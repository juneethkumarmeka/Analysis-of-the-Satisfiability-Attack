module basic_2000_20000_2500_10_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_767,In_409);
nand U1 (N_1,In_591,In_1651);
and U2 (N_2,In_1959,In_929);
and U3 (N_3,In_666,In_635);
nand U4 (N_4,In_489,In_320);
or U5 (N_5,In_382,In_1967);
and U6 (N_6,In_1220,In_1629);
nor U7 (N_7,In_1936,In_1970);
or U8 (N_8,In_1775,In_1460);
nand U9 (N_9,In_1957,In_390);
nand U10 (N_10,In_85,In_612);
or U11 (N_11,In_562,In_945);
and U12 (N_12,In_777,In_1781);
nand U13 (N_13,In_1178,In_810);
or U14 (N_14,In_616,In_374);
nand U15 (N_15,In_556,In_507);
nand U16 (N_16,In_1608,In_674);
nand U17 (N_17,In_903,In_1939);
nor U18 (N_18,In_1408,In_1848);
nand U19 (N_19,In_1382,In_1835);
nand U20 (N_20,In_1237,In_476);
and U21 (N_21,In_1779,In_1135);
and U22 (N_22,In_335,In_1155);
xor U23 (N_23,In_65,In_1963);
nor U24 (N_24,In_822,In_1710);
or U25 (N_25,In_8,In_1279);
nor U26 (N_26,In_1410,In_980);
nor U27 (N_27,In_1816,In_807);
and U28 (N_28,In_501,In_992);
and U29 (N_29,In_687,In_1977);
xor U30 (N_30,In_1482,In_1141);
xnor U31 (N_31,In_1873,In_1045);
or U32 (N_32,In_1513,In_473);
nor U33 (N_33,In_701,In_1298);
nand U34 (N_34,In_1769,In_295);
nand U35 (N_35,In_990,In_1346);
nor U36 (N_36,In_1707,In_716);
or U37 (N_37,In_1420,In_352);
or U38 (N_38,In_364,In_1744);
and U39 (N_39,In_1794,In_1945);
and U40 (N_40,In_289,In_1273);
or U41 (N_41,In_1789,In_244);
and U42 (N_42,In_1095,In_730);
and U43 (N_43,In_503,In_1714);
nor U44 (N_44,In_1191,In_1247);
xor U45 (N_45,In_422,In_359);
nand U46 (N_46,In_498,In_197);
and U47 (N_47,In_567,In_432);
and U48 (N_48,In_873,In_437);
xnor U49 (N_49,In_1209,In_392);
nor U50 (N_50,In_1469,In_1599);
nor U51 (N_51,In_1760,In_1260);
or U52 (N_52,In_494,In_1264);
or U53 (N_53,In_692,In_575);
and U54 (N_54,In_10,In_386);
nor U55 (N_55,In_1310,In_51);
nor U56 (N_56,In_1456,In_1948);
nand U57 (N_57,In_478,In_1767);
or U58 (N_58,In_54,In_1689);
nand U59 (N_59,In_1961,In_1532);
and U60 (N_60,In_869,In_7);
nor U61 (N_61,In_1227,In_310);
nor U62 (N_62,In_1242,In_319);
or U63 (N_63,In_1745,In_595);
or U64 (N_64,In_183,In_1907);
nor U65 (N_65,In_1331,In_754);
and U66 (N_66,In_1092,In_358);
and U67 (N_67,In_662,In_195);
nand U68 (N_68,In_941,In_1080);
nand U69 (N_69,In_632,In_1344);
or U70 (N_70,In_1366,In_761);
nor U71 (N_71,In_154,In_1684);
and U72 (N_72,In_337,In_203);
or U73 (N_73,In_1258,In_1069);
or U74 (N_74,In_1049,In_284);
or U75 (N_75,In_623,In_617);
and U76 (N_76,In_690,In_1051);
and U77 (N_77,In_1625,In_340);
and U78 (N_78,In_1859,In_1505);
or U79 (N_79,In_173,In_23);
nand U80 (N_80,In_238,In_518);
nand U81 (N_81,In_1063,In_1358);
nor U82 (N_82,In_539,In_1349);
or U83 (N_83,In_968,In_36);
nand U84 (N_84,In_1393,In_613);
or U85 (N_85,In_736,In_639);
nor U86 (N_86,In_469,In_788);
nor U87 (N_87,In_1960,In_893);
nor U88 (N_88,In_1971,In_651);
nor U89 (N_89,In_1404,In_144);
nor U90 (N_90,In_799,In_365);
xor U91 (N_91,In_520,In_830);
or U92 (N_92,In_78,In_574);
nand U93 (N_93,In_1206,In_602);
or U94 (N_94,In_1777,In_209);
nand U95 (N_95,In_544,In_738);
or U96 (N_96,In_1506,In_570);
and U97 (N_97,In_126,In_805);
nor U98 (N_98,In_845,In_1607);
and U99 (N_99,In_261,In_1475);
nand U100 (N_100,In_1565,In_69);
or U101 (N_101,In_668,In_649);
or U102 (N_102,In_673,In_491);
and U103 (N_103,In_1157,In_13);
nor U104 (N_104,In_418,In_597);
nor U105 (N_105,In_454,In_147);
and U106 (N_106,In_1337,In_1602);
and U107 (N_107,In_1172,In_1876);
xnor U108 (N_108,In_1706,In_973);
or U109 (N_109,In_603,In_578);
nand U110 (N_110,In_694,In_1418);
and U111 (N_111,In_447,In_633);
or U112 (N_112,In_940,In_908);
or U113 (N_113,In_317,In_224);
xnor U114 (N_114,In_379,In_1704);
or U115 (N_115,In_1234,In_1001);
nor U116 (N_116,In_551,In_824);
and U117 (N_117,In_1391,In_1383);
nand U118 (N_118,In_1664,In_555);
nor U119 (N_119,In_383,In_923);
and U120 (N_120,In_1119,In_1087);
or U121 (N_121,In_527,In_1526);
nand U122 (N_122,In_1484,In_506);
or U123 (N_123,In_1222,In_15);
nand U124 (N_124,In_1184,In_1831);
and U125 (N_125,In_1518,In_223);
and U126 (N_126,In_712,In_1660);
nor U127 (N_127,In_661,In_978);
nand U128 (N_128,In_1283,In_42);
and U129 (N_129,In_1177,In_1622);
nand U130 (N_130,In_168,In_1031);
nor U131 (N_131,In_1943,In_293);
nand U132 (N_132,In_466,In_1146);
and U133 (N_133,In_1500,In_1384);
and U134 (N_134,In_760,In_884);
and U135 (N_135,In_1009,In_1931);
or U136 (N_136,In_1200,In_142);
nand U137 (N_137,In_1357,In_324);
and U138 (N_138,In_1517,In_1807);
or U139 (N_139,In_1359,In_1373);
nand U140 (N_140,In_133,In_1604);
and U141 (N_141,In_667,In_1593);
or U142 (N_142,In_1034,In_637);
nor U143 (N_143,In_371,In_979);
and U144 (N_144,In_1434,In_937);
xor U145 (N_145,In_1403,In_1134);
or U146 (N_146,In_263,In_557);
or U147 (N_147,In_860,In_1474);
nand U148 (N_148,In_808,In_426);
or U149 (N_149,In_601,In_1730);
nand U150 (N_150,In_1309,In_1535);
and U151 (N_151,In_1569,In_160);
and U152 (N_152,In_1586,In_1877);
or U153 (N_153,In_1308,In_1468);
nor U154 (N_154,In_1056,In_172);
nor U155 (N_155,In_1496,In_1240);
nand U156 (N_156,In_1845,In_103);
xnor U157 (N_157,In_87,In_914);
nand U158 (N_158,In_1185,In_136);
or U159 (N_159,In_134,In_1100);
nand U160 (N_160,In_1552,In_1832);
xnor U161 (N_161,In_825,In_1296);
nor U162 (N_162,In_883,In_1551);
nor U163 (N_163,In_288,In_1052);
and U164 (N_164,In_823,In_746);
nor U165 (N_165,In_1720,In_1759);
nand U166 (N_166,In_151,In_1252);
nor U167 (N_167,In_1736,In_959);
nand U168 (N_168,In_786,In_1536);
or U169 (N_169,In_1028,In_1435);
nor U170 (N_170,In_975,In_1504);
nor U171 (N_171,In_1892,In_1508);
nand U172 (N_172,In_1424,In_566);
nand U173 (N_173,In_176,In_1840);
and U174 (N_174,In_1596,In_954);
and U175 (N_175,In_1074,In_251);
and U176 (N_176,In_1006,In_1020);
and U177 (N_177,In_1094,In_545);
nor U178 (N_178,In_665,In_1091);
or U179 (N_179,In_1969,In_486);
and U180 (N_180,In_707,In_1523);
and U181 (N_181,In_855,In_622);
or U182 (N_182,In_826,In_1849);
or U183 (N_183,In_1437,In_972);
or U184 (N_184,In_1464,In_983);
nor U185 (N_185,In_1547,In_888);
and U186 (N_186,In_113,In_107);
nor U187 (N_187,In_1335,In_1472);
and U188 (N_188,In_563,In_748);
nand U189 (N_189,In_47,In_170);
nand U190 (N_190,In_1495,In_419);
nor U191 (N_191,In_993,In_842);
nand U192 (N_192,In_1046,In_726);
xor U193 (N_193,In_309,In_119);
nand U194 (N_194,In_1215,In_1295);
or U195 (N_195,In_643,In_1639);
nor U196 (N_196,In_1755,In_1594);
nor U197 (N_197,In_1619,In_525);
nand U198 (N_198,In_408,In_453);
nand U199 (N_199,In_82,In_1365);
and U200 (N_200,In_1057,In_1966);
nor U201 (N_201,In_1728,In_1581);
or U202 (N_202,In_863,In_1617);
or U203 (N_203,In_833,In_262);
nand U204 (N_204,In_307,In_1842);
nor U205 (N_205,In_861,In_1114);
nor U206 (N_206,In_868,In_1352);
and U207 (N_207,In_135,In_1478);
nand U208 (N_208,In_225,In_1269);
nor U209 (N_209,In_5,In_179);
nand U210 (N_210,In_771,In_200);
or U211 (N_211,In_1897,In_1214);
nor U212 (N_212,In_1463,In_228);
nand U213 (N_213,In_129,In_1868);
nor U214 (N_214,In_1585,In_1803);
nand U215 (N_215,In_155,In_118);
or U216 (N_216,In_1400,In_290);
or U217 (N_217,In_1567,In_334);
nor U218 (N_218,In_1138,In_583);
and U219 (N_219,In_43,In_1187);
xnor U220 (N_220,In_1681,In_862);
nor U221 (N_221,In_1787,In_1224);
nand U222 (N_222,In_731,In_1678);
xnor U223 (N_223,In_504,In_1368);
and U224 (N_224,In_1416,In_1905);
xnor U225 (N_225,In_1415,In_30);
or U226 (N_226,In_1275,In_349);
or U227 (N_227,In_215,In_1053);
and U228 (N_228,In_894,In_721);
nand U229 (N_229,In_218,In_1439);
xor U230 (N_230,In_1205,In_360);
nand U231 (N_231,In_1661,In_165);
and U232 (N_232,In_1989,In_326);
nor U233 (N_233,In_306,In_363);
and U234 (N_234,In_483,In_400);
and U235 (N_235,In_158,In_1350);
and U236 (N_236,In_1659,In_1915);
and U237 (N_237,In_1412,In_531);
nand U238 (N_238,In_1318,In_1705);
and U239 (N_239,In_1904,In_373);
nand U240 (N_240,In_265,In_281);
nand U241 (N_241,In_161,In_1727);
or U242 (N_242,In_287,In_121);
nor U243 (N_243,In_1211,In_1314);
nand U244 (N_244,In_1498,In_1540);
and U245 (N_245,In_1733,In_1646);
and U246 (N_246,In_177,In_1583);
and U247 (N_247,In_267,In_401);
nor U248 (N_248,In_790,In_1159);
or U249 (N_249,In_76,In_1070);
nor U250 (N_250,In_272,In_21);
or U251 (N_251,In_615,In_528);
nand U252 (N_252,In_1324,In_598);
nand U253 (N_253,In_680,In_384);
and U254 (N_254,In_84,In_1470);
or U255 (N_255,In_770,In_977);
or U256 (N_256,In_485,In_463);
nor U257 (N_257,In_40,In_1347);
nor U258 (N_258,In_1255,In_96);
and U259 (N_259,In_1043,In_1993);
or U260 (N_260,In_1485,In_175);
nand U261 (N_261,In_1548,In_624);
xnor U262 (N_262,In_1825,In_1142);
nor U263 (N_263,In_1718,In_205);
nand U264 (N_264,In_459,In_111);
or U265 (N_265,In_1683,In_1738);
or U266 (N_266,In_604,In_282);
nand U267 (N_267,In_573,In_1562);
and U268 (N_268,In_547,In_1154);
and U269 (N_269,In_318,In_1898);
nand U270 (N_270,In_41,In_1951);
and U271 (N_271,In_1711,In_982);
nor U272 (N_272,In_1044,In_1919);
or U273 (N_273,In_1492,In_1797);
and U274 (N_274,In_369,In_1509);
or U275 (N_275,In_156,In_462);
nor U276 (N_276,In_1770,In_1407);
nand U277 (N_277,In_1421,In_1641);
and U278 (N_278,In_776,In_1870);
nand U279 (N_279,In_1988,In_211);
nand U280 (N_280,In_208,In_321);
and U281 (N_281,In_1457,In_377);
and U282 (N_282,In_875,In_339);
and U283 (N_283,In_1144,In_1979);
nor U284 (N_284,In_853,In_513);
or U285 (N_285,In_682,In_895);
xnor U286 (N_286,In_653,In_803);
and U287 (N_287,In_1944,In_274);
or U288 (N_288,In_782,In_468);
nand U289 (N_289,In_750,In_493);
nor U290 (N_290,In_1894,In_919);
or U291 (N_291,In_1522,In_1000);
or U292 (N_292,In_1941,In_1927);
nor U293 (N_293,In_1558,In_1645);
or U294 (N_294,In_542,In_1062);
nor U295 (N_295,In_1477,In_1232);
nand U296 (N_296,In_1414,In_1857);
nand U297 (N_297,In_74,In_1174);
and U298 (N_298,In_943,In_1731);
nand U299 (N_299,In_1480,In_1630);
nand U300 (N_300,In_1942,In_1925);
xnor U301 (N_301,In_1820,In_62);
nor U302 (N_302,In_1409,In_1102);
and U303 (N_303,In_32,In_193);
and U304 (N_304,In_204,In_1022);
nand U305 (N_305,In_343,In_1940);
nor U306 (N_306,In_1671,In_1503);
or U307 (N_307,In_1003,In_124);
xor U308 (N_308,In_1603,In_549);
nand U309 (N_309,In_350,In_458);
nand U310 (N_310,In_45,In_227);
or U311 (N_311,In_1106,In_98);
nand U312 (N_312,In_187,In_1766);
nor U313 (N_313,In_1918,In_210);
or U314 (N_314,In_1589,In_81);
or U315 (N_315,In_1855,In_735);
or U316 (N_316,In_1725,In_1345);
or U317 (N_317,In_588,In_564);
nor U318 (N_318,In_38,In_1489);
xnor U319 (N_319,In_778,In_1454);
nand U320 (N_320,In_1648,In_660);
or U321 (N_321,In_1542,In_471);
nor U322 (N_322,In_1635,In_97);
nor U323 (N_323,In_1124,In_792);
nand U324 (N_324,In_440,In_428);
or U325 (N_325,In_1566,In_1574);
or U326 (N_326,In_902,In_1348);
and U327 (N_327,In_681,In_1371);
nor U328 (N_328,In_715,In_1246);
or U329 (N_329,In_857,In_756);
or U330 (N_330,In_344,In_934);
nand U331 (N_331,In_1757,In_1055);
nor U332 (N_332,In_68,In_802);
xnor U333 (N_333,In_1018,In_609);
nand U334 (N_334,In_691,In_1427);
xor U335 (N_335,In_1450,In_877);
and U336 (N_336,In_1294,In_512);
and U337 (N_337,In_1229,In_1624);
nand U338 (N_338,In_1061,In_446);
and U339 (N_339,In_1101,In_37);
nor U340 (N_340,In_1890,In_734);
or U341 (N_341,In_1342,In_896);
nand U342 (N_342,In_449,In_693);
or U343 (N_343,In_1361,In_83);
xor U344 (N_344,In_890,In_1701);
and U345 (N_345,In_804,In_785);
or U346 (N_346,In_728,In_1654);
and U347 (N_347,In_1192,In_1559);
and U348 (N_348,In_1809,In_1375);
or U349 (N_349,In_232,In_850);
nand U350 (N_350,In_1013,In_1036);
or U351 (N_351,In_487,In_640);
and U352 (N_352,In_1311,In_559);
or U353 (N_353,In_137,In_216);
nand U354 (N_354,In_477,In_749);
and U355 (N_355,In_1529,In_672);
nor U356 (N_356,In_275,In_1449);
nand U357 (N_357,In_1600,In_387);
or U358 (N_358,In_1732,In_26);
nor U359 (N_359,In_380,In_1486);
nor U360 (N_360,In_904,In_1182);
nand U361 (N_361,In_429,In_72);
nand U362 (N_362,In_184,In_140);
nor U363 (N_363,In_152,In_1323);
nand U364 (N_364,In_1441,In_1995);
or U365 (N_365,In_61,In_1568);
xor U366 (N_366,In_565,In_354);
and U367 (N_367,In_273,In_1726);
nand U368 (N_368,In_733,In_519);
and U369 (N_369,In_55,In_546);
nor U370 (N_370,In_398,In_1555);
nand U371 (N_371,In_1886,In_296);
nand U372 (N_372,In_1634,In_1268);
and U373 (N_373,In_724,In_457);
or U374 (N_374,In_159,In_727);
nand U375 (N_375,In_592,In_1098);
xnor U376 (N_376,In_1047,In_912);
nor U377 (N_377,In_1306,In_1379);
nand U378 (N_378,In_1316,In_655);
and U379 (N_379,In_347,In_1871);
nor U380 (N_380,In_25,In_1204);
and U381 (N_381,In_1453,In_806);
and U382 (N_382,In_404,In_264);
and U383 (N_383,In_1016,In_1148);
xor U384 (N_384,In_1673,In_1773);
and U385 (N_385,In_1538,In_164);
nor U386 (N_386,In_1032,In_1367);
nand U387 (N_387,In_1244,In_1920);
nand U388 (N_388,In_663,In_817);
nand U389 (N_389,In_1992,In_259);
and U390 (N_390,In_1914,In_303);
nor U391 (N_391,In_106,In_571);
xnor U392 (N_392,In_241,In_743);
or U393 (N_393,In_1025,In_757);
xor U394 (N_394,In_798,In_679);
nor U395 (N_395,In_1436,In_1329);
nor U396 (N_396,In_1395,In_1241);
or U397 (N_397,In_1813,In_1462);
or U398 (N_398,In_1362,In_1642);
and U399 (N_399,In_255,In_1837);
and U400 (N_400,In_766,In_412);
nand U401 (N_401,In_1690,In_1250);
nand U402 (N_402,In_1280,In_1854);
and U403 (N_403,In_1259,In_1413);
or U404 (N_404,In_1734,In_1428);
and U405 (N_405,In_719,In_1067);
and U406 (N_406,In_327,In_1133);
nand U407 (N_407,In_1131,In_372);
or U408 (N_408,In_634,In_590);
nor U409 (N_409,In_1388,In_1029);
nand U410 (N_410,In_816,In_1305);
nor U411 (N_411,In_1719,In_1929);
or U412 (N_412,In_1411,In_201);
or U413 (N_413,In_787,In_1010);
nand U414 (N_414,In_1686,In_1334);
xor U415 (N_415,In_1312,In_1111);
and U416 (N_416,In_718,In_1355);
nor U417 (N_417,In_758,In_396);
or U418 (N_418,In_587,In_1390);
nand U419 (N_419,In_14,In_285);
or U420 (N_420,In_1923,In_1994);
xor U421 (N_421,In_252,In_191);
nand U422 (N_422,In_1169,In_219);
nor U423 (N_423,In_1575,In_509);
and U424 (N_424,In_948,In_1628);
and U425 (N_425,In_1483,In_1560);
xor U426 (N_426,In_1088,In_1175);
or U427 (N_427,In_844,In_190);
xor U428 (N_428,In_451,In_1153);
or U429 (N_429,In_1953,In_1805);
nor U430 (N_430,In_1399,In_1442);
nor U431 (N_431,In_1861,In_636);
nand U432 (N_432,In_1601,In_1328);
and U433 (N_433,In_1151,In_351);
or U434 (N_434,In_521,In_951);
and U435 (N_435,In_1254,In_1790);
xnor U436 (N_436,In_1620,In_1064);
or U437 (N_437,In_964,In_1037);
nor U438 (N_438,In_942,In_1864);
and U439 (N_439,In_1039,In_1702);
or U440 (N_440,In_1251,In_6);
nor U441 (N_441,In_648,In_1949);
xor U442 (N_442,In_1458,In_773);
nor U443 (N_443,In_93,In_1297);
and U444 (N_444,In_1377,In_759);
nor U445 (N_445,In_1054,In_1221);
nand U446 (N_446,In_314,In_530);
and U447 (N_447,In_28,In_1613);
nand U448 (N_448,In_646,In_969);
or U449 (N_449,In_1721,In_1595);
nand U450 (N_450,In_1304,In_866);
nor U451 (N_451,In_1360,In_811);
nand U452 (N_452,In_1655,In_1461);
nand U453 (N_453,In_809,In_797);
or U454 (N_454,In_1207,In_1007);
nor U455 (N_455,In_926,In_1746);
nor U456 (N_456,In_812,In_268);
nand U457 (N_457,In_801,In_417);
xnor U458 (N_458,In_461,In_465);
nor U459 (N_459,In_253,In_1445);
or U460 (N_460,In_77,In_1627);
and U461 (N_461,In_138,In_901);
nor U462 (N_462,In_1539,In_1479);
nand U463 (N_463,In_1005,In_1791);
nor U464 (N_464,In_1193,In_1014);
xor U465 (N_465,In_1433,In_1672);
and U466 (N_466,In_435,In_669);
nor U467 (N_467,In_146,In_1911);
and U468 (N_468,In_1800,In_772);
or U469 (N_469,In_558,In_1670);
nand U470 (N_470,In_1370,In_472);
and U471 (N_471,In_1423,In_952);
nand U472 (N_472,In_1156,In_1932);
nand U473 (N_473,In_1011,In_1652);
or U474 (N_474,In_1570,In_153);
nor U475 (N_475,In_1285,In_1287);
nor U476 (N_476,In_415,In_1120);
and U477 (N_477,In_1112,In_20);
nor U478 (N_478,In_1071,In_1284);
nor U479 (N_479,In_935,In_34);
nor U480 (N_480,In_90,In_876);
nand U481 (N_481,In_1050,In_1997);
nand U482 (N_482,In_552,In_1851);
nand U483 (N_483,In_171,In_927);
nor U484 (N_484,In_856,In_1606);
and U485 (N_485,In_357,In_1369);
nand U486 (N_486,In_66,In_1818);
or U487 (N_487,In_182,In_105);
nand U488 (N_488,In_1687,In_246);
nor U489 (N_489,In_385,In_741);
nor U490 (N_490,In_95,In_517);
nor U491 (N_491,In_596,In_600);
xor U492 (N_492,In_1650,In_1465);
xor U493 (N_493,In_1165,In_1040);
or U494 (N_494,In_832,In_1616);
nor U495 (N_495,In_481,In_1860);
or U496 (N_496,In_1924,In_995);
xor U497 (N_497,In_1888,In_774);
and U498 (N_498,In_925,In_1900);
nand U499 (N_499,In_1667,In_1700);
nand U500 (N_500,In_819,In_1179);
xor U501 (N_501,In_1488,In_924);
nor U502 (N_502,In_1947,In_515);
nand U503 (N_503,In_526,In_254);
or U504 (N_504,In_353,In_1722);
and U505 (N_505,In_1196,In_1743);
nor U506 (N_506,In_1965,In_1307);
and U507 (N_507,In_112,In_1521);
nor U508 (N_508,In_1230,In_1983);
or U509 (N_509,In_831,In_720);
and U510 (N_510,In_1163,In_12);
or U511 (N_511,In_1303,In_710);
xnor U512 (N_512,In_1398,In_405);
or U513 (N_513,In_73,In_1389);
nand U514 (N_514,In_1822,In_394);
and U515 (N_515,In_1281,In_1881);
or U516 (N_516,In_243,In_965);
and U517 (N_517,In_294,In_1249);
xnor U518 (N_518,In_1459,In_420);
or U519 (N_519,In_1293,In_1257);
nand U520 (N_520,In_1060,In_442);
and U521 (N_521,In_1194,In_706);
nor U522 (N_522,In_11,In_1024);
and U523 (N_523,In_186,In_207);
nor U524 (N_524,In_1161,In_1181);
and U525 (N_525,In_560,In_199);
or U526 (N_526,In_697,In_1691);
xor U527 (N_527,In_1109,In_611);
xor U528 (N_528,In_703,In_791);
or U529 (N_529,In_279,In_1615);
or U530 (N_530,In_1272,In_1330);
nor U531 (N_531,In_448,In_1675);
or U532 (N_532,In_1836,In_52);
nor U533 (N_533,In_577,In_441);
or U534 (N_534,In_108,In_1662);
or U535 (N_535,In_1072,In_1282);
xnor U536 (N_536,In_986,In_1089);
nor U537 (N_537,In_70,In_322);
or U538 (N_538,In_508,In_86);
nand U539 (N_539,In_1231,In_1802);
nand U540 (N_540,In_1640,In_920);
and U541 (N_541,In_899,In_242);
and U542 (N_542,In_331,In_1985);
nand U543 (N_543,In_533,In_538);
nand U544 (N_544,In_915,In_1592);
or U545 (N_545,In_657,In_2);
and U546 (N_546,In_1129,In_1618);
and U547 (N_547,In_1397,In_536);
nand U548 (N_548,In_1841,In_921);
nand U549 (N_549,In_936,In_1288);
nand U550 (N_550,In_452,In_1128);
or U551 (N_551,In_828,In_1333);
and U552 (N_552,In_714,In_416);
and U553 (N_553,In_328,In_411);
nand U554 (N_554,In_1019,In_1874);
and U555 (N_555,In_897,In_1545);
xnor U556 (N_556,In_1756,In_1846);
nor U557 (N_557,In_234,In_1497);
or U558 (N_558,In_1866,In_1764);
nand U559 (N_559,In_1754,In_1440);
and U560 (N_560,In_1833,In_1783);
and U561 (N_561,In_984,In_864);
and U562 (N_562,In_1826,In_654);
and U563 (N_563,In_1956,In_1422);
and U564 (N_564,In_188,In_614);
nor U565 (N_565,In_1811,In_1235);
xor U566 (N_566,In_1499,In_1170);
xnor U567 (N_567,In_1916,In_849);
and U568 (N_568,In_1302,In_367);
and U569 (N_569,In_747,In_1238);
or U570 (N_570,In_1315,In_1203);
or U571 (N_571,In_399,In_1784);
nor U572 (N_572,In_676,In_56);
and U573 (N_573,In_1557,In_887);
nand U574 (N_574,In_149,In_1313);
xnor U575 (N_575,In_1612,In_1819);
or U576 (N_576,In_1998,In_1685);
xnor U577 (N_577,In_1276,In_1609);
and U578 (N_578,In_1336,In_495);
or U579 (N_579,In_1473,In_480);
nor U580 (N_580,In_572,In_389);
or U581 (N_581,In_704,In_1210);
and U582 (N_582,In_16,In_301);
nand U583 (N_583,In_1341,In_9);
nand U584 (N_584,In_346,In_1443);
and U585 (N_585,In_258,In_1748);
or U586 (N_586,In_1708,In_1082);
nand U587 (N_587,In_532,In_239);
or U588 (N_588,In_641,In_1248);
xnor U589 (N_589,In_820,In_1038);
and U590 (N_590,In_568,In_342);
or U591 (N_591,In_1021,In_966);
and U592 (N_592,In_125,In_325);
and U593 (N_593,In_1623,In_996);
nand U594 (N_594,In_554,In_1137);
nand U595 (N_595,In_1208,In_167);
and U596 (N_596,In_1632,In_214);
and U597 (N_597,In_1768,In_1115);
nand U598 (N_598,In_605,In_1083);
nand U599 (N_599,In_1564,In_67);
and U600 (N_600,In_1017,In_256);
or U601 (N_601,In_1649,In_330);
nor U602 (N_602,In_49,In_762);
nor U603 (N_603,In_768,In_764);
nand U604 (N_604,In_1213,In_1875);
xnor U605 (N_605,In_1263,In_514);
and U606 (N_606,In_939,In_1059);
or U607 (N_607,In_1584,In_395);
xnor U608 (N_608,In_769,In_950);
and U609 (N_609,In_1834,In_874);
and U610 (N_610,In_1002,In_1147);
xor U611 (N_611,In_1527,In_1189);
xnor U612 (N_612,In_576,In_64);
nand U613 (N_613,In_1225,In_625);
or U614 (N_614,In_1127,In_230);
and U615 (N_615,In_1188,In_1891);
nor U616 (N_616,In_1430,In_1090);
xnor U617 (N_617,In_1494,In_1110);
nor U618 (N_618,In_953,In_425);
and U619 (N_619,In_961,In_92);
and U620 (N_620,In_1317,In_928);
nand U621 (N_621,In_1952,In_375);
nand U622 (N_622,In_1626,In_291);
nor U623 (N_623,In_599,In_523);
and U624 (N_624,In_742,In_1113);
and U625 (N_625,In_304,In_245);
xnor U626 (N_626,In_276,In_1872);
nor U627 (N_627,In_198,In_1325);
or U628 (N_628,In_1405,In_629);
xor U629 (N_629,In_17,In_713);
or U630 (N_630,In_1528,In_1291);
nor U631 (N_631,In_1270,In_1962);
nor U632 (N_632,In_407,In_1116);
nand U633 (N_633,In_450,In_886);
nor U634 (N_634,In_388,In_1909);
or U635 (N_635,In_102,In_1973);
nand U636 (N_636,In_1493,In_194);
nor U637 (N_637,In_932,In_1954);
and U638 (N_638,In_1561,In_1955);
nand U639 (N_639,In_1885,In_455);
nand U640 (N_640,In_795,In_1878);
and U641 (N_641,In_581,In_413);
nand U642 (N_642,In_1902,In_48);
xor U643 (N_643,In_1598,In_222);
or U644 (N_644,In_286,In_967);
and U645 (N_645,In_1798,In_1879);
and U646 (N_646,In_1321,In_579);
or U647 (N_647,In_628,In_427);
and U648 (N_648,In_1197,In_1926);
nand U649 (N_649,In_115,In_1201);
nor U650 (N_650,In_1749,In_1814);
nand U651 (N_651,In_1326,In_439);
and U652 (N_652,In_789,In_482);
nor U653 (N_653,In_841,In_192);
and U654 (N_654,In_1406,In_740);
or U655 (N_655,In_744,In_44);
nor U656 (N_656,In_499,In_702);
and U657 (N_657,In_1130,In_1621);
nand U658 (N_658,In_1804,In_89);
nand U659 (N_659,In_1827,In_700);
nand U660 (N_660,In_33,In_406);
nor U661 (N_661,In_166,In_1740);
or U662 (N_662,In_431,In_1858);
nor U663 (N_663,In_1431,In_1402);
and U664 (N_664,In_882,In_835);
and U665 (N_665,In_1162,In_178);
xor U666 (N_666,In_970,In_1446);
and U667 (N_667,In_1647,In_794);
nand U668 (N_668,In_1265,In_1578);
and U669 (N_669,In_836,In_1644);
nor U670 (N_670,In_1741,In_907);
and U671 (N_671,In_670,In_1742);
xor U672 (N_672,In_619,In_1356);
or U673 (N_673,In_582,In_779);
nand U674 (N_674,In_479,In_1844);
nor U675 (N_675,In_1928,In_1572);
nor U676 (N_676,In_1363,In_708);
nor U677 (N_677,In_280,In_1202);
and U678 (N_678,In_1739,In_1103);
and U679 (N_679,In_1553,In_341);
and U680 (N_680,In_626,In_1880);
or U681 (N_681,In_1636,In_1125);
nand U682 (N_682,In_27,In_421);
nor U683 (N_683,In_1376,In_104);
nor U684 (N_684,In_1587,In_1448);
nor U685 (N_685,In_1893,In_316);
nor U686 (N_686,In_561,In_467);
nor U687 (N_687,In_1763,In_1081);
nand U688 (N_688,In_537,In_1218);
and U689 (N_689,In_813,In_1066);
nor U690 (N_690,In_1392,In_1550);
nand U691 (N_691,In_127,In_956);
xnor U692 (N_692,In_445,In_1847);
or U693 (N_693,In_58,In_1882);
and U694 (N_694,In_586,In_236);
nor U695 (N_695,In_1981,In_658);
nand U696 (N_696,In_955,In_1676);
nor U697 (N_697,In_909,In_1571);
nor U698 (N_698,In_1516,In_1502);
nor U699 (N_699,In_1663,In_1674);
xor U700 (N_700,In_206,In_1788);
or U701 (N_701,In_283,In_1507);
nand U702 (N_702,In_765,In_1190);
xor U703 (N_703,In_918,In_1515);
xor U704 (N_704,In_1709,In_644);
nor U705 (N_705,In_1030,In_297);
nor U706 (N_706,In_717,In_838);
or U707 (N_707,In_196,In_1577);
or U708 (N_708,In_755,In_647);
nand U709 (N_709,In_821,In_1758);
or U710 (N_710,In_610,In_148);
nand U711 (N_711,In_510,In_1590);
nor U712 (N_712,In_1580,In_594);
nand U713 (N_713,In_1253,In_300);
and U714 (N_714,In_1139,In_1481);
nor U715 (N_715,In_1968,In_618);
nand U716 (N_716,In_1152,In_430);
and U717 (N_717,In_1656,In_1896);
nor U718 (N_718,In_1058,In_298);
nand U719 (N_719,In_695,In_1150);
nor U720 (N_720,In_645,In_139);
nor U721 (N_721,In_851,In_1982);
nor U722 (N_722,In_550,In_1122);
xor U723 (N_723,In_22,In_505);
and U724 (N_724,In_997,In_699);
nor U725 (N_725,In_1554,In_1394);
nor U726 (N_726,In_891,In_516);
and U727 (N_727,In_683,In_638);
nor U728 (N_728,In_723,In_858);
nor U729 (N_729,In_783,In_410);
or U730 (N_730,In_109,In_1104);
xor U731 (N_731,In_994,In_248);
nand U732 (N_732,In_827,In_345);
or U733 (N_733,In_1117,In_57);
nor U734 (N_734,In_1912,In_1934);
and U735 (N_735,In_75,In_145);
or U736 (N_736,In_88,In_35);
nand U737 (N_737,In_1300,In_308);
nor U738 (N_738,In_686,In_1697);
and U739 (N_739,In_1793,In_366);
nand U740 (N_740,In_1319,In_0);
nor U741 (N_741,In_889,In_1986);
nand U742 (N_742,In_910,In_1380);
xnor U743 (N_743,In_1476,In_50);
xor U744 (N_744,In_711,In_689);
and U745 (N_745,In_684,In_229);
xor U746 (N_746,In_1863,In_1677);
or U747 (N_747,In_745,In_1703);
nand U748 (N_748,In_116,In_991);
nor U749 (N_749,In_475,In_1716);
or U750 (N_750,In_502,In_424);
nand U751 (N_751,In_1320,In_1136);
nor U752 (N_752,In_585,In_233);
nor U753 (N_753,In_1865,In_260);
or U754 (N_754,In_329,In_1444);
or U755 (N_755,In_1027,In_1695);
or U756 (N_756,In_620,In_1883);
xnor U757 (N_757,In_217,In_1533);
or U758 (N_758,In_698,In_266);
nor U759 (N_759,In_1212,In_313);
and U760 (N_760,In_123,In_1901);
and U761 (N_761,In_739,In_608);
nand U762 (N_762,In_403,In_971);
xnor U763 (N_763,In_793,In_1862);
nand U764 (N_764,In_859,In_163);
xor U765 (N_765,In_212,In_1668);
and U766 (N_766,In_947,In_1167);
nand U767 (N_767,In_497,In_1610);
nand U768 (N_768,In_1729,In_1289);
and U769 (N_769,In_1747,In_31);
and U770 (N_770,In_1354,In_299);
nand U771 (N_771,In_1810,In_1750);
nand U772 (N_772,In_1830,In_1723);
or U773 (N_773,In_652,In_580);
or U774 (N_774,In_181,In_1339);
and U775 (N_775,In_240,In_100);
and U776 (N_776,In_725,In_1353);
xnor U777 (N_777,In_1277,In_1935);
or U778 (N_778,In_470,In_751);
and U779 (N_779,In_916,In_1591);
nand U780 (N_780,In_1543,In_1198);
or U781 (N_781,In_1950,In_1824);
nand U782 (N_782,In_1605,In_1682);
nand U783 (N_783,In_1512,In_1614);
and U784 (N_784,In_18,In_1823);
or U785 (N_785,In_1765,In_1075);
nor U786 (N_786,In_1236,In_226);
nor U787 (N_787,In_524,In_664);
xnor U788 (N_788,In_333,In_1762);
and U789 (N_789,In_1519,In_370);
or U790 (N_790,In_99,In_1843);
nor U791 (N_791,In_593,In_933);
nand U792 (N_792,In_1853,In_1364);
and U793 (N_793,In_987,In_1712);
or U794 (N_794,In_1425,In_1829);
and U795 (N_795,In_946,In_1869);
or U796 (N_796,In_906,In_356);
xor U797 (N_797,In_132,In_117);
nand U798 (N_798,In_1980,In_444);
and U799 (N_799,In_311,In_1799);
nor U800 (N_800,In_436,In_650);
or U801 (N_801,In_1839,In_110);
nand U802 (N_802,In_1176,In_362);
or U803 (N_803,In_627,In_361);
nor U804 (N_804,In_1597,In_1077);
xnor U805 (N_805,In_91,In_1821);
or U806 (N_806,In_1501,In_1);
nor U807 (N_807,In_94,In_1796);
nor U808 (N_808,In_1817,In_1976);
and U809 (N_809,In_705,In_1772);
or U810 (N_810,In_1713,In_292);
nor U811 (N_811,In_535,In_1452);
nand U812 (N_812,In_397,In_180);
nand U813 (N_813,In_917,In_202);
nand U814 (N_814,In_589,In_606);
and U815 (N_815,In_1160,In_1999);
xor U816 (N_816,In_957,In_985);
nand U817 (N_817,In_1401,In_1537);
nand U818 (N_818,In_1262,In_302);
nor U819 (N_819,In_931,In_250);
nor U820 (N_820,In_220,In_1266);
nand U821 (N_821,In_1785,In_938);
or U822 (N_822,In_1573,In_511);
nand U823 (N_823,In_1491,In_277);
or U824 (N_824,In_1079,In_39);
nand U825 (N_825,In_1372,In_1340);
nand U826 (N_826,In_840,In_1033);
or U827 (N_827,In_930,In_753);
and U828 (N_828,In_213,In_922);
or U829 (N_829,In_1026,In_1693);
or U830 (N_830,In_1556,In_114);
nand U831 (N_831,In_1381,In_722);
nor U832 (N_832,In_1426,In_732);
and U833 (N_833,In_1078,In_999);
or U834 (N_834,In_843,In_1895);
nand U835 (N_835,In_185,In_553);
nor U836 (N_836,In_269,In_150);
or U837 (N_837,In_1447,In_131);
or U838 (N_838,In_1261,In_1068);
nand U839 (N_839,In_780,In_1549);
nand U840 (N_840,In_529,In_128);
nand U841 (N_841,In_1653,In_1815);
nand U842 (N_842,In_1085,In_1908);
nor U843 (N_843,In_847,In_1086);
nor U844 (N_844,In_1884,In_1806);
nor U845 (N_845,In_1735,In_490);
nand U846 (N_846,In_355,In_141);
or U847 (N_847,In_913,In_1917);
nand U848 (N_848,In_1699,In_659);
xor U849 (N_849,In_443,In_1158);
or U850 (N_850,In_900,In_1792);
nor U851 (N_851,In_60,In_305);
nor U852 (N_852,In_1530,In_1987);
nor U853 (N_853,In_1795,In_737);
nand U854 (N_854,In_1145,In_162);
xor U855 (N_855,In_870,In_878);
nor U856 (N_856,In_1972,In_543);
and U857 (N_857,In_278,In_839);
nand U858 (N_858,In_1301,In_1171);
xor U859 (N_859,In_1808,In_1715);
nand U860 (N_860,In_414,In_1899);
nand U861 (N_861,In_1121,In_834);
and U862 (N_862,In_378,In_974);
nor U863 (N_863,In_976,In_1267);
or U864 (N_864,In_1338,In_880);
nand U865 (N_865,In_871,In_1782);
and U866 (N_866,In_1937,In_630);
nand U867 (N_867,In_1611,In_53);
nor U868 (N_868,In_1217,In_1698);
and U869 (N_869,In_1633,In_423);
nand U870 (N_870,In_1576,In_1271);
nor U871 (N_871,In_1780,In_1933);
nor U872 (N_872,In_1451,In_1097);
xor U873 (N_873,In_1012,In_1694);
and U874 (N_874,In_1386,In_1910);
nor U875 (N_875,In_221,In_1657);
xor U876 (N_876,In_892,In_24);
and U877 (N_877,In_784,In_885);
nor U878 (N_878,In_1374,In_642);
nand U879 (N_879,In_818,In_1471);
and U880 (N_880,In_752,In_949);
or U881 (N_881,In_1256,In_1290);
nand U882 (N_882,In_231,In_1186);
nor U883 (N_883,In_814,In_1867);
or U884 (N_884,In_675,In_1638);
or U885 (N_885,In_1990,In_1563);
xnor U886 (N_886,In_1974,In_1889);
nor U887 (N_887,In_1216,In_541);
nand U888 (N_888,In_1343,In_1076);
nor U889 (N_889,In_1938,In_1164);
or U890 (N_890,In_323,In_671);
nor U891 (N_891,In_1299,In_46);
or U892 (N_892,In_1432,In_898);
and U893 (N_893,In_1812,In_1510);
or U894 (N_894,In_1546,In_1438);
nor U895 (N_895,In_1008,In_962);
nor U896 (N_896,In_376,In_1455);
xor U897 (N_897,In_249,In_1579);
xor U898 (N_898,In_1093,In_1778);
nand U899 (N_899,In_19,In_998);
nor U900 (N_900,In_1351,In_1487);
nand U901 (N_901,In_101,In_846);
nor U902 (N_902,In_1042,In_1637);
nor U903 (N_903,In_1332,In_1233);
xor U904 (N_904,In_1761,In_338);
and U905 (N_905,In_1219,In_1099);
or U906 (N_906,In_696,In_1292);
nand U907 (N_907,In_1588,In_775);
nor U908 (N_908,In_500,In_460);
xnor U909 (N_909,In_79,In_1737);
nand U910 (N_910,In_800,In_1243);
and U911 (N_911,In_1525,In_402);
or U912 (N_912,In_71,In_1327);
and U913 (N_913,In_963,In_1239);
nand U914 (N_914,In_315,In_1922);
nand U915 (N_915,In_312,In_29);
nand U916 (N_916,In_368,In_1126);
nand U917 (N_917,In_631,In_1991);
nand U918 (N_918,In_1490,In_584);
or U919 (N_919,In_1887,In_1520);
or U920 (N_920,In_522,In_1168);
nand U921 (N_921,In_271,In_607);
nor U922 (N_922,In_1108,In_1511);
or U923 (N_923,In_1544,In_4);
or U924 (N_924,In_872,In_763);
and U925 (N_925,In_157,In_3);
xor U926 (N_926,In_1541,In_1669);
nor U927 (N_927,In_989,In_677);
nor U928 (N_928,In_1774,In_59);
or U929 (N_929,In_729,In_438);
or U930 (N_930,In_381,In_484);
and U931 (N_931,In_867,In_237);
xnor U932 (N_932,In_1679,In_247);
and U933 (N_933,In_1838,In_1226);
or U934 (N_934,In_1964,In_879);
nand U935 (N_935,In_1665,In_678);
nand U936 (N_936,In_656,In_1140);
nand U937 (N_937,In_1852,In_1771);
and U938 (N_938,In_685,In_1396);
or U939 (N_939,In_456,In_688);
nand U940 (N_940,In_911,In_1534);
or U941 (N_941,In_534,In_464);
nor U942 (N_942,In_1724,In_1048);
and U943 (N_943,In_1035,In_235);
nor U944 (N_944,In_474,In_434);
or U945 (N_945,In_1850,In_1696);
and U946 (N_946,In_1582,In_1322);
nor U947 (N_947,In_1913,In_332);
or U948 (N_948,In_1978,In_122);
nand U949 (N_949,In_1514,In_1996);
and U950 (N_950,In_1692,In_852);
nor U951 (N_951,In_540,In_1166);
nand U952 (N_952,In_1084,In_1751);
and U953 (N_953,In_169,In_1223);
nand U954 (N_954,In_1065,In_1387);
nor U955 (N_955,In_1105,In_960);
and U956 (N_956,In_1015,In_1975);
and U957 (N_957,In_1173,In_1776);
nor U958 (N_958,In_1274,In_1199);
or U959 (N_959,In_1419,In_1828);
or U960 (N_960,In_433,In_1073);
and U961 (N_961,In_1752,In_848);
nand U962 (N_962,In_1096,In_1004);
and U963 (N_963,In_1906,In_1195);
nor U964 (N_964,In_944,In_1023);
nand U965 (N_965,In_1688,In_1801);
nor U966 (N_966,In_1467,In_1856);
nor U967 (N_967,In_981,In_1531);
or U968 (N_968,In_1631,In_621);
nand U969 (N_969,In_1717,In_1524);
nor U970 (N_970,In_1107,In_1183);
or U971 (N_971,In_837,In_496);
and U972 (N_972,In_796,In_80);
or U973 (N_973,In_569,In_1041);
nor U974 (N_974,In_393,In_958);
xor U975 (N_975,In_829,In_1385);
nand U976 (N_976,In_130,In_1132);
xnor U977 (N_977,In_348,In_1149);
and U978 (N_978,In_1123,In_854);
or U979 (N_979,In_709,In_865);
nor U980 (N_980,In_815,In_1666);
and U981 (N_981,In_1118,In_1680);
nand U982 (N_982,In_1753,In_336);
or U983 (N_983,In_1378,In_1658);
xor U984 (N_984,In_174,In_120);
or U985 (N_985,In_63,In_391);
nand U986 (N_986,In_143,In_881);
and U987 (N_987,In_488,In_270);
or U988 (N_988,In_1466,In_1286);
nand U989 (N_989,In_1417,In_1429);
nor U990 (N_990,In_988,In_1786);
nor U991 (N_991,In_1143,In_1984);
nor U992 (N_992,In_1946,In_1930);
nand U993 (N_993,In_1245,In_1643);
nand U994 (N_994,In_189,In_257);
xor U995 (N_995,In_1278,In_1228);
and U996 (N_996,In_548,In_492);
or U997 (N_997,In_1921,In_905);
nor U998 (N_998,In_1903,In_1958);
or U999 (N_999,In_1180,In_781);
and U1000 (N_1000,In_1756,In_639);
or U1001 (N_1001,In_1303,In_1618);
nand U1002 (N_1002,In_1467,In_1487);
or U1003 (N_1003,In_364,In_354);
or U1004 (N_1004,In_1820,In_1525);
nor U1005 (N_1005,In_1152,In_53);
nand U1006 (N_1006,In_252,In_1027);
nor U1007 (N_1007,In_1873,In_1603);
or U1008 (N_1008,In_40,In_1764);
or U1009 (N_1009,In_1773,In_1202);
or U1010 (N_1010,In_1081,In_1436);
nand U1011 (N_1011,In_442,In_186);
nor U1012 (N_1012,In_92,In_1443);
or U1013 (N_1013,In_857,In_1498);
xor U1014 (N_1014,In_1226,In_731);
nand U1015 (N_1015,In_914,In_1899);
nor U1016 (N_1016,In_569,In_58);
nor U1017 (N_1017,In_1378,In_702);
and U1018 (N_1018,In_1128,In_1227);
xnor U1019 (N_1019,In_1654,In_725);
nor U1020 (N_1020,In_1377,In_218);
and U1021 (N_1021,In_550,In_386);
nand U1022 (N_1022,In_1338,In_1333);
nor U1023 (N_1023,In_166,In_1759);
nor U1024 (N_1024,In_929,In_1105);
nor U1025 (N_1025,In_87,In_1434);
or U1026 (N_1026,In_528,In_159);
and U1027 (N_1027,In_1541,In_1882);
xnor U1028 (N_1028,In_1837,In_1435);
and U1029 (N_1029,In_1095,In_657);
or U1030 (N_1030,In_1383,In_656);
and U1031 (N_1031,In_1094,In_1480);
and U1032 (N_1032,In_1536,In_927);
nor U1033 (N_1033,In_808,In_1881);
nand U1034 (N_1034,In_169,In_403);
nand U1035 (N_1035,In_1767,In_1967);
nand U1036 (N_1036,In_1817,In_801);
xor U1037 (N_1037,In_1228,In_840);
nand U1038 (N_1038,In_1321,In_877);
or U1039 (N_1039,In_539,In_82);
or U1040 (N_1040,In_620,In_1197);
and U1041 (N_1041,In_772,In_1008);
nor U1042 (N_1042,In_1056,In_1413);
and U1043 (N_1043,In_1987,In_249);
nor U1044 (N_1044,In_1392,In_96);
nor U1045 (N_1045,In_1154,In_1410);
nand U1046 (N_1046,In_928,In_1698);
nor U1047 (N_1047,In_307,In_1254);
or U1048 (N_1048,In_1484,In_40);
and U1049 (N_1049,In_520,In_883);
xnor U1050 (N_1050,In_1614,In_1228);
nor U1051 (N_1051,In_560,In_1213);
nand U1052 (N_1052,In_1102,In_1667);
and U1053 (N_1053,In_385,In_375);
xnor U1054 (N_1054,In_1025,In_1353);
and U1055 (N_1055,In_972,In_719);
or U1056 (N_1056,In_72,In_1678);
or U1057 (N_1057,In_1885,In_1077);
xnor U1058 (N_1058,In_797,In_156);
and U1059 (N_1059,In_1804,In_1967);
and U1060 (N_1060,In_129,In_609);
nand U1061 (N_1061,In_538,In_108);
or U1062 (N_1062,In_1644,In_1743);
or U1063 (N_1063,In_131,In_1252);
xnor U1064 (N_1064,In_1605,In_1228);
and U1065 (N_1065,In_513,In_494);
xnor U1066 (N_1066,In_449,In_1378);
nor U1067 (N_1067,In_1444,In_1305);
nor U1068 (N_1068,In_1816,In_749);
nor U1069 (N_1069,In_44,In_882);
nor U1070 (N_1070,In_737,In_1607);
nor U1071 (N_1071,In_1922,In_1693);
nand U1072 (N_1072,In_1236,In_1602);
nand U1073 (N_1073,In_335,In_738);
and U1074 (N_1074,In_301,In_1512);
or U1075 (N_1075,In_1420,In_1015);
nor U1076 (N_1076,In_491,In_1902);
nand U1077 (N_1077,In_1460,In_947);
nand U1078 (N_1078,In_626,In_1402);
nand U1079 (N_1079,In_1606,In_71);
nand U1080 (N_1080,In_196,In_1856);
nand U1081 (N_1081,In_11,In_1227);
xnor U1082 (N_1082,In_68,In_881);
nand U1083 (N_1083,In_59,In_1996);
or U1084 (N_1084,In_898,In_1093);
nor U1085 (N_1085,In_1929,In_1199);
or U1086 (N_1086,In_1767,In_883);
nor U1087 (N_1087,In_781,In_879);
xnor U1088 (N_1088,In_1353,In_1214);
and U1089 (N_1089,In_1403,In_1889);
or U1090 (N_1090,In_276,In_1236);
or U1091 (N_1091,In_202,In_934);
nand U1092 (N_1092,In_353,In_1394);
nand U1093 (N_1093,In_1912,In_763);
or U1094 (N_1094,In_1467,In_28);
nand U1095 (N_1095,In_1843,In_1348);
xnor U1096 (N_1096,In_1844,In_867);
nand U1097 (N_1097,In_1649,In_574);
or U1098 (N_1098,In_129,In_638);
or U1099 (N_1099,In_1975,In_407);
and U1100 (N_1100,In_1015,In_714);
nand U1101 (N_1101,In_1525,In_1211);
or U1102 (N_1102,In_581,In_465);
nand U1103 (N_1103,In_582,In_1193);
xnor U1104 (N_1104,In_943,In_1174);
or U1105 (N_1105,In_1128,In_123);
nand U1106 (N_1106,In_12,In_1580);
nor U1107 (N_1107,In_273,In_1596);
and U1108 (N_1108,In_1933,In_1554);
nor U1109 (N_1109,In_1391,In_1318);
nor U1110 (N_1110,In_1380,In_241);
or U1111 (N_1111,In_525,In_954);
nor U1112 (N_1112,In_348,In_1069);
nand U1113 (N_1113,In_1574,In_1118);
nor U1114 (N_1114,In_743,In_1451);
and U1115 (N_1115,In_1394,In_649);
nor U1116 (N_1116,In_978,In_437);
or U1117 (N_1117,In_1966,In_897);
or U1118 (N_1118,In_1470,In_887);
and U1119 (N_1119,In_1198,In_1864);
or U1120 (N_1120,In_1556,In_714);
nor U1121 (N_1121,In_1104,In_494);
nor U1122 (N_1122,In_1278,In_1998);
nor U1123 (N_1123,In_1554,In_1690);
and U1124 (N_1124,In_1887,In_41);
xnor U1125 (N_1125,In_1860,In_0);
nand U1126 (N_1126,In_1919,In_730);
nor U1127 (N_1127,In_1501,In_541);
nand U1128 (N_1128,In_1920,In_596);
or U1129 (N_1129,In_404,In_806);
and U1130 (N_1130,In_1571,In_594);
and U1131 (N_1131,In_119,In_581);
nor U1132 (N_1132,In_852,In_1447);
or U1133 (N_1133,In_1791,In_1295);
or U1134 (N_1134,In_1275,In_1650);
nand U1135 (N_1135,In_1344,In_1779);
and U1136 (N_1136,In_1599,In_711);
or U1137 (N_1137,In_1157,In_735);
nor U1138 (N_1138,In_1019,In_1061);
or U1139 (N_1139,In_588,In_1850);
nor U1140 (N_1140,In_708,In_636);
or U1141 (N_1141,In_1724,In_851);
nor U1142 (N_1142,In_1324,In_888);
and U1143 (N_1143,In_1174,In_1605);
nand U1144 (N_1144,In_825,In_468);
nor U1145 (N_1145,In_275,In_1034);
nand U1146 (N_1146,In_1961,In_678);
or U1147 (N_1147,In_1849,In_446);
and U1148 (N_1148,In_260,In_811);
nand U1149 (N_1149,In_712,In_239);
xor U1150 (N_1150,In_1390,In_538);
and U1151 (N_1151,In_1163,In_1458);
and U1152 (N_1152,In_758,In_1421);
nand U1153 (N_1153,In_497,In_1531);
and U1154 (N_1154,In_215,In_188);
and U1155 (N_1155,In_1925,In_508);
xnor U1156 (N_1156,In_394,In_1004);
and U1157 (N_1157,In_201,In_1285);
nand U1158 (N_1158,In_1427,In_249);
nand U1159 (N_1159,In_226,In_1711);
nand U1160 (N_1160,In_201,In_978);
nor U1161 (N_1161,In_1562,In_398);
nor U1162 (N_1162,In_595,In_611);
and U1163 (N_1163,In_699,In_54);
or U1164 (N_1164,In_372,In_1712);
or U1165 (N_1165,In_519,In_819);
and U1166 (N_1166,In_1225,In_414);
and U1167 (N_1167,In_379,In_1599);
or U1168 (N_1168,In_1303,In_430);
and U1169 (N_1169,In_262,In_1722);
nand U1170 (N_1170,In_5,In_1004);
nor U1171 (N_1171,In_558,In_1229);
or U1172 (N_1172,In_1246,In_578);
or U1173 (N_1173,In_448,In_1001);
or U1174 (N_1174,In_27,In_844);
and U1175 (N_1175,In_1294,In_928);
nand U1176 (N_1176,In_333,In_487);
nand U1177 (N_1177,In_466,In_1807);
or U1178 (N_1178,In_465,In_1882);
nor U1179 (N_1179,In_1692,In_1187);
or U1180 (N_1180,In_701,In_101);
nor U1181 (N_1181,In_376,In_457);
and U1182 (N_1182,In_723,In_1039);
nor U1183 (N_1183,In_262,In_612);
or U1184 (N_1184,In_675,In_137);
nor U1185 (N_1185,In_151,In_294);
nor U1186 (N_1186,In_458,In_959);
or U1187 (N_1187,In_813,In_427);
nand U1188 (N_1188,In_1523,In_1392);
and U1189 (N_1189,In_926,In_1166);
nand U1190 (N_1190,In_1170,In_739);
nand U1191 (N_1191,In_468,In_1027);
or U1192 (N_1192,In_381,In_5);
nand U1193 (N_1193,In_1748,In_610);
or U1194 (N_1194,In_1393,In_100);
nor U1195 (N_1195,In_1280,In_1935);
or U1196 (N_1196,In_164,In_1874);
nand U1197 (N_1197,In_1342,In_290);
or U1198 (N_1198,In_343,In_1014);
and U1199 (N_1199,In_1850,In_773);
or U1200 (N_1200,In_1738,In_297);
and U1201 (N_1201,In_367,In_376);
nand U1202 (N_1202,In_1108,In_620);
and U1203 (N_1203,In_1674,In_307);
nor U1204 (N_1204,In_100,In_1576);
nor U1205 (N_1205,In_632,In_1842);
nand U1206 (N_1206,In_304,In_1717);
or U1207 (N_1207,In_1635,In_1245);
or U1208 (N_1208,In_1181,In_1338);
nor U1209 (N_1209,In_1152,In_631);
nor U1210 (N_1210,In_55,In_970);
and U1211 (N_1211,In_432,In_1236);
nand U1212 (N_1212,In_90,In_1410);
nor U1213 (N_1213,In_1916,In_1761);
nor U1214 (N_1214,In_265,In_716);
nor U1215 (N_1215,In_345,In_1227);
xnor U1216 (N_1216,In_1740,In_1104);
or U1217 (N_1217,In_1804,In_1649);
nor U1218 (N_1218,In_949,In_551);
nor U1219 (N_1219,In_912,In_1733);
nand U1220 (N_1220,In_267,In_1378);
and U1221 (N_1221,In_76,In_1277);
nor U1222 (N_1222,In_1630,In_650);
nand U1223 (N_1223,In_1391,In_305);
and U1224 (N_1224,In_1799,In_1000);
and U1225 (N_1225,In_418,In_175);
or U1226 (N_1226,In_1822,In_1154);
or U1227 (N_1227,In_845,In_244);
nor U1228 (N_1228,In_23,In_1421);
or U1229 (N_1229,In_1461,In_468);
nor U1230 (N_1230,In_1291,In_395);
nand U1231 (N_1231,In_1729,In_1361);
and U1232 (N_1232,In_1624,In_706);
nor U1233 (N_1233,In_838,In_1618);
and U1234 (N_1234,In_1458,In_332);
or U1235 (N_1235,In_969,In_1263);
or U1236 (N_1236,In_1742,In_249);
or U1237 (N_1237,In_397,In_1886);
nor U1238 (N_1238,In_1885,In_1094);
nand U1239 (N_1239,In_1004,In_8);
xor U1240 (N_1240,In_1763,In_349);
and U1241 (N_1241,In_503,In_580);
or U1242 (N_1242,In_923,In_819);
or U1243 (N_1243,In_995,In_1939);
nor U1244 (N_1244,In_263,In_585);
nand U1245 (N_1245,In_806,In_1377);
nor U1246 (N_1246,In_932,In_325);
or U1247 (N_1247,In_205,In_1900);
nand U1248 (N_1248,In_330,In_1057);
nand U1249 (N_1249,In_1565,In_1431);
nand U1250 (N_1250,In_949,In_847);
nor U1251 (N_1251,In_875,In_1557);
xnor U1252 (N_1252,In_735,In_356);
and U1253 (N_1253,In_1107,In_201);
and U1254 (N_1254,In_1112,In_1847);
nand U1255 (N_1255,In_1571,In_400);
and U1256 (N_1256,In_1226,In_1011);
or U1257 (N_1257,In_416,In_368);
or U1258 (N_1258,In_537,In_315);
and U1259 (N_1259,In_1104,In_978);
or U1260 (N_1260,In_763,In_1449);
or U1261 (N_1261,In_1224,In_1989);
nor U1262 (N_1262,In_1057,In_615);
and U1263 (N_1263,In_1827,In_641);
nor U1264 (N_1264,In_109,In_192);
nor U1265 (N_1265,In_418,In_351);
or U1266 (N_1266,In_1351,In_1833);
nand U1267 (N_1267,In_429,In_1271);
and U1268 (N_1268,In_1906,In_709);
or U1269 (N_1269,In_1744,In_262);
nor U1270 (N_1270,In_696,In_201);
or U1271 (N_1271,In_405,In_919);
nand U1272 (N_1272,In_1547,In_1159);
nand U1273 (N_1273,In_959,In_1633);
nor U1274 (N_1274,In_1185,In_1424);
nand U1275 (N_1275,In_1219,In_920);
xnor U1276 (N_1276,In_260,In_1763);
and U1277 (N_1277,In_1429,In_654);
or U1278 (N_1278,In_1256,In_450);
nand U1279 (N_1279,In_770,In_200);
or U1280 (N_1280,In_319,In_1569);
and U1281 (N_1281,In_1278,In_508);
nor U1282 (N_1282,In_494,In_1693);
nand U1283 (N_1283,In_1289,In_678);
nand U1284 (N_1284,In_1069,In_129);
or U1285 (N_1285,In_309,In_204);
or U1286 (N_1286,In_362,In_1129);
and U1287 (N_1287,In_1655,In_1392);
or U1288 (N_1288,In_1906,In_978);
and U1289 (N_1289,In_1742,In_239);
nand U1290 (N_1290,In_916,In_1999);
and U1291 (N_1291,In_1986,In_29);
nand U1292 (N_1292,In_878,In_1795);
nand U1293 (N_1293,In_229,In_1207);
or U1294 (N_1294,In_227,In_931);
nor U1295 (N_1295,In_1831,In_997);
and U1296 (N_1296,In_1612,In_899);
and U1297 (N_1297,In_1798,In_890);
and U1298 (N_1298,In_1805,In_643);
and U1299 (N_1299,In_106,In_328);
and U1300 (N_1300,In_1391,In_682);
nand U1301 (N_1301,In_1109,In_1424);
nand U1302 (N_1302,In_1127,In_1142);
nor U1303 (N_1303,In_155,In_1843);
nor U1304 (N_1304,In_933,In_1555);
or U1305 (N_1305,In_754,In_240);
nand U1306 (N_1306,In_1306,In_244);
nand U1307 (N_1307,In_1422,In_393);
and U1308 (N_1308,In_1061,In_1320);
nand U1309 (N_1309,In_1444,In_1507);
or U1310 (N_1310,In_841,In_42);
xnor U1311 (N_1311,In_78,In_1804);
nor U1312 (N_1312,In_623,In_1492);
nand U1313 (N_1313,In_417,In_959);
xnor U1314 (N_1314,In_95,In_721);
or U1315 (N_1315,In_1712,In_1876);
nand U1316 (N_1316,In_663,In_1213);
nand U1317 (N_1317,In_127,In_318);
and U1318 (N_1318,In_1102,In_555);
nand U1319 (N_1319,In_1141,In_230);
nor U1320 (N_1320,In_1060,In_1502);
or U1321 (N_1321,In_1662,In_1145);
nand U1322 (N_1322,In_1915,In_1142);
or U1323 (N_1323,In_1101,In_1191);
and U1324 (N_1324,In_798,In_445);
nor U1325 (N_1325,In_358,In_657);
nor U1326 (N_1326,In_1340,In_31);
and U1327 (N_1327,In_1060,In_551);
nand U1328 (N_1328,In_307,In_887);
or U1329 (N_1329,In_1653,In_834);
nand U1330 (N_1330,In_961,In_454);
xor U1331 (N_1331,In_295,In_1168);
or U1332 (N_1332,In_848,In_292);
and U1333 (N_1333,In_1273,In_14);
nand U1334 (N_1334,In_773,In_237);
nor U1335 (N_1335,In_681,In_983);
nor U1336 (N_1336,In_1942,In_474);
or U1337 (N_1337,In_1860,In_1473);
and U1338 (N_1338,In_441,In_734);
and U1339 (N_1339,In_519,In_1457);
nor U1340 (N_1340,In_889,In_112);
nand U1341 (N_1341,In_340,In_162);
and U1342 (N_1342,In_1933,In_984);
nor U1343 (N_1343,In_1913,In_716);
and U1344 (N_1344,In_1266,In_102);
xnor U1345 (N_1345,In_1106,In_1496);
nand U1346 (N_1346,In_1143,In_1220);
or U1347 (N_1347,In_1085,In_1717);
and U1348 (N_1348,In_1246,In_304);
and U1349 (N_1349,In_890,In_5);
nand U1350 (N_1350,In_1119,In_313);
or U1351 (N_1351,In_374,In_1208);
and U1352 (N_1352,In_16,In_1079);
nand U1353 (N_1353,In_585,In_469);
xnor U1354 (N_1354,In_8,In_666);
nand U1355 (N_1355,In_531,In_328);
nand U1356 (N_1356,In_207,In_408);
nor U1357 (N_1357,In_385,In_529);
nor U1358 (N_1358,In_729,In_124);
and U1359 (N_1359,In_1973,In_394);
and U1360 (N_1360,In_1477,In_495);
xor U1361 (N_1361,In_570,In_817);
or U1362 (N_1362,In_627,In_681);
nor U1363 (N_1363,In_83,In_1398);
nor U1364 (N_1364,In_1294,In_1192);
nor U1365 (N_1365,In_1199,In_1575);
xor U1366 (N_1366,In_1045,In_1432);
nand U1367 (N_1367,In_1351,In_1048);
and U1368 (N_1368,In_887,In_503);
and U1369 (N_1369,In_1966,In_1106);
or U1370 (N_1370,In_1602,In_621);
or U1371 (N_1371,In_458,In_1100);
nor U1372 (N_1372,In_290,In_925);
and U1373 (N_1373,In_820,In_918);
nand U1374 (N_1374,In_114,In_1543);
nand U1375 (N_1375,In_1093,In_1671);
or U1376 (N_1376,In_1480,In_1603);
nand U1377 (N_1377,In_1790,In_359);
nor U1378 (N_1378,In_847,In_894);
or U1379 (N_1379,In_1777,In_1263);
and U1380 (N_1380,In_1220,In_1703);
nor U1381 (N_1381,In_903,In_880);
nor U1382 (N_1382,In_728,In_1934);
xor U1383 (N_1383,In_309,In_1101);
and U1384 (N_1384,In_1916,In_179);
xor U1385 (N_1385,In_1695,In_249);
nand U1386 (N_1386,In_957,In_1330);
and U1387 (N_1387,In_1407,In_63);
nand U1388 (N_1388,In_629,In_411);
or U1389 (N_1389,In_1741,In_1712);
and U1390 (N_1390,In_420,In_1659);
or U1391 (N_1391,In_1406,In_1227);
xnor U1392 (N_1392,In_377,In_1452);
nor U1393 (N_1393,In_924,In_1279);
or U1394 (N_1394,In_886,In_252);
nand U1395 (N_1395,In_151,In_1483);
nand U1396 (N_1396,In_546,In_1440);
or U1397 (N_1397,In_1871,In_764);
nor U1398 (N_1398,In_1935,In_388);
nand U1399 (N_1399,In_1488,In_1130);
nand U1400 (N_1400,In_533,In_1063);
nand U1401 (N_1401,In_1226,In_691);
or U1402 (N_1402,In_991,In_1154);
xor U1403 (N_1403,In_844,In_768);
or U1404 (N_1404,In_1618,In_77);
or U1405 (N_1405,In_1226,In_829);
or U1406 (N_1406,In_897,In_90);
or U1407 (N_1407,In_239,In_818);
xnor U1408 (N_1408,In_658,In_292);
or U1409 (N_1409,In_1924,In_632);
nand U1410 (N_1410,In_881,In_653);
and U1411 (N_1411,In_711,In_1608);
and U1412 (N_1412,In_1518,In_1679);
nor U1413 (N_1413,In_175,In_115);
or U1414 (N_1414,In_1660,In_1423);
nand U1415 (N_1415,In_1315,In_944);
or U1416 (N_1416,In_1325,In_216);
and U1417 (N_1417,In_1524,In_1519);
or U1418 (N_1418,In_765,In_1644);
or U1419 (N_1419,In_1855,In_1684);
and U1420 (N_1420,In_112,In_641);
nand U1421 (N_1421,In_1225,In_1091);
nand U1422 (N_1422,In_1647,In_14);
nand U1423 (N_1423,In_858,In_617);
nor U1424 (N_1424,In_376,In_1011);
and U1425 (N_1425,In_1931,In_749);
nand U1426 (N_1426,In_558,In_400);
or U1427 (N_1427,In_1424,In_633);
nand U1428 (N_1428,In_262,In_1696);
or U1429 (N_1429,In_1499,In_518);
nand U1430 (N_1430,In_1006,In_905);
or U1431 (N_1431,In_1561,In_1743);
nand U1432 (N_1432,In_1496,In_1630);
nor U1433 (N_1433,In_939,In_1782);
or U1434 (N_1434,In_1748,In_703);
or U1435 (N_1435,In_1210,In_950);
and U1436 (N_1436,In_1573,In_1048);
nor U1437 (N_1437,In_712,In_1355);
and U1438 (N_1438,In_699,In_689);
xor U1439 (N_1439,In_181,In_71);
nand U1440 (N_1440,In_1181,In_682);
or U1441 (N_1441,In_613,In_1944);
or U1442 (N_1442,In_686,In_562);
nand U1443 (N_1443,In_653,In_1445);
nor U1444 (N_1444,In_443,In_1251);
or U1445 (N_1445,In_187,In_1629);
and U1446 (N_1446,In_203,In_1468);
nor U1447 (N_1447,In_1946,In_1829);
and U1448 (N_1448,In_1375,In_1633);
or U1449 (N_1449,In_94,In_176);
and U1450 (N_1450,In_354,In_3);
and U1451 (N_1451,In_1017,In_1660);
nand U1452 (N_1452,In_1476,In_1793);
nor U1453 (N_1453,In_791,In_1665);
nand U1454 (N_1454,In_1709,In_1509);
nor U1455 (N_1455,In_380,In_269);
nor U1456 (N_1456,In_168,In_1217);
or U1457 (N_1457,In_960,In_311);
nand U1458 (N_1458,In_1570,In_1328);
nor U1459 (N_1459,In_1894,In_1787);
or U1460 (N_1460,In_1847,In_1868);
nor U1461 (N_1461,In_3,In_1691);
nand U1462 (N_1462,In_1006,In_217);
xor U1463 (N_1463,In_529,In_119);
and U1464 (N_1464,In_398,In_202);
or U1465 (N_1465,In_1209,In_678);
or U1466 (N_1466,In_909,In_754);
and U1467 (N_1467,In_241,In_218);
or U1468 (N_1468,In_1147,In_821);
xor U1469 (N_1469,In_102,In_1704);
and U1470 (N_1470,In_960,In_863);
nor U1471 (N_1471,In_583,In_124);
nor U1472 (N_1472,In_1765,In_846);
nor U1473 (N_1473,In_828,In_1640);
nor U1474 (N_1474,In_1116,In_1339);
or U1475 (N_1475,In_527,In_1061);
nand U1476 (N_1476,In_928,In_1411);
or U1477 (N_1477,In_874,In_1981);
nor U1478 (N_1478,In_149,In_1801);
and U1479 (N_1479,In_218,In_1874);
or U1480 (N_1480,In_146,In_1718);
nand U1481 (N_1481,In_208,In_1224);
or U1482 (N_1482,In_16,In_1263);
or U1483 (N_1483,In_1590,In_1190);
and U1484 (N_1484,In_1418,In_404);
nor U1485 (N_1485,In_1957,In_415);
and U1486 (N_1486,In_132,In_1906);
xnor U1487 (N_1487,In_553,In_398);
xor U1488 (N_1488,In_795,In_1124);
xor U1489 (N_1489,In_13,In_558);
xor U1490 (N_1490,In_1146,In_435);
or U1491 (N_1491,In_362,In_329);
nand U1492 (N_1492,In_1177,In_1160);
or U1493 (N_1493,In_1343,In_841);
nand U1494 (N_1494,In_1941,In_570);
nor U1495 (N_1495,In_737,In_198);
or U1496 (N_1496,In_1981,In_650);
or U1497 (N_1497,In_1357,In_1313);
and U1498 (N_1498,In_1007,In_568);
xnor U1499 (N_1499,In_1743,In_1689);
or U1500 (N_1500,In_1434,In_120);
or U1501 (N_1501,In_839,In_1734);
and U1502 (N_1502,In_68,In_1055);
nor U1503 (N_1503,In_649,In_464);
nor U1504 (N_1504,In_984,In_1498);
xor U1505 (N_1505,In_323,In_328);
and U1506 (N_1506,In_525,In_1459);
nor U1507 (N_1507,In_1629,In_230);
nand U1508 (N_1508,In_1891,In_248);
nand U1509 (N_1509,In_681,In_101);
or U1510 (N_1510,In_262,In_684);
nand U1511 (N_1511,In_1422,In_1683);
nor U1512 (N_1512,In_139,In_651);
xor U1513 (N_1513,In_1893,In_98);
and U1514 (N_1514,In_550,In_1201);
nor U1515 (N_1515,In_631,In_692);
nor U1516 (N_1516,In_883,In_545);
nand U1517 (N_1517,In_222,In_1940);
nor U1518 (N_1518,In_432,In_675);
nand U1519 (N_1519,In_1994,In_389);
and U1520 (N_1520,In_755,In_1453);
nand U1521 (N_1521,In_504,In_1392);
nand U1522 (N_1522,In_101,In_1964);
nand U1523 (N_1523,In_475,In_1128);
nor U1524 (N_1524,In_1031,In_339);
and U1525 (N_1525,In_1234,In_1332);
and U1526 (N_1526,In_51,In_1104);
nand U1527 (N_1527,In_961,In_271);
nand U1528 (N_1528,In_584,In_113);
nor U1529 (N_1529,In_1410,In_52);
nand U1530 (N_1530,In_816,In_1258);
or U1531 (N_1531,In_1045,In_1583);
or U1532 (N_1532,In_30,In_1473);
nor U1533 (N_1533,In_1955,In_324);
and U1534 (N_1534,In_40,In_128);
xnor U1535 (N_1535,In_1754,In_1181);
and U1536 (N_1536,In_1390,In_1465);
nor U1537 (N_1537,In_1533,In_996);
and U1538 (N_1538,In_337,In_1056);
nor U1539 (N_1539,In_963,In_1757);
nor U1540 (N_1540,In_707,In_559);
or U1541 (N_1541,In_1900,In_1532);
and U1542 (N_1542,In_1108,In_1106);
and U1543 (N_1543,In_63,In_1139);
and U1544 (N_1544,In_947,In_918);
nor U1545 (N_1545,In_1898,In_394);
or U1546 (N_1546,In_449,In_247);
nor U1547 (N_1547,In_1802,In_1483);
nor U1548 (N_1548,In_1718,In_1165);
and U1549 (N_1549,In_370,In_77);
nor U1550 (N_1550,In_1177,In_196);
nand U1551 (N_1551,In_723,In_1876);
nand U1552 (N_1552,In_0,In_1047);
nor U1553 (N_1553,In_54,In_1508);
nor U1554 (N_1554,In_1143,In_1180);
and U1555 (N_1555,In_1719,In_950);
or U1556 (N_1556,In_1266,In_1432);
nand U1557 (N_1557,In_478,In_416);
and U1558 (N_1558,In_59,In_811);
nand U1559 (N_1559,In_562,In_1160);
and U1560 (N_1560,In_251,In_151);
nor U1561 (N_1561,In_1720,In_1184);
nor U1562 (N_1562,In_1751,In_80);
or U1563 (N_1563,In_1484,In_1719);
or U1564 (N_1564,In_1999,In_1993);
nand U1565 (N_1565,In_1545,In_473);
and U1566 (N_1566,In_628,In_1891);
nor U1567 (N_1567,In_1835,In_765);
nand U1568 (N_1568,In_339,In_1967);
nand U1569 (N_1569,In_531,In_1794);
and U1570 (N_1570,In_337,In_657);
or U1571 (N_1571,In_1987,In_1148);
or U1572 (N_1572,In_118,In_1156);
nor U1573 (N_1573,In_1399,In_792);
or U1574 (N_1574,In_867,In_412);
and U1575 (N_1575,In_1757,In_188);
or U1576 (N_1576,In_113,In_220);
or U1577 (N_1577,In_162,In_1354);
nand U1578 (N_1578,In_653,In_125);
nor U1579 (N_1579,In_1816,In_945);
or U1580 (N_1580,In_1091,In_1206);
nand U1581 (N_1581,In_1987,In_1153);
nand U1582 (N_1582,In_1841,In_0);
nand U1583 (N_1583,In_9,In_1932);
xor U1584 (N_1584,In_1312,In_249);
nor U1585 (N_1585,In_1019,In_1975);
nand U1586 (N_1586,In_1181,In_942);
and U1587 (N_1587,In_1492,In_1134);
xnor U1588 (N_1588,In_685,In_1804);
nor U1589 (N_1589,In_817,In_637);
nor U1590 (N_1590,In_637,In_246);
nand U1591 (N_1591,In_626,In_1167);
or U1592 (N_1592,In_1101,In_975);
and U1593 (N_1593,In_1333,In_1989);
and U1594 (N_1594,In_726,In_1205);
or U1595 (N_1595,In_360,In_363);
and U1596 (N_1596,In_1745,In_226);
or U1597 (N_1597,In_469,In_517);
xnor U1598 (N_1598,In_667,In_1127);
nor U1599 (N_1599,In_1680,In_210);
nand U1600 (N_1600,In_1066,In_52);
nor U1601 (N_1601,In_1558,In_1285);
nand U1602 (N_1602,In_1577,In_827);
or U1603 (N_1603,In_1826,In_1820);
and U1604 (N_1604,In_555,In_36);
nand U1605 (N_1605,In_1810,In_864);
nor U1606 (N_1606,In_1567,In_659);
nand U1607 (N_1607,In_640,In_94);
xnor U1608 (N_1608,In_1840,In_578);
nor U1609 (N_1609,In_1109,In_1512);
nand U1610 (N_1610,In_1395,In_1994);
or U1611 (N_1611,In_1938,In_273);
xnor U1612 (N_1612,In_342,In_235);
nor U1613 (N_1613,In_1432,In_940);
nand U1614 (N_1614,In_1213,In_510);
and U1615 (N_1615,In_1756,In_303);
nor U1616 (N_1616,In_1681,In_622);
and U1617 (N_1617,In_1208,In_1340);
and U1618 (N_1618,In_961,In_1184);
nor U1619 (N_1619,In_1483,In_1280);
nand U1620 (N_1620,In_56,In_905);
and U1621 (N_1621,In_1338,In_73);
or U1622 (N_1622,In_1379,In_989);
nand U1623 (N_1623,In_411,In_578);
nor U1624 (N_1624,In_1890,In_1488);
nor U1625 (N_1625,In_408,In_1908);
nand U1626 (N_1626,In_997,In_1459);
or U1627 (N_1627,In_1380,In_1043);
and U1628 (N_1628,In_510,In_1091);
nand U1629 (N_1629,In_335,In_594);
nor U1630 (N_1630,In_1879,In_928);
and U1631 (N_1631,In_1609,In_1752);
or U1632 (N_1632,In_508,In_1424);
nand U1633 (N_1633,In_321,In_478);
or U1634 (N_1634,In_433,In_394);
nand U1635 (N_1635,In_1252,In_1675);
and U1636 (N_1636,In_245,In_79);
nor U1637 (N_1637,In_388,In_536);
and U1638 (N_1638,In_1481,In_1189);
and U1639 (N_1639,In_215,In_867);
nor U1640 (N_1640,In_129,In_1356);
and U1641 (N_1641,In_673,In_1333);
nor U1642 (N_1642,In_594,In_971);
nand U1643 (N_1643,In_1244,In_479);
or U1644 (N_1644,In_976,In_667);
xnor U1645 (N_1645,In_1238,In_1571);
and U1646 (N_1646,In_1774,In_856);
or U1647 (N_1647,In_1879,In_963);
and U1648 (N_1648,In_738,In_1624);
and U1649 (N_1649,In_767,In_212);
and U1650 (N_1650,In_840,In_470);
nor U1651 (N_1651,In_1506,In_1430);
nor U1652 (N_1652,In_704,In_190);
xnor U1653 (N_1653,In_1424,In_1263);
nor U1654 (N_1654,In_292,In_1884);
nand U1655 (N_1655,In_1680,In_312);
nor U1656 (N_1656,In_1228,In_672);
xnor U1657 (N_1657,In_1766,In_1915);
or U1658 (N_1658,In_1812,In_1203);
nand U1659 (N_1659,In_442,In_710);
nand U1660 (N_1660,In_672,In_1851);
or U1661 (N_1661,In_1689,In_247);
nand U1662 (N_1662,In_1047,In_1290);
nand U1663 (N_1663,In_1740,In_1058);
and U1664 (N_1664,In_411,In_1351);
nand U1665 (N_1665,In_1914,In_408);
and U1666 (N_1666,In_347,In_997);
nor U1667 (N_1667,In_1041,In_1107);
and U1668 (N_1668,In_374,In_329);
or U1669 (N_1669,In_1628,In_204);
nor U1670 (N_1670,In_1857,In_1383);
nor U1671 (N_1671,In_1732,In_375);
nor U1672 (N_1672,In_1674,In_296);
nor U1673 (N_1673,In_556,In_1358);
nand U1674 (N_1674,In_1353,In_30);
and U1675 (N_1675,In_995,In_1213);
nor U1676 (N_1676,In_369,In_177);
and U1677 (N_1677,In_125,In_938);
or U1678 (N_1678,In_1208,In_56);
or U1679 (N_1679,In_1280,In_544);
or U1680 (N_1680,In_114,In_1796);
nor U1681 (N_1681,In_1556,In_1324);
and U1682 (N_1682,In_1304,In_658);
and U1683 (N_1683,In_1059,In_1482);
or U1684 (N_1684,In_250,In_1802);
and U1685 (N_1685,In_729,In_294);
and U1686 (N_1686,In_167,In_1729);
or U1687 (N_1687,In_1577,In_1669);
or U1688 (N_1688,In_1138,In_1441);
xnor U1689 (N_1689,In_1118,In_1518);
and U1690 (N_1690,In_1822,In_894);
or U1691 (N_1691,In_1606,In_1906);
and U1692 (N_1692,In_1645,In_1588);
xor U1693 (N_1693,In_736,In_1076);
nand U1694 (N_1694,In_1563,In_552);
nand U1695 (N_1695,In_1025,In_566);
or U1696 (N_1696,In_1694,In_1191);
nor U1697 (N_1697,In_1925,In_296);
or U1698 (N_1698,In_1536,In_826);
and U1699 (N_1699,In_1259,In_40);
xor U1700 (N_1700,In_491,In_1298);
and U1701 (N_1701,In_565,In_1984);
nand U1702 (N_1702,In_156,In_1467);
nand U1703 (N_1703,In_834,In_1793);
and U1704 (N_1704,In_581,In_138);
and U1705 (N_1705,In_1073,In_1302);
nand U1706 (N_1706,In_1589,In_58);
and U1707 (N_1707,In_1471,In_765);
and U1708 (N_1708,In_1526,In_968);
nand U1709 (N_1709,In_1249,In_1707);
nor U1710 (N_1710,In_1712,In_1218);
xor U1711 (N_1711,In_394,In_1547);
nor U1712 (N_1712,In_1250,In_1354);
nand U1713 (N_1713,In_1362,In_1562);
and U1714 (N_1714,In_1456,In_763);
and U1715 (N_1715,In_961,In_1851);
xor U1716 (N_1716,In_1007,In_1107);
nor U1717 (N_1717,In_1383,In_276);
or U1718 (N_1718,In_1143,In_1939);
nand U1719 (N_1719,In_1223,In_15);
and U1720 (N_1720,In_1585,In_1307);
nand U1721 (N_1721,In_8,In_1721);
and U1722 (N_1722,In_1461,In_1850);
and U1723 (N_1723,In_1599,In_1121);
xnor U1724 (N_1724,In_1285,In_1340);
nor U1725 (N_1725,In_1727,In_1868);
xor U1726 (N_1726,In_1865,In_798);
nor U1727 (N_1727,In_605,In_1779);
and U1728 (N_1728,In_1627,In_159);
nor U1729 (N_1729,In_1610,In_451);
xor U1730 (N_1730,In_1567,In_1823);
and U1731 (N_1731,In_524,In_1104);
and U1732 (N_1732,In_552,In_226);
nand U1733 (N_1733,In_1720,In_483);
nand U1734 (N_1734,In_498,In_1752);
or U1735 (N_1735,In_785,In_1344);
or U1736 (N_1736,In_796,In_759);
nor U1737 (N_1737,In_432,In_345);
xnor U1738 (N_1738,In_1002,In_1414);
or U1739 (N_1739,In_866,In_1422);
xor U1740 (N_1740,In_130,In_588);
or U1741 (N_1741,In_109,In_1018);
and U1742 (N_1742,In_749,In_357);
and U1743 (N_1743,In_591,In_1638);
nand U1744 (N_1744,In_1671,In_1550);
nand U1745 (N_1745,In_1229,In_1517);
and U1746 (N_1746,In_632,In_728);
nand U1747 (N_1747,In_1341,In_1710);
nand U1748 (N_1748,In_1432,In_831);
nand U1749 (N_1749,In_1022,In_906);
nor U1750 (N_1750,In_226,In_994);
nor U1751 (N_1751,In_430,In_19);
and U1752 (N_1752,In_1115,In_500);
nor U1753 (N_1753,In_46,In_1853);
nand U1754 (N_1754,In_1341,In_881);
nand U1755 (N_1755,In_1133,In_1098);
nand U1756 (N_1756,In_1184,In_1522);
xnor U1757 (N_1757,In_1330,In_1707);
nand U1758 (N_1758,In_153,In_1217);
or U1759 (N_1759,In_1590,In_106);
and U1760 (N_1760,In_1700,In_1549);
nand U1761 (N_1761,In_1691,In_1048);
nor U1762 (N_1762,In_1182,In_1514);
nor U1763 (N_1763,In_1934,In_1207);
nor U1764 (N_1764,In_833,In_465);
and U1765 (N_1765,In_1697,In_1416);
or U1766 (N_1766,In_499,In_1947);
nand U1767 (N_1767,In_407,In_953);
and U1768 (N_1768,In_249,In_1571);
nand U1769 (N_1769,In_1309,In_620);
nor U1770 (N_1770,In_346,In_1521);
or U1771 (N_1771,In_838,In_1985);
nand U1772 (N_1772,In_28,In_1704);
nand U1773 (N_1773,In_964,In_293);
nand U1774 (N_1774,In_1098,In_1733);
nor U1775 (N_1775,In_1571,In_954);
and U1776 (N_1776,In_1916,In_1546);
nand U1777 (N_1777,In_554,In_1533);
nand U1778 (N_1778,In_1711,In_546);
xor U1779 (N_1779,In_189,In_1478);
xnor U1780 (N_1780,In_1754,In_1350);
and U1781 (N_1781,In_1073,In_195);
nand U1782 (N_1782,In_1844,In_1393);
nand U1783 (N_1783,In_1036,In_1980);
nor U1784 (N_1784,In_1084,In_1139);
nor U1785 (N_1785,In_1387,In_669);
xor U1786 (N_1786,In_1849,In_147);
and U1787 (N_1787,In_374,In_294);
and U1788 (N_1788,In_1107,In_1196);
xor U1789 (N_1789,In_1566,In_1180);
xor U1790 (N_1790,In_1564,In_328);
and U1791 (N_1791,In_1593,In_1562);
xnor U1792 (N_1792,In_680,In_308);
nor U1793 (N_1793,In_1513,In_148);
or U1794 (N_1794,In_681,In_1334);
nor U1795 (N_1795,In_1470,In_1202);
nand U1796 (N_1796,In_719,In_1483);
nor U1797 (N_1797,In_1745,In_1904);
nor U1798 (N_1798,In_783,In_356);
and U1799 (N_1799,In_819,In_1869);
or U1800 (N_1800,In_448,In_1271);
nand U1801 (N_1801,In_1830,In_502);
or U1802 (N_1802,In_1551,In_940);
xor U1803 (N_1803,In_29,In_1604);
nor U1804 (N_1804,In_1051,In_437);
xor U1805 (N_1805,In_344,In_1006);
nor U1806 (N_1806,In_13,In_590);
nor U1807 (N_1807,In_1032,In_266);
and U1808 (N_1808,In_1552,In_25);
nand U1809 (N_1809,In_1381,In_441);
or U1810 (N_1810,In_1532,In_1479);
or U1811 (N_1811,In_740,In_1885);
xor U1812 (N_1812,In_794,In_1013);
xnor U1813 (N_1813,In_102,In_634);
nand U1814 (N_1814,In_47,In_1462);
or U1815 (N_1815,In_1679,In_1648);
xnor U1816 (N_1816,In_42,In_470);
xor U1817 (N_1817,In_623,In_1420);
nor U1818 (N_1818,In_1028,In_334);
xnor U1819 (N_1819,In_1496,In_1863);
nand U1820 (N_1820,In_1099,In_1018);
or U1821 (N_1821,In_29,In_1873);
and U1822 (N_1822,In_840,In_1642);
and U1823 (N_1823,In_1559,In_127);
or U1824 (N_1824,In_176,In_535);
and U1825 (N_1825,In_246,In_1416);
or U1826 (N_1826,In_1480,In_1506);
xnor U1827 (N_1827,In_52,In_444);
nand U1828 (N_1828,In_1180,In_88);
or U1829 (N_1829,In_860,In_1729);
nor U1830 (N_1830,In_1312,In_169);
and U1831 (N_1831,In_1489,In_164);
or U1832 (N_1832,In_103,In_1531);
nor U1833 (N_1833,In_929,In_894);
nand U1834 (N_1834,In_783,In_1457);
xor U1835 (N_1835,In_250,In_1698);
nand U1836 (N_1836,In_1480,In_929);
and U1837 (N_1837,In_1677,In_512);
xnor U1838 (N_1838,In_1734,In_504);
and U1839 (N_1839,In_1274,In_1177);
and U1840 (N_1840,In_768,In_1765);
and U1841 (N_1841,In_653,In_139);
and U1842 (N_1842,In_1353,In_1789);
and U1843 (N_1843,In_146,In_739);
nor U1844 (N_1844,In_19,In_702);
nand U1845 (N_1845,In_1733,In_1630);
and U1846 (N_1846,In_1332,In_958);
nand U1847 (N_1847,In_1549,In_255);
nor U1848 (N_1848,In_1262,In_1526);
nor U1849 (N_1849,In_1388,In_137);
or U1850 (N_1850,In_616,In_349);
and U1851 (N_1851,In_177,In_1289);
nor U1852 (N_1852,In_884,In_184);
nor U1853 (N_1853,In_1853,In_199);
or U1854 (N_1854,In_1386,In_259);
nand U1855 (N_1855,In_1067,In_166);
nand U1856 (N_1856,In_929,In_1551);
nor U1857 (N_1857,In_1804,In_1983);
nand U1858 (N_1858,In_924,In_1280);
nor U1859 (N_1859,In_977,In_166);
and U1860 (N_1860,In_56,In_1512);
or U1861 (N_1861,In_1023,In_895);
nor U1862 (N_1862,In_1713,In_1739);
xnor U1863 (N_1863,In_1041,In_1245);
nand U1864 (N_1864,In_682,In_1412);
nand U1865 (N_1865,In_1996,In_359);
or U1866 (N_1866,In_1313,In_43);
nand U1867 (N_1867,In_363,In_1592);
nand U1868 (N_1868,In_16,In_1122);
and U1869 (N_1869,In_1917,In_369);
nand U1870 (N_1870,In_307,In_331);
and U1871 (N_1871,In_1862,In_1895);
and U1872 (N_1872,In_312,In_1329);
xnor U1873 (N_1873,In_1303,In_379);
and U1874 (N_1874,In_81,In_659);
xnor U1875 (N_1875,In_1401,In_1421);
nor U1876 (N_1876,In_1155,In_351);
nand U1877 (N_1877,In_1849,In_404);
or U1878 (N_1878,In_819,In_1514);
nand U1879 (N_1879,In_234,In_140);
and U1880 (N_1880,In_760,In_1466);
nand U1881 (N_1881,In_1809,In_1794);
xnor U1882 (N_1882,In_25,In_529);
xor U1883 (N_1883,In_1839,In_1975);
nor U1884 (N_1884,In_1631,In_75);
and U1885 (N_1885,In_911,In_700);
or U1886 (N_1886,In_126,In_587);
nand U1887 (N_1887,In_716,In_135);
nor U1888 (N_1888,In_1569,In_1725);
nand U1889 (N_1889,In_220,In_195);
xnor U1890 (N_1890,In_658,In_1389);
nor U1891 (N_1891,In_1242,In_1082);
or U1892 (N_1892,In_1386,In_616);
or U1893 (N_1893,In_1722,In_1023);
nand U1894 (N_1894,In_12,In_63);
nor U1895 (N_1895,In_1582,In_466);
nand U1896 (N_1896,In_1232,In_60);
nor U1897 (N_1897,In_1299,In_1024);
or U1898 (N_1898,In_1141,In_1309);
or U1899 (N_1899,In_845,In_1378);
or U1900 (N_1900,In_909,In_1417);
and U1901 (N_1901,In_1758,In_1513);
nor U1902 (N_1902,In_1402,In_1665);
or U1903 (N_1903,In_1898,In_393);
nor U1904 (N_1904,In_63,In_969);
nor U1905 (N_1905,In_54,In_1458);
and U1906 (N_1906,In_585,In_1821);
or U1907 (N_1907,In_1212,In_916);
and U1908 (N_1908,In_1619,In_648);
and U1909 (N_1909,In_1330,In_1073);
and U1910 (N_1910,In_785,In_1264);
nand U1911 (N_1911,In_1170,In_1663);
xnor U1912 (N_1912,In_1072,In_117);
nor U1913 (N_1913,In_474,In_1433);
or U1914 (N_1914,In_386,In_1796);
nand U1915 (N_1915,In_281,In_419);
nand U1916 (N_1916,In_1732,In_1966);
xor U1917 (N_1917,In_1235,In_1439);
nand U1918 (N_1918,In_1956,In_1320);
and U1919 (N_1919,In_1496,In_1809);
and U1920 (N_1920,In_1101,In_1105);
nor U1921 (N_1921,In_1574,In_1805);
nor U1922 (N_1922,In_1035,In_1039);
nor U1923 (N_1923,In_1384,In_1931);
nand U1924 (N_1924,In_1648,In_552);
and U1925 (N_1925,In_1600,In_982);
and U1926 (N_1926,In_753,In_387);
nand U1927 (N_1927,In_1407,In_211);
nor U1928 (N_1928,In_1752,In_1740);
and U1929 (N_1929,In_277,In_579);
or U1930 (N_1930,In_78,In_729);
xor U1931 (N_1931,In_228,In_555);
or U1932 (N_1932,In_1277,In_1164);
nand U1933 (N_1933,In_1610,In_1319);
nand U1934 (N_1934,In_416,In_621);
nand U1935 (N_1935,In_1598,In_542);
nor U1936 (N_1936,In_429,In_1822);
or U1937 (N_1937,In_1052,In_489);
and U1938 (N_1938,In_612,In_1241);
nand U1939 (N_1939,In_729,In_630);
or U1940 (N_1940,In_143,In_1205);
nand U1941 (N_1941,In_617,In_1719);
nor U1942 (N_1942,In_1980,In_1658);
or U1943 (N_1943,In_820,In_221);
or U1944 (N_1944,In_747,In_542);
nor U1945 (N_1945,In_512,In_481);
xor U1946 (N_1946,In_1471,In_1213);
nor U1947 (N_1947,In_1169,In_1150);
nand U1948 (N_1948,In_1953,In_1666);
and U1949 (N_1949,In_1094,In_597);
nor U1950 (N_1950,In_715,In_1967);
xnor U1951 (N_1951,In_180,In_1328);
or U1952 (N_1952,In_1355,In_1605);
nand U1953 (N_1953,In_269,In_933);
or U1954 (N_1954,In_927,In_346);
nand U1955 (N_1955,In_1845,In_1169);
and U1956 (N_1956,In_337,In_1975);
or U1957 (N_1957,In_1267,In_1703);
nand U1958 (N_1958,In_485,In_1464);
xor U1959 (N_1959,In_1387,In_1608);
nand U1960 (N_1960,In_403,In_123);
nand U1961 (N_1961,In_1945,In_1422);
and U1962 (N_1962,In_1807,In_1532);
and U1963 (N_1963,In_1250,In_988);
or U1964 (N_1964,In_1056,In_1076);
or U1965 (N_1965,In_546,In_1116);
nand U1966 (N_1966,In_1164,In_1756);
or U1967 (N_1967,In_771,In_597);
or U1968 (N_1968,In_793,In_1892);
nand U1969 (N_1969,In_1173,In_322);
and U1970 (N_1970,In_480,In_208);
and U1971 (N_1971,In_1919,In_362);
and U1972 (N_1972,In_1885,In_1520);
or U1973 (N_1973,In_1281,In_635);
xor U1974 (N_1974,In_4,In_1525);
xor U1975 (N_1975,In_1865,In_1661);
xor U1976 (N_1976,In_448,In_1427);
nand U1977 (N_1977,In_585,In_1473);
and U1978 (N_1978,In_1902,In_1442);
xor U1979 (N_1979,In_712,In_677);
or U1980 (N_1980,In_536,In_1014);
nand U1981 (N_1981,In_381,In_1469);
and U1982 (N_1982,In_277,In_1048);
nor U1983 (N_1983,In_1919,In_274);
nand U1984 (N_1984,In_248,In_1237);
or U1985 (N_1985,In_403,In_1758);
xor U1986 (N_1986,In_994,In_614);
or U1987 (N_1987,In_53,In_942);
or U1988 (N_1988,In_1995,In_647);
xnor U1989 (N_1989,In_1828,In_1921);
xnor U1990 (N_1990,In_281,In_1865);
or U1991 (N_1991,In_932,In_1676);
nand U1992 (N_1992,In_1544,In_1234);
or U1993 (N_1993,In_1843,In_1018);
or U1994 (N_1994,In_140,In_1321);
or U1995 (N_1995,In_905,In_109);
nor U1996 (N_1996,In_447,In_919);
xor U1997 (N_1997,In_1461,In_1886);
or U1998 (N_1998,In_1389,In_1106);
nor U1999 (N_1999,In_729,In_769);
xnor U2000 (N_2000,N_894,N_896);
nor U2001 (N_2001,N_1436,N_715);
and U2002 (N_2002,N_392,N_1660);
nand U2003 (N_2003,N_1937,N_615);
or U2004 (N_2004,N_599,N_1276);
or U2005 (N_2005,N_1770,N_1040);
and U2006 (N_2006,N_1594,N_1457);
nand U2007 (N_2007,N_1719,N_954);
and U2008 (N_2008,N_220,N_1603);
and U2009 (N_2009,N_1073,N_1613);
nor U2010 (N_2010,N_613,N_516);
and U2011 (N_2011,N_274,N_1991);
nand U2012 (N_2012,N_1110,N_306);
and U2013 (N_2013,N_247,N_1864);
and U2014 (N_2014,N_1575,N_101);
and U2015 (N_2015,N_1897,N_85);
xnor U2016 (N_2016,N_175,N_1776);
nand U2017 (N_2017,N_1096,N_77);
nor U2018 (N_2018,N_332,N_1044);
nand U2019 (N_2019,N_610,N_1086);
or U2020 (N_2020,N_366,N_1549);
or U2021 (N_2021,N_916,N_1765);
nor U2022 (N_2022,N_1692,N_1414);
nand U2023 (N_2023,N_1103,N_1329);
nor U2024 (N_2024,N_857,N_539);
and U2025 (N_2025,N_1139,N_1172);
and U2026 (N_2026,N_700,N_526);
or U2027 (N_2027,N_1905,N_1989);
and U2028 (N_2028,N_237,N_915);
and U2029 (N_2029,N_483,N_36);
or U2030 (N_2030,N_675,N_722);
or U2031 (N_2031,N_417,N_126);
nand U2032 (N_2032,N_787,N_64);
nor U2033 (N_2033,N_618,N_148);
nand U2034 (N_2034,N_1479,N_863);
or U2035 (N_2035,N_1188,N_714);
nor U2036 (N_2036,N_1595,N_1304);
nand U2037 (N_2037,N_1543,N_1358);
nand U2038 (N_2038,N_969,N_1015);
or U2039 (N_2039,N_405,N_1762);
or U2040 (N_2040,N_1957,N_345);
and U2041 (N_2041,N_1419,N_665);
or U2042 (N_2042,N_1371,N_119);
and U2043 (N_2043,N_1145,N_962);
or U2044 (N_2044,N_671,N_234);
nor U2045 (N_2045,N_472,N_1437);
and U2046 (N_2046,N_377,N_534);
nand U2047 (N_2047,N_1944,N_1552);
or U2048 (N_2048,N_1798,N_1085);
nand U2049 (N_2049,N_1287,N_606);
and U2050 (N_2050,N_1882,N_1931);
or U2051 (N_2051,N_433,N_543);
or U2052 (N_2052,N_308,N_1300);
and U2053 (N_2053,N_1727,N_1713);
or U2054 (N_2054,N_994,N_1749);
xor U2055 (N_2055,N_963,N_1097);
or U2056 (N_2056,N_359,N_435);
or U2057 (N_2057,N_872,N_1498);
or U2058 (N_2058,N_1837,N_533);
and U2059 (N_2059,N_1914,N_136);
or U2060 (N_2060,N_1639,N_1126);
or U2061 (N_2061,N_1334,N_737);
nand U2062 (N_2062,N_222,N_769);
or U2063 (N_2063,N_1791,N_1602);
nand U2064 (N_2064,N_745,N_1232);
nor U2065 (N_2065,N_42,N_1452);
and U2066 (N_2066,N_1638,N_321);
or U2067 (N_2067,N_114,N_348);
nand U2068 (N_2068,N_1652,N_725);
nand U2069 (N_2069,N_997,N_132);
or U2070 (N_2070,N_1783,N_1305);
or U2071 (N_2071,N_303,N_307);
or U2072 (N_2072,N_1078,N_1506);
nor U2073 (N_2073,N_649,N_133);
or U2074 (N_2074,N_463,N_1490);
nor U2075 (N_2075,N_1885,N_129);
and U2076 (N_2076,N_981,N_458);
nor U2077 (N_2077,N_1376,N_1855);
nor U2078 (N_2078,N_477,N_1683);
nor U2079 (N_2079,N_1546,N_960);
nand U2080 (N_2080,N_1737,N_1259);
xor U2081 (N_2081,N_447,N_1102);
or U2082 (N_2082,N_1813,N_595);
or U2083 (N_2083,N_556,N_1104);
or U2084 (N_2084,N_1434,N_445);
nand U2085 (N_2085,N_1654,N_1065);
xor U2086 (N_2086,N_1558,N_811);
nand U2087 (N_2087,N_741,N_1384);
and U2088 (N_2088,N_1442,N_1563);
or U2089 (N_2089,N_10,N_900);
nand U2090 (N_2090,N_198,N_494);
and U2091 (N_2091,N_632,N_1385);
or U2092 (N_2092,N_727,N_1889);
xor U2093 (N_2093,N_421,N_1938);
nor U2094 (N_2094,N_1890,N_780);
or U2095 (N_2095,N_596,N_322);
and U2096 (N_2096,N_621,N_668);
nor U2097 (N_2097,N_1845,N_1087);
nand U2098 (N_2098,N_1444,N_117);
and U2099 (N_2099,N_1165,N_1069);
and U2100 (N_2100,N_1386,N_1331);
and U2101 (N_2101,N_1243,N_1083);
and U2102 (N_2102,N_182,N_217);
nor U2103 (N_2103,N_868,N_235);
xor U2104 (N_2104,N_536,N_886);
and U2105 (N_2105,N_513,N_1904);
nor U2106 (N_2106,N_834,N_221);
nand U2107 (N_2107,N_210,N_992);
or U2108 (N_2108,N_196,N_407);
or U2109 (N_2109,N_1461,N_1545);
nand U2110 (N_2110,N_1251,N_853);
and U2111 (N_2111,N_1239,N_24);
and U2112 (N_2112,N_1676,N_1289);
nand U2113 (N_2113,N_1609,N_1057);
nor U2114 (N_2114,N_1034,N_1042);
nor U2115 (N_2115,N_1906,N_1803);
or U2116 (N_2116,N_1001,N_818);
nor U2117 (N_2117,N_1663,N_509);
and U2118 (N_2118,N_1075,N_1834);
and U2119 (N_2119,N_866,N_1651);
nor U2120 (N_2120,N_1159,N_468);
xor U2121 (N_2121,N_1012,N_1051);
or U2122 (N_2122,N_891,N_1659);
nor U2123 (N_2123,N_1818,N_1759);
xnor U2124 (N_2124,N_1895,N_1875);
or U2125 (N_2125,N_201,N_80);
and U2126 (N_2126,N_652,N_1050);
xor U2127 (N_2127,N_1828,N_1495);
and U2128 (N_2128,N_1880,N_643);
xor U2129 (N_2129,N_71,N_429);
nand U2130 (N_2130,N_1614,N_1);
nand U2131 (N_2131,N_1715,N_1965);
nor U2132 (N_2132,N_1560,N_940);
and U2133 (N_2133,N_1152,N_258);
nor U2134 (N_2134,N_289,N_920);
nor U2135 (N_2135,N_326,N_515);
and U2136 (N_2136,N_678,N_419);
or U2137 (N_2137,N_1747,N_1868);
xnor U2138 (N_2138,N_1852,N_1134);
and U2139 (N_2139,N_194,N_1084);
nand U2140 (N_2140,N_1425,N_487);
nand U2141 (N_2141,N_346,N_575);
nor U2142 (N_2142,N_1292,N_1650);
and U2143 (N_2143,N_319,N_197);
and U2144 (N_2144,N_440,N_1847);
and U2145 (N_2145,N_96,N_1548);
or U2146 (N_2146,N_1666,N_859);
and U2147 (N_2147,N_1951,N_1678);
nor U2148 (N_2148,N_4,N_58);
nor U2149 (N_2149,N_1841,N_43);
or U2150 (N_2150,N_687,N_1205);
or U2151 (N_2151,N_1094,N_1148);
or U2152 (N_2152,N_651,N_22);
or U2153 (N_2153,N_985,N_1234);
and U2154 (N_2154,N_967,N_420);
or U2155 (N_2155,N_479,N_318);
and U2156 (N_2156,N_1675,N_827);
and U2157 (N_2157,N_1522,N_1285);
nor U2158 (N_2158,N_152,N_638);
or U2159 (N_2159,N_1815,N_282);
nand U2160 (N_2160,N_977,N_734);
and U2161 (N_2161,N_1345,N_1181);
and U2162 (N_2162,N_735,N_709);
and U2163 (N_2163,N_1916,N_945);
and U2164 (N_2164,N_157,N_802);
nand U2165 (N_2165,N_78,N_1992);
nand U2166 (N_2166,N_1374,N_1248);
nor U2167 (N_2167,N_953,N_848);
nor U2168 (N_2168,N_1827,N_1272);
and U2169 (N_2169,N_1954,N_328);
and U2170 (N_2170,N_823,N_1218);
xor U2171 (N_2171,N_1821,N_1252);
nand U2172 (N_2172,N_1597,N_623);
or U2173 (N_2173,N_1910,N_887);
nor U2174 (N_2174,N_1691,N_1409);
and U2175 (N_2175,N_154,N_1557);
nor U2176 (N_2176,N_206,N_7);
xor U2177 (N_2177,N_386,N_1987);
nor U2178 (N_2178,N_1439,N_1564);
nand U2179 (N_2179,N_1736,N_288);
xnor U2180 (N_2180,N_211,N_1567);
and U2181 (N_2181,N_497,N_841);
nand U2182 (N_2182,N_246,N_171);
and U2183 (N_2183,N_213,N_391);
and U2184 (N_2184,N_100,N_545);
nand U2185 (N_2185,N_1127,N_1831);
or U2186 (N_2186,N_984,N_1198);
and U2187 (N_2187,N_973,N_1316);
and U2188 (N_2188,N_48,N_1279);
or U2189 (N_2189,N_824,N_1298);
nand U2190 (N_2190,N_243,N_1220);
or U2191 (N_2191,N_1222,N_67);
and U2192 (N_2192,N_1108,N_401);
or U2193 (N_2193,N_411,N_1014);
nor U2194 (N_2194,N_695,N_370);
and U2195 (N_2195,N_121,N_958);
and U2196 (N_2196,N_1440,N_1157);
and U2197 (N_2197,N_955,N_1227);
and U2198 (N_2198,N_1793,N_442);
or U2199 (N_2199,N_1350,N_1048);
nand U2200 (N_2200,N_1618,N_555);
or U2201 (N_2201,N_1915,N_600);
xor U2202 (N_2202,N_1738,N_1147);
and U2203 (N_2203,N_791,N_1854);
xnor U2204 (N_2204,N_972,N_876);
xnor U2205 (N_2205,N_209,N_885);
nor U2206 (N_2206,N_1799,N_1422);
and U2207 (N_2207,N_598,N_736);
nand U2208 (N_2208,N_507,N_1728);
and U2209 (N_2209,N_1664,N_1542);
nor U2210 (N_2210,N_290,N_1309);
or U2211 (N_2211,N_460,N_1607);
xor U2212 (N_2212,N_1777,N_1610);
or U2213 (N_2213,N_1608,N_1066);
or U2214 (N_2214,N_25,N_1346);
nor U2215 (N_2215,N_1514,N_949);
nand U2216 (N_2216,N_1231,N_1168);
nor U2217 (N_2217,N_858,N_219);
or U2218 (N_2218,N_699,N_12);
nor U2219 (N_2219,N_1076,N_53);
nor U2220 (N_2220,N_1337,N_1459);
xnor U2221 (N_2221,N_1007,N_1744);
and U2222 (N_2222,N_517,N_776);
nor U2223 (N_2223,N_11,N_1822);
and U2224 (N_2224,N_227,N_764);
nor U2225 (N_2225,N_1681,N_490);
and U2226 (N_2226,N_1537,N_1341);
nor U2227 (N_2227,N_69,N_1474);
xnor U2228 (N_2228,N_214,N_944);
nor U2229 (N_2229,N_1020,N_233);
nor U2230 (N_2230,N_1361,N_29);
or U2231 (N_2231,N_1934,N_612);
or U2232 (N_2232,N_943,N_1369);
xor U2233 (N_2233,N_719,N_204);
nor U2234 (N_2234,N_1708,N_188);
or U2235 (N_2235,N_1993,N_883);
or U2236 (N_2236,N_1859,N_1673);
nor U2237 (N_2237,N_200,N_167);
and U2238 (N_2238,N_603,N_35);
and U2239 (N_2239,N_1930,N_646);
nor U2240 (N_2240,N_1214,N_1039);
or U2241 (N_2241,N_1448,N_817);
xor U2242 (N_2242,N_1118,N_99);
and U2243 (N_2243,N_1997,N_1809);
nand U2244 (N_2244,N_1478,N_1959);
xnor U2245 (N_2245,N_554,N_1454);
or U2246 (N_2246,N_1806,N_284);
nand U2247 (N_2247,N_1842,N_1949);
or U2248 (N_2248,N_833,N_942);
nand U2249 (N_2249,N_557,N_1596);
nand U2250 (N_2250,N_1355,N_1401);
xor U2251 (N_2251,N_1184,N_1872);
nor U2252 (N_2252,N_1687,N_1253);
nand U2253 (N_2253,N_125,N_647);
nor U2254 (N_2254,N_1962,N_23);
and U2255 (N_2255,N_320,N_139);
or U2256 (N_2256,N_1458,N_783);
nand U2257 (N_2257,N_1632,N_1477);
and U2258 (N_2258,N_399,N_1990);
nor U2259 (N_2259,N_410,N_430);
nor U2260 (N_2260,N_843,N_910);
xor U2261 (N_2261,N_1843,N_295);
nand U2262 (N_2262,N_1463,N_131);
xnor U2263 (N_2263,N_939,N_1473);
and U2264 (N_2264,N_1698,N_796);
nor U2265 (N_2265,N_1848,N_1840);
or U2266 (N_2266,N_1812,N_1123);
and U2267 (N_2267,N_1344,N_1411);
nand U2268 (N_2268,N_1619,N_1208);
xnor U2269 (N_2269,N_1353,N_1233);
and U2270 (N_2270,N_1176,N_382);
or U2271 (N_2271,N_331,N_452);
or U2272 (N_2272,N_1981,N_1417);
and U2273 (N_2273,N_1964,N_323);
nand U2274 (N_2274,N_344,N_1296);
and U2275 (N_2275,N_164,N_1431);
or U2276 (N_2276,N_726,N_1695);
nand U2277 (N_2277,N_1271,N_1158);
or U2278 (N_2278,N_432,N_547);
or U2279 (N_2279,N_1499,N_1899);
or U2280 (N_2280,N_696,N_917);
and U2281 (N_2281,N_1515,N_913);
nor U2282 (N_2282,N_580,N_1430);
or U2283 (N_2283,N_1961,N_203);
and U2284 (N_2284,N_572,N_1927);
nor U2285 (N_2285,N_1013,N_94);
nand U2286 (N_2286,N_1213,N_1922);
or U2287 (N_2287,N_716,N_1186);
or U2288 (N_2288,N_74,N_1760);
or U2289 (N_2289,N_897,N_670);
xor U2290 (N_2290,N_1555,N_1811);
or U2291 (N_2291,N_241,N_679);
or U2292 (N_2292,N_1657,N_672);
or U2293 (N_2293,N_888,N_466);
and U2294 (N_2294,N_1443,N_814);
and U2295 (N_2295,N_1117,N_680);
and U2296 (N_2296,N_297,N_1447);
nand U2297 (N_2297,N_88,N_1162);
or U2298 (N_2298,N_847,N_865);
nor U2299 (N_2299,N_1041,N_496);
xor U2300 (N_2300,N_436,N_1299);
or U2301 (N_2301,N_861,N_128);
and U2302 (N_2302,N_845,N_146);
nor U2303 (N_2303,N_881,N_352);
nor U2304 (N_2304,N_564,N_180);
and U2305 (N_2305,N_1166,N_1701);
and U2306 (N_2306,N_1518,N_1779);
or U2307 (N_2307,N_1464,N_998);
or U2308 (N_2308,N_1153,N_1336);
nor U2309 (N_2309,N_609,N_1591);
xnor U2310 (N_2310,N_1260,N_601);
or U2311 (N_2311,N_1946,N_1326);
and U2312 (N_2312,N_110,N_89);
xor U2313 (N_2313,N_1704,N_1672);
and U2314 (N_2314,N_820,N_1753);
or U2315 (N_2315,N_768,N_505);
or U2316 (N_2316,N_1378,N_1128);
and U2317 (N_2317,N_427,N_995);
nand U2318 (N_2318,N_338,N_588);
nand U2319 (N_2319,N_1112,N_448);
xnor U2320 (N_2320,N_1058,N_717);
or U2321 (N_2321,N_1768,N_1052);
nand U2322 (N_2322,N_1342,N_1901);
or U2323 (N_2323,N_577,N_333);
and U2324 (N_2324,N_770,N_232);
xnor U2325 (N_2325,N_1590,N_251);
or U2326 (N_2326,N_761,N_974);
nor U2327 (N_2327,N_1772,N_1405);
and U2328 (N_2328,N_1982,N_461);
nand U2329 (N_2329,N_1343,N_927);
and U2330 (N_2330,N_816,N_383);
or U2331 (N_2331,N_1649,N_192);
nand U2332 (N_2332,N_926,N_971);
or U2333 (N_2333,N_830,N_1714);
nand U2334 (N_2334,N_1696,N_1160);
and U2335 (N_2335,N_1739,N_82);
and U2336 (N_2336,N_937,N_661);
xor U2337 (N_2337,N_1393,N_98);
nand U2338 (N_2338,N_895,N_1505);
and U2339 (N_2339,N_1053,N_62);
or U2340 (N_2340,N_395,N_1351);
nand U2341 (N_2341,N_1228,N_499);
or U2342 (N_2342,N_1623,N_1365);
nand U2343 (N_2343,N_1832,N_302);
or U2344 (N_2344,N_353,N_952);
nand U2345 (N_2345,N_1508,N_753);
xor U2346 (N_2346,N_1674,N_712);
nand U2347 (N_2347,N_1945,N_766);
and U2348 (N_2348,N_642,N_1970);
or U2349 (N_2349,N_660,N_403);
and U2350 (N_2350,N_772,N_1229);
nor U2351 (N_2351,N_1317,N_263);
nor U2352 (N_2352,N_842,N_238);
or U2353 (N_2353,N_819,N_226);
or U2354 (N_2354,N_456,N_676);
nor U2355 (N_2355,N_1028,N_677);
xor U2356 (N_2356,N_118,N_223);
nor U2357 (N_2357,N_549,N_558);
or U2358 (N_2358,N_1491,N_835);
or U2359 (N_2359,N_1426,N_376);
xor U2360 (N_2360,N_1113,N_1535);
or U2361 (N_2361,N_1503,N_1559);
or U2362 (N_2362,N_1870,N_65);
nor U2363 (N_2363,N_1242,N_270);
nor U2364 (N_2364,N_1284,N_1561);
nor U2365 (N_2365,N_805,N_629);
nor U2366 (N_2366,N_825,N_1235);
nor U2367 (N_2367,N_1022,N_1658);
nand U2368 (N_2368,N_1348,N_1423);
or U2369 (N_2369,N_627,N_228);
nand U2370 (N_2370,N_1534,N_1908);
nand U2371 (N_2371,N_708,N_86);
and U2372 (N_2372,N_160,N_546);
nor U2373 (N_2373,N_1070,N_1641);
or U2374 (N_2374,N_862,N_225);
xor U2375 (N_2375,N_1340,N_831);
nor U2376 (N_2376,N_1313,N_141);
or U2377 (N_2377,N_1400,N_1170);
and U2378 (N_2378,N_527,N_1725);
and U2379 (N_2379,N_70,N_611);
and U2380 (N_2380,N_1307,N_1138);
xnor U2381 (N_2381,N_537,N_855);
and U2382 (N_2382,N_1399,N_1270);
nor U2383 (N_2383,N_1199,N_1311);
or U2384 (N_2384,N_1390,N_1577);
or U2385 (N_2385,N_1903,N_570);
or U2386 (N_2386,N_925,N_1757);
and U2387 (N_2387,N_275,N_683);
nand U2388 (N_2388,N_449,N_854);
nand U2389 (N_2389,N_1119,N_339);
nand U2390 (N_2390,N_933,N_538);
or U2391 (N_2391,N_57,N_262);
or U2392 (N_2392,N_1403,N_1769);
nor U2393 (N_2393,N_648,N_1860);
xnor U2394 (N_2394,N_525,N_1178);
or U2395 (N_2395,N_1105,N_908);
nand U2396 (N_2396,N_590,N_46);
and U2397 (N_2397,N_16,N_159);
and U2398 (N_2398,N_155,N_552);
xor U2399 (N_2399,N_1986,N_47);
or U2400 (N_2400,N_1523,N_1866);
or U2401 (N_2401,N_1758,N_1064);
or U2402 (N_2402,N_1114,N_193);
nand U2403 (N_2403,N_898,N_1670);
nor U2404 (N_2404,N_578,N_1814);
nor U2405 (N_2405,N_1297,N_199);
nor U2406 (N_2406,N_1470,N_387);
and U2407 (N_2407,N_83,N_511);
xnor U2408 (N_2408,N_1718,N_298);
nor U2409 (N_2409,N_1653,N_907);
nor U2410 (N_2410,N_1942,N_1468);
or U2411 (N_2411,N_68,N_1204);
and U2412 (N_2412,N_1453,N_1116);
and U2413 (N_2413,N_743,N_1838);
nor U2414 (N_2414,N_1249,N_1356);
nand U2415 (N_2415,N_1767,N_437);
and U2416 (N_2416,N_1394,N_1211);
nor U2417 (N_2417,N_455,N_1969);
or U2418 (N_2418,N_1617,N_351);
or U2419 (N_2419,N_305,N_1129);
or U2420 (N_2420,N_356,N_636);
or U2421 (N_2421,N_373,N_1244);
xor U2422 (N_2422,N_1900,N_1634);
and U2423 (N_2423,N_1517,N_1643);
nor U2424 (N_2424,N_703,N_1258);
or U2425 (N_2425,N_187,N_697);
and U2426 (N_2426,N_828,N_1684);
xnor U2427 (N_2427,N_255,N_337);
nand U2428 (N_2428,N_271,N_1846);
nand U2429 (N_2429,N_49,N_1263);
and U2430 (N_2430,N_1068,N_240);
nor U2431 (N_2431,N_1869,N_357);
or U2432 (N_2432,N_574,N_113);
or U2433 (N_2433,N_143,N_1230);
xor U2434 (N_2434,N_287,N_1290);
or U2435 (N_2435,N_690,N_1541);
nor U2436 (N_2436,N_1741,N_807);
and U2437 (N_2437,N_684,N_424);
nor U2438 (N_2438,N_1709,N_312);
and U2439 (N_2439,N_173,N_987);
nor U2440 (N_2440,N_892,N_1295);
xor U2441 (N_2441,N_1631,N_1932);
and U2442 (N_2442,N_1045,N_81);
or U2443 (N_2443,N_1513,N_327);
nand U2444 (N_2444,N_711,N_1573);
nor U2445 (N_2445,N_573,N_1988);
and U2446 (N_2446,N_84,N_1000);
or U2447 (N_2447,N_1339,N_428);
xor U2448 (N_2448,N_1375,N_1533);
and U2449 (N_2449,N_1494,N_889);
and U2450 (N_2450,N_1389,N_1628);
xor U2451 (N_2451,N_1735,N_107);
and U2452 (N_2452,N_1861,N_374);
and U2453 (N_2453,N_1983,N_1876);
or U2454 (N_2454,N_309,N_1668);
nand U2455 (N_2455,N_362,N_721);
nor U2456 (N_2456,N_1929,N_626);
or U2457 (N_2457,N_1187,N_585);
xnor U2458 (N_2458,N_485,N_641);
nor U2459 (N_2459,N_581,N_1151);
and U2460 (N_2460,N_1850,N_947);
xnor U2461 (N_2461,N_60,N_1267);
and U2462 (N_2462,N_31,N_1286);
nor U2463 (N_2463,N_781,N_1140);
nand U2464 (N_2464,N_478,N_1497);
nor U2465 (N_2465,N_236,N_1584);
and U2466 (N_2466,N_457,N_681);
nand U2467 (N_2467,N_1200,N_354);
or U2468 (N_2468,N_1694,N_571);
xor U2469 (N_2469,N_304,N_170);
and U2470 (N_2470,N_1016,N_733);
nand U2471 (N_2471,N_1685,N_608);
or U2472 (N_2472,N_625,N_1382);
nor U2473 (N_2473,N_936,N_1245);
and U2474 (N_2474,N_1433,N_870);
or U2475 (N_2475,N_922,N_502);
or U2476 (N_2476,N_1268,N_195);
or U2477 (N_2477,N_1182,N_950);
xor U2478 (N_2478,N_1137,N_1817);
nor U2479 (N_2479,N_1554,N_1926);
xnor U2480 (N_2480,N_1174,N_1314);
xnor U2481 (N_2481,N_231,N_1894);
nand U2482 (N_2482,N_358,N_1720);
xor U2483 (N_2483,N_1291,N_1572);
or U2484 (N_2484,N_1892,N_912);
nand U2485 (N_2485,N_656,N_1773);
or U2486 (N_2486,N_1955,N_801);
and U2487 (N_2487,N_630,N_1125);
xor U2488 (N_2488,N_1027,N_1319);
nand U2489 (N_2489,N_1450,N_1540);
nor U2490 (N_2490,N_1082,N_142);
or U2491 (N_2491,N_518,N_1863);
nand U2492 (N_2492,N_909,N_1857);
nor U2493 (N_2493,N_207,N_257);
nor U2494 (N_2494,N_521,N_1621);
and U2495 (N_2495,N_1193,N_446);
nor U2496 (N_2496,N_718,N_1418);
nor U2497 (N_2497,N_786,N_1755);
and U2498 (N_2498,N_597,N_1702);
nor U2499 (N_2499,N_408,N_1080);
nor U2500 (N_2500,N_832,N_1787);
and U2501 (N_2501,N_33,N_970);
or U2502 (N_2502,N_692,N_1958);
xor U2503 (N_2503,N_694,N_1952);
or U2504 (N_2504,N_758,N_1451);
nor U2505 (N_2505,N_1221,N_591);
nor U2506 (N_2506,N_653,N_1330);
nor U2507 (N_2507,N_340,N_846);
nand U2508 (N_2508,N_280,N_105);
or U2509 (N_2509,N_1169,N_530);
and U2510 (N_2510,N_283,N_1033);
and U2511 (N_2511,N_1516,N_1079);
and U2512 (N_2512,N_32,N_324);
and U2513 (N_2513,N_1667,N_961);
or U2514 (N_2514,N_1636,N_1333);
nor U2515 (N_2515,N_1067,N_1574);
or U2516 (N_2516,N_594,N_821);
nand U2517 (N_2517,N_1500,N_839);
xor U2518 (N_2518,N_144,N_957);
nand U2519 (N_2519,N_431,N_882);
nor U2520 (N_2520,N_1359,N_750);
or U2521 (N_2521,N_617,N_6);
and U2522 (N_2522,N_249,N_720);
or U2523 (N_2523,N_542,N_1512);
or U2524 (N_2524,N_930,N_335);
nand U2525 (N_2525,N_434,N_903);
nand U2526 (N_2526,N_901,N_932);
nor U2527 (N_2527,N_464,N_762);
and U2528 (N_2528,N_1920,N_1784);
nor U2529 (N_2529,N_1164,N_474);
nand U2530 (N_2530,N_253,N_519);
and U2531 (N_2531,N_1726,N_122);
nor U2532 (N_2532,N_1911,N_1308);
nor U2533 (N_2533,N_176,N_1212);
nand U2534 (N_2534,N_1449,N_704);
nor U2535 (N_2535,N_1797,N_28);
or U2536 (N_2536,N_1018,N_93);
nand U2537 (N_2537,N_1829,N_166);
and U2538 (N_2538,N_1792,N_614);
nor U2539 (N_2539,N_562,N_550);
nand U2540 (N_2540,N_385,N_582);
nor U2541 (N_2541,N_264,N_278);
nand U2542 (N_2542,N_27,N_1115);
nand U2543 (N_2543,N_829,N_1420);
xnor U2544 (N_2544,N_145,N_1397);
nor U2545 (N_2545,N_622,N_414);
nand U2546 (N_2546,N_1141,N_568);
or U2547 (N_2547,N_347,N_644);
and U2548 (N_2548,N_277,N_1038);
and U2549 (N_2549,N_778,N_137);
and U2550 (N_2550,N_1917,N_938);
or U2551 (N_2551,N_1074,N_465);
nor U2552 (N_2552,N_425,N_1871);
and U2553 (N_2553,N_1238,N_13);
and U2554 (N_2554,N_968,N_242);
or U2555 (N_2555,N_837,N_1281);
and U2556 (N_2556,N_1009,N_946);
xor U2557 (N_2557,N_97,N_38);
xnor U2558 (N_2558,N_1975,N_1412);
or U2559 (N_2559,N_1862,N_918);
and U2560 (N_2560,N_808,N_760);
or U2561 (N_2561,N_1923,N_1132);
xor U2562 (N_2562,N_1255,N_795);
and U2563 (N_2563,N_1524,N_1665);
or U2564 (N_2564,N_1081,N_548);
nor U2565 (N_2565,N_106,N_1578);
nor U2566 (N_2566,N_1586,N_415);
or U2567 (N_2567,N_1644,N_1730);
nor U2568 (N_2568,N_873,N_404);
nand U2569 (N_2569,N_806,N_640);
xnor U2570 (N_2570,N_701,N_1700);
or U2571 (N_2571,N_397,N_1977);
nand U2572 (N_2572,N_1810,N_398);
and U2573 (N_2573,N_844,N_1858);
nand U2574 (N_2574,N_1312,N_1032);
nor U2575 (N_2575,N_746,N_61);
nand U2576 (N_2576,N_1604,N_310);
and U2577 (N_2577,N_1156,N_1963);
or U2578 (N_2578,N_1527,N_1531);
xnor U2579 (N_2579,N_1024,N_1802);
nor U2580 (N_2580,N_329,N_710);
nand U2581 (N_2581,N_663,N_1250);
nand U2582 (N_2582,N_1177,N_1998);
and U2583 (N_2583,N_239,N_1824);
and U2584 (N_2584,N_975,N_1471);
nand U2585 (N_2585,N_1324,N_1480);
and U2586 (N_2586,N_394,N_147);
nor U2587 (N_2587,N_619,N_1794);
and U2588 (N_2588,N_528,N_1202);
and U2589 (N_2589,N_951,N_473);
nor U2590 (N_2590,N_1192,N_1492);
xor U2591 (N_2591,N_1780,N_1950);
and U2592 (N_2592,N_797,N_1215);
and U2593 (N_2593,N_1724,N_1481);
or U2594 (N_2594,N_111,N_637);
nor U2595 (N_2595,N_956,N_645);
nand U2596 (N_2596,N_1947,N_1269);
nor U2597 (N_2597,N_254,N_1732);
nand U2598 (N_2598,N_822,N_1428);
or U2599 (N_2599,N_1778,N_1801);
nor U2600 (N_2600,N_1598,N_300);
and U2601 (N_2601,N_39,N_1960);
xnor U2602 (N_2602,N_8,N_1530);
and U2603 (N_2603,N_444,N_867);
or U2604 (N_2604,N_205,N_393);
xnor U2605 (N_2605,N_931,N_1421);
or U2606 (N_2606,N_109,N_1893);
nor U2607 (N_2607,N_349,N_112);
or U2608 (N_2608,N_1835,N_1568);
and U2609 (N_2609,N_174,N_639);
nor U2610 (N_2610,N_1370,N_1722);
nor U2611 (N_2611,N_230,N_1354);
nor U2612 (N_2612,N_212,N_755);
nor U2613 (N_2613,N_481,N_1122);
or U2614 (N_2614,N_384,N_838);
xor U2615 (N_2615,N_261,N_79);
nor U2616 (N_2616,N_1774,N_1367);
nand U2617 (N_2617,N_875,N_1179);
nor U2618 (N_2618,N_45,N_1576);
xor U2619 (N_2619,N_579,N_979);
and U2620 (N_2620,N_104,N_864);
nor U2621 (N_2621,N_21,N_739);
xor U2622 (N_2622,N_799,N_1967);
or U2623 (N_2623,N_1465,N_731);
and U2624 (N_2624,N_740,N_1569);
and U2625 (N_2625,N_269,N_602);
or U2626 (N_2626,N_905,N_1823);
nor U2627 (N_2627,N_1550,N_1553);
and U2628 (N_2628,N_1133,N_489);
or U2629 (N_2629,N_1130,N_658);
or U2630 (N_2630,N_1839,N_350);
or U2631 (N_2631,N_501,N_1844);
nand U2632 (N_2632,N_1690,N_1788);
and U2633 (N_2633,N_30,N_506);
and U2634 (N_2634,N_948,N_299);
or U2635 (N_2635,N_1410,N_52);
and U2636 (N_2636,N_1381,N_544);
and U2637 (N_2637,N_1750,N_706);
and U2638 (N_2638,N_467,N_779);
and U2639 (N_2639,N_73,N_1413);
or U2640 (N_2640,N_662,N_1913);
nor U2641 (N_2641,N_1335,N_422);
or U2642 (N_2642,N_1183,N_1438);
nor U2643 (N_2643,N_1098,N_798);
nor U2644 (N_2644,N_1120,N_1049);
nor U2645 (N_2645,N_1520,N_1763);
and U2646 (N_2646,N_1647,N_1936);
or U2647 (N_2647,N_890,N_161);
nand U2648 (N_2648,N_1746,N_524);
or U2649 (N_2649,N_364,N_1710);
or U2650 (N_2650,N_1320,N_934);
xnor U2651 (N_2651,N_771,N_921);
nor U2652 (N_2652,N_978,N_1404);
nand U2653 (N_2653,N_1571,N_878);
nor U2654 (N_2654,N_1010,N_869);
or U2655 (N_2655,N_732,N_0);
or U2656 (N_2656,N_495,N_279);
or U2657 (N_2657,N_782,N_1790);
nor U2658 (N_2658,N_1655,N_792);
and U2659 (N_2659,N_982,N_773);
nand U2660 (N_2660,N_1195,N_765);
nor U2661 (N_2661,N_560,N_1379);
or U2662 (N_2662,N_812,N_412);
nand U2663 (N_2663,N_1529,N_367);
or U2664 (N_2664,N_149,N_1240);
nand U2665 (N_2665,N_165,N_1146);
and U2666 (N_2666,N_1486,N_1912);
or U2667 (N_2667,N_95,N_744);
or U2668 (N_2668,N_1754,N_532);
or U2669 (N_2669,N_1600,N_1507);
or U2670 (N_2670,N_1940,N_1154);
nand U2671 (N_2671,N_1482,N_1462);
nor U2672 (N_2672,N_793,N_1743);
nand U2673 (N_2673,N_1008,N_162);
and U2674 (N_2674,N_1971,N_1306);
or U2675 (N_2675,N_1616,N_1424);
or U2676 (N_2676,N_1721,N_512);
nor U2677 (N_2677,N_1264,N_1246);
and U2678 (N_2678,N_1669,N_1974);
nor U2679 (N_2679,N_1985,N_1939);
nand U2680 (N_2680,N_1979,N_705);
or U2681 (N_2681,N_693,N_87);
or U2682 (N_2682,N_686,N_1364);
xor U2683 (N_2683,N_923,N_757);
or U2684 (N_2684,N_655,N_1677);
or U2685 (N_2685,N_454,N_120);
xor U2686 (N_2686,N_1999,N_1031);
nand U2687 (N_2687,N_902,N_1484);
and U2688 (N_2688,N_1216,N_1888);
nor U2689 (N_2689,N_1223,N_1606);
or U2690 (N_2690,N_1217,N_1310);
and U2691 (N_2691,N_291,N_1539);
nand U2692 (N_2692,N_1782,N_1100);
nor U2693 (N_2693,N_1460,N_728);
or U2694 (N_2694,N_169,N_569);
nor U2695 (N_2695,N_1101,N_342);
nor U2696 (N_2696,N_650,N_1662);
and U2697 (N_2697,N_1011,N_748);
or U2698 (N_2698,N_1037,N_1622);
xor U2699 (N_2699,N_1036,N_1489);
and U2700 (N_2700,N_1825,N_1435);
nor U2701 (N_2701,N_566,N_576);
xor U2702 (N_2702,N_1090,N_1338);
xnor U2703 (N_2703,N_124,N_135);
xor U2704 (N_2704,N_988,N_1973);
and U2705 (N_2705,N_1088,N_1761);
nand U2706 (N_2706,N_698,N_1836);
nor U2707 (N_2707,N_1771,N_482);
or U2708 (N_2708,N_1475,N_216);
nor U2709 (N_2709,N_685,N_453);
nand U2710 (N_2710,N_1237,N_19);
and U2711 (N_2711,N_1347,N_423);
or U2712 (N_2712,N_1149,N_1826);
or U2713 (N_2713,N_1630,N_368);
nor U2714 (N_2714,N_1633,N_1071);
nand U2715 (N_2715,N_664,N_871);
or U2716 (N_2716,N_1867,N_294);
or U2717 (N_2717,N_1171,N_1785);
xnor U2718 (N_2718,N_92,N_470);
nand U2719 (N_2719,N_252,N_1175);
and U2720 (N_2720,N_229,N_369);
nand U2721 (N_2721,N_666,N_1392);
xor U2722 (N_2722,N_738,N_1611);
and U2723 (N_2723,N_586,N_1257);
xnor U2724 (N_2724,N_1795,N_1328);
or U2725 (N_2725,N_488,N_265);
nand U2726 (N_2726,N_1196,N_713);
nand U2727 (N_2727,N_475,N_691);
or U2728 (N_2728,N_1878,N_996);
and U2729 (N_2729,N_965,N_535);
nand U2730 (N_2730,N_742,N_1136);
and U2731 (N_2731,N_669,N_1642);
nor U2732 (N_2732,N_788,N_1055);
nor U2733 (N_2733,N_498,N_378);
xor U2734 (N_2734,N_1620,N_5);
and U2735 (N_2735,N_462,N_1256);
or U2736 (N_2736,N_1775,N_116);
nand U2737 (N_2737,N_1109,N_1807);
xor U2738 (N_2738,N_1005,N_1483);
xnor U2739 (N_2739,N_1124,N_813);
and U2740 (N_2740,N_775,N_1883);
nor U2741 (N_2741,N_899,N_1427);
or U2742 (N_2742,N_2,N_190);
or U2743 (N_2743,N_365,N_729);
xnor U2744 (N_2744,N_1302,N_520);
and U2745 (N_2745,N_1717,N_1501);
nor U2746 (N_2746,N_1887,N_1646);
nand U2747 (N_2747,N_1003,N_1407);
nand U2748 (N_2748,N_1197,N_1191);
and U2749 (N_2749,N_1030,N_1830);
and U2750 (N_2750,N_1388,N_50);
or U2751 (N_2751,N_1808,N_1173);
nor U2752 (N_2752,N_1266,N_72);
nor U2753 (N_2753,N_153,N_1487);
or U2754 (N_2754,N_1368,N_1521);
and U2755 (N_2755,N_1656,N_1697);
nor U2756 (N_2756,N_1396,N_259);
or U2757 (N_2757,N_409,N_1093);
xor U2758 (N_2758,N_1274,N_76);
or U2759 (N_2759,N_450,N_15);
or U2760 (N_2760,N_1789,N_1275);
or U2761 (N_2761,N_1601,N_286);
nor U2762 (N_2762,N_439,N_674);
nand U2763 (N_2763,N_245,N_1980);
xnor U2764 (N_2764,N_631,N_1023);
nand U2765 (N_2765,N_1391,N_1092);
nor U2766 (N_2766,N_123,N_268);
nor U2767 (N_2767,N_1360,N_784);
nand U2768 (N_2768,N_959,N_1321);
xnor U2769 (N_2769,N_789,N_707);
nand U2770 (N_2770,N_593,N_754);
and U2771 (N_2771,N_1851,N_471);
or U2772 (N_2772,N_379,N_1740);
and U2773 (N_2773,N_999,N_983);
or U2774 (N_2774,N_273,N_880);
nand U2775 (N_2775,N_1416,N_514);
and U2776 (N_2776,N_809,N_156);
or U2777 (N_2777,N_1538,N_325);
or U2778 (N_2778,N_635,N_906);
nor U2779 (N_2779,N_311,N_102);
nor U2780 (N_2780,N_1476,N_1377);
nor U2781 (N_2781,N_272,N_1363);
or U2782 (N_2782,N_1043,N_1896);
nand U2783 (N_2783,N_1587,N_1224);
or U2784 (N_2784,N_1210,N_1472);
nor U2785 (N_2785,N_1645,N_1318);
or U2786 (N_2786,N_1303,N_1509);
or U2787 (N_2787,N_438,N_1060);
and U2788 (N_2788,N_371,N_1994);
and U2789 (N_2789,N_790,N_285);
or U2790 (N_2790,N_1976,N_1054);
or U2791 (N_2791,N_924,N_1699);
nand U2792 (N_2792,N_37,N_1978);
or U2793 (N_2793,N_1029,N_1624);
nor U2794 (N_2794,N_1599,N_1671);
nor U2795 (N_2795,N_1693,N_1711);
nand U2796 (N_2796,N_1532,N_1941);
and U2797 (N_2797,N_877,N_1918);
and U2798 (N_2798,N_522,N_1528);
nand U2799 (N_2799,N_1956,N_17);
or U2800 (N_2800,N_1581,N_1398);
or U2801 (N_2801,N_218,N_1167);
or U2802 (N_2802,N_59,N_1155);
nand U2803 (N_2803,N_1781,N_749);
and U2804 (N_2804,N_55,N_1731);
nor U2805 (N_2805,N_1706,N_1592);
nand U2806 (N_2806,N_1705,N_1025);
nand U2807 (N_2807,N_1547,N_1061);
and U2808 (N_2808,N_1881,N_1349);
xor U2809 (N_2809,N_767,N_1322);
or U2810 (N_2810,N_1021,N_565);
or U2811 (N_2811,N_1362,N_9);
or U2812 (N_2812,N_314,N_301);
and U2813 (N_2813,N_1456,N_1686);
xor U2814 (N_2814,N_1002,N_375);
nor U2815 (N_2815,N_14,N_1247);
and U2816 (N_2816,N_108,N_250);
or U2817 (N_2817,N_929,N_1886);
or U2818 (N_2818,N_476,N_1019);
or U2819 (N_2819,N_604,N_163);
nor U2820 (N_2820,N_1948,N_724);
nand U2821 (N_2821,N_266,N_1161);
nand U2822 (N_2822,N_1583,N_654);
and U2823 (N_2823,N_1469,N_34);
nor U2824 (N_2824,N_583,N_563);
nand U2825 (N_2825,N_904,N_1261);
xor U2826 (N_2826,N_40,N_1579);
nor U2827 (N_2827,N_1226,N_1063);
nand U2828 (N_2828,N_202,N_1919);
nor U2829 (N_2829,N_151,N_1637);
or U2830 (N_2830,N_1383,N_1745);
nor U2831 (N_2831,N_659,N_18);
xor U2832 (N_2832,N_1849,N_508);
and U2833 (N_2833,N_689,N_1907);
and U2834 (N_2834,N_1877,N_1194);
nor U2835 (N_2835,N_567,N_1357);
or U2836 (N_2836,N_1688,N_860);
nor U2837 (N_2837,N_1996,N_1924);
xor U2838 (N_2838,N_966,N_990);
nor U2839 (N_2839,N_26,N_1689);
or U2840 (N_2840,N_850,N_51);
and U2841 (N_2841,N_991,N_1640);
nand U2842 (N_2842,N_1163,N_1626);
and U2843 (N_2843,N_244,N_1536);
or U2844 (N_2844,N_134,N_361);
nor U2845 (N_2845,N_1589,N_529);
or U2846 (N_2846,N_531,N_179);
nand U2847 (N_2847,N_1106,N_1395);
nor U2848 (N_2848,N_1280,N_667);
nand U2849 (N_2849,N_1301,N_66);
nand U2850 (N_2850,N_140,N_1593);
nor U2851 (N_2851,N_1294,N_1995);
and U2852 (N_2852,N_1062,N_150);
or U2853 (N_2853,N_1820,N_1928);
and U2854 (N_2854,N_1455,N_702);
xor U2855 (N_2855,N_1099,N_589);
nor U2856 (N_2856,N_1415,N_390);
nand U2857 (N_2857,N_774,N_1766);
xor U2858 (N_2858,N_1466,N_1921);
and U2859 (N_2859,N_804,N_1441);
and U2860 (N_2860,N_682,N_54);
or U2861 (N_2861,N_541,N_1277);
and U2862 (N_2862,N_1077,N_1510);
and U2863 (N_2863,N_281,N_1733);
nor U2864 (N_2864,N_620,N_158);
nor U2865 (N_2865,N_1485,N_1059);
nand U2866 (N_2866,N_986,N_1627);
nor U2867 (N_2867,N_1006,N_360);
nand U2868 (N_2868,N_1089,N_673);
or U2869 (N_2869,N_292,N_752);
nand U2870 (N_2870,N_815,N_316);
xor U2871 (N_2871,N_1467,N_747);
xor U2872 (N_2872,N_1953,N_1935);
and U2873 (N_2873,N_1046,N_759);
nor U2874 (N_2874,N_372,N_1209);
nor U2875 (N_2875,N_1805,N_402);
nor U2876 (N_2876,N_1723,N_1366);
or U2877 (N_2877,N_849,N_914);
and U2878 (N_2878,N_451,N_396);
nor U2879 (N_2879,N_551,N_91);
and U2880 (N_2880,N_587,N_1853);
nor U2881 (N_2881,N_1504,N_363);
xnor U2882 (N_2882,N_1189,N_491);
nor U2883 (N_2883,N_191,N_1800);
nand U2884 (N_2884,N_260,N_484);
nand U2885 (N_2885,N_1135,N_1445);
xnor U2886 (N_2886,N_1190,N_1756);
nand U2887 (N_2887,N_248,N_172);
nand U2888 (N_2888,N_413,N_336);
nor U2889 (N_2889,N_1873,N_168);
xor U2890 (N_2890,N_1909,N_317);
nand U2891 (N_2891,N_1432,N_503);
or U2892 (N_2892,N_1612,N_330);
xor U2893 (N_2893,N_1107,N_785);
nor U2894 (N_2894,N_592,N_1751);
or U2895 (N_2895,N_400,N_980);
xor U2896 (N_2896,N_1833,N_803);
nor U2897 (N_2897,N_63,N_1387);
nand U2898 (N_2898,N_836,N_3);
nand U2899 (N_2899,N_810,N_186);
and U2900 (N_2900,N_127,N_874);
and U2901 (N_2901,N_469,N_1017);
or U2902 (N_2902,N_1236,N_1648);
nand U2903 (N_2903,N_1283,N_388);
or U2904 (N_2904,N_177,N_1680);
or U2905 (N_2905,N_181,N_935);
or U2906 (N_2906,N_1615,N_928);
nand U2907 (N_2907,N_879,N_1712);
nor U2908 (N_2908,N_1588,N_1185);
nand U2909 (N_2909,N_1629,N_1004);
or U2910 (N_2910,N_657,N_1488);
and U2911 (N_2911,N_426,N_1373);
and U2912 (N_2912,N_1925,N_561);
or U2913 (N_2913,N_763,N_138);
and U2914 (N_2914,N_130,N_1716);
or U2915 (N_2915,N_224,N_756);
nand U2916 (N_2916,N_1585,N_41);
and U2917 (N_2917,N_293,N_852);
nand U2918 (N_2918,N_1902,N_1526);
nand U2919 (N_2919,N_1293,N_380);
or U2920 (N_2920,N_459,N_44);
or U2921 (N_2921,N_1446,N_1874);
nor U2922 (N_2922,N_315,N_178);
and U2923 (N_2923,N_256,N_1091);
nor U2924 (N_2924,N_1131,N_1144);
nand U2925 (N_2925,N_628,N_1968);
and U2926 (N_2926,N_634,N_688);
or U2927 (N_2927,N_911,N_1327);
and U2928 (N_2928,N_1142,N_215);
nand U2929 (N_2929,N_1493,N_1273);
nor U2930 (N_2930,N_1219,N_1544);
nand U2931 (N_2931,N_334,N_1729);
and U2932 (N_2932,N_1072,N_1966);
or U2933 (N_2933,N_75,N_1150);
nand U2934 (N_2934,N_964,N_1734);
nor U2935 (N_2935,N_441,N_584);
nand U2936 (N_2936,N_510,N_1819);
and U2937 (N_2937,N_1325,N_1262);
and U2938 (N_2938,N_884,N_976);
xor U2939 (N_2939,N_1429,N_406);
nand U2940 (N_2940,N_826,N_1816);
nand U2941 (N_2941,N_486,N_1203);
nor U2942 (N_2942,N_1315,N_1519);
or U2943 (N_2943,N_343,N_492);
nor U2944 (N_2944,N_1352,N_1582);
or U2945 (N_2945,N_1323,N_1972);
xnor U2946 (N_2946,N_1884,N_1278);
and U2947 (N_2947,N_1703,N_20);
xnor U2948 (N_2948,N_1933,N_840);
nand U2949 (N_2949,N_1551,N_1865);
and U2950 (N_2950,N_1796,N_276);
or U2951 (N_2951,N_1143,N_1047);
xor U2952 (N_2952,N_800,N_1682);
nor U2953 (N_2953,N_115,N_1201);
and U2954 (N_2954,N_1570,N_493);
or U2955 (N_2955,N_1111,N_1748);
nor U2956 (N_2956,N_1265,N_553);
xor U2957 (N_2957,N_267,N_1408);
or U2958 (N_2958,N_1254,N_418);
or U2959 (N_2959,N_993,N_1402);
and U2960 (N_2960,N_208,N_90);
xor U2961 (N_2961,N_1891,N_777);
nor U2962 (N_2962,N_989,N_1225);
or U2963 (N_2963,N_480,N_1380);
or U2964 (N_2964,N_1625,N_504);
nand U2965 (N_2965,N_751,N_633);
nor U2966 (N_2966,N_1661,N_1511);
or U2967 (N_2967,N_1707,N_1943);
or U2968 (N_2968,N_443,N_341);
or U2969 (N_2969,N_1406,N_559);
or U2970 (N_2970,N_389,N_1206);
or U2971 (N_2971,N_1856,N_1984);
or U2972 (N_2972,N_1742,N_1288);
or U2973 (N_2973,N_1566,N_1496);
or U2974 (N_2974,N_1282,N_1502);
or U2975 (N_2975,N_103,N_1372);
and U2976 (N_2976,N_56,N_184);
xor U2977 (N_2977,N_893,N_616);
nand U2978 (N_2978,N_856,N_523);
and U2979 (N_2979,N_1556,N_607);
xor U2980 (N_2980,N_296,N_1605);
nand U2981 (N_2981,N_1679,N_1562);
nand U2982 (N_2982,N_1026,N_1764);
nand U2983 (N_2983,N_1035,N_919);
nand U2984 (N_2984,N_1056,N_624);
xnor U2985 (N_2985,N_1879,N_1095);
nor U2986 (N_2986,N_851,N_185);
nor U2987 (N_2987,N_1565,N_313);
or U2988 (N_2988,N_355,N_1241);
nand U2989 (N_2989,N_794,N_183);
or U2990 (N_2990,N_605,N_1332);
or U2991 (N_2991,N_189,N_1525);
nand U2992 (N_2992,N_540,N_1786);
xor U2993 (N_2993,N_1121,N_416);
nor U2994 (N_2994,N_730,N_1898);
nor U2995 (N_2995,N_381,N_1752);
nor U2996 (N_2996,N_1207,N_1804);
nand U2997 (N_2997,N_941,N_500);
nor U2998 (N_2998,N_1635,N_1580);
or U2999 (N_2999,N_1180,N_723);
xor U3000 (N_3000,N_1237,N_1661);
or U3001 (N_3001,N_948,N_1952);
nor U3002 (N_3002,N_1794,N_330);
or U3003 (N_3003,N_1086,N_1129);
nand U3004 (N_3004,N_1636,N_1907);
and U3005 (N_3005,N_448,N_1835);
xor U3006 (N_3006,N_494,N_302);
nand U3007 (N_3007,N_1579,N_304);
and U3008 (N_3008,N_762,N_525);
and U3009 (N_3009,N_1262,N_776);
and U3010 (N_3010,N_208,N_498);
and U3011 (N_3011,N_31,N_1242);
or U3012 (N_3012,N_1721,N_441);
or U3013 (N_3013,N_1044,N_1875);
nor U3014 (N_3014,N_36,N_1060);
xor U3015 (N_3015,N_816,N_1244);
or U3016 (N_3016,N_561,N_405);
nand U3017 (N_3017,N_154,N_853);
nand U3018 (N_3018,N_1879,N_1273);
nor U3019 (N_3019,N_796,N_1898);
nor U3020 (N_3020,N_1481,N_171);
nor U3021 (N_3021,N_484,N_792);
or U3022 (N_3022,N_954,N_1023);
or U3023 (N_3023,N_1893,N_1239);
or U3024 (N_3024,N_813,N_1660);
or U3025 (N_3025,N_1935,N_454);
nor U3026 (N_3026,N_825,N_1068);
nand U3027 (N_3027,N_64,N_646);
xor U3028 (N_3028,N_862,N_671);
or U3029 (N_3029,N_602,N_342);
nor U3030 (N_3030,N_1432,N_1719);
and U3031 (N_3031,N_531,N_1536);
and U3032 (N_3032,N_1593,N_995);
and U3033 (N_3033,N_850,N_186);
nor U3034 (N_3034,N_1596,N_1373);
nand U3035 (N_3035,N_323,N_1409);
nor U3036 (N_3036,N_437,N_679);
nor U3037 (N_3037,N_1810,N_734);
nor U3038 (N_3038,N_1814,N_866);
and U3039 (N_3039,N_1561,N_222);
and U3040 (N_3040,N_56,N_117);
xor U3041 (N_3041,N_1618,N_1999);
and U3042 (N_3042,N_1771,N_15);
or U3043 (N_3043,N_56,N_1203);
and U3044 (N_3044,N_58,N_117);
or U3045 (N_3045,N_1395,N_934);
or U3046 (N_3046,N_1761,N_893);
or U3047 (N_3047,N_628,N_177);
nand U3048 (N_3048,N_1070,N_1707);
and U3049 (N_3049,N_1066,N_1897);
or U3050 (N_3050,N_1980,N_193);
or U3051 (N_3051,N_1361,N_1608);
and U3052 (N_3052,N_379,N_28);
nand U3053 (N_3053,N_1539,N_849);
and U3054 (N_3054,N_412,N_1529);
nor U3055 (N_3055,N_1774,N_968);
and U3056 (N_3056,N_1191,N_1281);
or U3057 (N_3057,N_694,N_243);
and U3058 (N_3058,N_513,N_528);
and U3059 (N_3059,N_1254,N_958);
or U3060 (N_3060,N_1314,N_153);
and U3061 (N_3061,N_1426,N_1955);
or U3062 (N_3062,N_16,N_1690);
or U3063 (N_3063,N_898,N_932);
or U3064 (N_3064,N_219,N_1923);
or U3065 (N_3065,N_601,N_187);
nand U3066 (N_3066,N_495,N_1997);
and U3067 (N_3067,N_810,N_147);
nand U3068 (N_3068,N_1301,N_394);
and U3069 (N_3069,N_1222,N_829);
nand U3070 (N_3070,N_347,N_432);
and U3071 (N_3071,N_1482,N_1718);
or U3072 (N_3072,N_1121,N_542);
or U3073 (N_3073,N_354,N_993);
nand U3074 (N_3074,N_1910,N_1983);
nor U3075 (N_3075,N_905,N_983);
or U3076 (N_3076,N_1309,N_1103);
nor U3077 (N_3077,N_1925,N_533);
nor U3078 (N_3078,N_1218,N_624);
nor U3079 (N_3079,N_259,N_440);
or U3080 (N_3080,N_1546,N_98);
or U3081 (N_3081,N_367,N_1435);
nor U3082 (N_3082,N_1414,N_1685);
nand U3083 (N_3083,N_580,N_1485);
nand U3084 (N_3084,N_577,N_1760);
or U3085 (N_3085,N_389,N_920);
nand U3086 (N_3086,N_327,N_783);
and U3087 (N_3087,N_303,N_1431);
xor U3088 (N_3088,N_276,N_1399);
nor U3089 (N_3089,N_1198,N_1526);
nand U3090 (N_3090,N_1322,N_1136);
and U3091 (N_3091,N_610,N_85);
nor U3092 (N_3092,N_1836,N_1042);
and U3093 (N_3093,N_981,N_1321);
and U3094 (N_3094,N_1961,N_1379);
or U3095 (N_3095,N_1018,N_663);
and U3096 (N_3096,N_51,N_1097);
or U3097 (N_3097,N_19,N_587);
nand U3098 (N_3098,N_1246,N_745);
nor U3099 (N_3099,N_1874,N_832);
nor U3100 (N_3100,N_443,N_1255);
and U3101 (N_3101,N_82,N_1125);
and U3102 (N_3102,N_1062,N_1339);
nand U3103 (N_3103,N_1860,N_1039);
nand U3104 (N_3104,N_1695,N_1946);
nor U3105 (N_3105,N_1804,N_927);
nor U3106 (N_3106,N_1002,N_1728);
nand U3107 (N_3107,N_1083,N_638);
nor U3108 (N_3108,N_1891,N_168);
or U3109 (N_3109,N_73,N_1929);
nand U3110 (N_3110,N_723,N_1385);
nor U3111 (N_3111,N_476,N_1225);
or U3112 (N_3112,N_1292,N_193);
xnor U3113 (N_3113,N_1583,N_144);
and U3114 (N_3114,N_955,N_65);
and U3115 (N_3115,N_264,N_1473);
or U3116 (N_3116,N_363,N_1686);
or U3117 (N_3117,N_720,N_912);
or U3118 (N_3118,N_1164,N_1776);
and U3119 (N_3119,N_1296,N_146);
nand U3120 (N_3120,N_774,N_107);
nor U3121 (N_3121,N_737,N_1690);
nor U3122 (N_3122,N_1962,N_536);
or U3123 (N_3123,N_285,N_1247);
and U3124 (N_3124,N_303,N_1079);
and U3125 (N_3125,N_281,N_1148);
nand U3126 (N_3126,N_266,N_1977);
nor U3127 (N_3127,N_1480,N_1190);
or U3128 (N_3128,N_40,N_407);
nor U3129 (N_3129,N_426,N_589);
and U3130 (N_3130,N_560,N_1059);
or U3131 (N_3131,N_1747,N_1394);
or U3132 (N_3132,N_378,N_1874);
nor U3133 (N_3133,N_1212,N_708);
nand U3134 (N_3134,N_1082,N_1200);
or U3135 (N_3135,N_283,N_1825);
nand U3136 (N_3136,N_1059,N_283);
and U3137 (N_3137,N_604,N_1938);
nand U3138 (N_3138,N_1971,N_12);
nor U3139 (N_3139,N_1713,N_821);
or U3140 (N_3140,N_657,N_1491);
nand U3141 (N_3141,N_50,N_1344);
nand U3142 (N_3142,N_278,N_305);
xor U3143 (N_3143,N_1230,N_592);
nand U3144 (N_3144,N_1975,N_1941);
nor U3145 (N_3145,N_1718,N_1120);
nor U3146 (N_3146,N_1125,N_1986);
and U3147 (N_3147,N_923,N_67);
or U3148 (N_3148,N_1485,N_65);
nand U3149 (N_3149,N_1682,N_1198);
nor U3150 (N_3150,N_391,N_38);
or U3151 (N_3151,N_1151,N_618);
nor U3152 (N_3152,N_1512,N_672);
and U3153 (N_3153,N_1989,N_138);
or U3154 (N_3154,N_255,N_925);
nand U3155 (N_3155,N_298,N_207);
and U3156 (N_3156,N_1136,N_542);
or U3157 (N_3157,N_102,N_71);
nor U3158 (N_3158,N_217,N_1597);
and U3159 (N_3159,N_1257,N_1496);
nand U3160 (N_3160,N_1330,N_1427);
nand U3161 (N_3161,N_1193,N_921);
nand U3162 (N_3162,N_44,N_62);
nand U3163 (N_3163,N_1450,N_1932);
xnor U3164 (N_3164,N_1782,N_1093);
or U3165 (N_3165,N_1997,N_39);
and U3166 (N_3166,N_111,N_47);
and U3167 (N_3167,N_1093,N_1521);
and U3168 (N_3168,N_1242,N_1239);
nor U3169 (N_3169,N_357,N_1513);
nand U3170 (N_3170,N_1933,N_916);
xor U3171 (N_3171,N_1924,N_1785);
nor U3172 (N_3172,N_871,N_1661);
and U3173 (N_3173,N_1242,N_1613);
and U3174 (N_3174,N_778,N_234);
xor U3175 (N_3175,N_484,N_1153);
or U3176 (N_3176,N_1648,N_1363);
or U3177 (N_3177,N_709,N_1076);
nand U3178 (N_3178,N_385,N_234);
nand U3179 (N_3179,N_935,N_1693);
or U3180 (N_3180,N_1131,N_804);
nor U3181 (N_3181,N_1231,N_1321);
nand U3182 (N_3182,N_1799,N_46);
xor U3183 (N_3183,N_1073,N_134);
and U3184 (N_3184,N_1787,N_302);
and U3185 (N_3185,N_1480,N_1548);
or U3186 (N_3186,N_637,N_1578);
nand U3187 (N_3187,N_1804,N_728);
nand U3188 (N_3188,N_233,N_1829);
nand U3189 (N_3189,N_362,N_1661);
nand U3190 (N_3190,N_1326,N_1332);
xor U3191 (N_3191,N_1890,N_1463);
and U3192 (N_3192,N_258,N_1908);
and U3193 (N_3193,N_256,N_1038);
xor U3194 (N_3194,N_932,N_977);
or U3195 (N_3195,N_901,N_1016);
xnor U3196 (N_3196,N_555,N_887);
nor U3197 (N_3197,N_724,N_1352);
xor U3198 (N_3198,N_172,N_1737);
xnor U3199 (N_3199,N_912,N_1754);
nor U3200 (N_3200,N_867,N_420);
nand U3201 (N_3201,N_1423,N_969);
and U3202 (N_3202,N_1229,N_332);
and U3203 (N_3203,N_412,N_707);
or U3204 (N_3204,N_1068,N_455);
and U3205 (N_3205,N_577,N_414);
and U3206 (N_3206,N_325,N_588);
xor U3207 (N_3207,N_1276,N_1566);
nand U3208 (N_3208,N_197,N_227);
or U3209 (N_3209,N_436,N_1016);
or U3210 (N_3210,N_665,N_91);
nand U3211 (N_3211,N_549,N_317);
nor U3212 (N_3212,N_950,N_995);
and U3213 (N_3213,N_1931,N_1481);
and U3214 (N_3214,N_1560,N_1147);
xor U3215 (N_3215,N_1633,N_1563);
nor U3216 (N_3216,N_1695,N_1515);
and U3217 (N_3217,N_506,N_1304);
xor U3218 (N_3218,N_90,N_197);
or U3219 (N_3219,N_296,N_204);
nor U3220 (N_3220,N_1221,N_1984);
or U3221 (N_3221,N_476,N_1071);
nand U3222 (N_3222,N_1217,N_1876);
nor U3223 (N_3223,N_718,N_1542);
nor U3224 (N_3224,N_1375,N_644);
nand U3225 (N_3225,N_164,N_1608);
nor U3226 (N_3226,N_122,N_1012);
or U3227 (N_3227,N_288,N_833);
nor U3228 (N_3228,N_726,N_1510);
nand U3229 (N_3229,N_71,N_947);
nand U3230 (N_3230,N_602,N_1561);
nor U3231 (N_3231,N_1775,N_1684);
or U3232 (N_3232,N_479,N_1816);
or U3233 (N_3233,N_1870,N_249);
and U3234 (N_3234,N_613,N_231);
xor U3235 (N_3235,N_812,N_930);
and U3236 (N_3236,N_181,N_1601);
nand U3237 (N_3237,N_371,N_1131);
nand U3238 (N_3238,N_1980,N_1402);
nand U3239 (N_3239,N_761,N_557);
nor U3240 (N_3240,N_650,N_63);
and U3241 (N_3241,N_962,N_417);
and U3242 (N_3242,N_1581,N_947);
or U3243 (N_3243,N_1351,N_367);
nand U3244 (N_3244,N_929,N_640);
nor U3245 (N_3245,N_1716,N_1409);
and U3246 (N_3246,N_522,N_333);
nor U3247 (N_3247,N_49,N_181);
nor U3248 (N_3248,N_1811,N_869);
or U3249 (N_3249,N_1255,N_198);
xor U3250 (N_3250,N_1656,N_1748);
and U3251 (N_3251,N_981,N_1475);
and U3252 (N_3252,N_1733,N_1122);
or U3253 (N_3253,N_24,N_490);
or U3254 (N_3254,N_1716,N_1097);
or U3255 (N_3255,N_1845,N_1519);
or U3256 (N_3256,N_991,N_777);
and U3257 (N_3257,N_315,N_571);
or U3258 (N_3258,N_1689,N_368);
xnor U3259 (N_3259,N_1872,N_1717);
and U3260 (N_3260,N_1910,N_1794);
and U3261 (N_3261,N_1402,N_1240);
and U3262 (N_3262,N_1705,N_1564);
or U3263 (N_3263,N_961,N_1993);
or U3264 (N_3264,N_1305,N_1394);
and U3265 (N_3265,N_18,N_1855);
and U3266 (N_3266,N_1812,N_721);
nand U3267 (N_3267,N_580,N_1167);
nand U3268 (N_3268,N_1063,N_494);
and U3269 (N_3269,N_702,N_1336);
or U3270 (N_3270,N_1553,N_1383);
nand U3271 (N_3271,N_1165,N_1826);
nor U3272 (N_3272,N_862,N_1812);
or U3273 (N_3273,N_941,N_1456);
nand U3274 (N_3274,N_484,N_1128);
nor U3275 (N_3275,N_415,N_32);
nor U3276 (N_3276,N_551,N_330);
and U3277 (N_3277,N_1822,N_628);
and U3278 (N_3278,N_513,N_543);
and U3279 (N_3279,N_536,N_104);
and U3280 (N_3280,N_955,N_1583);
and U3281 (N_3281,N_1448,N_26);
nand U3282 (N_3282,N_1387,N_1829);
xor U3283 (N_3283,N_1451,N_1863);
nand U3284 (N_3284,N_1684,N_672);
and U3285 (N_3285,N_1394,N_324);
or U3286 (N_3286,N_578,N_1366);
or U3287 (N_3287,N_377,N_844);
nor U3288 (N_3288,N_1087,N_1112);
or U3289 (N_3289,N_1319,N_1671);
and U3290 (N_3290,N_1038,N_281);
and U3291 (N_3291,N_1946,N_491);
nand U3292 (N_3292,N_1698,N_732);
nor U3293 (N_3293,N_358,N_873);
or U3294 (N_3294,N_1197,N_27);
nor U3295 (N_3295,N_1332,N_455);
nor U3296 (N_3296,N_788,N_1397);
nand U3297 (N_3297,N_1128,N_1246);
nor U3298 (N_3298,N_948,N_1751);
nand U3299 (N_3299,N_292,N_1961);
and U3300 (N_3300,N_88,N_1396);
and U3301 (N_3301,N_1401,N_1208);
or U3302 (N_3302,N_511,N_515);
and U3303 (N_3303,N_345,N_1611);
or U3304 (N_3304,N_1688,N_1255);
nor U3305 (N_3305,N_1906,N_500);
nor U3306 (N_3306,N_1932,N_823);
nor U3307 (N_3307,N_816,N_133);
or U3308 (N_3308,N_549,N_197);
xnor U3309 (N_3309,N_1345,N_1938);
and U3310 (N_3310,N_883,N_1379);
or U3311 (N_3311,N_1693,N_983);
or U3312 (N_3312,N_224,N_210);
nor U3313 (N_3313,N_206,N_167);
or U3314 (N_3314,N_736,N_1825);
xnor U3315 (N_3315,N_984,N_1740);
or U3316 (N_3316,N_845,N_921);
nand U3317 (N_3317,N_206,N_1205);
xnor U3318 (N_3318,N_200,N_1880);
and U3319 (N_3319,N_1986,N_935);
and U3320 (N_3320,N_1284,N_943);
nor U3321 (N_3321,N_474,N_1146);
nor U3322 (N_3322,N_348,N_1843);
and U3323 (N_3323,N_1537,N_720);
and U3324 (N_3324,N_1243,N_289);
or U3325 (N_3325,N_821,N_1067);
nor U3326 (N_3326,N_212,N_1740);
xor U3327 (N_3327,N_1809,N_1932);
nor U3328 (N_3328,N_46,N_1852);
xnor U3329 (N_3329,N_163,N_586);
nand U3330 (N_3330,N_1979,N_306);
xnor U3331 (N_3331,N_1332,N_61);
and U3332 (N_3332,N_989,N_1326);
nand U3333 (N_3333,N_78,N_1765);
nand U3334 (N_3334,N_1628,N_1138);
nor U3335 (N_3335,N_1121,N_713);
nor U3336 (N_3336,N_1982,N_1970);
and U3337 (N_3337,N_700,N_1803);
or U3338 (N_3338,N_43,N_414);
and U3339 (N_3339,N_903,N_1664);
xor U3340 (N_3340,N_1828,N_414);
nor U3341 (N_3341,N_110,N_1870);
or U3342 (N_3342,N_589,N_93);
nand U3343 (N_3343,N_1058,N_1800);
or U3344 (N_3344,N_61,N_1768);
or U3345 (N_3345,N_449,N_1371);
nand U3346 (N_3346,N_332,N_1404);
and U3347 (N_3347,N_1306,N_1763);
nand U3348 (N_3348,N_1793,N_1618);
nor U3349 (N_3349,N_814,N_867);
nand U3350 (N_3350,N_1786,N_1534);
and U3351 (N_3351,N_897,N_42);
nor U3352 (N_3352,N_1824,N_1717);
or U3353 (N_3353,N_530,N_1878);
xor U3354 (N_3354,N_842,N_912);
or U3355 (N_3355,N_126,N_502);
nor U3356 (N_3356,N_358,N_1452);
and U3357 (N_3357,N_1810,N_1155);
nor U3358 (N_3358,N_590,N_1266);
nor U3359 (N_3359,N_1502,N_770);
and U3360 (N_3360,N_1750,N_335);
and U3361 (N_3361,N_704,N_1776);
nor U3362 (N_3362,N_1155,N_1744);
xor U3363 (N_3363,N_1835,N_888);
and U3364 (N_3364,N_514,N_1865);
and U3365 (N_3365,N_579,N_543);
nand U3366 (N_3366,N_237,N_56);
and U3367 (N_3367,N_1605,N_1374);
nor U3368 (N_3368,N_584,N_560);
and U3369 (N_3369,N_935,N_1960);
or U3370 (N_3370,N_1240,N_720);
nand U3371 (N_3371,N_991,N_1811);
or U3372 (N_3372,N_209,N_1395);
or U3373 (N_3373,N_388,N_1233);
or U3374 (N_3374,N_1301,N_514);
or U3375 (N_3375,N_931,N_376);
nand U3376 (N_3376,N_1796,N_150);
xnor U3377 (N_3377,N_1666,N_657);
xnor U3378 (N_3378,N_611,N_1757);
and U3379 (N_3379,N_638,N_1276);
nand U3380 (N_3380,N_169,N_486);
nor U3381 (N_3381,N_1987,N_1833);
nand U3382 (N_3382,N_68,N_902);
nand U3383 (N_3383,N_1264,N_1);
nand U3384 (N_3384,N_785,N_1821);
nor U3385 (N_3385,N_1234,N_124);
xor U3386 (N_3386,N_1496,N_714);
or U3387 (N_3387,N_401,N_1762);
nor U3388 (N_3388,N_1290,N_111);
nor U3389 (N_3389,N_976,N_1462);
xor U3390 (N_3390,N_1179,N_1976);
or U3391 (N_3391,N_1980,N_1129);
nand U3392 (N_3392,N_781,N_184);
nand U3393 (N_3393,N_1550,N_1327);
and U3394 (N_3394,N_1566,N_1529);
or U3395 (N_3395,N_984,N_1530);
and U3396 (N_3396,N_1592,N_570);
nor U3397 (N_3397,N_1706,N_1992);
nor U3398 (N_3398,N_1273,N_832);
nor U3399 (N_3399,N_952,N_866);
xor U3400 (N_3400,N_1361,N_1290);
and U3401 (N_3401,N_838,N_210);
nor U3402 (N_3402,N_1,N_1608);
or U3403 (N_3403,N_89,N_1586);
or U3404 (N_3404,N_795,N_844);
xnor U3405 (N_3405,N_96,N_517);
or U3406 (N_3406,N_185,N_466);
and U3407 (N_3407,N_86,N_32);
or U3408 (N_3408,N_1477,N_313);
or U3409 (N_3409,N_316,N_1509);
nand U3410 (N_3410,N_1009,N_1385);
and U3411 (N_3411,N_863,N_1539);
or U3412 (N_3412,N_712,N_974);
nand U3413 (N_3413,N_509,N_1060);
or U3414 (N_3414,N_181,N_182);
and U3415 (N_3415,N_1694,N_1881);
nand U3416 (N_3416,N_1431,N_1458);
or U3417 (N_3417,N_1899,N_1868);
or U3418 (N_3418,N_875,N_1271);
nor U3419 (N_3419,N_871,N_338);
or U3420 (N_3420,N_685,N_1066);
nor U3421 (N_3421,N_45,N_1193);
or U3422 (N_3422,N_1114,N_38);
nor U3423 (N_3423,N_1201,N_1808);
nand U3424 (N_3424,N_36,N_2);
or U3425 (N_3425,N_150,N_1421);
xor U3426 (N_3426,N_602,N_704);
and U3427 (N_3427,N_452,N_832);
nand U3428 (N_3428,N_1936,N_1530);
nand U3429 (N_3429,N_642,N_1182);
or U3430 (N_3430,N_1482,N_514);
and U3431 (N_3431,N_1406,N_1120);
nor U3432 (N_3432,N_1508,N_1721);
nor U3433 (N_3433,N_1396,N_376);
and U3434 (N_3434,N_1487,N_237);
and U3435 (N_3435,N_864,N_1543);
or U3436 (N_3436,N_802,N_400);
or U3437 (N_3437,N_1460,N_29);
xor U3438 (N_3438,N_17,N_1516);
and U3439 (N_3439,N_1293,N_490);
and U3440 (N_3440,N_400,N_695);
nand U3441 (N_3441,N_1621,N_1738);
nand U3442 (N_3442,N_225,N_974);
nor U3443 (N_3443,N_1992,N_1345);
or U3444 (N_3444,N_338,N_703);
xnor U3445 (N_3445,N_796,N_1299);
and U3446 (N_3446,N_156,N_1837);
nand U3447 (N_3447,N_1008,N_639);
nor U3448 (N_3448,N_1067,N_1216);
nor U3449 (N_3449,N_711,N_429);
and U3450 (N_3450,N_1626,N_1915);
nand U3451 (N_3451,N_89,N_1967);
nand U3452 (N_3452,N_1865,N_428);
nand U3453 (N_3453,N_1600,N_37);
nand U3454 (N_3454,N_140,N_539);
and U3455 (N_3455,N_1713,N_1244);
or U3456 (N_3456,N_1927,N_1944);
or U3457 (N_3457,N_788,N_1015);
xnor U3458 (N_3458,N_792,N_1601);
xnor U3459 (N_3459,N_872,N_195);
nand U3460 (N_3460,N_1365,N_1630);
nor U3461 (N_3461,N_549,N_1538);
nand U3462 (N_3462,N_677,N_1030);
and U3463 (N_3463,N_322,N_1709);
and U3464 (N_3464,N_898,N_349);
xnor U3465 (N_3465,N_187,N_559);
nand U3466 (N_3466,N_723,N_515);
or U3467 (N_3467,N_930,N_1782);
and U3468 (N_3468,N_733,N_335);
and U3469 (N_3469,N_1048,N_910);
xnor U3470 (N_3470,N_351,N_225);
and U3471 (N_3471,N_1019,N_1100);
nand U3472 (N_3472,N_1644,N_1159);
nand U3473 (N_3473,N_202,N_719);
or U3474 (N_3474,N_1339,N_32);
or U3475 (N_3475,N_1737,N_1050);
or U3476 (N_3476,N_612,N_518);
and U3477 (N_3477,N_1397,N_1531);
and U3478 (N_3478,N_938,N_1228);
nand U3479 (N_3479,N_147,N_605);
nand U3480 (N_3480,N_137,N_832);
nand U3481 (N_3481,N_196,N_152);
and U3482 (N_3482,N_1619,N_1596);
and U3483 (N_3483,N_1044,N_1484);
or U3484 (N_3484,N_593,N_552);
nor U3485 (N_3485,N_1185,N_1310);
nor U3486 (N_3486,N_926,N_1035);
nor U3487 (N_3487,N_1886,N_899);
nor U3488 (N_3488,N_663,N_1661);
nor U3489 (N_3489,N_1684,N_480);
nand U3490 (N_3490,N_40,N_1114);
and U3491 (N_3491,N_1986,N_1639);
and U3492 (N_3492,N_1714,N_851);
nor U3493 (N_3493,N_1131,N_1845);
or U3494 (N_3494,N_1531,N_1728);
nor U3495 (N_3495,N_1628,N_1666);
xor U3496 (N_3496,N_8,N_985);
nand U3497 (N_3497,N_815,N_1646);
or U3498 (N_3498,N_1748,N_1424);
and U3499 (N_3499,N_1749,N_1576);
nand U3500 (N_3500,N_750,N_41);
xnor U3501 (N_3501,N_1960,N_1838);
nand U3502 (N_3502,N_1924,N_595);
and U3503 (N_3503,N_1245,N_959);
nand U3504 (N_3504,N_1714,N_1708);
or U3505 (N_3505,N_1789,N_1037);
nand U3506 (N_3506,N_1547,N_1839);
nand U3507 (N_3507,N_852,N_715);
nand U3508 (N_3508,N_1489,N_219);
or U3509 (N_3509,N_1313,N_1488);
nand U3510 (N_3510,N_1011,N_131);
or U3511 (N_3511,N_1313,N_1455);
nor U3512 (N_3512,N_1766,N_788);
nor U3513 (N_3513,N_1220,N_1466);
nand U3514 (N_3514,N_528,N_660);
nor U3515 (N_3515,N_766,N_563);
and U3516 (N_3516,N_216,N_314);
xor U3517 (N_3517,N_1038,N_1757);
nor U3518 (N_3518,N_291,N_717);
nor U3519 (N_3519,N_1673,N_372);
nor U3520 (N_3520,N_1949,N_483);
or U3521 (N_3521,N_318,N_1940);
or U3522 (N_3522,N_1600,N_1755);
nor U3523 (N_3523,N_1045,N_1202);
or U3524 (N_3524,N_1220,N_1202);
or U3525 (N_3525,N_128,N_370);
and U3526 (N_3526,N_1771,N_1167);
and U3527 (N_3527,N_94,N_656);
and U3528 (N_3528,N_390,N_877);
nand U3529 (N_3529,N_164,N_82);
and U3530 (N_3530,N_797,N_1491);
nor U3531 (N_3531,N_935,N_114);
and U3532 (N_3532,N_487,N_1242);
nand U3533 (N_3533,N_358,N_500);
and U3534 (N_3534,N_55,N_987);
xor U3535 (N_3535,N_967,N_195);
nand U3536 (N_3536,N_401,N_1587);
nor U3537 (N_3537,N_1335,N_1520);
or U3538 (N_3538,N_460,N_1798);
xnor U3539 (N_3539,N_1010,N_222);
xor U3540 (N_3540,N_1641,N_1272);
and U3541 (N_3541,N_549,N_171);
and U3542 (N_3542,N_1537,N_262);
and U3543 (N_3543,N_1746,N_1727);
nand U3544 (N_3544,N_379,N_1700);
and U3545 (N_3545,N_351,N_1685);
nand U3546 (N_3546,N_366,N_357);
nor U3547 (N_3547,N_1898,N_1480);
and U3548 (N_3548,N_1114,N_521);
nor U3549 (N_3549,N_369,N_220);
and U3550 (N_3550,N_1335,N_1968);
nand U3551 (N_3551,N_1096,N_1148);
nand U3552 (N_3552,N_1495,N_781);
nor U3553 (N_3553,N_211,N_1393);
or U3554 (N_3554,N_1381,N_1491);
nor U3555 (N_3555,N_389,N_747);
nand U3556 (N_3556,N_1547,N_1989);
nand U3557 (N_3557,N_1393,N_1923);
nor U3558 (N_3558,N_567,N_1853);
nor U3559 (N_3559,N_1532,N_1067);
or U3560 (N_3560,N_700,N_1186);
xor U3561 (N_3561,N_1541,N_208);
or U3562 (N_3562,N_653,N_1883);
nor U3563 (N_3563,N_387,N_540);
nand U3564 (N_3564,N_985,N_580);
nand U3565 (N_3565,N_1797,N_459);
or U3566 (N_3566,N_1536,N_1806);
nand U3567 (N_3567,N_943,N_883);
nor U3568 (N_3568,N_301,N_1219);
or U3569 (N_3569,N_868,N_292);
or U3570 (N_3570,N_647,N_1541);
xor U3571 (N_3571,N_1317,N_1230);
nand U3572 (N_3572,N_1921,N_1878);
nor U3573 (N_3573,N_1514,N_1181);
nor U3574 (N_3574,N_1565,N_682);
or U3575 (N_3575,N_607,N_1787);
nand U3576 (N_3576,N_1739,N_889);
or U3577 (N_3577,N_91,N_952);
xnor U3578 (N_3578,N_128,N_1682);
and U3579 (N_3579,N_594,N_26);
xnor U3580 (N_3580,N_1594,N_990);
or U3581 (N_3581,N_94,N_1054);
or U3582 (N_3582,N_1713,N_1473);
and U3583 (N_3583,N_1776,N_1284);
nor U3584 (N_3584,N_217,N_1561);
nand U3585 (N_3585,N_596,N_631);
xor U3586 (N_3586,N_1504,N_460);
nor U3587 (N_3587,N_581,N_687);
and U3588 (N_3588,N_651,N_473);
nor U3589 (N_3589,N_1217,N_327);
nor U3590 (N_3590,N_1556,N_1799);
xnor U3591 (N_3591,N_12,N_920);
nand U3592 (N_3592,N_1938,N_133);
xnor U3593 (N_3593,N_911,N_1074);
or U3594 (N_3594,N_272,N_1430);
and U3595 (N_3595,N_228,N_607);
and U3596 (N_3596,N_1874,N_1042);
nor U3597 (N_3597,N_617,N_1603);
or U3598 (N_3598,N_104,N_1037);
nand U3599 (N_3599,N_23,N_1299);
nor U3600 (N_3600,N_1930,N_143);
nand U3601 (N_3601,N_1394,N_1399);
and U3602 (N_3602,N_351,N_503);
or U3603 (N_3603,N_752,N_577);
nand U3604 (N_3604,N_802,N_1964);
or U3605 (N_3605,N_1941,N_233);
and U3606 (N_3606,N_1571,N_1298);
nand U3607 (N_3607,N_900,N_551);
xor U3608 (N_3608,N_808,N_1014);
or U3609 (N_3609,N_1106,N_157);
and U3610 (N_3610,N_1784,N_74);
nor U3611 (N_3611,N_419,N_1302);
and U3612 (N_3612,N_1767,N_1146);
nor U3613 (N_3613,N_902,N_189);
xnor U3614 (N_3614,N_874,N_644);
nand U3615 (N_3615,N_380,N_905);
or U3616 (N_3616,N_900,N_1051);
nor U3617 (N_3617,N_335,N_544);
nor U3618 (N_3618,N_1192,N_1175);
and U3619 (N_3619,N_1779,N_407);
nand U3620 (N_3620,N_1460,N_948);
nand U3621 (N_3621,N_1259,N_1195);
or U3622 (N_3622,N_110,N_1344);
nand U3623 (N_3623,N_51,N_1404);
xnor U3624 (N_3624,N_358,N_621);
xnor U3625 (N_3625,N_266,N_141);
nand U3626 (N_3626,N_880,N_74);
nor U3627 (N_3627,N_1116,N_1978);
nor U3628 (N_3628,N_946,N_399);
nand U3629 (N_3629,N_1194,N_1262);
nor U3630 (N_3630,N_726,N_1795);
nor U3631 (N_3631,N_843,N_533);
and U3632 (N_3632,N_1267,N_1279);
nor U3633 (N_3633,N_719,N_1200);
nor U3634 (N_3634,N_1487,N_1030);
xnor U3635 (N_3635,N_1462,N_1781);
nor U3636 (N_3636,N_1131,N_1051);
nor U3637 (N_3637,N_1134,N_647);
nand U3638 (N_3638,N_683,N_84);
or U3639 (N_3639,N_571,N_1197);
or U3640 (N_3640,N_372,N_1560);
nand U3641 (N_3641,N_1256,N_410);
or U3642 (N_3642,N_1257,N_14);
nand U3643 (N_3643,N_219,N_1298);
nand U3644 (N_3644,N_699,N_771);
or U3645 (N_3645,N_1406,N_389);
nand U3646 (N_3646,N_245,N_1274);
nand U3647 (N_3647,N_1219,N_1941);
or U3648 (N_3648,N_1917,N_421);
nand U3649 (N_3649,N_636,N_915);
nand U3650 (N_3650,N_571,N_1638);
or U3651 (N_3651,N_1282,N_1224);
nor U3652 (N_3652,N_1505,N_827);
nand U3653 (N_3653,N_1179,N_487);
nor U3654 (N_3654,N_1341,N_1909);
nor U3655 (N_3655,N_539,N_1901);
or U3656 (N_3656,N_1084,N_364);
or U3657 (N_3657,N_1481,N_873);
nor U3658 (N_3658,N_1723,N_177);
nor U3659 (N_3659,N_853,N_299);
nor U3660 (N_3660,N_1132,N_1936);
and U3661 (N_3661,N_1498,N_83);
and U3662 (N_3662,N_1606,N_1202);
or U3663 (N_3663,N_1682,N_484);
and U3664 (N_3664,N_1882,N_1714);
or U3665 (N_3665,N_943,N_996);
xor U3666 (N_3666,N_575,N_471);
nand U3667 (N_3667,N_741,N_1262);
and U3668 (N_3668,N_1074,N_556);
nor U3669 (N_3669,N_1570,N_387);
and U3670 (N_3670,N_78,N_531);
nor U3671 (N_3671,N_1266,N_494);
and U3672 (N_3672,N_645,N_60);
nor U3673 (N_3673,N_285,N_132);
or U3674 (N_3674,N_261,N_854);
and U3675 (N_3675,N_675,N_1672);
nor U3676 (N_3676,N_323,N_1581);
and U3677 (N_3677,N_114,N_1800);
and U3678 (N_3678,N_1985,N_585);
xor U3679 (N_3679,N_1820,N_904);
and U3680 (N_3680,N_1742,N_1743);
nand U3681 (N_3681,N_1088,N_808);
xnor U3682 (N_3682,N_1594,N_1261);
nor U3683 (N_3683,N_1500,N_1383);
and U3684 (N_3684,N_1680,N_1701);
nand U3685 (N_3685,N_1559,N_1048);
and U3686 (N_3686,N_1602,N_300);
or U3687 (N_3687,N_1116,N_482);
xor U3688 (N_3688,N_1156,N_96);
nor U3689 (N_3689,N_375,N_609);
nand U3690 (N_3690,N_903,N_1332);
and U3691 (N_3691,N_1052,N_1221);
and U3692 (N_3692,N_118,N_1099);
and U3693 (N_3693,N_1385,N_1307);
nand U3694 (N_3694,N_895,N_1279);
nor U3695 (N_3695,N_611,N_845);
and U3696 (N_3696,N_1711,N_1902);
or U3697 (N_3697,N_1686,N_1423);
or U3698 (N_3698,N_1366,N_1649);
and U3699 (N_3699,N_1495,N_1396);
nand U3700 (N_3700,N_523,N_1837);
nand U3701 (N_3701,N_224,N_1753);
or U3702 (N_3702,N_1244,N_481);
nor U3703 (N_3703,N_1888,N_365);
nor U3704 (N_3704,N_890,N_1982);
or U3705 (N_3705,N_1382,N_1434);
and U3706 (N_3706,N_1696,N_1550);
and U3707 (N_3707,N_213,N_1016);
nor U3708 (N_3708,N_1167,N_941);
nand U3709 (N_3709,N_1895,N_1652);
xnor U3710 (N_3710,N_299,N_198);
xor U3711 (N_3711,N_1768,N_382);
or U3712 (N_3712,N_422,N_131);
nand U3713 (N_3713,N_479,N_410);
or U3714 (N_3714,N_1810,N_1593);
nand U3715 (N_3715,N_1234,N_1013);
nor U3716 (N_3716,N_1991,N_947);
and U3717 (N_3717,N_1869,N_1273);
nand U3718 (N_3718,N_891,N_1766);
nand U3719 (N_3719,N_96,N_1889);
or U3720 (N_3720,N_37,N_1559);
or U3721 (N_3721,N_1050,N_1419);
nand U3722 (N_3722,N_1512,N_1567);
or U3723 (N_3723,N_1042,N_409);
and U3724 (N_3724,N_750,N_1199);
or U3725 (N_3725,N_1017,N_702);
nor U3726 (N_3726,N_1372,N_461);
nor U3727 (N_3727,N_367,N_867);
or U3728 (N_3728,N_515,N_1608);
and U3729 (N_3729,N_1485,N_1056);
or U3730 (N_3730,N_656,N_739);
and U3731 (N_3731,N_1025,N_1239);
nand U3732 (N_3732,N_1067,N_1399);
nand U3733 (N_3733,N_549,N_1493);
nand U3734 (N_3734,N_1094,N_1874);
and U3735 (N_3735,N_454,N_1275);
or U3736 (N_3736,N_1169,N_1902);
or U3737 (N_3737,N_1684,N_870);
nor U3738 (N_3738,N_1081,N_144);
nor U3739 (N_3739,N_1591,N_710);
nor U3740 (N_3740,N_556,N_1780);
xor U3741 (N_3741,N_1417,N_78);
or U3742 (N_3742,N_1523,N_1152);
or U3743 (N_3743,N_1751,N_355);
nor U3744 (N_3744,N_1748,N_38);
nand U3745 (N_3745,N_902,N_191);
nor U3746 (N_3746,N_1487,N_1877);
xor U3747 (N_3747,N_1869,N_255);
nor U3748 (N_3748,N_990,N_1188);
or U3749 (N_3749,N_97,N_1568);
xnor U3750 (N_3750,N_1350,N_1772);
and U3751 (N_3751,N_556,N_683);
xnor U3752 (N_3752,N_1981,N_649);
nand U3753 (N_3753,N_1657,N_1090);
xor U3754 (N_3754,N_1971,N_1834);
and U3755 (N_3755,N_571,N_1884);
nor U3756 (N_3756,N_1544,N_1253);
and U3757 (N_3757,N_725,N_1935);
nand U3758 (N_3758,N_123,N_1232);
nor U3759 (N_3759,N_1480,N_1172);
or U3760 (N_3760,N_49,N_433);
or U3761 (N_3761,N_768,N_1760);
and U3762 (N_3762,N_388,N_1061);
and U3763 (N_3763,N_1563,N_757);
nand U3764 (N_3764,N_1355,N_709);
nor U3765 (N_3765,N_24,N_404);
and U3766 (N_3766,N_1528,N_1593);
or U3767 (N_3767,N_1330,N_1086);
or U3768 (N_3768,N_1370,N_1852);
and U3769 (N_3769,N_1622,N_1245);
and U3770 (N_3770,N_517,N_1029);
nand U3771 (N_3771,N_1214,N_534);
nand U3772 (N_3772,N_1298,N_1845);
and U3773 (N_3773,N_1491,N_19);
or U3774 (N_3774,N_89,N_1805);
or U3775 (N_3775,N_1486,N_832);
and U3776 (N_3776,N_1335,N_929);
or U3777 (N_3777,N_1499,N_954);
and U3778 (N_3778,N_1133,N_1589);
or U3779 (N_3779,N_1051,N_788);
nand U3780 (N_3780,N_1596,N_226);
and U3781 (N_3781,N_1558,N_967);
xnor U3782 (N_3782,N_1966,N_1069);
nand U3783 (N_3783,N_1705,N_1598);
or U3784 (N_3784,N_556,N_247);
nand U3785 (N_3785,N_890,N_1829);
or U3786 (N_3786,N_1370,N_1777);
nand U3787 (N_3787,N_1600,N_704);
nand U3788 (N_3788,N_1644,N_565);
xor U3789 (N_3789,N_773,N_1178);
or U3790 (N_3790,N_797,N_753);
nor U3791 (N_3791,N_1019,N_662);
or U3792 (N_3792,N_1526,N_1391);
or U3793 (N_3793,N_836,N_1013);
or U3794 (N_3794,N_672,N_26);
nor U3795 (N_3795,N_1007,N_973);
or U3796 (N_3796,N_333,N_1281);
nor U3797 (N_3797,N_1686,N_701);
nand U3798 (N_3798,N_586,N_882);
xnor U3799 (N_3799,N_1569,N_1217);
nor U3800 (N_3800,N_619,N_1874);
xor U3801 (N_3801,N_895,N_1021);
xnor U3802 (N_3802,N_130,N_1375);
and U3803 (N_3803,N_587,N_603);
nor U3804 (N_3804,N_365,N_841);
and U3805 (N_3805,N_1400,N_1819);
nand U3806 (N_3806,N_758,N_1512);
and U3807 (N_3807,N_1640,N_945);
nor U3808 (N_3808,N_873,N_647);
or U3809 (N_3809,N_1932,N_1376);
xnor U3810 (N_3810,N_525,N_1288);
or U3811 (N_3811,N_1090,N_129);
xor U3812 (N_3812,N_1596,N_849);
and U3813 (N_3813,N_178,N_1959);
nand U3814 (N_3814,N_948,N_684);
nand U3815 (N_3815,N_1327,N_1790);
nor U3816 (N_3816,N_1827,N_1294);
or U3817 (N_3817,N_340,N_978);
xor U3818 (N_3818,N_1285,N_1937);
nor U3819 (N_3819,N_475,N_494);
and U3820 (N_3820,N_1735,N_1823);
xor U3821 (N_3821,N_1969,N_1509);
and U3822 (N_3822,N_952,N_396);
nor U3823 (N_3823,N_628,N_1297);
or U3824 (N_3824,N_1579,N_617);
nor U3825 (N_3825,N_1131,N_1086);
nand U3826 (N_3826,N_1059,N_1687);
or U3827 (N_3827,N_1540,N_1253);
nor U3828 (N_3828,N_351,N_659);
xnor U3829 (N_3829,N_111,N_709);
nor U3830 (N_3830,N_1705,N_639);
nor U3831 (N_3831,N_574,N_1547);
nor U3832 (N_3832,N_175,N_607);
nand U3833 (N_3833,N_1034,N_1079);
xor U3834 (N_3834,N_1800,N_302);
and U3835 (N_3835,N_700,N_1313);
nand U3836 (N_3836,N_1345,N_726);
xor U3837 (N_3837,N_1370,N_1122);
or U3838 (N_3838,N_64,N_800);
or U3839 (N_3839,N_967,N_1430);
nand U3840 (N_3840,N_1499,N_1014);
nand U3841 (N_3841,N_527,N_617);
xnor U3842 (N_3842,N_142,N_1599);
nor U3843 (N_3843,N_1595,N_736);
or U3844 (N_3844,N_1878,N_1867);
or U3845 (N_3845,N_1150,N_1971);
and U3846 (N_3846,N_1643,N_142);
nand U3847 (N_3847,N_1061,N_1747);
nor U3848 (N_3848,N_914,N_1678);
and U3849 (N_3849,N_941,N_891);
nor U3850 (N_3850,N_1075,N_1609);
nor U3851 (N_3851,N_487,N_1115);
nor U3852 (N_3852,N_1346,N_367);
or U3853 (N_3853,N_1540,N_32);
xor U3854 (N_3854,N_8,N_210);
nor U3855 (N_3855,N_925,N_1901);
nand U3856 (N_3856,N_1482,N_1887);
nand U3857 (N_3857,N_355,N_1581);
nand U3858 (N_3858,N_1555,N_118);
and U3859 (N_3859,N_1118,N_1562);
or U3860 (N_3860,N_1202,N_1718);
xnor U3861 (N_3861,N_1778,N_1948);
nor U3862 (N_3862,N_1452,N_1374);
and U3863 (N_3863,N_444,N_1723);
nand U3864 (N_3864,N_224,N_1185);
xnor U3865 (N_3865,N_1785,N_679);
and U3866 (N_3866,N_703,N_480);
nand U3867 (N_3867,N_182,N_124);
and U3868 (N_3868,N_894,N_877);
nor U3869 (N_3869,N_1495,N_237);
or U3870 (N_3870,N_569,N_1765);
or U3871 (N_3871,N_1735,N_761);
xnor U3872 (N_3872,N_15,N_1237);
nor U3873 (N_3873,N_359,N_674);
or U3874 (N_3874,N_1822,N_151);
nand U3875 (N_3875,N_9,N_1724);
nand U3876 (N_3876,N_783,N_896);
nand U3877 (N_3877,N_1660,N_761);
nor U3878 (N_3878,N_455,N_1991);
and U3879 (N_3879,N_1227,N_1477);
xor U3880 (N_3880,N_989,N_174);
and U3881 (N_3881,N_1550,N_49);
or U3882 (N_3882,N_105,N_984);
and U3883 (N_3883,N_659,N_557);
or U3884 (N_3884,N_1035,N_1257);
nand U3885 (N_3885,N_1064,N_1069);
and U3886 (N_3886,N_1265,N_77);
nand U3887 (N_3887,N_685,N_647);
and U3888 (N_3888,N_908,N_62);
nand U3889 (N_3889,N_173,N_1108);
or U3890 (N_3890,N_1925,N_855);
or U3891 (N_3891,N_259,N_727);
nand U3892 (N_3892,N_926,N_1543);
and U3893 (N_3893,N_668,N_1196);
and U3894 (N_3894,N_754,N_946);
nand U3895 (N_3895,N_1862,N_1603);
nand U3896 (N_3896,N_467,N_237);
xor U3897 (N_3897,N_1839,N_1067);
and U3898 (N_3898,N_1533,N_671);
or U3899 (N_3899,N_946,N_796);
nand U3900 (N_3900,N_1108,N_1472);
and U3901 (N_3901,N_1809,N_574);
or U3902 (N_3902,N_1781,N_280);
and U3903 (N_3903,N_976,N_801);
or U3904 (N_3904,N_1473,N_376);
xnor U3905 (N_3905,N_181,N_415);
or U3906 (N_3906,N_1449,N_570);
and U3907 (N_3907,N_608,N_464);
nand U3908 (N_3908,N_1039,N_1462);
nor U3909 (N_3909,N_1560,N_1199);
nor U3910 (N_3910,N_72,N_40);
nand U3911 (N_3911,N_1752,N_86);
nor U3912 (N_3912,N_741,N_1887);
xor U3913 (N_3913,N_361,N_1202);
or U3914 (N_3914,N_1376,N_174);
nand U3915 (N_3915,N_1535,N_1873);
nor U3916 (N_3916,N_941,N_1613);
and U3917 (N_3917,N_736,N_851);
nand U3918 (N_3918,N_148,N_725);
xor U3919 (N_3919,N_126,N_425);
and U3920 (N_3920,N_1127,N_1882);
or U3921 (N_3921,N_1489,N_1480);
nand U3922 (N_3922,N_958,N_1542);
nor U3923 (N_3923,N_590,N_627);
nand U3924 (N_3924,N_1810,N_1565);
or U3925 (N_3925,N_1180,N_1820);
xnor U3926 (N_3926,N_78,N_1120);
xnor U3927 (N_3927,N_1637,N_1489);
and U3928 (N_3928,N_262,N_1436);
nand U3929 (N_3929,N_1807,N_387);
or U3930 (N_3930,N_1273,N_13);
nor U3931 (N_3931,N_1850,N_1844);
nand U3932 (N_3932,N_8,N_1228);
nand U3933 (N_3933,N_1161,N_14);
nor U3934 (N_3934,N_334,N_373);
and U3935 (N_3935,N_747,N_600);
nand U3936 (N_3936,N_426,N_1347);
and U3937 (N_3937,N_1422,N_1004);
nand U3938 (N_3938,N_672,N_584);
nand U3939 (N_3939,N_717,N_508);
and U3940 (N_3940,N_1606,N_786);
xor U3941 (N_3941,N_610,N_1229);
nor U3942 (N_3942,N_955,N_719);
nand U3943 (N_3943,N_295,N_768);
and U3944 (N_3944,N_1297,N_1633);
nor U3945 (N_3945,N_329,N_4);
nand U3946 (N_3946,N_143,N_686);
and U3947 (N_3947,N_82,N_979);
nand U3948 (N_3948,N_873,N_301);
and U3949 (N_3949,N_1950,N_932);
nand U3950 (N_3950,N_377,N_1090);
or U3951 (N_3951,N_1864,N_1476);
and U3952 (N_3952,N_823,N_909);
or U3953 (N_3953,N_1132,N_1260);
nor U3954 (N_3954,N_760,N_753);
xnor U3955 (N_3955,N_819,N_148);
nor U3956 (N_3956,N_721,N_1731);
nor U3957 (N_3957,N_1379,N_1926);
or U3958 (N_3958,N_442,N_763);
and U3959 (N_3959,N_1927,N_1643);
or U3960 (N_3960,N_1293,N_1334);
nor U3961 (N_3961,N_917,N_1172);
or U3962 (N_3962,N_1114,N_684);
nand U3963 (N_3963,N_741,N_1152);
or U3964 (N_3964,N_1863,N_1974);
nand U3965 (N_3965,N_888,N_1347);
xor U3966 (N_3966,N_600,N_1204);
nor U3967 (N_3967,N_1391,N_1605);
nor U3968 (N_3968,N_1613,N_1397);
or U3969 (N_3969,N_498,N_1169);
nor U3970 (N_3970,N_1508,N_1995);
and U3971 (N_3971,N_1986,N_1160);
nand U3972 (N_3972,N_1788,N_1211);
and U3973 (N_3973,N_71,N_600);
xor U3974 (N_3974,N_1130,N_635);
or U3975 (N_3975,N_680,N_811);
and U3976 (N_3976,N_1464,N_444);
and U3977 (N_3977,N_382,N_1540);
nor U3978 (N_3978,N_591,N_1684);
xnor U3979 (N_3979,N_1994,N_623);
and U3980 (N_3980,N_84,N_1515);
or U3981 (N_3981,N_1646,N_1647);
and U3982 (N_3982,N_969,N_1625);
nor U3983 (N_3983,N_1053,N_471);
and U3984 (N_3984,N_152,N_319);
xnor U3985 (N_3985,N_825,N_1360);
xnor U3986 (N_3986,N_1719,N_1502);
nor U3987 (N_3987,N_427,N_680);
or U3988 (N_3988,N_177,N_773);
nor U3989 (N_3989,N_1016,N_1495);
and U3990 (N_3990,N_1839,N_1541);
or U3991 (N_3991,N_501,N_1463);
or U3992 (N_3992,N_518,N_186);
and U3993 (N_3993,N_961,N_1384);
or U3994 (N_3994,N_1595,N_1599);
and U3995 (N_3995,N_1953,N_919);
xor U3996 (N_3996,N_1398,N_956);
nor U3997 (N_3997,N_1135,N_100);
nor U3998 (N_3998,N_1939,N_966);
xnor U3999 (N_3999,N_489,N_1898);
or U4000 (N_4000,N_3015,N_2095);
nand U4001 (N_4001,N_3336,N_3436);
xor U4002 (N_4002,N_2011,N_2090);
and U4003 (N_4003,N_2573,N_2805);
or U4004 (N_4004,N_2294,N_3018);
and U4005 (N_4005,N_3920,N_2923);
nand U4006 (N_4006,N_3598,N_2393);
or U4007 (N_4007,N_3719,N_2466);
nor U4008 (N_4008,N_3533,N_2258);
nand U4009 (N_4009,N_2539,N_2665);
and U4010 (N_4010,N_3371,N_3618);
nor U4011 (N_4011,N_3069,N_3343);
and U4012 (N_4012,N_3833,N_3315);
nand U4013 (N_4013,N_2333,N_2528);
xnor U4014 (N_4014,N_3965,N_2626);
or U4015 (N_4015,N_2203,N_3638);
and U4016 (N_4016,N_3269,N_2775);
nor U4017 (N_4017,N_3035,N_2536);
and U4018 (N_4018,N_3189,N_3379);
nor U4019 (N_4019,N_3161,N_2318);
and U4020 (N_4020,N_2839,N_2083);
nand U4021 (N_4021,N_2050,N_3448);
nand U4022 (N_4022,N_3107,N_3478);
nand U4023 (N_4023,N_3001,N_2413);
or U4024 (N_4024,N_2981,N_3687);
nand U4025 (N_4025,N_3990,N_2568);
xor U4026 (N_4026,N_3144,N_2708);
and U4027 (N_4027,N_3134,N_2340);
or U4028 (N_4028,N_3435,N_2409);
and U4029 (N_4029,N_3308,N_2969);
or U4030 (N_4030,N_3845,N_2717);
and U4031 (N_4031,N_3510,N_2404);
or U4032 (N_4032,N_3779,N_3546);
nor U4033 (N_4033,N_2062,N_3658);
xor U4034 (N_4034,N_3917,N_3378);
and U4035 (N_4035,N_2281,N_3317);
or U4036 (N_4036,N_2591,N_2799);
and U4037 (N_4037,N_3162,N_3762);
or U4038 (N_4038,N_2423,N_2540);
nor U4039 (N_4039,N_3079,N_2209);
nand U4040 (N_4040,N_3670,N_2368);
or U4041 (N_4041,N_2977,N_2102);
and U4042 (N_4042,N_2779,N_3333);
or U4043 (N_4043,N_2054,N_3178);
and U4044 (N_4044,N_3212,N_2504);
and U4045 (N_4045,N_3485,N_2984);
xnor U4046 (N_4046,N_3787,N_2342);
or U4047 (N_4047,N_3587,N_2713);
and U4048 (N_4048,N_3856,N_3733);
or U4049 (N_4049,N_2986,N_2718);
nor U4050 (N_4050,N_3483,N_2214);
nor U4051 (N_4051,N_2444,N_2639);
nand U4052 (N_4052,N_3053,N_2110);
nand U4053 (N_4053,N_3661,N_3950);
xnor U4054 (N_4054,N_2651,N_3443);
nor U4055 (N_4055,N_2921,N_3802);
nand U4056 (N_4056,N_3398,N_3303);
nand U4057 (N_4057,N_2558,N_2937);
nand U4058 (N_4058,N_2046,N_2467);
nand U4059 (N_4059,N_2350,N_3803);
xnor U4060 (N_4060,N_3260,N_2111);
nand U4061 (N_4061,N_3791,N_2885);
xnor U4062 (N_4062,N_2551,N_3342);
or U4063 (N_4063,N_2786,N_3637);
nor U4064 (N_4064,N_3849,N_3326);
nand U4065 (N_4065,N_3111,N_3578);
nand U4066 (N_4066,N_3931,N_2594);
nand U4067 (N_4067,N_2190,N_3384);
or U4068 (N_4068,N_2360,N_2223);
xor U4069 (N_4069,N_3701,N_2187);
nand U4070 (N_4070,N_3657,N_3365);
nor U4071 (N_4071,N_3408,N_3044);
and U4072 (N_4072,N_3594,N_3309);
xor U4073 (N_4073,N_3356,N_3520);
or U4074 (N_4074,N_3771,N_2668);
and U4075 (N_4075,N_3686,N_3962);
nor U4076 (N_4076,N_3496,N_2972);
nand U4077 (N_4077,N_2048,N_3539);
or U4078 (N_4078,N_2869,N_3997);
and U4079 (N_4079,N_3509,N_2850);
or U4080 (N_4080,N_2553,N_2823);
nand U4081 (N_4081,N_3293,N_2679);
and U4082 (N_4082,N_2566,N_3900);
or U4083 (N_4083,N_3160,N_2402);
or U4084 (N_4084,N_2186,N_3066);
xor U4085 (N_4085,N_3146,N_2240);
nand U4086 (N_4086,N_3766,N_3486);
xnor U4087 (N_4087,N_3428,N_3334);
or U4088 (N_4088,N_3964,N_2367);
or U4089 (N_4089,N_3763,N_3050);
nor U4090 (N_4090,N_3251,N_2925);
or U4091 (N_4091,N_3767,N_2653);
xor U4092 (N_4092,N_3185,N_2552);
and U4093 (N_4093,N_2341,N_2815);
and U4094 (N_4094,N_2509,N_2139);
nand U4095 (N_4095,N_2579,N_2947);
nor U4096 (N_4096,N_3707,N_3959);
xnor U4097 (N_4097,N_2629,N_3799);
or U4098 (N_4098,N_3005,N_2785);
or U4099 (N_4099,N_2895,N_2464);
xor U4100 (N_4100,N_2960,N_2018);
nor U4101 (N_4101,N_3873,N_2141);
xnor U4102 (N_4102,N_2765,N_2230);
and U4103 (N_4103,N_2771,N_3324);
nor U4104 (N_4104,N_2273,N_2748);
nor U4105 (N_4105,N_2267,N_3591);
nor U4106 (N_4106,N_2491,N_2122);
nand U4107 (N_4107,N_2479,N_3499);
and U4108 (N_4108,N_2429,N_3535);
xnor U4109 (N_4109,N_3278,N_2495);
nand U4110 (N_4110,N_2917,N_2037);
nand U4111 (N_4111,N_2487,N_3217);
nor U4112 (N_4112,N_3240,N_3983);
or U4113 (N_4113,N_2452,N_2218);
nor U4114 (N_4114,N_2189,N_3930);
nand U4115 (N_4115,N_3331,N_3459);
nand U4116 (N_4116,N_3416,N_3447);
or U4117 (N_4117,N_2118,N_3122);
and U4118 (N_4118,N_2681,N_2123);
or U4119 (N_4119,N_2134,N_3070);
nor U4120 (N_4120,N_3912,N_3453);
or U4121 (N_4121,N_2430,N_3903);
and U4122 (N_4122,N_3057,N_3726);
xnor U4123 (N_4123,N_3671,N_3387);
or U4124 (N_4124,N_3798,N_2891);
nor U4125 (N_4125,N_3713,N_2978);
nand U4126 (N_4126,N_3742,N_3809);
nand U4127 (N_4127,N_3274,N_2656);
nor U4128 (N_4128,N_2535,N_3038);
nor U4129 (N_4129,N_2843,N_2389);
and U4130 (N_4130,N_2262,N_2329);
xor U4131 (N_4131,N_2688,N_3471);
nor U4132 (N_4132,N_2147,N_3033);
nand U4133 (N_4133,N_3346,N_2761);
and U4134 (N_4134,N_3233,N_3624);
and U4135 (N_4135,N_3581,N_2352);
nor U4136 (N_4136,N_2928,N_3734);
or U4137 (N_4137,N_3355,N_2967);
nand U4138 (N_4138,N_2956,N_2778);
and U4139 (N_4139,N_3115,N_3630);
nor U4140 (N_4140,N_2531,N_2047);
or U4141 (N_4141,N_2655,N_2988);
nand U4142 (N_4142,N_2414,N_2069);
nor U4143 (N_4143,N_2072,N_2798);
nand U4144 (N_4144,N_3544,N_3414);
nand U4145 (N_4145,N_3706,N_2354);
xnor U4146 (N_4146,N_3330,N_2683);
nor U4147 (N_4147,N_2330,N_2879);
nand U4148 (N_4148,N_2968,N_3463);
xnor U4149 (N_4149,N_2517,N_3222);
nand U4150 (N_4150,N_3316,N_3773);
or U4151 (N_4151,N_2399,N_2445);
and U4152 (N_4152,N_3700,N_3261);
nand U4153 (N_4153,N_3511,N_2345);
or U4154 (N_4154,N_2001,N_2058);
or U4155 (N_4155,N_3602,N_3036);
or U4156 (N_4156,N_2266,N_2161);
nand U4157 (N_4157,N_2982,N_3148);
or U4158 (N_4158,N_3277,N_3548);
or U4159 (N_4159,N_3305,N_2720);
nor U4160 (N_4160,N_2637,N_3027);
and U4161 (N_4161,N_3825,N_3560);
nand U4162 (N_4162,N_2555,N_3826);
or U4163 (N_4163,N_3968,N_2938);
and U4164 (N_4164,N_3221,N_2261);
nor U4165 (N_4165,N_3009,N_3527);
nor U4166 (N_4166,N_2227,N_2888);
nor U4167 (N_4167,N_2313,N_3859);
xnor U4168 (N_4168,N_2620,N_3603);
nand U4169 (N_4169,N_2622,N_3655);
nand U4170 (N_4170,N_3926,N_2632);
or U4171 (N_4171,N_2115,N_2783);
nor U4172 (N_4172,N_3074,N_2385);
xor U4173 (N_4173,N_3270,N_2569);
xor U4174 (N_4174,N_3385,N_2634);
and U4175 (N_4175,N_3494,N_3302);
nand U4176 (N_4176,N_2840,N_3649);
nand U4177 (N_4177,N_3828,N_2678);
and U4178 (N_4178,N_2315,N_2074);
nand U4179 (N_4179,N_3597,N_2661);
and U4180 (N_4180,N_2019,N_2098);
or U4181 (N_4181,N_3982,N_2347);
and U4182 (N_4182,N_2201,N_2195);
nand U4183 (N_4183,N_3444,N_2480);
or U4184 (N_4184,N_3257,N_3176);
nand U4185 (N_4185,N_2392,N_2924);
nand U4186 (N_4186,N_2225,N_3789);
or U4187 (N_4187,N_2600,N_3208);
and U4188 (N_4188,N_2314,N_2416);
or U4189 (N_4189,N_3613,N_3285);
xor U4190 (N_4190,N_2763,N_2983);
nor U4191 (N_4191,N_3061,N_2127);
nand U4192 (N_4192,N_3490,N_3557);
nor U4193 (N_4193,N_2507,N_3939);
or U4194 (N_4194,N_3843,N_3164);
nand U4195 (N_4195,N_3023,N_3413);
or U4196 (N_4196,N_2476,N_2739);
nand U4197 (N_4197,N_2207,N_3423);
nor U4198 (N_4198,N_2343,N_2899);
nand U4199 (N_4199,N_2269,N_2515);
or U4200 (N_4200,N_3238,N_2338);
nor U4201 (N_4201,N_3039,N_3646);
nand U4202 (N_4202,N_2485,N_3392);
or U4203 (N_4203,N_2420,N_2232);
nor U4204 (N_4204,N_2469,N_2846);
or U4205 (N_4205,N_2370,N_2824);
nor U4206 (N_4206,N_2725,N_3476);
xor U4207 (N_4207,N_3916,N_2893);
or U4208 (N_4208,N_2819,N_3190);
nor U4209 (N_4209,N_2962,N_2930);
nand U4210 (N_4210,N_3446,N_2167);
and U4211 (N_4211,N_2870,N_2541);
or U4212 (N_4212,N_3580,N_2386);
nor U4213 (N_4213,N_2880,N_2035);
or U4214 (N_4214,N_3163,N_2081);
nand U4215 (N_4215,N_3690,N_3155);
or U4216 (N_4216,N_2913,N_2120);
nand U4217 (N_4217,N_3932,N_3362);
or U4218 (N_4218,N_2835,N_3821);
and U4219 (N_4219,N_3521,N_3996);
nor U4220 (N_4220,N_2822,N_2245);
or U4221 (N_4221,N_2138,N_3054);
nor U4222 (N_4222,N_2987,N_3994);
and U4223 (N_4223,N_3263,N_2135);
and U4224 (N_4224,N_2009,N_2669);
and U4225 (N_4225,N_2890,N_2132);
nor U4226 (N_4226,N_3663,N_2272);
xnor U4227 (N_4227,N_3808,N_2670);
xnor U4228 (N_4228,N_2897,N_3680);
nand U4229 (N_4229,N_3220,N_2715);
nor U4230 (N_4230,N_2070,N_3820);
and U4231 (N_4231,N_3367,N_3518);
and U4232 (N_4232,N_2997,N_3505);
nor U4233 (N_4233,N_3427,N_3174);
or U4234 (N_4234,N_3345,N_2442);
or U4235 (N_4235,N_3712,N_3940);
or U4236 (N_4236,N_3858,N_3695);
nor U4237 (N_4237,N_3745,N_2176);
or U4238 (N_4238,N_2649,N_3377);
xor U4239 (N_4239,N_3052,N_2421);
nor U4240 (N_4240,N_3542,N_3851);
and U4241 (N_4241,N_2825,N_3210);
or U4242 (N_4242,N_3438,N_2797);
nor U4243 (N_4243,N_2658,N_2304);
nor U4244 (N_4244,N_2813,N_2296);
nand U4245 (N_4245,N_2690,N_3375);
nand U4246 (N_4246,N_2680,N_2355);
nand U4247 (N_4247,N_2441,N_3314);
nand U4248 (N_4248,N_2605,N_2438);
nor U4249 (N_4249,N_2571,N_2397);
nor U4250 (N_4250,N_3249,N_3410);
nor U4251 (N_4251,N_2321,N_2630);
or U4252 (N_4252,N_2547,N_2929);
nand U4253 (N_4253,N_3106,N_2538);
nand U4254 (N_4254,N_2625,N_3622);
or U4255 (N_4255,N_2185,N_2933);
nor U4256 (N_4256,N_3457,N_3643);
and U4257 (N_4257,N_2896,N_3230);
nand U4258 (N_4258,N_3801,N_3906);
nor U4259 (N_4259,N_3306,N_3525);
xnor U4260 (N_4260,N_2631,N_3216);
nor U4261 (N_4261,N_3236,N_2503);
or U4262 (N_4262,N_3454,N_3697);
nor U4263 (N_4263,N_2596,N_3517);
nor U4264 (N_4264,N_2744,N_2288);
nor U4265 (N_4265,N_2006,N_3123);
nand U4266 (N_4266,N_2801,N_2702);
nand U4267 (N_4267,N_2082,N_3065);
nand U4268 (N_4268,N_2124,N_2534);
or U4269 (N_4269,N_2436,N_2807);
nor U4270 (N_4270,N_2506,N_3855);
xnor U4271 (N_4271,N_3328,N_2970);
and U4272 (N_4272,N_3970,N_3895);
xnor U4273 (N_4273,N_3609,N_2184);
nor U4274 (N_4274,N_3685,N_2999);
and U4275 (N_4275,N_2092,N_2085);
nor U4276 (N_4276,N_3307,N_3831);
nor U4277 (N_4277,N_2532,N_2474);
and U4278 (N_4278,N_3172,N_3340);
or U4279 (N_4279,N_3567,N_3758);
nor U4280 (N_4280,N_2745,N_2060);
nand U4281 (N_4281,N_3089,N_3899);
xnor U4282 (N_4282,N_3313,N_2107);
and U4283 (N_4283,N_2121,N_3691);
nand U4284 (N_4284,N_2914,N_2494);
or U4285 (N_4285,N_2864,N_3938);
nand U4286 (N_4286,N_2434,N_3013);
or U4287 (N_4287,N_3749,N_3049);
nand U4288 (N_4288,N_3312,N_3402);
nand U4289 (N_4289,N_3639,N_2998);
nor U4290 (N_4290,N_3225,N_3275);
nand U4291 (N_4291,N_3272,N_3862);
nand U4292 (N_4292,N_2836,N_3359);
nor U4293 (N_4293,N_2295,N_2915);
nand U4294 (N_4294,N_2910,N_2738);
nor U4295 (N_4295,N_2348,N_3586);
and U4296 (N_4296,N_3894,N_2671);
nand U4297 (N_4297,N_2527,N_3287);
or U4298 (N_4298,N_2471,N_2278);
nand U4299 (N_4299,N_2640,N_3677);
nor U4300 (N_4300,N_3118,N_3610);
and U4301 (N_4301,N_3783,N_2781);
nor U4302 (N_4302,N_3806,N_3228);
or U4303 (N_4303,N_2165,N_2156);
nand U4304 (N_4304,N_2382,N_3688);
xor U4305 (N_4305,N_2390,N_3088);
and U4306 (N_4306,N_2465,N_3605);
nor U4307 (N_4307,N_2212,N_2950);
nand U4308 (N_4308,N_3759,N_2621);
or U4309 (N_4309,N_3874,N_2061);
nor U4310 (N_4310,N_2422,N_2034);
nand U4311 (N_4311,N_3987,N_3750);
or U4312 (N_4312,N_3589,N_2312);
nor U4313 (N_4313,N_3473,N_3226);
nand U4314 (N_4314,N_2618,N_3197);
nor U4315 (N_4315,N_2084,N_2437);
xnor U4316 (N_4316,N_2387,N_2829);
nor U4317 (N_4317,N_2130,N_2769);
nand U4318 (N_4318,N_2756,N_3563);
nor U4319 (N_4319,N_3376,N_3642);
and U4320 (N_4320,N_2777,N_2433);
and U4321 (N_4321,N_3246,N_2335);
nand U4322 (N_4322,N_2286,N_2667);
or U4323 (N_4323,N_3844,N_3028);
and U4324 (N_4324,N_3883,N_3516);
or U4325 (N_4325,N_2707,N_2451);
and U4326 (N_4326,N_2361,N_3692);
and U4327 (N_4327,N_3421,N_3479);
and U4328 (N_4328,N_3999,N_2307);
nand U4329 (N_4329,N_2758,N_3682);
nand U4330 (N_4330,N_3433,N_3540);
and U4331 (N_4331,N_2908,N_2719);
or U4332 (N_4332,N_2692,N_3031);
nor U4333 (N_4333,N_3370,N_2216);
nor U4334 (N_4334,N_2652,N_3952);
and U4335 (N_4335,N_3046,N_2821);
nor U4336 (N_4336,N_2577,N_2619);
and U4337 (N_4337,N_2643,N_2776);
or U4338 (N_4338,N_2832,N_2816);
nor U4339 (N_4339,N_2844,N_3656);
or U4340 (N_4340,N_2627,N_3056);
and U4341 (N_4341,N_3924,N_2511);
nand U4342 (N_4342,N_3588,N_3592);
nand U4343 (N_4343,N_3425,N_3788);
or U4344 (N_4344,N_2255,N_3877);
or U4345 (N_4345,N_2737,N_2066);
nand U4346 (N_4346,N_3953,N_3757);
nor U4347 (N_4347,N_2375,N_2991);
nand U4348 (N_4348,N_2965,N_2525);
or U4349 (N_4349,N_2331,N_2391);
xor U4350 (N_4350,N_3623,N_3439);
or U4351 (N_4351,N_2181,N_2337);
nand U4352 (N_4352,N_3577,N_3565);
or U4353 (N_4353,N_3528,N_3321);
and U4354 (N_4354,N_3011,N_3575);
xnor U4355 (N_4355,N_3149,N_2704);
nand U4356 (N_4356,N_2410,N_3583);
or U4357 (N_4357,N_3295,N_3645);
nand U4358 (N_4358,N_2767,N_3409);
and U4359 (N_4359,N_2936,N_2570);
xnor U4360 (N_4360,N_2689,N_2016);
xor U4361 (N_4361,N_3718,N_2543);
nand U4362 (N_4362,N_2332,N_3519);
and U4363 (N_4363,N_3668,N_2664);
nor U4364 (N_4364,N_3019,N_3523);
or U4365 (N_4365,N_3395,N_2125);
and U4366 (N_4366,N_3404,N_3291);
and U4367 (N_4367,N_2530,N_2500);
and U4368 (N_4368,N_3142,N_2323);
and U4369 (N_4369,N_2654,N_3672);
and U4370 (N_4370,N_3202,N_3529);
or U4371 (N_4371,N_2202,N_3441);
or U4372 (N_4372,N_3048,N_2700);
nor U4373 (N_4373,N_2100,N_3256);
and U4374 (N_4374,N_2894,N_3555);
or U4375 (N_4375,N_3465,N_3841);
or U4376 (N_4376,N_3886,N_2126);
nor U4377 (N_4377,N_2523,N_2136);
or U4378 (N_4378,N_2542,N_3524);
nand U4379 (N_4379,N_3286,N_2754);
nand U4380 (N_4380,N_3770,N_2475);
or U4381 (N_4381,N_2306,N_2992);
xnor U4382 (N_4382,N_3568,N_2007);
nand U4383 (N_4383,N_3390,N_3374);
nand U4384 (N_4384,N_2254,N_2563);
or U4385 (N_4385,N_3727,N_2927);
nor U4386 (N_4386,N_3360,N_2488);
and U4387 (N_4387,N_2979,N_2882);
or U4388 (N_4388,N_3635,N_2460);
nor U4389 (N_4389,N_2320,N_2633);
nand U4390 (N_4390,N_3991,N_2898);
and U4391 (N_4391,N_3461,N_2602);
and U4392 (N_4392,N_3449,N_2097);
nor U4393 (N_4393,N_3258,N_2157);
nor U4394 (N_4394,N_2153,N_3949);
nor U4395 (N_4395,N_3021,N_2903);
nor U4396 (N_4396,N_3195,N_2610);
and U4397 (N_4397,N_3292,N_3937);
and U4398 (N_4398,N_3405,N_3248);
and U4399 (N_4399,N_2440,N_2714);
and U4400 (N_4400,N_3971,N_2635);
and U4401 (N_4401,N_2379,N_3958);
nor U4402 (N_4402,N_2663,N_3017);
nand U4403 (N_4403,N_3218,N_2583);
or U4404 (N_4404,N_2265,N_2883);
nand U4405 (N_4405,N_2952,N_3393);
xnor U4406 (N_4406,N_2709,N_2473);
or U4407 (N_4407,N_2900,N_3902);
or U4408 (N_4408,N_2662,N_2855);
nand U4409 (N_4409,N_3353,N_3863);
and U4410 (N_4410,N_2966,N_3244);
nand U4411 (N_4411,N_3945,N_3403);
nor U4412 (N_4412,N_3495,N_3412);
nor U4413 (N_4413,N_2114,N_2164);
nor U4414 (N_4414,N_2453,N_2857);
nor U4415 (N_4415,N_2484,N_2468);
or U4416 (N_4416,N_2400,N_3304);
nand U4417 (N_4417,N_3103,N_2526);
nand U4418 (N_4418,N_2148,N_2863);
and U4419 (N_4419,N_2291,N_2067);
nor U4420 (N_4420,N_3811,N_2012);
and U4421 (N_4421,N_3191,N_2064);
nand U4422 (N_4422,N_3870,N_3364);
and U4423 (N_4423,N_2376,N_2311);
or U4424 (N_4424,N_3710,N_3929);
nor U4425 (N_4425,N_3612,N_2943);
or U4426 (N_4426,N_3878,N_3711);
nor U4427 (N_4427,N_2743,N_3299);
and U4428 (N_4428,N_3797,N_2310);
nand U4429 (N_4429,N_3110,N_3325);
or U4430 (N_4430,N_3865,N_2219);
nor U4431 (N_4431,N_3179,N_3332);
and U4432 (N_4432,N_3606,N_2705);
and U4433 (N_4433,N_3265,N_2706);
nor U4434 (N_4434,N_2106,N_3349);
nand U4435 (N_4435,N_3867,N_2172);
and U4436 (N_4436,N_3171,N_3098);
and U4437 (N_4437,N_2193,N_2224);
nor U4438 (N_4438,N_3232,N_3782);
nor U4439 (N_4439,N_2076,N_3747);
and U4440 (N_4440,N_3678,N_3193);
or U4441 (N_4441,N_2033,N_3255);
nand U4442 (N_4442,N_3008,N_2684);
or U4443 (N_4443,N_2886,N_2065);
or U4444 (N_4444,N_2008,N_2431);
and U4445 (N_4445,N_2996,N_3175);
nor U4446 (N_4446,N_2757,N_2727);
xor U4447 (N_4447,N_3060,N_3834);
or U4448 (N_4448,N_2283,N_2806);
and U4449 (N_4449,N_3761,N_3474);
nor U4450 (N_4450,N_2617,N_3957);
or U4451 (N_4451,N_3501,N_3201);
nor U4452 (N_4452,N_3918,N_3319);
nand U4453 (N_4453,N_2359,N_3633);
or U4454 (N_4454,N_2398,N_2772);
and U4455 (N_4455,N_3729,N_3016);
nor U4456 (N_4456,N_3925,N_3401);
nor U4457 (N_4457,N_3116,N_2450);
or U4458 (N_4458,N_2292,N_2584);
xnor U4459 (N_4459,N_3062,N_3621);
or U4460 (N_4460,N_3754,N_3660);
nor U4461 (N_4461,N_3810,N_2567);
nand U4462 (N_4462,N_3105,N_2169);
nor U4463 (N_4463,N_2023,N_3892);
and U4464 (N_4464,N_3041,N_3076);
and U4465 (N_4465,N_3815,N_3599);
and U4466 (N_4466,N_3085,N_2319);
nand U4467 (N_4467,N_2588,N_2934);
or U4468 (N_4468,N_3124,N_2834);
and U4469 (N_4469,N_3662,N_3531);
nor U4470 (N_4470,N_3620,N_2149);
and U4471 (N_4471,N_2694,N_3984);
and U4472 (N_4472,N_3430,N_3864);
nor U4473 (N_4473,N_3667,N_3978);
xnor U4474 (N_4474,N_3003,N_2580);
xnor U4475 (N_4475,N_3536,N_3145);
and U4476 (N_4476,N_2145,N_3616);
or U4477 (N_4477,N_3007,N_3989);
or U4478 (N_4478,N_2673,N_3167);
xor U4479 (N_4479,N_2792,N_3653);
nor U4480 (N_4480,N_3960,N_3000);
or U4481 (N_4481,N_3135,N_2247);
xor U4482 (N_4482,N_2809,N_2191);
or U4483 (N_4483,N_2603,N_3716);
nor U4484 (N_4484,N_2803,N_2211);
and U4485 (N_4485,N_2795,N_2875);
nand U4486 (N_4486,N_2143,N_3629);
or U4487 (N_4487,N_3147,N_3186);
nor U4488 (N_4488,N_2078,N_3852);
xnor U4489 (N_4489,N_3659,N_3466);
nand U4490 (N_4490,N_2736,N_2217);
nor U4491 (N_4491,N_2194,N_3868);
or U4492 (N_4492,N_2305,N_3652);
nand U4493 (N_4493,N_3551,N_3506);
nor U4494 (N_4494,N_3824,N_2682);
or U4495 (N_4495,N_3114,N_2648);
nand U4496 (N_4496,N_2647,N_3676);
nand U4497 (N_4497,N_2802,N_2325);
and U4498 (N_4498,N_2514,N_3698);
or U4499 (N_4499,N_3322,N_2188);
nor U4500 (N_4500,N_2729,N_2592);
or U4501 (N_4501,N_3361,N_3823);
nor U4502 (N_4502,N_2545,N_3338);
and U4503 (N_4503,N_2179,N_3566);
or U4504 (N_4504,N_2365,N_2582);
or U4505 (N_4505,N_3814,N_2884);
nor U4506 (N_4506,N_3552,N_3569);
or U4507 (N_4507,N_2274,N_3470);
nand U4508 (N_4508,N_3976,N_2140);
nand U4509 (N_4509,N_2942,N_3120);
and U4510 (N_4510,N_3032,N_2287);
nand U4511 (N_4511,N_2449,N_3481);
nor U4512 (N_4512,N_2470,N_2578);
and U4513 (N_4513,N_2939,N_2038);
nor U4514 (N_4514,N_3608,N_3252);
nor U4515 (N_4515,N_3647,N_3150);
nor U4516 (N_4516,N_2259,N_3813);
nor U4517 (N_4517,N_2871,N_2443);
or U4518 (N_4518,N_2456,N_3012);
and U4519 (N_4519,N_3790,N_2119);
and U4520 (N_4520,N_3836,N_3590);
nand U4521 (N_4521,N_3857,N_3879);
xor U4522 (N_4522,N_2206,N_3966);
or U4523 (N_4523,N_2773,N_3354);
nor U4524 (N_4524,N_3961,N_3775);
or U4525 (N_4525,N_2103,N_2171);
and U4526 (N_4526,N_2113,N_3804);
nand U4527 (N_4527,N_3132,N_2830);
xor U4528 (N_4528,N_2782,N_3627);
nor U4529 (N_4529,N_3480,N_3717);
xnor U4530 (N_4530,N_3383,N_2353);
nor U4531 (N_4531,N_3556,N_2482);
nand U4532 (N_4532,N_2056,N_3723);
or U4533 (N_4533,N_2235,N_2024);
xnor U4534 (N_4534,N_2215,N_2749);
and U4535 (N_4535,N_2685,N_3250);
or U4536 (N_4536,N_3995,N_2876);
and U4537 (N_4537,N_2976,N_3204);
and U4538 (N_4538,N_3290,N_3876);
nand U4539 (N_4539,N_2277,N_3604);
and U4540 (N_4540,N_2344,N_2808);
nor U4541 (N_4541,N_3993,N_3188);
and U4542 (N_4542,N_3184,N_3909);
nor U4543 (N_4543,N_3777,N_2182);
nand U4544 (N_4544,N_3830,N_3203);
nand U4545 (N_4545,N_3206,N_2520);
and U4546 (N_4546,N_3358,N_3477);
xnor U4547 (N_4547,N_3822,N_2959);
and U4548 (N_4548,N_3936,N_3547);
nand U4549 (N_4549,N_3077,N_3998);
or U4550 (N_4550,N_3708,N_3484);
xnor U4551 (N_4551,N_2221,N_2406);
and U4552 (N_4552,N_3755,N_2152);
nand U4553 (N_4553,N_3399,N_3211);
and U4554 (N_4554,N_3615,N_2862);
nand U4555 (N_4555,N_2901,N_3200);
nor U4556 (N_4556,N_2595,N_2096);
and U4557 (N_4557,N_2613,N_3915);
xor U4558 (N_4558,N_3273,N_2297);
nor U4559 (N_4559,N_3288,N_2384);
or U4560 (N_4560,N_3545,N_2660);
xor U4561 (N_4561,N_3180,N_3407);
and U4562 (N_4562,N_3975,N_3559);
nor U4563 (N_4563,N_3239,N_2053);
or U4564 (N_4564,N_2693,N_3366);
and U4565 (N_4565,N_3406,N_3942);
nand U4566 (N_4566,N_3297,N_2606);
nand U4567 (N_4567,N_3666,N_3784);
and U4568 (N_4568,N_2590,N_3764);
nor U4569 (N_4569,N_3386,N_2837);
and U4570 (N_4570,N_2116,N_2233);
and U4571 (N_4571,N_3795,N_3271);
nand U4572 (N_4572,N_2838,N_2010);
nand U4573 (N_4573,N_2574,N_2205);
nor U4574 (N_4574,N_3102,N_2089);
nor U4575 (N_4575,N_2512,N_3337);
nor U4576 (N_4576,N_3224,N_2162);
nor U4577 (N_4577,N_3838,N_2612);
or U4578 (N_4578,N_3986,N_3796);
or U4579 (N_4579,N_3928,N_2874);
and U4580 (N_4580,N_3735,N_3094);
or U4581 (N_4581,N_2303,N_2213);
and U4582 (N_4582,N_2133,N_2128);
nand U4583 (N_4583,N_2251,N_2377);
or U4584 (N_4584,N_2753,N_2963);
nand U4585 (N_4585,N_3237,N_2021);
nor U4586 (N_4586,N_3158,N_2636);
xor U4587 (N_4587,N_3347,N_3679);
and U4588 (N_4588,N_3829,N_2015);
or U4589 (N_4589,N_3869,N_3985);
nand U4590 (N_4590,N_3242,N_3159);
nor U4591 (N_4591,N_2242,N_3748);
nor U4592 (N_4592,N_3890,N_3381);
or U4593 (N_4593,N_2746,N_2154);
xor U4594 (N_4594,N_3429,N_2137);
nand U4595 (N_4595,N_2764,N_2740);
or U4596 (N_4596,N_3935,N_2614);
nor U4597 (N_4597,N_2159,N_2833);
or U4598 (N_4598,N_2505,N_2432);
nand U4599 (N_4599,N_3919,N_3561);
or U4600 (N_4600,N_2866,N_3006);
nand U4601 (N_4601,N_3884,N_2183);
nor U4602 (N_4602,N_3318,N_2794);
or U4603 (N_4603,N_2094,N_3097);
or U4604 (N_4604,N_3756,N_2395);
nor U4605 (N_4605,N_3840,N_2253);
xnor U4606 (N_4606,N_3654,N_2293);
or U4607 (N_4607,N_2868,N_3571);
or U4608 (N_4608,N_3253,N_3772);
nand U4609 (N_4609,N_3963,N_3946);
nor U4610 (N_4610,N_3455,N_3199);
nor U4611 (N_4611,N_2151,N_2529);
xor U4612 (N_4612,N_3640,N_2887);
or U4613 (N_4613,N_2659,N_2246);
and U4614 (N_4614,N_3681,N_2025);
xnor U4615 (N_4615,N_2498,N_2336);
nand U4616 (N_4616,N_2766,N_2916);
nor U4617 (N_4617,N_3327,N_3730);
or U4618 (N_4618,N_3973,N_2623);
nor U4619 (N_4619,N_2051,N_3907);
nor U4620 (N_4620,N_2284,N_3010);
and U4621 (N_4621,N_2645,N_3357);
xor U4622 (N_4622,N_3927,N_2747);
nand U4623 (N_4623,N_2075,N_3266);
and U4624 (N_4624,N_2810,N_3140);
xnor U4625 (N_4625,N_3391,N_3047);
and U4626 (N_4626,N_2881,N_2522);
nor U4627 (N_4627,N_3847,N_2572);
nor U4628 (N_4628,N_3778,N_3445);
and U4629 (N_4629,N_3722,N_2175);
xnor U4630 (N_4630,N_3948,N_3914);
nand U4631 (N_4631,N_2285,N_3980);
or U4632 (N_4632,N_2150,N_2774);
or U4633 (N_4633,N_3153,N_3411);
and U4634 (N_4634,N_2755,N_2701);
and U4635 (N_4635,N_3732,N_3117);
and U4636 (N_4636,N_2405,N_2827);
nand U4637 (N_4637,N_2741,N_2905);
and U4638 (N_4638,N_2079,N_3744);
xor U4639 (N_4639,N_2666,N_3507);
or U4640 (N_4640,N_3450,N_3380);
nand U4641 (N_4641,N_3078,N_3166);
nor U4642 (N_4642,N_2497,N_2985);
or U4643 (N_4643,N_2537,N_3600);
nor U4644 (N_4644,N_3254,N_3839);
or U4645 (N_4645,N_2461,N_3515);
or U4646 (N_4646,N_2585,N_2299);
and U4647 (N_4647,N_2057,N_3805);
xnor U4648 (N_4648,N_2279,N_3329);
nor U4649 (N_4649,N_3794,N_3241);
xor U4650 (N_4650,N_3452,N_3245);
and U4651 (N_4651,N_3296,N_3786);
nor U4652 (N_4652,N_2818,N_3848);
or U4653 (N_4653,N_3702,N_2424);
or U4654 (N_4654,N_3101,N_2328);
nor U4655 (N_4655,N_3626,N_2200);
or U4656 (N_4656,N_3231,N_2142);
or U4657 (N_4657,N_2462,N_2000);
nand U4658 (N_4658,N_2519,N_2131);
nor U4659 (N_4659,N_3064,N_3243);
and U4660 (N_4660,N_3100,N_3651);
nand U4661 (N_4661,N_3944,N_3699);
nand U4662 (N_4662,N_3492,N_2691);
nor U4663 (N_4663,N_3572,N_3720);
nor U4664 (N_4664,N_3703,N_3636);
nor U4665 (N_4665,N_3125,N_3689);
and U4666 (N_4666,N_2447,N_2080);
and U4667 (N_4667,N_3675,N_2044);
or U4668 (N_4668,N_2403,N_3550);
xnor U4669 (N_4669,N_2351,N_3553);
and U4670 (N_4670,N_2814,N_3151);
nor U4671 (N_4671,N_2516,N_3832);
nand U4672 (N_4672,N_3067,N_3619);
or U4673 (N_4673,N_3921,N_3344);
or U4674 (N_4674,N_3800,N_2364);
xnor U4675 (N_4675,N_3705,N_3860);
or U4676 (N_4676,N_2940,N_3152);
nand U4677 (N_4677,N_3974,N_2220);
or U4678 (N_4678,N_2013,N_2091);
nor U4679 (N_4679,N_3034,N_2931);
or U4680 (N_4680,N_3363,N_3534);
or U4681 (N_4681,N_3055,N_3170);
or U4682 (N_4682,N_3099,N_2027);
and U4683 (N_4683,N_2964,N_3896);
or U4684 (N_4684,N_3276,N_3893);
and U4685 (N_4685,N_2040,N_3768);
or U4686 (N_4686,N_2260,N_2904);
or U4687 (N_4687,N_2724,N_2731);
or U4688 (N_4688,N_3508,N_2146);
and U4689 (N_4689,N_2995,N_3072);
and U4690 (N_4690,N_3714,N_3866);
nand U4691 (N_4691,N_3025,N_3564);
xor U4692 (N_4692,N_2641,N_2878);
and U4693 (N_4693,N_2811,N_2556);
nand U4694 (N_4694,N_2672,N_2463);
or U4695 (N_4695,N_3875,N_3596);
nor U4696 (N_4696,N_3259,N_2372);
nand U4697 (N_4697,N_3214,N_3093);
or U4698 (N_4698,N_2728,N_3223);
and U4699 (N_4699,N_2454,N_2676);
or U4700 (N_4700,N_2426,N_3045);
or U4701 (N_4701,N_3526,N_2177);
and U4702 (N_4702,N_2907,N_2383);
or U4703 (N_4703,N_2155,N_2349);
nand U4704 (N_4704,N_3264,N_3382);
nor U4705 (N_4705,N_2581,N_2270);
nor U4706 (N_4706,N_2817,N_3601);
xor U4707 (N_4707,N_2088,N_3650);
or U4708 (N_4708,N_2112,N_3614);
nor U4709 (N_4709,N_3108,N_3488);
nand U4710 (N_4710,N_2586,N_2280);
nor U4711 (N_4711,N_2036,N_3954);
nand U4712 (N_4712,N_3497,N_2687);
nand U4713 (N_4713,N_3282,N_3644);
or U4714 (N_4714,N_2178,N_3209);
nor U4715 (N_4715,N_2854,N_3284);
nand U4716 (N_4716,N_3709,N_3502);
and U4717 (N_4717,N_3030,N_3187);
nor U4718 (N_4718,N_2222,N_2650);
nor U4719 (N_4719,N_2282,N_3051);
nor U4720 (N_4720,N_3493,N_3368);
or U4721 (N_4721,N_2401,N_3522);
nand U4722 (N_4722,N_2363,N_2841);
and U4723 (N_4723,N_3475,N_3351);
nand U4724 (N_4724,N_2922,N_3584);
nor U4725 (N_4725,N_3503,N_3951);
and U4726 (N_4726,N_3424,N_3126);
and U4727 (N_4727,N_3113,N_2919);
nor U4728 (N_4728,N_2521,N_2020);
and U4729 (N_4729,N_3415,N_3388);
nor U4730 (N_4730,N_2858,N_2334);
nand U4731 (N_4731,N_3063,N_2954);
nor U4732 (N_4732,N_3981,N_2860);
xor U4733 (N_4733,N_2918,N_3059);
or U4734 (N_4734,N_3020,N_3607);
nor U4735 (N_4735,N_2760,N_3737);
nor U4736 (N_4736,N_3817,N_3121);
or U4737 (N_4737,N_3369,N_3913);
nor U4738 (N_4738,N_3882,N_2624);
or U4739 (N_4739,N_2902,N_2356);
and U4740 (N_4740,N_2546,N_3139);
nor U4741 (N_4741,N_2243,N_2486);
or U4742 (N_4742,N_3469,N_2073);
or U4743 (N_4743,N_3904,N_3769);
or U4744 (N_4744,N_3871,N_2446);
or U4745 (N_4745,N_3129,N_3091);
nand U4746 (N_4746,N_2415,N_2003);
or U4747 (N_4747,N_3842,N_2851);
nor U4748 (N_4748,N_2435,N_2239);
or U4749 (N_4749,N_3664,N_2768);
or U4750 (N_4750,N_2457,N_3641);
nor U4751 (N_4751,N_2099,N_2231);
and U4752 (N_4752,N_2524,N_2324);
nor U4753 (N_4753,N_2990,N_2550);
or U4754 (N_4754,N_2492,N_2039);
or U4755 (N_4755,N_3372,N_3611);
nand U4756 (N_4756,N_3934,N_3498);
or U4757 (N_4757,N_3753,N_3514);
nor U4758 (N_4758,N_3739,N_3897);
nor U4759 (N_4759,N_2608,N_3979);
nor U4760 (N_4760,N_3977,N_3715);
nor U4761 (N_4761,N_3487,N_3154);
or U4762 (N_4762,N_2309,N_3437);
nand U4763 (N_4763,N_2865,N_2948);
nand U4764 (N_4764,N_3765,N_2852);
nor U4765 (N_4765,N_2249,N_2077);
nor U4766 (N_4766,N_3431,N_3137);
or U4767 (N_4767,N_3472,N_3310);
or U4768 (N_4768,N_3417,N_2828);
or U4769 (N_4769,N_2859,N_2941);
xor U4770 (N_4770,N_2380,N_3394);
xor U4771 (N_4771,N_3969,N_2174);
and U4772 (N_4772,N_2298,N_3022);
or U4773 (N_4773,N_3819,N_3543);
and U4774 (N_4774,N_2101,N_2049);
or U4775 (N_4775,N_2750,N_2052);
and U4776 (N_4776,N_2842,N_2716);
nor U4777 (N_4777,N_2502,N_3182);
nand U4778 (N_4778,N_3704,N_3348);
nand U4779 (N_4779,N_2759,N_3156);
nand U4780 (N_4780,N_3213,N_3339);
nor U4781 (N_4781,N_2926,N_3992);
nand U4782 (N_4782,N_2607,N_3911);
or U4783 (N_4783,N_3458,N_2710);
nand U4784 (N_4784,N_3835,N_3026);
or U4785 (N_4785,N_2872,N_3268);
and U4786 (N_4786,N_2369,N_2791);
or U4787 (N_4787,N_3092,N_3235);
nor U4788 (N_4788,N_3141,N_2501);
and U4789 (N_4789,N_3133,N_3731);
nor U4790 (N_4790,N_3227,N_3593);
nor U4791 (N_4791,N_3058,N_2339);
nand U4792 (N_4792,N_2697,N_2346);
nand U4793 (N_4793,N_2848,N_2975);
nand U4794 (N_4794,N_2173,N_2322);
nand U4795 (N_4795,N_3434,N_2417);
nor U4796 (N_4796,N_2117,N_3632);
nand U4797 (N_4797,N_3504,N_2071);
nor U4798 (N_4798,N_2770,N_3451);
and U4799 (N_4799,N_2548,N_2168);
or U4800 (N_4800,N_2017,N_3693);
nor U4801 (N_4801,N_3736,N_2686);
or U4802 (N_4802,N_3910,N_2252);
and U4803 (N_4803,N_3683,N_3891);
nor U4804 (N_4804,N_2004,N_3323);
and U4805 (N_4805,N_3947,N_2257);
nor U4806 (N_4806,N_2598,N_2597);
nand U4807 (N_4807,N_3192,N_2411);
and U4808 (N_4808,N_2002,N_2508);
nand U4809 (N_4809,N_2703,N_3549);
xnor U4810 (N_4810,N_3420,N_3086);
nand U4811 (N_4811,N_3943,N_2093);
and U4812 (N_4812,N_2419,N_3760);
nand U4813 (N_4813,N_2289,N_3082);
and U4814 (N_4814,N_2055,N_2428);
and U4815 (N_4815,N_2533,N_3955);
or U4816 (N_4816,N_3684,N_2477);
nor U4817 (N_4817,N_3885,N_3574);
or U4818 (N_4818,N_3743,N_2198);
nand U4819 (N_4819,N_3442,N_3837);
or U4820 (N_4820,N_2108,N_3558);
nand U4821 (N_4821,N_3262,N_3538);
nor U4822 (N_4822,N_2459,N_3617);
or U4823 (N_4823,N_2412,N_2366);
nand U4824 (N_4824,N_3422,N_2751);
xor U4825 (N_4825,N_2712,N_2722);
and U4826 (N_4826,N_3579,N_3207);
or U4827 (N_4827,N_2562,N_2373);
and U4828 (N_4828,N_3037,N_3827);
nor U4829 (N_4829,N_3922,N_2849);
and U4830 (N_4830,N_3198,N_2032);
and U4831 (N_4831,N_3513,N_2166);
nand U4832 (N_4832,N_2993,N_2557);
nand U4833 (N_4833,N_2256,N_2109);
and U4834 (N_4834,N_3298,N_2787);
and U4835 (N_4835,N_2788,N_3194);
nand U4836 (N_4836,N_2086,N_3774);
and U4837 (N_4837,N_3462,N_2378);
nand U4838 (N_4838,N_3776,N_3173);
nor U4839 (N_4839,N_3923,N_2911);
nor U4840 (N_4840,N_3905,N_2326);
and U4841 (N_4841,N_3267,N_2180);
or U4842 (N_4842,N_2554,N_3740);
nor U4843 (N_4843,N_2593,N_2793);
nand U4844 (N_4844,N_2616,N_3872);
or U4845 (N_4845,N_3090,N_3491);
nor U4846 (N_4846,N_3084,N_3096);
nand U4847 (N_4847,N_2129,N_2644);
nor U4848 (N_4848,N_2784,N_2263);
nor U4849 (N_4849,N_3080,N_3071);
nor U4850 (N_4850,N_2439,N_3042);
and U4851 (N_4851,N_3460,N_2980);
nor U4852 (N_4852,N_2638,N_2576);
xnor U4853 (N_4853,N_3229,N_3941);
and U4854 (N_4854,N_3793,N_3247);
and U4855 (N_4855,N_2812,N_3988);
nor U4856 (N_4856,N_3281,N_2244);
xnor U4857 (N_4857,N_3541,N_3818);
or U4858 (N_4858,N_2906,N_2721);
and U4859 (N_4859,N_2831,N_2973);
nand U4860 (N_4860,N_2742,N_2268);
nand U4861 (N_4861,N_3850,N_2711);
nand U4862 (N_4862,N_2301,N_2276);
or U4863 (N_4863,N_2726,N_3888);
xnor U4864 (N_4864,N_3136,N_2264);
nor U4865 (N_4865,N_3109,N_2199);
nor U4866 (N_4866,N_3746,N_3280);
nor U4867 (N_4867,N_2455,N_3396);
and U4868 (N_4868,N_3024,N_2068);
nor U4869 (N_4869,N_2513,N_2951);
and U4870 (N_4870,N_2796,N_3389);
and U4871 (N_4871,N_2396,N_2043);
nor U4872 (N_4872,N_2104,N_2873);
nand U4873 (N_4873,N_3648,N_2026);
nor U4874 (N_4874,N_2856,N_2238);
and U4875 (N_4875,N_3751,N_3816);
nor U4876 (N_4876,N_3972,N_2642);
nor U4877 (N_4877,N_3081,N_2628);
or U4878 (N_4878,N_2561,N_3582);
nor U4879 (N_4879,N_2565,N_3482);
or U4880 (N_4880,N_3350,N_3352);
nand U4881 (N_4881,N_2611,N_2601);
nor U4882 (N_4882,N_3812,N_2362);
nor U4883 (N_4883,N_2022,N_3530);
or U4884 (N_4884,N_3068,N_2820);
and U4885 (N_4885,N_2944,N_2489);
nand U4886 (N_4886,N_2699,N_3785);
or U4887 (N_4887,N_2425,N_2974);
and U4888 (N_4888,N_2063,N_3489);
nor U4889 (N_4889,N_2472,N_2674);
or U4890 (N_4890,N_3807,N_2945);
or U4891 (N_4891,N_3889,N_3724);
or U4892 (N_4892,N_3373,N_3112);
nand U4893 (N_4893,N_3301,N_2029);
nor U4894 (N_4894,N_3397,N_3537);
nor U4895 (N_4895,N_2483,N_3512);
or U4896 (N_4896,N_2158,N_3418);
xor U4897 (N_4897,N_2789,N_2144);
or U4898 (N_4898,N_2518,N_3127);
nand U4899 (N_4899,N_2427,N_3665);
nand U4900 (N_4900,N_2228,N_3846);
nor U4901 (N_4901,N_3311,N_2374);
or U4902 (N_4902,N_2028,N_3087);
nand U4903 (N_4903,N_2458,N_3500);
or U4904 (N_4904,N_2358,N_2675);
and U4905 (N_4905,N_2407,N_2609);
nor U4906 (N_4906,N_3157,N_2041);
nor U4907 (N_4907,N_3130,N_3440);
or U4908 (N_4908,N_3741,N_2045);
and U4909 (N_4909,N_3887,N_2935);
nand U4910 (N_4910,N_3721,N_3234);
nor U4911 (N_4911,N_3694,N_3083);
or U4912 (N_4912,N_2853,N_3792);
xor U4913 (N_4913,N_2448,N_3468);
or U4914 (N_4914,N_2241,N_3570);
and U4915 (N_4915,N_2657,N_2408);
and U4916 (N_4916,N_2615,N_2735);
or U4917 (N_4917,N_3554,N_2949);
and U4918 (N_4918,N_3432,N_2560);
xor U4919 (N_4919,N_2867,N_2290);
or U4920 (N_4920,N_2210,N_2300);
or U4921 (N_4921,N_2734,N_2957);
nor U4922 (N_4922,N_3165,N_3674);
xor U4923 (N_4923,N_3573,N_3183);
nor U4924 (N_4924,N_3854,N_3029);
and U4925 (N_4925,N_3752,N_3075);
or U4926 (N_4926,N_2499,N_3631);
xor U4927 (N_4927,N_2971,N_2559);
and U4928 (N_4928,N_3908,N_3004);
nor U4929 (N_4929,N_2695,N_2826);
nor U4930 (N_4930,N_3040,N_2912);
nor U4931 (N_4931,N_2418,N_2961);
or U4932 (N_4932,N_3881,N_2790);
nand U4933 (N_4933,N_3215,N_2250);
or U4934 (N_4934,N_3002,N_2388);
nor U4935 (N_4935,N_3131,N_3576);
and U4936 (N_4936,N_3673,N_3696);
nor U4937 (N_4937,N_3853,N_2909);
nand U4938 (N_4938,N_3320,N_3219);
nand U4939 (N_4939,N_2271,N_3861);
nor U4940 (N_4940,N_2847,N_2234);
and U4941 (N_4941,N_2160,N_2589);
and U4942 (N_4942,N_2989,N_2394);
and U4943 (N_4943,N_2696,N_2031);
or U4944 (N_4944,N_2732,N_2030);
xor U4945 (N_4945,N_2920,N_2308);
and U4946 (N_4946,N_2845,N_2698);
and U4947 (N_4947,N_2197,N_3104);
xor U4948 (N_4948,N_2762,N_2604);
nor U4949 (N_4949,N_2804,N_2204);
and U4950 (N_4950,N_3933,N_3532);
nor U4951 (N_4951,N_2752,N_2677);
nor U4952 (N_4952,N_2248,N_2564);
nand U4953 (N_4953,N_2317,N_2236);
nor U4954 (N_4954,N_2237,N_3341);
and U4955 (N_4955,N_2196,N_2861);
nand U4956 (N_4956,N_2510,N_2478);
nor U4957 (N_4957,N_3585,N_3119);
or U4958 (N_4958,N_3283,N_3289);
nand U4959 (N_4959,N_2208,N_2229);
nand U4960 (N_4960,N_2730,N_3294);
and U4961 (N_4961,N_3128,N_2490);
nor U4962 (N_4962,N_3967,N_2275);
and U4963 (N_4963,N_3456,N_2493);
nor U4964 (N_4964,N_3625,N_2496);
nor U4965 (N_4965,N_3138,N_2005);
or U4966 (N_4966,N_3669,N_2723);
nand U4967 (N_4967,N_2587,N_2226);
and U4968 (N_4968,N_3738,N_3464);
nand U4969 (N_4969,N_2780,N_2599);
and U4970 (N_4970,N_3956,N_3901);
and U4971 (N_4971,N_2357,N_3467);
nor U4972 (N_4972,N_2105,N_2042);
or U4973 (N_4973,N_3335,N_3177);
and U4974 (N_4974,N_3725,N_2994);
and U4975 (N_4975,N_2646,N_2327);
nor U4976 (N_4976,N_3880,N_2544);
and U4977 (N_4977,N_2575,N_2087);
and U4978 (N_4978,N_3196,N_2163);
xor U4979 (N_4979,N_2302,N_2481);
or U4980 (N_4980,N_3562,N_2733);
nand U4981 (N_4981,N_2877,N_2932);
nand U4982 (N_4982,N_2800,N_3143);
and U4983 (N_4983,N_2549,N_3595);
nor U4984 (N_4984,N_3205,N_2889);
and U4985 (N_4985,N_2892,N_2953);
nand U4986 (N_4986,N_2192,N_2371);
or U4987 (N_4987,N_3169,N_3628);
nor U4988 (N_4988,N_3780,N_2958);
xnor U4989 (N_4989,N_2316,N_2955);
nor U4990 (N_4990,N_2014,N_2059);
nand U4991 (N_4991,N_3426,N_3043);
nand U4992 (N_4992,N_3095,N_3168);
or U4993 (N_4993,N_3634,N_3300);
nand U4994 (N_4994,N_3400,N_3898);
xor U4995 (N_4995,N_3728,N_3073);
and U4996 (N_4996,N_2381,N_3419);
xnor U4997 (N_4997,N_2170,N_3781);
and U4998 (N_4998,N_2946,N_3279);
nand U4999 (N_4999,N_3014,N_3181);
and U5000 (N_5000,N_3755,N_2966);
or U5001 (N_5001,N_2936,N_3299);
or U5002 (N_5002,N_2115,N_3110);
nor U5003 (N_5003,N_2790,N_3258);
and U5004 (N_5004,N_3136,N_3314);
and U5005 (N_5005,N_2564,N_3095);
and U5006 (N_5006,N_3784,N_2842);
or U5007 (N_5007,N_3069,N_2302);
nor U5008 (N_5008,N_2379,N_2503);
nand U5009 (N_5009,N_3220,N_2952);
and U5010 (N_5010,N_2676,N_3121);
or U5011 (N_5011,N_2360,N_3994);
nand U5012 (N_5012,N_2546,N_2684);
nor U5013 (N_5013,N_3913,N_2315);
and U5014 (N_5014,N_2510,N_2613);
nand U5015 (N_5015,N_2366,N_3458);
and U5016 (N_5016,N_3515,N_3402);
xor U5017 (N_5017,N_2770,N_2685);
and U5018 (N_5018,N_3082,N_2266);
or U5019 (N_5019,N_2618,N_3671);
nand U5020 (N_5020,N_2324,N_2432);
and U5021 (N_5021,N_2050,N_2332);
and U5022 (N_5022,N_2523,N_3544);
or U5023 (N_5023,N_2256,N_3965);
nand U5024 (N_5024,N_2418,N_3674);
nand U5025 (N_5025,N_2094,N_3731);
nand U5026 (N_5026,N_2085,N_3793);
nor U5027 (N_5027,N_2330,N_3361);
and U5028 (N_5028,N_2696,N_3326);
nand U5029 (N_5029,N_2307,N_2107);
xnor U5030 (N_5030,N_3961,N_3931);
nand U5031 (N_5031,N_2039,N_3428);
and U5032 (N_5032,N_2480,N_2935);
and U5033 (N_5033,N_3871,N_3626);
nor U5034 (N_5034,N_3249,N_2069);
and U5035 (N_5035,N_3804,N_2032);
or U5036 (N_5036,N_2079,N_2953);
or U5037 (N_5037,N_2399,N_3804);
or U5038 (N_5038,N_2605,N_2905);
nand U5039 (N_5039,N_2881,N_3359);
xnor U5040 (N_5040,N_2479,N_2833);
or U5041 (N_5041,N_3349,N_2554);
and U5042 (N_5042,N_2490,N_3736);
nand U5043 (N_5043,N_3621,N_3484);
nand U5044 (N_5044,N_2739,N_3077);
nor U5045 (N_5045,N_3999,N_2586);
nor U5046 (N_5046,N_3790,N_2718);
nor U5047 (N_5047,N_3910,N_2613);
or U5048 (N_5048,N_3225,N_2190);
nor U5049 (N_5049,N_2326,N_2524);
nand U5050 (N_5050,N_2489,N_3523);
or U5051 (N_5051,N_2174,N_3411);
or U5052 (N_5052,N_3173,N_3038);
xnor U5053 (N_5053,N_3126,N_2720);
nor U5054 (N_5054,N_2848,N_2603);
nor U5055 (N_5055,N_3015,N_2595);
or U5056 (N_5056,N_3073,N_2813);
nor U5057 (N_5057,N_2365,N_3126);
xnor U5058 (N_5058,N_2278,N_2355);
xor U5059 (N_5059,N_3609,N_3820);
nand U5060 (N_5060,N_2972,N_2833);
nor U5061 (N_5061,N_2120,N_2894);
and U5062 (N_5062,N_3264,N_2269);
nand U5063 (N_5063,N_2900,N_2018);
and U5064 (N_5064,N_3505,N_3558);
or U5065 (N_5065,N_2569,N_2274);
or U5066 (N_5066,N_2146,N_2944);
nor U5067 (N_5067,N_3800,N_3680);
and U5068 (N_5068,N_2543,N_2256);
or U5069 (N_5069,N_2837,N_3088);
or U5070 (N_5070,N_3584,N_3804);
nand U5071 (N_5071,N_3173,N_2066);
nand U5072 (N_5072,N_3377,N_3896);
or U5073 (N_5073,N_3108,N_3467);
or U5074 (N_5074,N_3328,N_2664);
and U5075 (N_5075,N_3729,N_3774);
nand U5076 (N_5076,N_2379,N_3709);
and U5077 (N_5077,N_3727,N_3773);
or U5078 (N_5078,N_3743,N_3541);
nor U5079 (N_5079,N_2129,N_2053);
nor U5080 (N_5080,N_2663,N_2375);
nand U5081 (N_5081,N_3079,N_2526);
xnor U5082 (N_5082,N_2239,N_3832);
nand U5083 (N_5083,N_3759,N_2411);
nand U5084 (N_5084,N_3174,N_2012);
nor U5085 (N_5085,N_2275,N_3754);
and U5086 (N_5086,N_2154,N_2709);
nor U5087 (N_5087,N_3046,N_3121);
and U5088 (N_5088,N_2184,N_3749);
and U5089 (N_5089,N_2733,N_2644);
and U5090 (N_5090,N_3819,N_2066);
nor U5091 (N_5091,N_3658,N_2451);
and U5092 (N_5092,N_3836,N_3714);
or U5093 (N_5093,N_2981,N_3486);
or U5094 (N_5094,N_2089,N_2621);
nand U5095 (N_5095,N_2389,N_3547);
or U5096 (N_5096,N_3885,N_3206);
xor U5097 (N_5097,N_3448,N_2669);
nor U5098 (N_5098,N_3135,N_2799);
and U5099 (N_5099,N_3197,N_2462);
nor U5100 (N_5100,N_2209,N_3232);
and U5101 (N_5101,N_2692,N_2372);
and U5102 (N_5102,N_3286,N_2963);
nor U5103 (N_5103,N_2805,N_3710);
nor U5104 (N_5104,N_3074,N_2989);
nor U5105 (N_5105,N_2138,N_3384);
xor U5106 (N_5106,N_2270,N_2645);
or U5107 (N_5107,N_2501,N_2664);
xor U5108 (N_5108,N_2424,N_2018);
or U5109 (N_5109,N_2655,N_2087);
nand U5110 (N_5110,N_3458,N_3120);
or U5111 (N_5111,N_2853,N_2891);
nand U5112 (N_5112,N_3410,N_3159);
or U5113 (N_5113,N_3696,N_2921);
nand U5114 (N_5114,N_3749,N_2224);
and U5115 (N_5115,N_3113,N_2946);
nand U5116 (N_5116,N_2657,N_3941);
nand U5117 (N_5117,N_2686,N_3060);
and U5118 (N_5118,N_2200,N_3303);
or U5119 (N_5119,N_2173,N_2781);
xor U5120 (N_5120,N_2058,N_3951);
or U5121 (N_5121,N_2445,N_3065);
and U5122 (N_5122,N_2833,N_3660);
and U5123 (N_5123,N_2590,N_3966);
xnor U5124 (N_5124,N_3722,N_3592);
nor U5125 (N_5125,N_3805,N_3774);
nand U5126 (N_5126,N_3453,N_3687);
nand U5127 (N_5127,N_3917,N_3474);
nand U5128 (N_5128,N_3990,N_3606);
nand U5129 (N_5129,N_3166,N_2601);
or U5130 (N_5130,N_2160,N_2817);
nand U5131 (N_5131,N_2296,N_2891);
or U5132 (N_5132,N_3649,N_3740);
or U5133 (N_5133,N_3090,N_3875);
nand U5134 (N_5134,N_2661,N_2015);
nor U5135 (N_5135,N_3897,N_3662);
or U5136 (N_5136,N_2528,N_2064);
and U5137 (N_5137,N_3719,N_2975);
nand U5138 (N_5138,N_2044,N_3772);
and U5139 (N_5139,N_3951,N_2111);
nand U5140 (N_5140,N_2563,N_2526);
and U5141 (N_5141,N_3579,N_2915);
or U5142 (N_5142,N_2716,N_2189);
nor U5143 (N_5143,N_3173,N_3399);
nor U5144 (N_5144,N_3051,N_2035);
and U5145 (N_5145,N_2140,N_3219);
nand U5146 (N_5146,N_3699,N_2578);
nand U5147 (N_5147,N_2677,N_3405);
and U5148 (N_5148,N_2656,N_3882);
nor U5149 (N_5149,N_2034,N_3621);
or U5150 (N_5150,N_2093,N_3144);
nand U5151 (N_5151,N_3078,N_3547);
or U5152 (N_5152,N_2950,N_2004);
or U5153 (N_5153,N_3210,N_2519);
xor U5154 (N_5154,N_2538,N_2218);
nand U5155 (N_5155,N_2833,N_2678);
nor U5156 (N_5156,N_2728,N_2896);
nor U5157 (N_5157,N_2950,N_2308);
nor U5158 (N_5158,N_3142,N_3607);
and U5159 (N_5159,N_3725,N_2538);
xor U5160 (N_5160,N_2843,N_3428);
xnor U5161 (N_5161,N_3170,N_2702);
nor U5162 (N_5162,N_2186,N_3914);
nand U5163 (N_5163,N_3632,N_2581);
nand U5164 (N_5164,N_2274,N_2008);
and U5165 (N_5165,N_3505,N_3967);
and U5166 (N_5166,N_2441,N_2538);
and U5167 (N_5167,N_3287,N_3610);
nand U5168 (N_5168,N_3213,N_3389);
nand U5169 (N_5169,N_2458,N_2762);
nand U5170 (N_5170,N_2277,N_2160);
nand U5171 (N_5171,N_3190,N_2605);
and U5172 (N_5172,N_2167,N_3022);
nand U5173 (N_5173,N_2597,N_2430);
nor U5174 (N_5174,N_2515,N_3127);
or U5175 (N_5175,N_3972,N_2724);
or U5176 (N_5176,N_2362,N_2829);
nand U5177 (N_5177,N_3075,N_3337);
or U5178 (N_5178,N_2406,N_3065);
nor U5179 (N_5179,N_3097,N_3847);
nand U5180 (N_5180,N_2631,N_3739);
nand U5181 (N_5181,N_3527,N_3505);
and U5182 (N_5182,N_3046,N_3875);
or U5183 (N_5183,N_2290,N_3003);
nor U5184 (N_5184,N_2662,N_3585);
nand U5185 (N_5185,N_3755,N_3345);
nand U5186 (N_5186,N_3454,N_2494);
or U5187 (N_5187,N_2881,N_2088);
nor U5188 (N_5188,N_2176,N_2041);
or U5189 (N_5189,N_3034,N_3649);
nand U5190 (N_5190,N_3395,N_2404);
and U5191 (N_5191,N_3791,N_2161);
xor U5192 (N_5192,N_3851,N_2434);
and U5193 (N_5193,N_2816,N_2320);
nor U5194 (N_5194,N_3610,N_3361);
nand U5195 (N_5195,N_3343,N_2542);
nand U5196 (N_5196,N_3588,N_3255);
and U5197 (N_5197,N_2960,N_2052);
and U5198 (N_5198,N_3798,N_2365);
nor U5199 (N_5199,N_3339,N_3861);
nand U5200 (N_5200,N_2747,N_3717);
nor U5201 (N_5201,N_2187,N_3361);
xnor U5202 (N_5202,N_2614,N_3770);
nor U5203 (N_5203,N_3655,N_3400);
or U5204 (N_5204,N_3703,N_3477);
nor U5205 (N_5205,N_3966,N_2982);
nand U5206 (N_5206,N_2926,N_2238);
or U5207 (N_5207,N_3381,N_3736);
xnor U5208 (N_5208,N_2680,N_3636);
and U5209 (N_5209,N_2037,N_2154);
and U5210 (N_5210,N_2566,N_3594);
nand U5211 (N_5211,N_2679,N_3213);
and U5212 (N_5212,N_3755,N_3779);
nand U5213 (N_5213,N_3173,N_3773);
or U5214 (N_5214,N_2930,N_3774);
or U5215 (N_5215,N_2955,N_2011);
or U5216 (N_5216,N_2900,N_3319);
or U5217 (N_5217,N_3329,N_2734);
nor U5218 (N_5218,N_3114,N_3169);
nand U5219 (N_5219,N_3794,N_3971);
or U5220 (N_5220,N_2402,N_3325);
or U5221 (N_5221,N_3817,N_3052);
and U5222 (N_5222,N_3009,N_2532);
or U5223 (N_5223,N_3585,N_2958);
nor U5224 (N_5224,N_2800,N_2206);
and U5225 (N_5225,N_2458,N_3446);
nor U5226 (N_5226,N_2233,N_3573);
or U5227 (N_5227,N_2315,N_2053);
nor U5228 (N_5228,N_3149,N_3967);
and U5229 (N_5229,N_3095,N_3740);
or U5230 (N_5230,N_3889,N_3604);
xnor U5231 (N_5231,N_2920,N_3567);
xnor U5232 (N_5232,N_2312,N_2215);
nand U5233 (N_5233,N_3905,N_3219);
nand U5234 (N_5234,N_2969,N_2778);
or U5235 (N_5235,N_3010,N_3872);
or U5236 (N_5236,N_3886,N_2386);
and U5237 (N_5237,N_2297,N_3594);
or U5238 (N_5238,N_2769,N_2660);
nand U5239 (N_5239,N_3963,N_2147);
or U5240 (N_5240,N_2001,N_2936);
nor U5241 (N_5241,N_2327,N_3325);
and U5242 (N_5242,N_3738,N_3244);
and U5243 (N_5243,N_2403,N_3765);
or U5244 (N_5244,N_3378,N_2207);
xor U5245 (N_5245,N_3197,N_2907);
nand U5246 (N_5246,N_2245,N_3794);
nand U5247 (N_5247,N_2665,N_2946);
xor U5248 (N_5248,N_3916,N_2276);
nand U5249 (N_5249,N_3149,N_2104);
nor U5250 (N_5250,N_3542,N_3663);
nor U5251 (N_5251,N_2365,N_3746);
nor U5252 (N_5252,N_2255,N_3295);
nand U5253 (N_5253,N_3916,N_2820);
and U5254 (N_5254,N_3499,N_2053);
nor U5255 (N_5255,N_3029,N_2592);
nor U5256 (N_5256,N_2195,N_3564);
or U5257 (N_5257,N_2131,N_2239);
xnor U5258 (N_5258,N_3161,N_2959);
nor U5259 (N_5259,N_3431,N_2139);
or U5260 (N_5260,N_3335,N_3458);
nor U5261 (N_5261,N_2548,N_3056);
or U5262 (N_5262,N_3819,N_3296);
nand U5263 (N_5263,N_2477,N_2009);
nand U5264 (N_5264,N_2825,N_2042);
nor U5265 (N_5265,N_3693,N_3332);
nand U5266 (N_5266,N_2621,N_2942);
and U5267 (N_5267,N_2519,N_2932);
and U5268 (N_5268,N_2816,N_2298);
and U5269 (N_5269,N_3133,N_3138);
and U5270 (N_5270,N_3559,N_2517);
nand U5271 (N_5271,N_3340,N_2021);
and U5272 (N_5272,N_3383,N_2875);
nor U5273 (N_5273,N_3428,N_3814);
nor U5274 (N_5274,N_2850,N_2041);
nand U5275 (N_5275,N_2201,N_3422);
nand U5276 (N_5276,N_2481,N_3783);
and U5277 (N_5277,N_3296,N_2610);
or U5278 (N_5278,N_2469,N_3906);
or U5279 (N_5279,N_3460,N_3025);
nand U5280 (N_5280,N_3254,N_3979);
nor U5281 (N_5281,N_2545,N_2659);
or U5282 (N_5282,N_2663,N_3844);
and U5283 (N_5283,N_2713,N_2076);
or U5284 (N_5284,N_3822,N_3702);
nor U5285 (N_5285,N_3585,N_3215);
and U5286 (N_5286,N_3498,N_3131);
or U5287 (N_5287,N_3406,N_2334);
nor U5288 (N_5288,N_3204,N_3745);
nor U5289 (N_5289,N_2892,N_3598);
or U5290 (N_5290,N_2476,N_3150);
nand U5291 (N_5291,N_2934,N_2868);
and U5292 (N_5292,N_3949,N_3229);
or U5293 (N_5293,N_2252,N_3610);
xnor U5294 (N_5294,N_2039,N_3507);
nor U5295 (N_5295,N_2671,N_3405);
or U5296 (N_5296,N_3755,N_2271);
and U5297 (N_5297,N_2209,N_3495);
xor U5298 (N_5298,N_2494,N_2936);
nand U5299 (N_5299,N_2517,N_2633);
and U5300 (N_5300,N_3877,N_2468);
and U5301 (N_5301,N_2160,N_3121);
nand U5302 (N_5302,N_2594,N_3816);
and U5303 (N_5303,N_2094,N_3319);
nand U5304 (N_5304,N_3481,N_3367);
and U5305 (N_5305,N_2610,N_3970);
xnor U5306 (N_5306,N_2668,N_3781);
or U5307 (N_5307,N_2390,N_3116);
and U5308 (N_5308,N_3252,N_3840);
nor U5309 (N_5309,N_3025,N_2754);
nor U5310 (N_5310,N_2506,N_3637);
and U5311 (N_5311,N_2075,N_2130);
nor U5312 (N_5312,N_3210,N_3337);
or U5313 (N_5313,N_2518,N_2796);
xor U5314 (N_5314,N_2450,N_2140);
nand U5315 (N_5315,N_2260,N_2361);
and U5316 (N_5316,N_2922,N_3767);
and U5317 (N_5317,N_2784,N_2353);
or U5318 (N_5318,N_2793,N_3303);
or U5319 (N_5319,N_2809,N_2334);
and U5320 (N_5320,N_3935,N_3715);
and U5321 (N_5321,N_2810,N_2061);
nand U5322 (N_5322,N_2899,N_2970);
xnor U5323 (N_5323,N_3902,N_3849);
or U5324 (N_5324,N_3140,N_3460);
nand U5325 (N_5325,N_2904,N_3235);
or U5326 (N_5326,N_3111,N_3608);
or U5327 (N_5327,N_3117,N_3254);
or U5328 (N_5328,N_2023,N_2459);
nand U5329 (N_5329,N_2046,N_2391);
and U5330 (N_5330,N_3016,N_2333);
xnor U5331 (N_5331,N_3254,N_3236);
or U5332 (N_5332,N_2617,N_3181);
or U5333 (N_5333,N_2500,N_3911);
or U5334 (N_5334,N_2429,N_3303);
and U5335 (N_5335,N_3367,N_3033);
nor U5336 (N_5336,N_2576,N_3628);
xor U5337 (N_5337,N_2462,N_2613);
nor U5338 (N_5338,N_3935,N_2643);
or U5339 (N_5339,N_3512,N_3785);
and U5340 (N_5340,N_3471,N_3107);
nand U5341 (N_5341,N_2528,N_3297);
nand U5342 (N_5342,N_2441,N_3828);
nor U5343 (N_5343,N_3449,N_2810);
nand U5344 (N_5344,N_3101,N_2922);
or U5345 (N_5345,N_2899,N_2647);
or U5346 (N_5346,N_3370,N_2437);
xnor U5347 (N_5347,N_2684,N_2089);
xor U5348 (N_5348,N_3238,N_2854);
or U5349 (N_5349,N_2909,N_2317);
and U5350 (N_5350,N_3306,N_3426);
xnor U5351 (N_5351,N_3749,N_2297);
or U5352 (N_5352,N_3961,N_2853);
nand U5353 (N_5353,N_3969,N_2240);
and U5354 (N_5354,N_3716,N_2016);
and U5355 (N_5355,N_3728,N_2640);
nand U5356 (N_5356,N_2190,N_2012);
nor U5357 (N_5357,N_2237,N_2984);
nor U5358 (N_5358,N_2904,N_3943);
or U5359 (N_5359,N_2811,N_3432);
or U5360 (N_5360,N_3157,N_2603);
nand U5361 (N_5361,N_3209,N_2421);
nand U5362 (N_5362,N_3112,N_3113);
nor U5363 (N_5363,N_2625,N_3525);
xor U5364 (N_5364,N_3548,N_3310);
or U5365 (N_5365,N_3963,N_3340);
nand U5366 (N_5366,N_3173,N_3604);
or U5367 (N_5367,N_2478,N_2138);
xor U5368 (N_5368,N_2074,N_2914);
and U5369 (N_5369,N_2223,N_2808);
and U5370 (N_5370,N_2004,N_3772);
nor U5371 (N_5371,N_2209,N_3150);
and U5372 (N_5372,N_2403,N_3463);
nor U5373 (N_5373,N_2945,N_2481);
nand U5374 (N_5374,N_2208,N_2862);
xnor U5375 (N_5375,N_3936,N_3952);
and U5376 (N_5376,N_3264,N_3543);
nand U5377 (N_5377,N_2104,N_2496);
and U5378 (N_5378,N_2567,N_2712);
xor U5379 (N_5379,N_2460,N_2346);
nand U5380 (N_5380,N_3488,N_2502);
nor U5381 (N_5381,N_2366,N_3959);
nor U5382 (N_5382,N_2772,N_3972);
and U5383 (N_5383,N_3701,N_3919);
and U5384 (N_5384,N_3796,N_3784);
and U5385 (N_5385,N_2174,N_2324);
or U5386 (N_5386,N_3377,N_3671);
nand U5387 (N_5387,N_2288,N_2485);
nor U5388 (N_5388,N_3769,N_2479);
and U5389 (N_5389,N_2686,N_3282);
or U5390 (N_5390,N_2985,N_2460);
or U5391 (N_5391,N_3124,N_3943);
and U5392 (N_5392,N_2015,N_3668);
nand U5393 (N_5393,N_2343,N_3782);
xnor U5394 (N_5394,N_2527,N_3245);
nand U5395 (N_5395,N_3450,N_3927);
or U5396 (N_5396,N_3111,N_3009);
and U5397 (N_5397,N_2437,N_3836);
nor U5398 (N_5398,N_2498,N_3300);
and U5399 (N_5399,N_2976,N_3938);
and U5400 (N_5400,N_2037,N_3176);
xnor U5401 (N_5401,N_2721,N_3048);
nor U5402 (N_5402,N_3935,N_3218);
and U5403 (N_5403,N_2631,N_3510);
or U5404 (N_5404,N_3068,N_2444);
nor U5405 (N_5405,N_2751,N_2912);
or U5406 (N_5406,N_3647,N_2482);
nand U5407 (N_5407,N_3171,N_2583);
and U5408 (N_5408,N_2366,N_2064);
xnor U5409 (N_5409,N_3273,N_3354);
or U5410 (N_5410,N_2141,N_2502);
nor U5411 (N_5411,N_2239,N_2293);
or U5412 (N_5412,N_3305,N_2938);
and U5413 (N_5413,N_3391,N_3891);
or U5414 (N_5414,N_2703,N_2662);
xor U5415 (N_5415,N_2574,N_2432);
nor U5416 (N_5416,N_2024,N_3067);
or U5417 (N_5417,N_3230,N_2663);
or U5418 (N_5418,N_3865,N_2652);
or U5419 (N_5419,N_2512,N_3390);
nand U5420 (N_5420,N_2183,N_2375);
xnor U5421 (N_5421,N_2308,N_3583);
and U5422 (N_5422,N_3616,N_2430);
nor U5423 (N_5423,N_3594,N_3293);
or U5424 (N_5424,N_3173,N_3897);
nor U5425 (N_5425,N_2895,N_2517);
or U5426 (N_5426,N_3190,N_3106);
or U5427 (N_5427,N_2139,N_2930);
or U5428 (N_5428,N_2079,N_2954);
nor U5429 (N_5429,N_2171,N_3731);
nand U5430 (N_5430,N_3765,N_2188);
xor U5431 (N_5431,N_3822,N_3845);
and U5432 (N_5432,N_2170,N_3826);
and U5433 (N_5433,N_3613,N_3885);
nor U5434 (N_5434,N_3477,N_2367);
and U5435 (N_5435,N_3102,N_3899);
nor U5436 (N_5436,N_2321,N_2497);
or U5437 (N_5437,N_2001,N_3524);
and U5438 (N_5438,N_2305,N_3376);
xnor U5439 (N_5439,N_3029,N_3622);
xnor U5440 (N_5440,N_3984,N_2837);
nand U5441 (N_5441,N_3188,N_3391);
nor U5442 (N_5442,N_2299,N_2561);
nand U5443 (N_5443,N_3941,N_3181);
nand U5444 (N_5444,N_2782,N_2359);
nand U5445 (N_5445,N_2690,N_2520);
and U5446 (N_5446,N_2529,N_2676);
or U5447 (N_5447,N_2243,N_2132);
xor U5448 (N_5448,N_2327,N_2403);
nor U5449 (N_5449,N_2713,N_3517);
nor U5450 (N_5450,N_3652,N_3356);
nor U5451 (N_5451,N_3700,N_3304);
or U5452 (N_5452,N_3216,N_2009);
or U5453 (N_5453,N_2538,N_2213);
nand U5454 (N_5454,N_3890,N_3645);
nor U5455 (N_5455,N_2159,N_3593);
or U5456 (N_5456,N_3941,N_3657);
or U5457 (N_5457,N_3645,N_3338);
and U5458 (N_5458,N_3240,N_3231);
or U5459 (N_5459,N_3972,N_3458);
or U5460 (N_5460,N_2204,N_2696);
nand U5461 (N_5461,N_3310,N_3307);
or U5462 (N_5462,N_2688,N_3649);
nand U5463 (N_5463,N_3843,N_3036);
nand U5464 (N_5464,N_2755,N_3969);
and U5465 (N_5465,N_2171,N_2163);
or U5466 (N_5466,N_3727,N_2237);
xor U5467 (N_5467,N_3041,N_2034);
and U5468 (N_5468,N_2174,N_3527);
nand U5469 (N_5469,N_3842,N_2770);
nand U5470 (N_5470,N_3684,N_2128);
nand U5471 (N_5471,N_2434,N_2210);
nand U5472 (N_5472,N_2013,N_2651);
xnor U5473 (N_5473,N_2123,N_3084);
nor U5474 (N_5474,N_3340,N_2325);
or U5475 (N_5475,N_3276,N_3863);
nor U5476 (N_5476,N_3464,N_3242);
nand U5477 (N_5477,N_2823,N_2694);
and U5478 (N_5478,N_2359,N_2447);
nand U5479 (N_5479,N_3924,N_3786);
or U5480 (N_5480,N_3351,N_2544);
and U5481 (N_5481,N_3560,N_2597);
nand U5482 (N_5482,N_2655,N_3640);
nand U5483 (N_5483,N_2585,N_3370);
nor U5484 (N_5484,N_2916,N_2279);
or U5485 (N_5485,N_3691,N_3031);
nand U5486 (N_5486,N_3547,N_3518);
and U5487 (N_5487,N_2791,N_2831);
xor U5488 (N_5488,N_2854,N_3571);
xnor U5489 (N_5489,N_2991,N_3991);
and U5490 (N_5490,N_3765,N_2595);
and U5491 (N_5491,N_2645,N_2237);
or U5492 (N_5492,N_3167,N_2604);
nand U5493 (N_5493,N_3400,N_2245);
and U5494 (N_5494,N_2952,N_2874);
xor U5495 (N_5495,N_2290,N_3324);
and U5496 (N_5496,N_3952,N_2694);
nor U5497 (N_5497,N_3851,N_2026);
xnor U5498 (N_5498,N_3659,N_2995);
nor U5499 (N_5499,N_2637,N_3684);
xnor U5500 (N_5500,N_2681,N_3846);
and U5501 (N_5501,N_3805,N_2712);
nor U5502 (N_5502,N_2626,N_3245);
nand U5503 (N_5503,N_3543,N_2970);
nand U5504 (N_5504,N_2138,N_3365);
nand U5505 (N_5505,N_3172,N_3619);
nand U5506 (N_5506,N_3507,N_2056);
or U5507 (N_5507,N_3281,N_2995);
and U5508 (N_5508,N_2651,N_2625);
nor U5509 (N_5509,N_3785,N_2776);
and U5510 (N_5510,N_2401,N_2175);
nor U5511 (N_5511,N_3094,N_3126);
nor U5512 (N_5512,N_2002,N_2601);
and U5513 (N_5513,N_2566,N_3599);
nand U5514 (N_5514,N_3569,N_2860);
nor U5515 (N_5515,N_3098,N_2758);
or U5516 (N_5516,N_2699,N_3655);
nor U5517 (N_5517,N_3011,N_3916);
or U5518 (N_5518,N_2480,N_2120);
or U5519 (N_5519,N_2099,N_3811);
and U5520 (N_5520,N_3493,N_3470);
nor U5521 (N_5521,N_2780,N_3248);
or U5522 (N_5522,N_2455,N_3523);
nor U5523 (N_5523,N_2186,N_3580);
and U5524 (N_5524,N_2769,N_2389);
and U5525 (N_5525,N_2626,N_3265);
or U5526 (N_5526,N_2442,N_2787);
nor U5527 (N_5527,N_3521,N_2414);
and U5528 (N_5528,N_2797,N_3350);
and U5529 (N_5529,N_3903,N_2944);
nor U5530 (N_5530,N_2841,N_2884);
or U5531 (N_5531,N_2661,N_3375);
or U5532 (N_5532,N_3839,N_2333);
nor U5533 (N_5533,N_2879,N_2100);
and U5534 (N_5534,N_2173,N_2552);
nand U5535 (N_5535,N_3716,N_3599);
or U5536 (N_5536,N_2757,N_3144);
and U5537 (N_5537,N_3474,N_3985);
or U5538 (N_5538,N_2079,N_2442);
nor U5539 (N_5539,N_3508,N_3120);
xor U5540 (N_5540,N_2065,N_2438);
nor U5541 (N_5541,N_2255,N_3457);
and U5542 (N_5542,N_3403,N_2121);
nor U5543 (N_5543,N_2014,N_2538);
or U5544 (N_5544,N_2166,N_3527);
nand U5545 (N_5545,N_2428,N_3289);
nand U5546 (N_5546,N_3937,N_2748);
nor U5547 (N_5547,N_2491,N_2444);
or U5548 (N_5548,N_2747,N_2517);
nor U5549 (N_5549,N_3724,N_3606);
nand U5550 (N_5550,N_3725,N_2268);
and U5551 (N_5551,N_3124,N_3129);
nand U5552 (N_5552,N_3260,N_2187);
nor U5553 (N_5553,N_3497,N_3089);
or U5554 (N_5554,N_2220,N_2050);
xor U5555 (N_5555,N_2849,N_2572);
or U5556 (N_5556,N_3684,N_3529);
and U5557 (N_5557,N_3603,N_3895);
or U5558 (N_5558,N_3887,N_3481);
nor U5559 (N_5559,N_2686,N_3558);
nand U5560 (N_5560,N_2618,N_3764);
nand U5561 (N_5561,N_2086,N_3198);
nor U5562 (N_5562,N_3024,N_2761);
xor U5563 (N_5563,N_2976,N_3998);
xor U5564 (N_5564,N_3303,N_2034);
nand U5565 (N_5565,N_3381,N_3497);
and U5566 (N_5566,N_2328,N_2522);
or U5567 (N_5567,N_2512,N_3596);
nor U5568 (N_5568,N_2375,N_3144);
nor U5569 (N_5569,N_3725,N_3410);
and U5570 (N_5570,N_2825,N_3203);
nand U5571 (N_5571,N_2941,N_2917);
nor U5572 (N_5572,N_3863,N_2025);
or U5573 (N_5573,N_3629,N_3051);
nand U5574 (N_5574,N_2437,N_2061);
nor U5575 (N_5575,N_3571,N_2881);
and U5576 (N_5576,N_2525,N_3622);
and U5577 (N_5577,N_2154,N_2603);
xnor U5578 (N_5578,N_3432,N_3791);
or U5579 (N_5579,N_2948,N_3864);
xor U5580 (N_5580,N_3873,N_3243);
nand U5581 (N_5581,N_3403,N_2777);
or U5582 (N_5582,N_3698,N_2603);
nand U5583 (N_5583,N_3903,N_2495);
nand U5584 (N_5584,N_3858,N_2759);
or U5585 (N_5585,N_2985,N_2098);
or U5586 (N_5586,N_3637,N_3936);
and U5587 (N_5587,N_2077,N_3751);
nand U5588 (N_5588,N_3555,N_2416);
nand U5589 (N_5589,N_3371,N_3709);
nor U5590 (N_5590,N_3235,N_3667);
nand U5591 (N_5591,N_2541,N_2536);
and U5592 (N_5592,N_2014,N_2551);
nor U5593 (N_5593,N_2592,N_3086);
nor U5594 (N_5594,N_3754,N_2890);
or U5595 (N_5595,N_3553,N_2839);
nand U5596 (N_5596,N_2863,N_2261);
nor U5597 (N_5597,N_2071,N_3127);
nor U5598 (N_5598,N_2998,N_3434);
nand U5599 (N_5599,N_2763,N_2382);
nor U5600 (N_5600,N_3045,N_3640);
or U5601 (N_5601,N_3745,N_3805);
and U5602 (N_5602,N_3333,N_3175);
nor U5603 (N_5603,N_3982,N_3068);
nand U5604 (N_5604,N_2090,N_3356);
or U5605 (N_5605,N_2308,N_2600);
xor U5606 (N_5606,N_3747,N_3801);
nand U5607 (N_5607,N_3485,N_3878);
nor U5608 (N_5608,N_3363,N_3853);
and U5609 (N_5609,N_2629,N_3594);
and U5610 (N_5610,N_3044,N_3685);
nor U5611 (N_5611,N_2359,N_3654);
or U5612 (N_5612,N_3061,N_2451);
and U5613 (N_5613,N_3999,N_2142);
xor U5614 (N_5614,N_3626,N_2402);
and U5615 (N_5615,N_3238,N_3175);
or U5616 (N_5616,N_3044,N_3882);
nand U5617 (N_5617,N_2673,N_2465);
and U5618 (N_5618,N_2959,N_2280);
nor U5619 (N_5619,N_3535,N_2196);
nor U5620 (N_5620,N_3946,N_3552);
and U5621 (N_5621,N_2230,N_3023);
or U5622 (N_5622,N_2197,N_2390);
and U5623 (N_5623,N_2561,N_2765);
nor U5624 (N_5624,N_2087,N_2737);
nor U5625 (N_5625,N_2499,N_3288);
or U5626 (N_5626,N_2535,N_3471);
or U5627 (N_5627,N_2235,N_3387);
nor U5628 (N_5628,N_2664,N_2818);
nor U5629 (N_5629,N_3572,N_3031);
and U5630 (N_5630,N_2574,N_3495);
or U5631 (N_5631,N_2450,N_2732);
and U5632 (N_5632,N_3975,N_2034);
nor U5633 (N_5633,N_3239,N_3031);
and U5634 (N_5634,N_3181,N_2598);
or U5635 (N_5635,N_2123,N_2853);
xor U5636 (N_5636,N_2781,N_3419);
nor U5637 (N_5637,N_2116,N_3114);
and U5638 (N_5638,N_3018,N_2481);
nand U5639 (N_5639,N_2729,N_2251);
xor U5640 (N_5640,N_2205,N_2061);
nand U5641 (N_5641,N_3297,N_2064);
and U5642 (N_5642,N_3512,N_3100);
xor U5643 (N_5643,N_2867,N_2006);
nor U5644 (N_5644,N_3707,N_2586);
xnor U5645 (N_5645,N_3659,N_2391);
nand U5646 (N_5646,N_3634,N_2945);
and U5647 (N_5647,N_3232,N_3623);
or U5648 (N_5648,N_2921,N_3753);
or U5649 (N_5649,N_3264,N_2942);
nand U5650 (N_5650,N_2388,N_2409);
xor U5651 (N_5651,N_2960,N_2971);
or U5652 (N_5652,N_2719,N_3135);
or U5653 (N_5653,N_3755,N_2839);
nand U5654 (N_5654,N_2057,N_2132);
nor U5655 (N_5655,N_3484,N_2824);
or U5656 (N_5656,N_2254,N_2890);
nand U5657 (N_5657,N_3221,N_2348);
and U5658 (N_5658,N_3134,N_3473);
xor U5659 (N_5659,N_3787,N_2619);
xor U5660 (N_5660,N_3297,N_3326);
nand U5661 (N_5661,N_3880,N_3233);
or U5662 (N_5662,N_3049,N_3316);
nor U5663 (N_5663,N_3493,N_2619);
xor U5664 (N_5664,N_2269,N_2745);
and U5665 (N_5665,N_2998,N_3873);
nor U5666 (N_5666,N_3744,N_2061);
and U5667 (N_5667,N_3989,N_3911);
and U5668 (N_5668,N_2958,N_2016);
or U5669 (N_5669,N_2213,N_2444);
and U5670 (N_5670,N_2721,N_2383);
xor U5671 (N_5671,N_3958,N_3927);
and U5672 (N_5672,N_2991,N_3270);
or U5673 (N_5673,N_2922,N_2340);
xor U5674 (N_5674,N_3274,N_3934);
and U5675 (N_5675,N_2762,N_2454);
xor U5676 (N_5676,N_2312,N_2421);
nand U5677 (N_5677,N_3321,N_3550);
or U5678 (N_5678,N_2401,N_3374);
xnor U5679 (N_5679,N_2495,N_3053);
and U5680 (N_5680,N_2448,N_3868);
or U5681 (N_5681,N_2659,N_2157);
and U5682 (N_5682,N_3662,N_2124);
nand U5683 (N_5683,N_3130,N_2370);
nand U5684 (N_5684,N_3319,N_2279);
or U5685 (N_5685,N_2377,N_3458);
nand U5686 (N_5686,N_2466,N_2958);
nor U5687 (N_5687,N_3783,N_2973);
xnor U5688 (N_5688,N_2603,N_2020);
nand U5689 (N_5689,N_3473,N_3147);
and U5690 (N_5690,N_3504,N_2145);
and U5691 (N_5691,N_2463,N_3021);
nand U5692 (N_5692,N_3393,N_2435);
xnor U5693 (N_5693,N_2520,N_3839);
or U5694 (N_5694,N_2167,N_2388);
or U5695 (N_5695,N_2134,N_3432);
nor U5696 (N_5696,N_3955,N_3287);
and U5697 (N_5697,N_2948,N_2709);
nor U5698 (N_5698,N_3786,N_3411);
xnor U5699 (N_5699,N_2902,N_3919);
nand U5700 (N_5700,N_2260,N_3293);
and U5701 (N_5701,N_2414,N_3035);
nand U5702 (N_5702,N_2584,N_2652);
nor U5703 (N_5703,N_2395,N_2663);
nand U5704 (N_5704,N_3222,N_3494);
and U5705 (N_5705,N_2035,N_3954);
or U5706 (N_5706,N_2567,N_3389);
nor U5707 (N_5707,N_3153,N_3817);
or U5708 (N_5708,N_2403,N_2834);
or U5709 (N_5709,N_3438,N_2815);
xnor U5710 (N_5710,N_2559,N_2637);
and U5711 (N_5711,N_3869,N_3125);
and U5712 (N_5712,N_2935,N_3257);
nand U5713 (N_5713,N_3161,N_2136);
nand U5714 (N_5714,N_3815,N_2626);
xnor U5715 (N_5715,N_2369,N_3292);
or U5716 (N_5716,N_2116,N_3472);
xor U5717 (N_5717,N_3673,N_3890);
and U5718 (N_5718,N_2299,N_2490);
nor U5719 (N_5719,N_2587,N_3421);
and U5720 (N_5720,N_3025,N_3492);
or U5721 (N_5721,N_2529,N_2089);
and U5722 (N_5722,N_3695,N_2627);
nor U5723 (N_5723,N_2897,N_3588);
nand U5724 (N_5724,N_3035,N_3902);
nand U5725 (N_5725,N_2956,N_2005);
or U5726 (N_5726,N_2002,N_3734);
nor U5727 (N_5727,N_2286,N_2864);
nand U5728 (N_5728,N_3045,N_3603);
or U5729 (N_5729,N_2590,N_2330);
nor U5730 (N_5730,N_3006,N_2466);
nor U5731 (N_5731,N_2250,N_3195);
and U5732 (N_5732,N_3183,N_3674);
nand U5733 (N_5733,N_3738,N_2834);
xnor U5734 (N_5734,N_2702,N_3799);
nor U5735 (N_5735,N_3099,N_3741);
nand U5736 (N_5736,N_2958,N_2743);
or U5737 (N_5737,N_2110,N_3385);
xnor U5738 (N_5738,N_2494,N_3282);
xor U5739 (N_5739,N_3844,N_2364);
xor U5740 (N_5740,N_3611,N_3116);
or U5741 (N_5741,N_2874,N_2479);
nor U5742 (N_5742,N_2581,N_2155);
nand U5743 (N_5743,N_2244,N_2092);
and U5744 (N_5744,N_2615,N_3709);
and U5745 (N_5745,N_3028,N_2614);
nand U5746 (N_5746,N_3195,N_3772);
nand U5747 (N_5747,N_2712,N_3102);
and U5748 (N_5748,N_3153,N_2799);
or U5749 (N_5749,N_2363,N_2743);
xor U5750 (N_5750,N_3472,N_2653);
nor U5751 (N_5751,N_3682,N_3065);
nand U5752 (N_5752,N_2717,N_3154);
nand U5753 (N_5753,N_2246,N_2302);
and U5754 (N_5754,N_3129,N_2782);
xor U5755 (N_5755,N_2325,N_3865);
or U5756 (N_5756,N_2132,N_3614);
nand U5757 (N_5757,N_3246,N_3371);
xor U5758 (N_5758,N_3452,N_3307);
nor U5759 (N_5759,N_2265,N_3430);
nor U5760 (N_5760,N_2951,N_2602);
nor U5761 (N_5761,N_3209,N_3321);
nand U5762 (N_5762,N_2166,N_2888);
nor U5763 (N_5763,N_2398,N_3601);
and U5764 (N_5764,N_2537,N_3863);
or U5765 (N_5765,N_2868,N_3795);
or U5766 (N_5766,N_3715,N_3592);
xnor U5767 (N_5767,N_3071,N_2007);
and U5768 (N_5768,N_2618,N_3597);
and U5769 (N_5769,N_2065,N_2263);
nand U5770 (N_5770,N_2319,N_2619);
nor U5771 (N_5771,N_2732,N_3564);
and U5772 (N_5772,N_2912,N_2786);
nor U5773 (N_5773,N_2727,N_3151);
and U5774 (N_5774,N_2792,N_2623);
nand U5775 (N_5775,N_2531,N_2441);
nor U5776 (N_5776,N_2848,N_3538);
or U5777 (N_5777,N_3177,N_3804);
or U5778 (N_5778,N_2490,N_2733);
and U5779 (N_5779,N_3965,N_3212);
and U5780 (N_5780,N_3190,N_2336);
and U5781 (N_5781,N_2127,N_2566);
nor U5782 (N_5782,N_2961,N_2052);
xor U5783 (N_5783,N_3634,N_2168);
xor U5784 (N_5784,N_2375,N_2256);
and U5785 (N_5785,N_2637,N_3117);
or U5786 (N_5786,N_3497,N_3191);
nor U5787 (N_5787,N_2147,N_2969);
nor U5788 (N_5788,N_2253,N_2891);
or U5789 (N_5789,N_3656,N_2786);
nor U5790 (N_5790,N_3969,N_3473);
xnor U5791 (N_5791,N_3837,N_2662);
nand U5792 (N_5792,N_2881,N_3765);
nor U5793 (N_5793,N_2375,N_2760);
or U5794 (N_5794,N_2565,N_3724);
nor U5795 (N_5795,N_3700,N_2096);
and U5796 (N_5796,N_3654,N_3192);
and U5797 (N_5797,N_2308,N_2655);
xor U5798 (N_5798,N_3026,N_2114);
and U5799 (N_5799,N_2233,N_3913);
or U5800 (N_5800,N_3458,N_2675);
nor U5801 (N_5801,N_2260,N_2402);
and U5802 (N_5802,N_2587,N_2107);
and U5803 (N_5803,N_2144,N_2329);
and U5804 (N_5804,N_2982,N_2937);
and U5805 (N_5805,N_3075,N_2872);
nand U5806 (N_5806,N_2330,N_2807);
and U5807 (N_5807,N_2216,N_3399);
and U5808 (N_5808,N_3716,N_3872);
or U5809 (N_5809,N_2987,N_3004);
or U5810 (N_5810,N_3404,N_2143);
nor U5811 (N_5811,N_3236,N_3926);
nand U5812 (N_5812,N_2875,N_2902);
xor U5813 (N_5813,N_3675,N_2852);
or U5814 (N_5814,N_3984,N_2873);
nand U5815 (N_5815,N_2616,N_2387);
and U5816 (N_5816,N_2227,N_2266);
or U5817 (N_5817,N_2511,N_2917);
nor U5818 (N_5818,N_3743,N_3738);
or U5819 (N_5819,N_3817,N_2094);
or U5820 (N_5820,N_2919,N_2830);
xnor U5821 (N_5821,N_3697,N_3832);
nor U5822 (N_5822,N_3184,N_3043);
or U5823 (N_5823,N_2110,N_3886);
or U5824 (N_5824,N_2578,N_3157);
nand U5825 (N_5825,N_3043,N_2372);
nand U5826 (N_5826,N_2420,N_2558);
or U5827 (N_5827,N_3017,N_3400);
nand U5828 (N_5828,N_2653,N_3459);
or U5829 (N_5829,N_3356,N_3760);
nor U5830 (N_5830,N_3845,N_3998);
and U5831 (N_5831,N_3399,N_2594);
or U5832 (N_5832,N_3099,N_2539);
nand U5833 (N_5833,N_3467,N_2562);
or U5834 (N_5834,N_3310,N_3504);
xor U5835 (N_5835,N_3884,N_2015);
nand U5836 (N_5836,N_2544,N_3790);
nor U5837 (N_5837,N_2449,N_2538);
nand U5838 (N_5838,N_2272,N_2788);
and U5839 (N_5839,N_2536,N_2604);
nor U5840 (N_5840,N_3791,N_3086);
or U5841 (N_5841,N_3619,N_2578);
or U5842 (N_5842,N_2344,N_2103);
xor U5843 (N_5843,N_2072,N_3933);
and U5844 (N_5844,N_2913,N_3017);
xor U5845 (N_5845,N_3408,N_3386);
or U5846 (N_5846,N_2169,N_3400);
nor U5847 (N_5847,N_3676,N_3801);
nor U5848 (N_5848,N_3628,N_2085);
xor U5849 (N_5849,N_2453,N_3982);
and U5850 (N_5850,N_2972,N_2549);
and U5851 (N_5851,N_2873,N_2721);
and U5852 (N_5852,N_3402,N_2845);
nand U5853 (N_5853,N_2332,N_3923);
nand U5854 (N_5854,N_3227,N_3660);
or U5855 (N_5855,N_3875,N_2153);
xnor U5856 (N_5856,N_2931,N_3105);
nor U5857 (N_5857,N_3010,N_2251);
nor U5858 (N_5858,N_3336,N_2026);
nand U5859 (N_5859,N_3954,N_2863);
nand U5860 (N_5860,N_2715,N_3432);
nand U5861 (N_5861,N_2656,N_3182);
xnor U5862 (N_5862,N_3772,N_3312);
or U5863 (N_5863,N_2392,N_3980);
and U5864 (N_5864,N_2390,N_2219);
nand U5865 (N_5865,N_2749,N_3477);
and U5866 (N_5866,N_2159,N_3846);
or U5867 (N_5867,N_2611,N_3834);
xor U5868 (N_5868,N_3003,N_3890);
nand U5869 (N_5869,N_3236,N_2383);
nor U5870 (N_5870,N_3423,N_3174);
or U5871 (N_5871,N_2870,N_2217);
nand U5872 (N_5872,N_2563,N_2428);
and U5873 (N_5873,N_2177,N_2129);
or U5874 (N_5874,N_3044,N_2731);
or U5875 (N_5875,N_2478,N_2551);
nor U5876 (N_5876,N_3872,N_3958);
and U5877 (N_5877,N_3916,N_2164);
nor U5878 (N_5878,N_2446,N_3875);
and U5879 (N_5879,N_2503,N_2532);
or U5880 (N_5880,N_3170,N_3158);
or U5881 (N_5881,N_2206,N_3594);
nor U5882 (N_5882,N_2667,N_3579);
and U5883 (N_5883,N_3301,N_3394);
nand U5884 (N_5884,N_2949,N_2825);
nor U5885 (N_5885,N_3060,N_3049);
and U5886 (N_5886,N_3508,N_3213);
or U5887 (N_5887,N_3046,N_3546);
nand U5888 (N_5888,N_2507,N_3584);
nor U5889 (N_5889,N_2771,N_3001);
nor U5890 (N_5890,N_3325,N_2169);
nand U5891 (N_5891,N_2551,N_3949);
or U5892 (N_5892,N_2130,N_3397);
and U5893 (N_5893,N_2555,N_2579);
or U5894 (N_5894,N_3800,N_2994);
nand U5895 (N_5895,N_2539,N_2975);
and U5896 (N_5896,N_2405,N_2843);
nor U5897 (N_5897,N_2092,N_2961);
nand U5898 (N_5898,N_2458,N_3191);
and U5899 (N_5899,N_2564,N_3492);
xnor U5900 (N_5900,N_2864,N_3022);
nor U5901 (N_5901,N_3666,N_3369);
nor U5902 (N_5902,N_2025,N_2206);
or U5903 (N_5903,N_2254,N_3458);
nor U5904 (N_5904,N_2216,N_2728);
nor U5905 (N_5905,N_3892,N_2875);
nand U5906 (N_5906,N_3192,N_2504);
and U5907 (N_5907,N_3840,N_2592);
or U5908 (N_5908,N_2625,N_2075);
and U5909 (N_5909,N_2664,N_2191);
xor U5910 (N_5910,N_2790,N_2070);
or U5911 (N_5911,N_3906,N_3580);
and U5912 (N_5912,N_3532,N_2002);
nand U5913 (N_5913,N_2087,N_3580);
nor U5914 (N_5914,N_2017,N_2112);
nand U5915 (N_5915,N_2616,N_2832);
nor U5916 (N_5916,N_2557,N_3503);
nor U5917 (N_5917,N_3976,N_3719);
nor U5918 (N_5918,N_3667,N_2826);
xnor U5919 (N_5919,N_2953,N_3769);
and U5920 (N_5920,N_2663,N_2995);
nor U5921 (N_5921,N_3626,N_3273);
xnor U5922 (N_5922,N_3077,N_3837);
or U5923 (N_5923,N_2051,N_2487);
nand U5924 (N_5924,N_3563,N_2300);
or U5925 (N_5925,N_3935,N_2210);
or U5926 (N_5926,N_2119,N_2182);
nor U5927 (N_5927,N_2719,N_3626);
nor U5928 (N_5928,N_2741,N_3771);
nand U5929 (N_5929,N_3334,N_2011);
xnor U5930 (N_5930,N_3526,N_2010);
xnor U5931 (N_5931,N_3043,N_3297);
xor U5932 (N_5932,N_3958,N_2350);
nor U5933 (N_5933,N_3119,N_2492);
and U5934 (N_5934,N_3438,N_3375);
nand U5935 (N_5935,N_3050,N_3551);
xor U5936 (N_5936,N_2913,N_3768);
and U5937 (N_5937,N_2804,N_2883);
xor U5938 (N_5938,N_3285,N_3361);
or U5939 (N_5939,N_3653,N_2582);
or U5940 (N_5940,N_3594,N_2936);
or U5941 (N_5941,N_2222,N_3460);
xnor U5942 (N_5942,N_3113,N_3771);
or U5943 (N_5943,N_2040,N_2313);
and U5944 (N_5944,N_3385,N_3572);
or U5945 (N_5945,N_3975,N_3301);
xnor U5946 (N_5946,N_2542,N_3774);
nand U5947 (N_5947,N_3023,N_2508);
nand U5948 (N_5948,N_3604,N_3771);
nor U5949 (N_5949,N_2726,N_3954);
nand U5950 (N_5950,N_2684,N_2378);
xnor U5951 (N_5951,N_3778,N_3605);
nand U5952 (N_5952,N_3226,N_2247);
or U5953 (N_5953,N_3432,N_3457);
or U5954 (N_5954,N_3082,N_2511);
nor U5955 (N_5955,N_2216,N_2423);
nand U5956 (N_5956,N_3400,N_3455);
or U5957 (N_5957,N_2289,N_2196);
and U5958 (N_5958,N_3294,N_2450);
or U5959 (N_5959,N_2426,N_2791);
or U5960 (N_5960,N_2364,N_3593);
xnor U5961 (N_5961,N_2905,N_3718);
nand U5962 (N_5962,N_2760,N_2602);
or U5963 (N_5963,N_3770,N_2137);
or U5964 (N_5964,N_3615,N_3790);
nor U5965 (N_5965,N_3628,N_2004);
and U5966 (N_5966,N_2474,N_2216);
xnor U5967 (N_5967,N_2053,N_3156);
nand U5968 (N_5968,N_2716,N_2387);
nand U5969 (N_5969,N_2517,N_3564);
and U5970 (N_5970,N_2605,N_3390);
nor U5971 (N_5971,N_2295,N_3568);
xnor U5972 (N_5972,N_2623,N_3333);
nand U5973 (N_5973,N_3370,N_3670);
nand U5974 (N_5974,N_3021,N_3031);
or U5975 (N_5975,N_3126,N_2587);
and U5976 (N_5976,N_3873,N_2694);
nor U5977 (N_5977,N_3513,N_3996);
or U5978 (N_5978,N_2570,N_2528);
nor U5979 (N_5979,N_2094,N_3545);
nor U5980 (N_5980,N_3753,N_3279);
and U5981 (N_5981,N_3530,N_2982);
or U5982 (N_5982,N_3137,N_3299);
nor U5983 (N_5983,N_3355,N_2729);
xnor U5984 (N_5984,N_3038,N_3776);
nor U5985 (N_5985,N_3178,N_2398);
nand U5986 (N_5986,N_2713,N_3521);
xor U5987 (N_5987,N_2883,N_3477);
nor U5988 (N_5988,N_3538,N_3212);
nand U5989 (N_5989,N_2047,N_3939);
nand U5990 (N_5990,N_2403,N_2124);
and U5991 (N_5991,N_2306,N_2644);
xor U5992 (N_5992,N_3120,N_2459);
and U5993 (N_5993,N_2938,N_3212);
or U5994 (N_5994,N_3074,N_3232);
nand U5995 (N_5995,N_2936,N_3643);
or U5996 (N_5996,N_3885,N_2498);
nor U5997 (N_5997,N_2353,N_3104);
or U5998 (N_5998,N_3843,N_3570);
nor U5999 (N_5999,N_3214,N_2436);
or U6000 (N_6000,N_5527,N_5092);
and U6001 (N_6001,N_5535,N_4995);
or U6002 (N_6002,N_5890,N_5095);
nor U6003 (N_6003,N_4239,N_4007);
or U6004 (N_6004,N_4884,N_4607);
nor U6005 (N_6005,N_5748,N_5870);
nand U6006 (N_6006,N_5462,N_4271);
nor U6007 (N_6007,N_4197,N_5503);
or U6008 (N_6008,N_4925,N_4045);
nor U6009 (N_6009,N_4701,N_4377);
nor U6010 (N_6010,N_4026,N_5582);
nand U6011 (N_6011,N_4190,N_5264);
nand U6012 (N_6012,N_4285,N_5616);
nand U6013 (N_6013,N_5229,N_5162);
xnor U6014 (N_6014,N_4895,N_4466);
nand U6015 (N_6015,N_5836,N_5041);
nand U6016 (N_6016,N_4100,N_4678);
and U6017 (N_6017,N_5115,N_4220);
xnor U6018 (N_6018,N_4738,N_5546);
and U6019 (N_6019,N_5165,N_4296);
and U6020 (N_6020,N_5654,N_4522);
and U6021 (N_6021,N_4828,N_5333);
and U6022 (N_6022,N_4796,N_4155);
nor U6023 (N_6023,N_4105,N_5119);
or U6024 (N_6024,N_4689,N_5519);
or U6025 (N_6025,N_4160,N_5743);
and U6026 (N_6026,N_5400,N_5130);
and U6027 (N_6027,N_5925,N_4668);
or U6028 (N_6028,N_4735,N_5966);
xor U6029 (N_6029,N_5219,N_5822);
nor U6030 (N_6030,N_4347,N_5961);
or U6031 (N_6031,N_5094,N_4438);
nand U6032 (N_6032,N_5117,N_5929);
nand U6033 (N_6033,N_4393,N_4443);
nor U6034 (N_6034,N_4742,N_4502);
nand U6035 (N_6035,N_5956,N_4189);
nand U6036 (N_6036,N_5808,N_4059);
nor U6037 (N_6037,N_5177,N_5817);
nor U6038 (N_6038,N_5413,N_4693);
and U6039 (N_6039,N_4875,N_4496);
or U6040 (N_6040,N_5238,N_5834);
or U6041 (N_6041,N_4099,N_4856);
nor U6042 (N_6042,N_4208,N_4988);
nand U6043 (N_6043,N_4450,N_5526);
nor U6044 (N_6044,N_5901,N_5428);
nand U6045 (N_6045,N_5299,N_5957);
nand U6046 (N_6046,N_5416,N_4052);
nor U6047 (N_6047,N_5068,N_5626);
and U6048 (N_6048,N_4010,N_4696);
and U6049 (N_6049,N_4919,N_4817);
and U6050 (N_6050,N_5309,N_4824);
nor U6051 (N_6051,N_4511,N_5632);
or U6052 (N_6052,N_5676,N_5829);
nand U6053 (N_6053,N_4628,N_4241);
or U6054 (N_6054,N_5980,N_5935);
nor U6055 (N_6055,N_4287,N_5417);
nor U6056 (N_6056,N_4161,N_4226);
nor U6057 (N_6057,N_4282,N_4308);
and U6058 (N_6058,N_4143,N_5279);
xnor U6059 (N_6059,N_5543,N_5859);
xor U6060 (N_6060,N_4908,N_5713);
nor U6061 (N_6061,N_4156,N_5769);
nor U6062 (N_6062,N_5157,N_4711);
nor U6063 (N_6063,N_5110,N_4371);
nor U6064 (N_6064,N_5927,N_5953);
or U6065 (N_6065,N_4372,N_5537);
and U6066 (N_6066,N_5287,N_4539);
nand U6067 (N_6067,N_4107,N_4993);
or U6068 (N_6068,N_5833,N_4953);
nand U6069 (N_6069,N_5215,N_5572);
and U6070 (N_6070,N_5320,N_4872);
or U6071 (N_6071,N_5058,N_5600);
nor U6072 (N_6072,N_4302,N_5650);
xnor U6073 (N_6073,N_5906,N_5342);
nand U6074 (N_6074,N_4719,N_5647);
and U6075 (N_6075,N_4986,N_4427);
nand U6076 (N_6076,N_4721,N_4391);
or U6077 (N_6077,N_4221,N_4482);
nand U6078 (N_6078,N_5217,N_5746);
or U6079 (N_6079,N_4619,N_5666);
nand U6080 (N_6080,N_4829,N_4848);
and U6081 (N_6081,N_4041,N_4124);
nand U6082 (N_6082,N_4493,N_5168);
and U6083 (N_6083,N_4236,N_4057);
or U6084 (N_6084,N_4228,N_4526);
xor U6085 (N_6085,N_4853,N_4334);
nand U6086 (N_6086,N_4501,N_4690);
and U6087 (N_6087,N_4558,N_4777);
nand U6088 (N_6088,N_4675,N_4900);
xor U6089 (N_6089,N_4821,N_4487);
nor U6090 (N_6090,N_5576,N_4219);
nand U6091 (N_6091,N_5096,N_5951);
and U6092 (N_6092,N_4996,N_5545);
and U6093 (N_6093,N_4399,N_5077);
or U6094 (N_6094,N_4645,N_5153);
or U6095 (N_6095,N_5685,N_4048);
nand U6096 (N_6096,N_4449,N_5160);
and U6097 (N_6097,N_4576,N_4209);
or U6098 (N_6098,N_5203,N_5263);
nand U6099 (N_6099,N_4431,N_5126);
and U6100 (N_6100,N_4398,N_4704);
or U6101 (N_6101,N_4213,N_5774);
and U6102 (N_6102,N_5924,N_5023);
xnor U6103 (N_6103,N_5878,N_5381);
or U6104 (N_6104,N_4773,N_4808);
nand U6105 (N_6105,N_4553,N_5761);
and U6106 (N_6106,N_5234,N_4113);
nor U6107 (N_6107,N_5628,N_4842);
and U6108 (N_6108,N_5670,N_5105);
nand U6109 (N_6109,N_4568,N_5308);
or U6110 (N_6110,N_5667,N_5864);
and U6111 (N_6111,N_4657,N_5069);
nor U6112 (N_6112,N_5766,N_5763);
or U6113 (N_6113,N_5211,N_4653);
nor U6114 (N_6114,N_4660,N_4561);
nand U6115 (N_6115,N_5196,N_5240);
nand U6116 (N_6116,N_5163,N_4823);
xor U6117 (N_6117,N_4638,N_5845);
or U6118 (N_6118,N_4877,N_4676);
or U6119 (N_6119,N_4646,N_4324);
nor U6120 (N_6120,N_5158,N_5262);
or U6121 (N_6121,N_5866,N_5590);
and U6122 (N_6122,N_5410,N_4980);
or U6123 (N_6123,N_4977,N_5648);
nor U6124 (N_6124,N_4467,N_5018);
nand U6125 (N_6125,N_5129,N_4374);
nor U6126 (N_6126,N_5950,N_5180);
or U6127 (N_6127,N_5361,N_4182);
nand U6128 (N_6128,N_4267,N_5179);
nor U6129 (N_6129,N_5137,N_5594);
or U6130 (N_6130,N_5249,N_4663);
nand U6131 (N_6131,N_4506,N_5491);
nand U6132 (N_6132,N_4330,N_4290);
nand U6133 (N_6133,N_4178,N_5093);
or U6134 (N_6134,N_5445,N_4637);
nor U6135 (N_6135,N_4193,N_4035);
xnor U6136 (N_6136,N_5990,N_5181);
xnor U6137 (N_6137,N_5700,N_5634);
and U6138 (N_6138,N_5208,N_4751);
xnor U6139 (N_6139,N_4061,N_5668);
nor U6140 (N_6140,N_5882,N_4661);
nor U6141 (N_6141,N_4076,N_5938);
nand U6142 (N_6142,N_5300,N_4433);
or U6143 (N_6143,N_4771,N_5359);
nor U6144 (N_6144,N_5268,N_4176);
nor U6145 (N_6145,N_5360,N_4327);
or U6146 (N_6146,N_5290,N_5236);
or U6147 (N_6147,N_5529,N_4020);
or U6148 (N_6148,N_4713,N_4886);
or U6149 (N_6149,N_4303,N_5678);
and U6150 (N_6150,N_4888,N_4613);
nand U6151 (N_6151,N_5450,N_5739);
nand U6152 (N_6152,N_5827,N_4830);
or U6153 (N_6153,N_5188,N_5837);
xor U6154 (N_6154,N_4958,N_4086);
or U6155 (N_6155,N_4695,N_5948);
nand U6156 (N_6156,N_4862,N_5496);
nor U6157 (N_6157,N_4602,N_5660);
and U6158 (N_6158,N_5765,N_4135);
nor U6159 (N_6159,N_4752,N_5880);
or U6160 (N_6160,N_4621,N_5116);
nor U6161 (N_6161,N_4357,N_5851);
and U6162 (N_6162,N_4520,N_4625);
xor U6163 (N_6163,N_4051,N_5454);
and U6164 (N_6164,N_5464,N_4688);
nor U6165 (N_6165,N_4874,N_4024);
nand U6166 (N_6166,N_4618,N_5191);
nand U6167 (N_6167,N_5883,N_5037);
or U6168 (N_6168,N_4928,N_4305);
nand U6169 (N_6169,N_4543,N_4232);
nand U6170 (N_6170,N_5371,N_4158);
nor U6171 (N_6171,N_4911,N_4034);
nor U6172 (N_6172,N_4974,N_5143);
nor U6173 (N_6173,N_5846,N_5858);
nand U6174 (N_6174,N_5348,N_5121);
nand U6175 (N_6175,N_4536,N_4011);
or U6176 (N_6176,N_4112,N_4710);
nor U6177 (N_6177,N_4110,N_4730);
xor U6178 (N_6178,N_5151,N_5710);
and U6179 (N_6179,N_4413,N_5427);
and U6180 (N_6180,N_5193,N_4906);
nor U6181 (N_6181,N_5050,N_5964);
or U6182 (N_6182,N_4707,N_4442);
or U6183 (N_6183,N_4692,N_5978);
and U6184 (N_6184,N_4832,N_4591);
or U6185 (N_6185,N_4192,N_4534);
nor U6186 (N_6186,N_4441,N_5909);
nand U6187 (N_6187,N_5708,N_5969);
or U6188 (N_6188,N_4163,N_4018);
nor U6189 (N_6189,N_5843,N_5610);
nor U6190 (N_6190,N_5782,N_4896);
nand U6191 (N_6191,N_5184,N_5122);
and U6192 (N_6192,N_4656,N_4074);
and U6193 (N_6193,N_4827,N_4437);
nand U6194 (N_6194,N_5794,N_5169);
nand U6195 (N_6195,N_5335,N_5391);
nand U6196 (N_6196,N_4328,N_5035);
nor U6197 (N_6197,N_4097,N_4078);
nand U6198 (N_6198,N_5141,N_5494);
or U6199 (N_6199,N_5718,N_4669);
nand U6200 (N_6200,N_4120,N_4781);
and U6201 (N_6201,N_5013,N_4352);
nand U6202 (N_6202,N_5759,N_4629);
nor U6203 (N_6203,N_5326,N_4902);
nand U6204 (N_6204,N_4849,N_4488);
nor U6205 (N_6205,N_5672,N_5479);
or U6206 (N_6206,N_5098,N_4293);
nor U6207 (N_6207,N_5271,N_5190);
and U6208 (N_6208,N_5656,N_4733);
nand U6209 (N_6209,N_4126,N_4595);
nor U6210 (N_6210,N_4434,N_5434);
or U6211 (N_6211,N_5532,N_4724);
and U6212 (N_6212,N_4639,N_5871);
nor U6213 (N_6213,N_5675,N_4168);
nand U6214 (N_6214,N_4108,N_4154);
nand U6215 (N_6215,N_5109,N_5011);
and U6216 (N_6216,N_5049,N_5051);
or U6217 (N_6217,N_5895,N_4535);
nor U6218 (N_6218,N_4942,N_4318);
nor U6219 (N_6219,N_5438,N_5226);
and U6220 (N_6220,N_4822,N_4150);
nor U6221 (N_6221,N_4789,N_4390);
nand U6222 (N_6222,N_4262,N_5079);
or U6223 (N_6223,N_4892,N_5892);
nor U6224 (N_6224,N_5235,N_4538);
nand U6225 (N_6225,N_4556,N_5664);
or U6226 (N_6226,N_5409,N_4869);
nor U6227 (N_6227,N_5056,N_5799);
nand U6228 (N_6228,N_5449,N_5558);
xnor U6229 (N_6229,N_5560,N_4409);
or U6230 (N_6230,N_5719,N_5912);
xnor U6231 (N_6231,N_4909,N_4764);
xor U6232 (N_6232,N_4174,N_5877);
nor U6233 (N_6233,N_4729,N_4366);
or U6234 (N_6234,N_5057,N_4732);
nor U6235 (N_6235,N_5317,N_5498);
or U6236 (N_6236,N_5596,N_5627);
nand U6237 (N_6237,N_5161,N_5198);
xnor U6238 (N_6238,N_5824,N_5606);
or U6239 (N_6239,N_4640,N_5362);
nor U6240 (N_6240,N_5974,N_5911);
and U6241 (N_6241,N_5915,N_5302);
or U6242 (N_6242,N_5021,N_5398);
xor U6243 (N_6243,N_4758,N_5237);
and U6244 (N_6244,N_4340,N_4382);
or U6245 (N_6245,N_4876,N_4720);
and U6246 (N_6246,N_5175,N_5478);
and U6247 (N_6247,N_4804,N_4134);
nor U6248 (N_6248,N_5195,N_4858);
and U6249 (N_6249,N_4141,N_4813);
xnor U6250 (N_6250,N_4944,N_4883);
nor U6251 (N_6251,N_5483,N_5727);
nand U6252 (N_6252,N_4799,N_4662);
and U6253 (N_6253,N_4123,N_5644);
nand U6254 (N_6254,N_5977,N_5844);
nor U6255 (N_6255,N_5762,N_5651);
nor U6256 (N_6256,N_5164,N_4300);
or U6257 (N_6257,N_4945,N_5301);
xnor U6258 (N_6258,N_5351,N_4106);
nor U6259 (N_6259,N_5749,N_5534);
nor U6260 (N_6260,N_5176,N_5073);
nor U6261 (N_6261,N_4866,N_4527);
or U6262 (N_6262,N_5455,N_4079);
nand U6263 (N_6263,N_4465,N_4363);
nand U6264 (N_6264,N_5370,N_5415);
and U6265 (N_6265,N_4354,N_5930);
nor U6266 (N_6266,N_4893,N_4857);
nor U6267 (N_6267,N_5541,N_4286);
or U6268 (N_6268,N_4489,N_5293);
xnor U6269 (N_6269,N_4791,N_5394);
xnor U6270 (N_6270,N_5233,N_5019);
nor U6271 (N_6271,N_5554,N_4064);
or U6272 (N_6272,N_4151,N_5500);
and U6273 (N_6273,N_5940,N_4270);
nand U6274 (N_6274,N_4991,N_4575);
and U6275 (N_6275,N_5083,N_5742);
nand U6276 (N_6276,N_4455,N_4075);
xnor U6277 (N_6277,N_5114,N_5559);
nand U6278 (N_6278,N_5745,N_4400);
and U6279 (N_6279,N_4524,N_5379);
nor U6280 (N_6280,N_4083,N_5477);
and U6281 (N_6281,N_4175,N_5783);
nor U6282 (N_6282,N_5932,N_5881);
nor U6283 (N_6283,N_4565,N_4708);
nor U6284 (N_6284,N_5078,N_5914);
nand U6285 (N_6285,N_5091,N_4424);
nor U6286 (N_6286,N_5006,N_5192);
or U6287 (N_6287,N_4985,N_5809);
nor U6288 (N_6288,N_5142,N_4321);
or U6289 (N_6289,N_5721,N_5276);
nor U6290 (N_6290,N_4109,N_4295);
and U6291 (N_6291,N_5828,N_4394);
nor U6292 (N_6292,N_5507,N_5508);
nor U6293 (N_6293,N_4860,N_4544);
xnor U6294 (N_6294,N_5680,N_5586);
nor U6295 (N_6295,N_4320,N_4573);
or U6296 (N_6296,N_4976,N_5777);
xnor U6297 (N_6297,N_5922,N_4005);
or U6298 (N_6298,N_4803,N_5431);
and U6299 (N_6299,N_4968,N_5889);
or U6300 (N_6300,N_5533,N_5459);
and U6301 (N_6301,N_5252,N_4307);
xor U6302 (N_6302,N_4844,N_4929);
xnor U6303 (N_6303,N_4040,N_5949);
nor U6304 (N_6304,N_5973,N_5753);
and U6305 (N_6305,N_4651,N_4338);
xnor U6306 (N_6306,N_4885,N_5820);
nand U6307 (N_6307,N_4187,N_5062);
nor U6308 (N_6308,N_4070,N_5885);
nor U6309 (N_6309,N_5767,N_5609);
or U6310 (N_6310,N_4339,N_4766);
nand U6311 (N_6311,N_5170,N_5599);
and U6312 (N_6312,N_4089,N_5045);
and U6313 (N_6313,N_5277,N_4420);
and U6314 (N_6314,N_4772,N_4463);
nand U6315 (N_6315,N_5256,N_4335);
nand U6316 (N_6316,N_5643,N_5819);
or U6317 (N_6317,N_4594,N_4117);
nand U6318 (N_6318,N_5486,N_5807);
or U6319 (N_6319,N_4947,N_5711);
and U6320 (N_6320,N_4631,N_4746);
or U6321 (N_6321,N_5009,N_4960);
and U6322 (N_6322,N_5404,N_4148);
xor U6323 (N_6323,N_4776,N_4468);
nor U6324 (N_6324,N_4432,N_5502);
nor U6325 (N_6325,N_5107,N_4998);
and U6326 (N_6326,N_4403,N_5795);
nor U6327 (N_6327,N_4627,N_5330);
and U6328 (N_6328,N_5352,N_5778);
nand U6329 (N_6329,N_4418,N_5206);
nor U6330 (N_6330,N_4205,N_4071);
xnor U6331 (N_6331,N_4248,N_5365);
and U6332 (N_6332,N_5801,N_4705);
nand U6333 (N_6333,N_5061,N_5564);
nor U6334 (N_6334,N_4261,N_5064);
and U6335 (N_6335,N_4053,N_5033);
nor U6336 (N_6336,N_5941,N_5364);
nand U6337 (N_6337,N_5341,N_4589);
or U6338 (N_6338,N_5812,N_5955);
xor U6339 (N_6339,N_4769,N_5182);
nor U6340 (N_6340,N_5954,N_4227);
and U6341 (N_6341,N_5460,N_5471);
and U6342 (N_6342,N_4770,N_5020);
nor U6343 (N_6343,N_5149,N_4940);
and U6344 (N_6344,N_4647,N_4727);
and U6345 (N_6345,N_5280,N_4650);
or U6346 (N_6346,N_5452,N_5891);
nand U6347 (N_6347,N_5806,N_5322);
and U6348 (N_6348,N_5108,N_4207);
and U6349 (N_6349,N_5228,N_4868);
nand U6350 (N_6350,N_5216,N_4564);
and U6351 (N_6351,N_4157,N_4069);
or U6352 (N_6352,N_4936,N_5888);
nand U6353 (N_6353,N_5910,N_4878);
or U6354 (N_6354,N_4127,N_4899);
nor U6355 (N_6355,N_5085,N_4412);
nand U6356 (N_6356,N_5592,N_5430);
or U6357 (N_6357,N_4578,N_4843);
xnor U6358 (N_6358,N_4571,N_4376);
and U6359 (N_6359,N_4454,N_5574);
or U6360 (N_6360,N_4211,N_4604);
nor U6361 (N_6361,N_5810,N_4952);
nor U6362 (N_6362,N_4459,N_4333);
or U6363 (N_6363,N_4028,N_4469);
or U6364 (N_6364,N_5875,N_5690);
and U6365 (N_6365,N_4581,N_4624);
or U6366 (N_6366,N_4084,N_5312);
nand U6367 (N_6367,N_4590,N_5306);
or U6368 (N_6368,N_5705,N_4072);
or U6369 (N_6369,N_5042,N_4956);
nor U6370 (N_6370,N_5552,N_4761);
and U6371 (N_6371,N_4782,N_5225);
or U6372 (N_6372,N_4025,N_4671);
xnor U6373 (N_6373,N_5630,N_4677);
nand U6374 (N_6374,N_4038,N_5484);
nand U6375 (N_6375,N_4723,N_5908);
or U6376 (N_6376,N_5612,N_5345);
nand U6377 (N_6377,N_5318,N_5470);
or U6378 (N_6378,N_4491,N_4850);
nand U6379 (N_6379,N_5097,N_4067);
and U6380 (N_6380,N_4898,N_4739);
xor U6381 (N_6381,N_5826,N_4181);
nand U6382 (N_6382,N_4421,N_5793);
nand U6383 (N_6383,N_4429,N_5201);
and U6384 (N_6384,N_5028,N_5729);
or U6385 (N_6385,N_4879,N_4013);
nor U6386 (N_6386,N_5304,N_5946);
nor U6387 (N_6387,N_5993,N_4370);
or U6388 (N_6388,N_5321,N_4255);
nor U6389 (N_6389,N_5038,N_4592);
or U6390 (N_6390,N_5231,N_5566);
nand U6391 (N_6391,N_5022,N_4983);
and U6392 (N_6392,N_4697,N_5084);
nor U6393 (N_6393,N_4448,N_5082);
nand U6394 (N_6394,N_5702,N_5336);
nor U6395 (N_6395,N_5703,N_4863);
nor U6396 (N_6396,N_4703,N_4358);
xor U6397 (N_6397,N_4430,N_4577);
or U6398 (N_6398,N_4180,N_4404);
nor U6399 (N_6399,N_5865,N_5723);
and U6400 (N_6400,N_5907,N_4254);
nor U6401 (N_6401,N_4243,N_5305);
nand U6402 (N_6402,N_5099,N_4445);
and U6403 (N_6403,N_4926,N_5573);
and U6404 (N_6404,N_5923,N_4294);
nor U6405 (N_6405,N_5076,N_5707);
or U6406 (N_6406,N_5232,N_4915);
xnor U6407 (N_6407,N_5601,N_5853);
nand U6408 (N_6408,N_4199,N_5048);
or U6409 (N_6409,N_5960,N_4674);
nand U6410 (N_6410,N_5677,N_4699);
xnor U6411 (N_6411,N_4768,N_5384);
nor U6412 (N_6412,N_5555,N_5147);
and U6413 (N_6413,N_5337,N_5551);
nor U6414 (N_6414,N_4179,N_4224);
nand U6415 (N_6415,N_5687,N_5625);
or U6416 (N_6416,N_4792,N_4162);
and U6417 (N_6417,N_4825,N_5442);
nand U6418 (N_6418,N_4805,N_4840);
or U6419 (N_6419,N_5005,N_4935);
nand U6420 (N_6420,N_5463,N_5372);
nor U6421 (N_6421,N_5135,N_4406);
nor U6422 (N_6422,N_5522,N_5492);
xor U6423 (N_6423,N_5081,N_5172);
or U6424 (N_6424,N_5007,N_4081);
xor U6425 (N_6425,N_4380,N_5619);
xor U6426 (N_6426,N_4289,N_5039);
and U6427 (N_6427,N_4559,N_5173);
xor U6428 (N_6428,N_4206,N_5145);
or U6429 (N_6429,N_5043,N_5367);
nor U6430 (N_6430,N_4615,N_4423);
xnor U6431 (N_6431,N_5608,N_5289);
nor U6432 (N_6432,N_4164,N_5896);
nor U6433 (N_6433,N_5242,N_4636);
nand U6434 (N_6434,N_4167,N_5821);
and U6435 (N_6435,N_4408,N_5303);
and U6436 (N_6436,N_4375,N_5046);
or U6437 (N_6437,N_5008,N_5712);
and U6438 (N_6438,N_4165,N_5433);
or U6439 (N_6439,N_5128,N_4684);
or U6440 (N_6440,N_4183,N_4835);
or U6441 (N_6441,N_4345,N_5520);
nor U6442 (N_6442,N_4683,N_5059);
and U6443 (N_6443,N_4125,N_4200);
and U6444 (N_6444,N_4111,N_4461);
or U6445 (N_6445,N_4278,N_4889);
nor U6446 (N_6446,N_4128,N_5649);
and U6447 (N_6447,N_4060,N_5916);
nor U6448 (N_6448,N_4000,N_5260);
and U6449 (N_6449,N_5358,N_5615);
nor U6450 (N_6450,N_5241,N_4331);
nand U6451 (N_6451,N_4353,N_4251);
nand U6452 (N_6452,N_5926,N_4485);
nand U6453 (N_6453,N_5025,N_5380);
xor U6454 (N_6454,N_5183,N_4475);
or U6455 (N_6455,N_4978,N_5787);
and U6456 (N_6456,N_5490,N_4129);
nor U6457 (N_6457,N_4687,N_4975);
and U6458 (N_6458,N_5611,N_5246);
nand U6459 (N_6459,N_4597,N_5016);
xor U6460 (N_6460,N_5474,N_4728);
and U6461 (N_6461,N_4149,N_4273);
nand U6462 (N_6462,N_4921,N_4519);
and U6463 (N_6463,N_4516,N_4030);
and U6464 (N_6464,N_5402,N_4999);
or U6465 (N_6465,N_5893,N_5512);
nand U6466 (N_6466,N_4685,N_4542);
and U6467 (N_6467,N_4039,N_4523);
nand U6468 (N_6468,N_5429,N_5988);
nand U6469 (N_6469,N_5425,N_4797);
nor U6470 (N_6470,N_5350,N_5257);
and U6471 (N_6471,N_5495,N_4966);
nor U6472 (N_6472,N_5735,N_5991);
and U6473 (N_6473,N_5839,N_4091);
xnor U6474 (N_6474,N_4379,N_4982);
nor U6475 (N_6475,N_5674,N_4009);
nor U6476 (N_6476,N_4541,N_5469);
or U6477 (N_6477,N_4159,N_5239);
nor U6478 (N_6478,N_4600,N_4924);
nor U6479 (N_6479,N_4507,N_5984);
and U6480 (N_6480,N_5602,N_4023);
or U6481 (N_6481,N_4306,N_4831);
xor U6482 (N_6482,N_5032,N_4917);
and U6483 (N_6483,N_5903,N_4140);
nand U6484 (N_6484,N_4166,N_5542);
and U6485 (N_6485,N_5849,N_5771);
and U6486 (N_6486,N_5869,N_5185);
or U6487 (N_6487,N_4029,N_5720);
or U6488 (N_6488,N_4740,N_5740);
xor U6489 (N_6489,N_5716,N_5465);
and U6490 (N_6490,N_5036,N_4044);
and U6491 (N_6491,N_4754,N_5489);
and U6492 (N_6492,N_5751,N_4341);
and U6493 (N_6493,N_4019,N_4880);
or U6494 (N_6494,N_4215,N_5325);
xor U6495 (N_6495,N_4116,N_5150);
nor U6496 (N_6496,N_4622,N_5259);
nand U6497 (N_6497,N_4492,N_4790);
xnor U6498 (N_6498,N_4649,N_5525);
or U6499 (N_6499,N_4686,N_4670);
nand U6500 (N_6500,N_5197,N_4562);
or U6501 (N_6501,N_5331,N_5420);
or U6502 (N_6502,N_4887,N_5186);
and U6503 (N_6503,N_4865,N_5120);
and U6504 (N_6504,N_4003,N_4839);
nor U6505 (N_6505,N_5475,N_4709);
and U6506 (N_6506,N_4043,N_5187);
nand U6507 (N_6507,N_5575,N_4932);
or U6508 (N_6508,N_5741,N_5080);
or U6509 (N_6509,N_4816,N_5657);
and U6510 (N_6510,N_5585,N_5692);
or U6511 (N_6511,N_4903,N_5368);
nand U6512 (N_6512,N_5593,N_4891);
or U6513 (N_6513,N_5298,N_4356);
nand U6514 (N_6514,N_4694,N_4812);
and U6515 (N_6515,N_5272,N_5517);
nor U6516 (N_6516,N_5311,N_5756);
nor U6517 (N_6517,N_4554,N_5204);
nand U6518 (N_6518,N_4195,N_5942);
nor U6519 (N_6519,N_4237,N_5737);
and U6520 (N_6520,N_4579,N_5688);
nor U6521 (N_6521,N_5665,N_5156);
nor U6522 (N_6522,N_4798,N_5562);
nor U6523 (N_6523,N_5734,N_5408);
or U6524 (N_6524,N_5802,N_4833);
and U6525 (N_6525,N_4297,N_4914);
nor U6526 (N_6526,N_4612,N_4731);
or U6527 (N_6527,N_5899,N_5768);
nand U6528 (N_6528,N_5003,N_5835);
nor U6529 (N_6529,N_5701,N_5212);
nor U6530 (N_6530,N_4951,N_5736);
nor U6531 (N_6531,N_5118,N_5291);
xor U6532 (N_6532,N_4806,N_4402);
nor U6533 (N_6533,N_4760,N_4836);
xor U6534 (N_6534,N_5825,N_5544);
nand U6535 (N_6535,N_4245,N_5944);
xnor U6536 (N_6536,N_4610,N_5523);
and U6537 (N_6537,N_5171,N_5933);
and U6538 (N_6538,N_5140,N_5531);
nor U6539 (N_6539,N_5514,N_4864);
and U6540 (N_6540,N_4311,N_4077);
nor U6541 (N_6541,N_5958,N_4006);
nor U6542 (N_6542,N_5111,N_5344);
xor U6543 (N_6543,N_5424,N_5509);
nor U6544 (N_6544,N_4550,N_4266);
nand U6545 (N_6545,N_5060,N_4800);
nand U6546 (N_6546,N_5343,N_5133);
nand U6547 (N_6547,N_4369,N_5653);
nor U6548 (N_6548,N_4419,N_4484);
nand U6549 (N_6549,N_4923,N_5635);
and U6550 (N_6550,N_5389,N_4967);
nand U6551 (N_6551,N_4185,N_4242);
and U6552 (N_6552,N_4389,N_4088);
nand U6553 (N_6553,N_4460,N_4172);
and U6554 (N_6554,N_4132,N_4984);
and U6555 (N_6555,N_5510,N_5072);
xnor U6556 (N_6556,N_4779,N_4349);
nor U6557 (N_6557,N_5178,N_4939);
xnor U6558 (N_6558,N_5658,N_4422);
nor U6559 (N_6559,N_5754,N_5987);
xnor U6560 (N_6560,N_5136,N_5999);
nand U6561 (N_6561,N_5265,N_4714);
and U6562 (N_6562,N_5403,N_4415);
or U6563 (N_6563,N_5587,N_5515);
and U6564 (N_6564,N_4905,N_4959);
nand U6565 (N_6565,N_4969,N_5724);
and U6566 (N_6566,N_4566,N_5591);
or U6567 (N_6567,N_5414,N_4841);
nand U6568 (N_6568,N_5457,N_5931);
nor U6569 (N_6569,N_5441,N_4749);
nor U6570 (N_6570,N_5505,N_4743);
or U6571 (N_6571,N_4802,N_5986);
nor U6572 (N_6572,N_5618,N_4788);
and U6573 (N_6573,N_5224,N_5419);
xor U6574 (N_6574,N_5770,N_5396);
and U6575 (N_6575,N_4722,N_4498);
and U6576 (N_6576,N_4194,N_5339);
nor U6577 (N_6577,N_5223,N_4648);
nand U6578 (N_6578,N_4250,N_4426);
nor U6579 (N_6579,N_4056,N_5620);
and U6580 (N_6580,N_4654,N_5354);
or U6581 (N_6581,N_5518,N_4362);
nor U6582 (N_6582,N_4337,N_4365);
nand U6583 (N_6583,N_5315,N_5790);
nor U6584 (N_6584,N_4546,N_4547);
nor U6585 (N_6585,N_5516,N_4963);
and U6586 (N_6586,N_5472,N_4563);
nand U6587 (N_6587,N_5613,N_5102);
nand U6588 (N_6588,N_5066,N_4476);
or U6589 (N_6589,N_5755,N_4855);
xnor U6590 (N_6590,N_5928,N_5758);
or U6591 (N_6591,N_5563,N_5521);
xor U6592 (N_6592,N_5316,N_5106);
and U6593 (N_6593,N_5528,N_4396);
nor U6594 (N_6594,N_4188,N_4177);
nand U6595 (N_6595,N_5904,N_5524);
xor U6596 (N_6596,N_4934,N_5034);
xnor U6597 (N_6597,N_4186,N_5453);
nand U6598 (N_6598,N_4173,N_4946);
nor U6599 (N_6599,N_4090,N_5788);
and U6600 (N_6600,N_5813,N_4774);
nor U6601 (N_6601,N_5435,N_4169);
nor U6602 (N_6602,N_4961,N_4490);
and U6603 (N_6603,N_4846,N_4994);
or U6604 (N_6604,N_5848,N_5919);
nand U6605 (N_6605,N_4313,N_5861);
and U6606 (N_6606,N_5962,N_4118);
nand U6607 (N_6607,N_4521,N_5730);
and U6608 (N_6608,N_5731,N_5947);
nand U6609 (N_6609,N_4252,N_4279);
nor U6610 (N_6610,N_5887,N_4665);
nand U6611 (N_6611,N_5139,N_5772);
xor U6612 (N_6612,N_4567,N_5934);
and U6613 (N_6613,N_4258,N_4473);
and U6614 (N_6614,N_4263,N_5055);
and U6615 (N_6615,N_4103,N_5636);
and U6616 (N_6616,N_4191,N_5673);
xor U6617 (N_6617,N_4225,N_5659);
nor U6618 (N_6618,N_5860,N_5779);
and U6619 (N_6619,N_4323,N_4170);
and U6620 (N_6620,N_4820,N_5637);
nand U6621 (N_6621,N_4304,N_5423);
nor U6622 (N_6622,N_4505,N_5230);
nand U6623 (N_6623,N_4001,N_5589);
or U6624 (N_6624,N_5965,N_4229);
and U6625 (N_6625,N_5487,N_5681);
and U6626 (N_6626,N_4838,N_4870);
and U6627 (N_6627,N_4322,N_4373);
and U6628 (N_6628,N_5785,N_4726);
and U6629 (N_6629,N_4759,N_4312);
and U6630 (N_6630,N_4316,N_5101);
or U6631 (N_6631,N_5538,N_5357);
nor U6632 (N_6632,N_5283,N_5561);
nor U6633 (N_6633,N_4214,N_5044);
nor U6634 (N_6634,N_5281,N_4047);
nor U6635 (N_6635,N_5972,N_4291);
or U6636 (N_6636,N_4367,N_4497);
nor U6637 (N_6637,N_5997,N_5750);
nand U6638 (N_6638,N_5553,N_5054);
nand U6639 (N_6639,N_4131,N_5661);
nand U6640 (N_6640,N_5967,N_4503);
and U6641 (N_6641,N_4508,N_5070);
nand U6642 (N_6642,N_5994,N_4659);
nand U6643 (N_6643,N_5189,N_5451);
and U6644 (N_6644,N_4301,N_5390);
nor U6645 (N_6645,N_5797,N_4184);
or U6646 (N_6646,N_4681,N_5791);
or U6647 (N_6647,N_5209,N_4231);
nor U6648 (N_6648,N_4809,N_5395);
nor U6649 (N_6649,N_5063,N_5884);
nor U6650 (N_6650,N_5671,N_4818);
nand U6651 (N_6651,N_4845,N_5152);
nand U6652 (N_6652,N_5569,N_4609);
and U6653 (N_6653,N_5565,N_5439);
and U6654 (N_6654,N_5662,N_4098);
or U6655 (N_6655,N_5227,N_5706);
or U6656 (N_6656,N_4203,N_4446);
nand U6657 (N_6657,N_4643,N_4068);
and U6658 (N_6658,N_4472,N_4515);
or U6659 (N_6659,N_5332,N_5982);
and U6660 (N_6660,N_5000,N_5513);
and U6661 (N_6661,N_5663,N_5485);
xor U6662 (N_6662,N_5437,N_4428);
nand U6663 (N_6663,N_4008,N_5399);
nand U6664 (N_6664,N_4269,N_4912);
or U6665 (N_6665,N_4381,N_5773);
nor U6666 (N_6666,N_4264,N_5090);
nor U6667 (N_6667,N_4680,N_4748);
and U6668 (N_6668,N_5579,N_5963);
nor U6669 (N_6669,N_4765,N_5030);
and U6670 (N_6670,N_4753,N_4317);
and U6671 (N_6671,N_5567,N_4588);
nor U6672 (N_6672,N_5728,N_4552);
and U6673 (N_6673,N_4457,N_5695);
nand U6674 (N_6674,N_4268,N_5818);
and U6675 (N_6675,N_5936,N_4210);
and U6676 (N_6676,N_5349,N_4606);
and U6677 (N_6677,N_5200,N_4658);
or U6678 (N_6678,N_4275,N_4032);
nor U6679 (N_6679,N_4778,N_4997);
and U6680 (N_6680,N_5086,N_4144);
nand U6681 (N_6681,N_4453,N_5412);
nand U6682 (N_6682,N_5814,N_5261);
or U6683 (N_6683,N_5571,N_5278);
nand U6684 (N_6684,N_4065,N_4387);
and U6685 (N_6685,N_4310,N_4837);
nor U6686 (N_6686,N_5388,N_5273);
nor U6687 (N_6687,N_5857,N_5346);
or U6688 (N_6688,N_4021,N_4933);
xor U6689 (N_6689,N_4329,N_5800);
or U6690 (N_6690,N_4309,N_5631);
xor U6691 (N_6691,N_4775,N_5131);
and U6692 (N_6692,N_5868,N_5879);
and U6693 (N_6693,N_5418,N_4979);
and U6694 (N_6694,N_4927,N_4031);
nand U6695 (N_6695,N_4901,N_5937);
or U6696 (N_6696,N_5155,N_5401);
nand U6697 (N_6697,N_4223,N_4635);
nor U6698 (N_6698,N_5275,N_4439);
xor U6699 (N_6699,N_4012,N_4212);
nor U6700 (N_6700,N_4259,N_5210);
xor U6701 (N_6701,N_4142,N_4922);
and U6702 (N_6702,N_5296,N_5220);
or U6703 (N_6703,N_5902,N_4957);
nor U6704 (N_6704,N_4583,N_4101);
and U6705 (N_6705,N_4702,N_5466);
or U6706 (N_6706,N_4073,N_5856);
and U6707 (N_6707,N_4634,N_4549);
and U6708 (N_6708,N_5992,N_5863);
nand U6709 (N_6709,N_5294,N_5468);
or U6710 (N_6710,N_4537,N_5598);
xnor U6711 (N_6711,N_4058,N_4509);
or U6712 (N_6712,N_4385,N_4655);
and U6713 (N_6713,N_4082,N_5898);
nand U6714 (N_6714,N_4283,N_4783);
nor U6715 (N_6715,N_5001,N_5319);
nor U6716 (N_6716,N_4626,N_4284);
nor U6717 (N_6717,N_4093,N_4002);
and U6718 (N_6718,N_5968,N_5075);
xnor U6719 (N_6719,N_5027,N_5709);
nand U6720 (N_6720,N_4037,N_4867);
nand U6721 (N_6721,N_4355,N_5269);
and U6722 (N_6722,N_4368,N_5983);
nor U6723 (N_6723,N_5641,N_5338);
nand U6724 (N_6724,N_5698,N_4616);
and U6725 (N_6725,N_5732,N_5780);
nor U6726 (N_6726,N_4277,N_4405);
nor U6727 (N_6727,N_5725,N_4725);
and U6728 (N_6728,N_4036,N_4314);
or U6729 (N_6729,N_4757,N_4943);
and U6730 (N_6730,N_5775,N_4747);
and U6731 (N_6731,N_4717,N_4672);
nand U6732 (N_6732,N_4528,N_4916);
and U6733 (N_6733,N_4990,N_5803);
nor U6734 (N_6734,N_5570,N_4054);
xnor U6735 (N_6735,N_5604,N_5205);
nand U6736 (N_6736,N_5547,N_5146);
and U6737 (N_6737,N_4027,N_4582);
and U6738 (N_6738,N_4533,N_4042);
and U6739 (N_6739,N_4570,N_5411);
xor U6740 (N_6740,N_4470,N_4767);
and U6741 (N_6741,N_5373,N_4055);
or U6742 (N_6742,N_5017,N_5642);
or U6743 (N_6743,N_4897,N_5029);
and U6744 (N_6744,N_5323,N_4096);
nand U6745 (N_6745,N_5623,N_4344);
xor U6746 (N_6746,N_4222,N_4756);
nand U6747 (N_6747,N_4218,N_5760);
nand U6748 (N_6748,N_4411,N_4481);
nor U6749 (N_6749,N_4907,N_5840);
nor U6750 (N_6750,N_5905,N_5697);
and U6751 (N_6751,N_4971,N_4620);
nor U6752 (N_6752,N_4786,N_4395);
or U6753 (N_6753,N_5816,N_5222);
and U6754 (N_6754,N_5733,N_4950);
nor U6755 (N_6755,N_5270,N_4795);
nand U6756 (N_6756,N_4859,N_5501);
xor U6757 (N_6757,N_4049,N_4004);
nand U6758 (N_6758,N_5557,N_5597);
xor U6759 (N_6759,N_5488,N_5577);
nor U6760 (N_6760,N_4585,N_5274);
nor U6761 (N_6761,N_5010,N_5166);
nand U6762 (N_6762,N_5786,N_4274);
or U6763 (N_6763,N_5266,N_5012);
or U6764 (N_6764,N_5148,N_5493);
nand U6765 (N_6765,N_5696,N_4931);
nand U6766 (N_6766,N_4871,N_4572);
or U6767 (N_6767,N_4452,N_5443);
nor U6768 (N_6768,N_5976,N_4826);
nand U6769 (N_6769,N_4346,N_4593);
nand U6770 (N_6770,N_4630,N_4989);
nand U6771 (N_6771,N_5202,N_5284);
nand U6772 (N_6772,N_4679,N_5694);
and U6773 (N_6773,N_5174,N_4930);
nor U6774 (N_6774,N_5481,N_5355);
and U6775 (N_6775,N_5796,N_5382);
or U6776 (N_6776,N_5781,N_4281);
or U6777 (N_6777,N_4632,N_4913);
nand U6778 (N_6778,N_4530,N_5556);
or U6779 (N_6779,N_4417,N_5248);
nor U6780 (N_6780,N_5679,N_5385);
or U6781 (N_6781,N_5805,N_4392);
nor U6782 (N_6782,N_4336,N_5838);
and U6783 (N_6783,N_5607,N_5113);
nand U6784 (N_6784,N_5392,N_5482);
or U6785 (N_6785,N_5683,N_5480);
nor U6786 (N_6786,N_5689,N_4325);
and U6787 (N_6787,N_4249,N_4596);
nand U6788 (N_6788,N_5047,N_5310);
and U6789 (N_6789,N_4234,N_5638);
nor U6790 (N_6790,N_4682,N_5253);
nor U6791 (N_6791,N_4763,N_4288);
nand U6792 (N_6792,N_4378,N_5244);
nand U6793 (N_6793,N_5536,N_5458);
and U6794 (N_6794,N_5832,N_4981);
and U6795 (N_6795,N_5622,N_5347);
or U6796 (N_6796,N_4513,N_5127);
nor U6797 (N_6797,N_5595,N_5314);
nand U6798 (N_6798,N_5581,N_4718);
nor U6799 (N_6799,N_4652,N_4910);
and U6800 (N_6800,N_4601,N_4941);
nor U6801 (N_6801,N_5461,N_5804);
or U6802 (N_6802,N_4949,N_5548);
and U6803 (N_6803,N_4332,N_4954);
and U6804 (N_6804,N_5747,N_5897);
nor U6805 (N_6805,N_5652,N_5920);
nand U6806 (N_6806,N_4608,N_5539);
nand U6807 (N_6807,N_5448,N_4276);
nor U6808 (N_6808,N_5921,N_5798);
or U6809 (N_6809,N_4716,N_5375);
or U6810 (N_6810,N_5530,N_5872);
or U6811 (N_6811,N_4094,N_5629);
nor U6812 (N_6812,N_4964,N_4642);
and U6813 (N_6813,N_4087,N_5847);
xor U6814 (N_6814,N_5250,N_4478);
or U6815 (N_6815,N_4499,N_5605);
nand U6816 (N_6816,N_4834,N_4202);
nor U6817 (N_6817,N_5504,N_4815);
xor U6818 (N_6818,N_4145,N_4750);
nor U6819 (N_6819,N_5421,N_4462);
and U6820 (N_6820,N_5134,N_5307);
and U6821 (N_6821,N_4046,N_4617);
and U6822 (N_6822,N_5945,N_4480);
nor U6823 (N_6823,N_4397,N_5088);
and U6824 (N_6824,N_5757,N_4580);
xor U6825 (N_6825,N_5873,N_4292);
or U6826 (N_6826,N_4486,N_4464);
nor U6827 (N_6827,N_5744,N_4315);
nand U6828 (N_6828,N_4873,N_4384);
nor U6829 (N_6829,N_5640,N_4667);
nor U6830 (N_6830,N_5144,N_5405);
or U6831 (N_6831,N_5862,N_4238);
nor U6832 (N_6832,N_5065,N_5406);
or U6833 (N_6833,N_5540,N_5313);
xor U6834 (N_6834,N_5998,N_5959);
nor U6835 (N_6835,N_4706,N_5811);
or U6836 (N_6836,N_4257,N_5444);
nor U6837 (N_6837,N_5024,N_4698);
nor U6838 (N_6838,N_5568,N_4122);
or U6839 (N_6839,N_4644,N_5614);
xnor U6840 (N_6840,N_5549,N_4881);
and U6841 (N_6841,N_4784,N_5194);
and U6842 (N_6842,N_4256,N_4280);
nor U6843 (N_6843,N_5167,N_5292);
or U6844 (N_6844,N_5717,N_5646);
and U6845 (N_6845,N_4904,N_5633);
xor U6846 (N_6846,N_5714,N_5900);
and U6847 (N_6847,N_4062,N_5715);
nand U6848 (N_6848,N_5089,N_4851);
nand U6849 (N_6849,N_5686,N_4965);
or U6850 (N_6850,N_5831,N_5376);
nand U6851 (N_6851,N_4364,N_4477);
or U6852 (N_6852,N_4479,N_4955);
nand U6853 (N_6853,N_4050,N_4092);
and U6854 (N_6854,N_4115,N_4973);
nor U6855 (N_6855,N_5436,N_4483);
nor U6856 (N_6856,N_4471,N_5255);
or U6857 (N_6857,N_5918,N_4474);
nand U6858 (N_6858,N_4745,N_5040);
nand U6859 (N_6859,N_5580,N_4514);
or U6860 (N_6860,N_5329,N_4201);
nand U6861 (N_6861,N_4504,N_4130);
or U6862 (N_6862,N_5913,N_4253);
or U6863 (N_6863,N_4970,N_4548);
xnor U6864 (N_6864,N_4987,N_5823);
xor U6865 (N_6865,N_5123,N_4586);
nand U6866 (N_6866,N_4712,N_4152);
nand U6867 (N_6867,N_5324,N_5764);
nand U6868 (N_6868,N_5199,N_4787);
nand U6869 (N_6869,N_5624,N_4085);
nand U6870 (N_6870,N_5067,N_4080);
nand U6871 (N_6871,N_5792,N_5841);
and U6872 (N_6872,N_5506,N_4810);
xnor U6873 (N_6873,N_4066,N_4937);
nand U6874 (N_6874,N_4033,N_4359);
and U6875 (N_6875,N_5588,N_4737);
and U6876 (N_6876,N_5125,N_4780);
nand U6877 (N_6877,N_4447,N_5221);
nand U6878 (N_6878,N_5699,N_5004);
and U6879 (N_6879,N_4265,N_5369);
or U6880 (N_6880,N_5267,N_4882);
or U6881 (N_6881,N_4551,N_5894);
and U6882 (N_6882,N_5874,N_4918);
or U6883 (N_6883,N_5655,N_5124);
nor U6884 (N_6884,N_4852,N_4574);
nor U6885 (N_6885,N_5014,N_4383);
and U6886 (N_6886,N_4785,N_5645);
or U6887 (N_6887,N_4235,N_4137);
or U6888 (N_6888,N_4360,N_4611);
or U6889 (N_6889,N_4962,N_4691);
and U6890 (N_6890,N_4014,N_5297);
nand U6891 (N_6891,N_5639,N_4133);
nand U6892 (N_6892,N_4102,N_4715);
xnor U6893 (N_6893,N_5952,N_5691);
nor U6894 (N_6894,N_5356,N_5446);
and U6895 (N_6895,N_4451,N_4440);
or U6896 (N_6896,N_5258,N_4494);
and U6897 (N_6897,N_4890,N_4948);
nor U6898 (N_6898,N_5340,N_5985);
nand U6899 (N_6899,N_4458,N_5876);
nor U6900 (N_6900,N_5989,N_4920);
nand U6901 (N_6901,N_4410,N_4666);
and U6902 (N_6902,N_5295,N_5584);
nor U6903 (N_6903,N_4560,N_4136);
and U6904 (N_6904,N_4138,N_4217);
and U6905 (N_6905,N_4153,N_4171);
or U6906 (N_6906,N_5511,N_5784);
nand U6907 (N_6907,N_5251,N_5074);
nand U6908 (N_6908,N_5981,N_4510);
or U6909 (N_6909,N_4762,N_4196);
or U6910 (N_6910,N_5617,N_5842);
nor U6911 (N_6911,N_5100,N_5327);
and U6912 (N_6912,N_4531,N_4198);
or U6913 (N_6913,N_4584,N_4139);
nand U6914 (N_6914,N_5363,N_5254);
and U6915 (N_6915,N_4319,N_5386);
or U6916 (N_6916,N_4741,N_5288);
nor U6917 (N_6917,N_5789,N_5476);
or U6918 (N_6918,N_5432,N_4744);
nand U6919 (N_6919,N_4495,N_4343);
or U6920 (N_6920,N_5621,N_5578);
nor U6921 (N_6921,N_5071,N_5970);
xnor U6922 (N_6922,N_5850,N_5726);
nand U6923 (N_6923,N_5378,N_5550);
nand U6924 (N_6924,N_4500,N_5467);
nor U6925 (N_6925,N_4348,N_5104);
nor U6926 (N_6926,N_4811,N_4518);
or U6927 (N_6927,N_4569,N_5154);
nor U6928 (N_6928,N_5917,N_4700);
or U6929 (N_6929,N_4095,N_5971);
nand U6930 (N_6930,N_4260,N_5684);
and U6931 (N_6931,N_4299,N_5245);
nand U6932 (N_6932,N_4326,N_5583);
nor U6933 (N_6933,N_5132,N_5407);
and U6934 (N_6934,N_4736,N_4121);
and U6935 (N_6935,N_4022,N_5422);
nand U6936 (N_6936,N_5855,N_4605);
nor U6937 (N_6937,N_4216,N_5752);
and U6938 (N_6938,N_4972,N_5247);
and U6939 (N_6939,N_4351,N_5426);
or U6940 (N_6940,N_4532,N_4529);
and U6941 (N_6941,N_5456,N_4847);
and U6942 (N_6942,N_5447,N_5603);
or U6943 (N_6943,N_4204,N_5213);
nand U6944 (N_6944,N_4425,N_4555);
xnor U6945 (N_6945,N_4342,N_4114);
nand U6946 (N_6946,N_5087,N_4146);
or U6947 (N_6947,N_4272,N_4119);
nor U6948 (N_6948,N_4233,N_5669);
and U6949 (N_6949,N_4388,N_4801);
nor U6950 (N_6950,N_4517,N_5693);
xnor U6951 (N_6951,N_5497,N_5031);
nor U6952 (N_6952,N_5704,N_5473);
xnor U6953 (N_6953,N_5682,N_4247);
and U6954 (N_6954,N_5397,N_4015);
nand U6955 (N_6955,N_4614,N_4623);
xor U6956 (N_6956,N_4545,N_4557);
xnor U6957 (N_6957,N_5285,N_4807);
and U6958 (N_6958,N_4361,N_5026);
nor U6959 (N_6959,N_5015,N_4386);
nand U6960 (N_6960,N_5002,N_5852);
nor U6961 (N_6961,N_5867,N_4641);
nor U6962 (N_6962,N_5103,N_5328);
and U6963 (N_6963,N_4992,N_4793);
or U6964 (N_6964,N_5815,N_4016);
nand U6965 (N_6965,N_5440,N_4244);
nand U6966 (N_6966,N_5979,N_5943);
nor U6967 (N_6967,N_4436,N_5159);
nand U6968 (N_6968,N_5393,N_5776);
or U6969 (N_6969,N_4603,N_5738);
nor U6970 (N_6970,N_4861,N_4414);
or U6971 (N_6971,N_4599,N_5830);
nor U6972 (N_6972,N_4633,N_4673);
or U6973 (N_6973,N_4525,N_5854);
or U6974 (N_6974,N_5377,N_4407);
xor U6975 (N_6975,N_5499,N_5214);
nor U6976 (N_6976,N_4814,N_5722);
and U6977 (N_6977,N_5112,N_5374);
nor U6978 (N_6978,N_5052,N_4938);
nor U6979 (N_6979,N_5996,N_4230);
nor U6980 (N_6980,N_4894,N_4664);
or U6981 (N_6981,N_4416,N_4794);
nand U6982 (N_6982,N_4104,N_4246);
or U6983 (N_6983,N_5334,N_4819);
and U6984 (N_6984,N_4350,N_5218);
or U6985 (N_6985,N_4017,N_4854);
nand U6986 (N_6986,N_5207,N_5995);
and U6987 (N_6987,N_5138,N_5243);
or U6988 (N_6988,N_4456,N_5383);
or U6989 (N_6989,N_4240,N_5353);
or U6990 (N_6990,N_4147,N_4435);
nand U6991 (N_6991,N_4598,N_4512);
and U6992 (N_6992,N_4755,N_4401);
nor U6993 (N_6993,N_5886,N_5387);
or U6994 (N_6994,N_5053,N_5975);
and U6995 (N_6995,N_4734,N_4587);
or U6996 (N_6996,N_5282,N_5286);
nand U6997 (N_6997,N_5366,N_4298);
nor U6998 (N_6998,N_4540,N_5939);
nand U6999 (N_6999,N_4444,N_4063);
and U7000 (N_7000,N_4720,N_5568);
xnor U7001 (N_7001,N_5659,N_5826);
nand U7002 (N_7002,N_5253,N_5348);
or U7003 (N_7003,N_4531,N_4499);
or U7004 (N_7004,N_4870,N_4474);
and U7005 (N_7005,N_5161,N_5522);
nand U7006 (N_7006,N_5189,N_5296);
nand U7007 (N_7007,N_5673,N_5424);
nor U7008 (N_7008,N_5383,N_4169);
nor U7009 (N_7009,N_5911,N_4454);
or U7010 (N_7010,N_4005,N_4017);
and U7011 (N_7011,N_4370,N_5645);
and U7012 (N_7012,N_5627,N_5975);
or U7013 (N_7013,N_4350,N_5902);
nor U7014 (N_7014,N_5680,N_5027);
or U7015 (N_7015,N_4730,N_4636);
nor U7016 (N_7016,N_5157,N_5196);
nor U7017 (N_7017,N_4621,N_5627);
and U7018 (N_7018,N_4869,N_4675);
and U7019 (N_7019,N_4465,N_5499);
nor U7020 (N_7020,N_4858,N_5949);
and U7021 (N_7021,N_4620,N_5436);
nand U7022 (N_7022,N_5404,N_4731);
xnor U7023 (N_7023,N_4414,N_5118);
nor U7024 (N_7024,N_4799,N_5872);
nand U7025 (N_7025,N_4446,N_5741);
and U7026 (N_7026,N_4597,N_5257);
or U7027 (N_7027,N_5766,N_4646);
nor U7028 (N_7028,N_5698,N_5500);
nor U7029 (N_7029,N_4154,N_5143);
and U7030 (N_7030,N_5766,N_5769);
and U7031 (N_7031,N_4324,N_5483);
nand U7032 (N_7032,N_5871,N_5887);
nor U7033 (N_7033,N_5670,N_5618);
nand U7034 (N_7034,N_5469,N_5827);
and U7035 (N_7035,N_4375,N_4858);
xor U7036 (N_7036,N_4417,N_4167);
xor U7037 (N_7037,N_5691,N_5777);
or U7038 (N_7038,N_4215,N_4012);
nor U7039 (N_7039,N_5685,N_5316);
nor U7040 (N_7040,N_5835,N_4335);
and U7041 (N_7041,N_5617,N_5972);
or U7042 (N_7042,N_5364,N_4812);
xnor U7043 (N_7043,N_4980,N_5032);
or U7044 (N_7044,N_5428,N_5541);
xnor U7045 (N_7045,N_4106,N_5108);
nand U7046 (N_7046,N_4354,N_5903);
and U7047 (N_7047,N_5317,N_4404);
or U7048 (N_7048,N_4582,N_5246);
and U7049 (N_7049,N_4079,N_5160);
nor U7050 (N_7050,N_4946,N_4183);
nor U7051 (N_7051,N_4882,N_5225);
nand U7052 (N_7052,N_4901,N_4953);
and U7053 (N_7053,N_5264,N_4336);
or U7054 (N_7054,N_5100,N_4594);
xnor U7055 (N_7055,N_4515,N_4316);
xor U7056 (N_7056,N_4706,N_5886);
nand U7057 (N_7057,N_4321,N_4504);
and U7058 (N_7058,N_5993,N_5699);
nand U7059 (N_7059,N_5719,N_5733);
nand U7060 (N_7060,N_5517,N_4241);
nand U7061 (N_7061,N_4330,N_5467);
nand U7062 (N_7062,N_4653,N_5042);
nor U7063 (N_7063,N_4615,N_5879);
xnor U7064 (N_7064,N_5357,N_4363);
and U7065 (N_7065,N_5585,N_4155);
nand U7066 (N_7066,N_5441,N_5094);
or U7067 (N_7067,N_4186,N_4875);
nor U7068 (N_7068,N_5701,N_5341);
or U7069 (N_7069,N_5780,N_5006);
nor U7070 (N_7070,N_4232,N_5199);
and U7071 (N_7071,N_5635,N_5541);
nor U7072 (N_7072,N_5836,N_5467);
nand U7073 (N_7073,N_5433,N_4480);
or U7074 (N_7074,N_4382,N_5647);
nor U7075 (N_7075,N_4965,N_4667);
nor U7076 (N_7076,N_4284,N_5619);
xor U7077 (N_7077,N_5181,N_4186);
nand U7078 (N_7078,N_5979,N_5289);
nor U7079 (N_7079,N_5322,N_5912);
nor U7080 (N_7080,N_5766,N_5991);
nor U7081 (N_7081,N_5714,N_4160);
xor U7082 (N_7082,N_5397,N_4288);
or U7083 (N_7083,N_4169,N_4117);
xnor U7084 (N_7084,N_4899,N_4826);
and U7085 (N_7085,N_4813,N_4783);
or U7086 (N_7086,N_4005,N_4218);
and U7087 (N_7087,N_5487,N_4930);
xnor U7088 (N_7088,N_4261,N_4591);
xor U7089 (N_7089,N_5964,N_4041);
or U7090 (N_7090,N_5579,N_5580);
and U7091 (N_7091,N_4090,N_5214);
nand U7092 (N_7092,N_5829,N_4229);
nor U7093 (N_7093,N_4088,N_4493);
xor U7094 (N_7094,N_4723,N_4815);
xnor U7095 (N_7095,N_4249,N_4439);
or U7096 (N_7096,N_4234,N_4306);
nand U7097 (N_7097,N_4605,N_5594);
and U7098 (N_7098,N_4203,N_5123);
xnor U7099 (N_7099,N_5265,N_4329);
or U7100 (N_7100,N_5543,N_5343);
or U7101 (N_7101,N_5553,N_4965);
and U7102 (N_7102,N_4830,N_4518);
and U7103 (N_7103,N_4255,N_4904);
nor U7104 (N_7104,N_4072,N_4524);
nor U7105 (N_7105,N_4382,N_5317);
xor U7106 (N_7106,N_5828,N_5469);
and U7107 (N_7107,N_5348,N_5182);
nand U7108 (N_7108,N_4781,N_4368);
nor U7109 (N_7109,N_4835,N_5940);
nand U7110 (N_7110,N_5939,N_4176);
or U7111 (N_7111,N_5897,N_5412);
and U7112 (N_7112,N_4219,N_4711);
nor U7113 (N_7113,N_5363,N_4859);
nand U7114 (N_7114,N_5702,N_4045);
nor U7115 (N_7115,N_4779,N_5399);
or U7116 (N_7116,N_5215,N_5509);
nand U7117 (N_7117,N_4522,N_5109);
nand U7118 (N_7118,N_5108,N_5112);
xnor U7119 (N_7119,N_4352,N_5487);
nor U7120 (N_7120,N_4904,N_5638);
and U7121 (N_7121,N_5169,N_5223);
xnor U7122 (N_7122,N_5985,N_4703);
and U7123 (N_7123,N_4787,N_5230);
or U7124 (N_7124,N_5759,N_4700);
or U7125 (N_7125,N_5059,N_5527);
and U7126 (N_7126,N_4558,N_5792);
nor U7127 (N_7127,N_4526,N_5545);
nand U7128 (N_7128,N_4819,N_4469);
or U7129 (N_7129,N_4024,N_4189);
or U7130 (N_7130,N_4378,N_4077);
and U7131 (N_7131,N_5572,N_5056);
or U7132 (N_7132,N_4067,N_5597);
xnor U7133 (N_7133,N_5367,N_4068);
nor U7134 (N_7134,N_4451,N_5287);
nor U7135 (N_7135,N_5975,N_5205);
and U7136 (N_7136,N_5409,N_5915);
nand U7137 (N_7137,N_4486,N_5060);
nor U7138 (N_7138,N_4824,N_5020);
and U7139 (N_7139,N_4735,N_5047);
and U7140 (N_7140,N_4707,N_5235);
or U7141 (N_7141,N_4983,N_4343);
xnor U7142 (N_7142,N_4856,N_5645);
nor U7143 (N_7143,N_5669,N_4348);
xnor U7144 (N_7144,N_4945,N_5245);
or U7145 (N_7145,N_5173,N_4152);
or U7146 (N_7146,N_4164,N_4307);
xnor U7147 (N_7147,N_5363,N_5376);
nor U7148 (N_7148,N_5465,N_5981);
nand U7149 (N_7149,N_4275,N_5906);
xor U7150 (N_7150,N_5271,N_5587);
and U7151 (N_7151,N_5689,N_4749);
or U7152 (N_7152,N_4036,N_5469);
nand U7153 (N_7153,N_4942,N_5538);
nor U7154 (N_7154,N_4763,N_4349);
nor U7155 (N_7155,N_4451,N_5976);
or U7156 (N_7156,N_4349,N_5583);
nor U7157 (N_7157,N_5700,N_4308);
or U7158 (N_7158,N_5823,N_5230);
or U7159 (N_7159,N_5545,N_5913);
xor U7160 (N_7160,N_5840,N_4013);
or U7161 (N_7161,N_4031,N_4628);
nor U7162 (N_7162,N_5699,N_5175);
nor U7163 (N_7163,N_5831,N_5939);
nand U7164 (N_7164,N_5675,N_5379);
nand U7165 (N_7165,N_4280,N_5844);
nor U7166 (N_7166,N_5069,N_4390);
and U7167 (N_7167,N_5928,N_5726);
and U7168 (N_7168,N_5383,N_4120);
and U7169 (N_7169,N_5071,N_4152);
or U7170 (N_7170,N_4543,N_5007);
and U7171 (N_7171,N_5131,N_4029);
nor U7172 (N_7172,N_4240,N_5624);
nor U7173 (N_7173,N_4683,N_4091);
nor U7174 (N_7174,N_5466,N_4268);
and U7175 (N_7175,N_4868,N_5130);
and U7176 (N_7176,N_5844,N_5253);
xnor U7177 (N_7177,N_5091,N_5173);
and U7178 (N_7178,N_4772,N_4404);
and U7179 (N_7179,N_5530,N_5765);
nand U7180 (N_7180,N_5945,N_4646);
and U7181 (N_7181,N_5420,N_4717);
or U7182 (N_7182,N_5585,N_5058);
or U7183 (N_7183,N_5654,N_4214);
and U7184 (N_7184,N_4760,N_4822);
or U7185 (N_7185,N_5053,N_5136);
nor U7186 (N_7186,N_5122,N_5778);
xor U7187 (N_7187,N_5768,N_5689);
nand U7188 (N_7188,N_4295,N_5666);
nand U7189 (N_7189,N_5744,N_5523);
and U7190 (N_7190,N_4370,N_4452);
xnor U7191 (N_7191,N_5691,N_5591);
nor U7192 (N_7192,N_5548,N_4193);
and U7193 (N_7193,N_4675,N_5291);
nor U7194 (N_7194,N_4335,N_5238);
or U7195 (N_7195,N_5941,N_5780);
and U7196 (N_7196,N_5077,N_5310);
xor U7197 (N_7197,N_5928,N_5197);
xor U7198 (N_7198,N_5963,N_5897);
nor U7199 (N_7199,N_5670,N_4919);
xor U7200 (N_7200,N_4648,N_4191);
nand U7201 (N_7201,N_4081,N_5321);
nor U7202 (N_7202,N_4803,N_5205);
nand U7203 (N_7203,N_5057,N_4806);
or U7204 (N_7204,N_4265,N_4581);
or U7205 (N_7205,N_5204,N_4000);
nor U7206 (N_7206,N_4703,N_4737);
nand U7207 (N_7207,N_5091,N_5295);
and U7208 (N_7208,N_5719,N_5934);
or U7209 (N_7209,N_4642,N_5156);
nand U7210 (N_7210,N_4495,N_5579);
or U7211 (N_7211,N_4984,N_4980);
or U7212 (N_7212,N_5354,N_5531);
nor U7213 (N_7213,N_5605,N_4812);
nor U7214 (N_7214,N_5103,N_5341);
or U7215 (N_7215,N_4172,N_5134);
nand U7216 (N_7216,N_5176,N_4623);
nand U7217 (N_7217,N_4952,N_4921);
or U7218 (N_7218,N_4910,N_5585);
and U7219 (N_7219,N_4645,N_4931);
nor U7220 (N_7220,N_5061,N_4147);
nand U7221 (N_7221,N_4354,N_5039);
nor U7222 (N_7222,N_4318,N_4439);
and U7223 (N_7223,N_5293,N_5762);
nand U7224 (N_7224,N_4858,N_5857);
nand U7225 (N_7225,N_5664,N_5911);
or U7226 (N_7226,N_5709,N_5524);
or U7227 (N_7227,N_4828,N_4783);
and U7228 (N_7228,N_4010,N_5969);
or U7229 (N_7229,N_4508,N_5458);
nand U7230 (N_7230,N_5534,N_5242);
or U7231 (N_7231,N_5721,N_5686);
xor U7232 (N_7232,N_4639,N_4902);
nor U7233 (N_7233,N_5798,N_4922);
and U7234 (N_7234,N_5263,N_4981);
and U7235 (N_7235,N_5861,N_5658);
nand U7236 (N_7236,N_5478,N_5284);
nor U7237 (N_7237,N_4908,N_4140);
nor U7238 (N_7238,N_4038,N_5142);
nor U7239 (N_7239,N_4869,N_4011);
or U7240 (N_7240,N_4633,N_5226);
or U7241 (N_7241,N_5416,N_4272);
nand U7242 (N_7242,N_4912,N_4154);
nor U7243 (N_7243,N_5363,N_4340);
or U7244 (N_7244,N_5928,N_4527);
or U7245 (N_7245,N_5312,N_5322);
or U7246 (N_7246,N_4592,N_5217);
or U7247 (N_7247,N_5977,N_5661);
nand U7248 (N_7248,N_5868,N_5617);
and U7249 (N_7249,N_5153,N_4832);
and U7250 (N_7250,N_4514,N_4719);
or U7251 (N_7251,N_5014,N_5769);
nand U7252 (N_7252,N_4708,N_5224);
and U7253 (N_7253,N_5101,N_5227);
nor U7254 (N_7254,N_5801,N_5561);
and U7255 (N_7255,N_5822,N_4026);
nor U7256 (N_7256,N_5923,N_4759);
xor U7257 (N_7257,N_5628,N_4409);
or U7258 (N_7258,N_5779,N_5682);
nor U7259 (N_7259,N_4844,N_5034);
or U7260 (N_7260,N_5161,N_5759);
nand U7261 (N_7261,N_5602,N_4120);
or U7262 (N_7262,N_4288,N_5146);
or U7263 (N_7263,N_4595,N_5774);
nor U7264 (N_7264,N_5762,N_4260);
nand U7265 (N_7265,N_5573,N_5051);
xor U7266 (N_7266,N_4184,N_5823);
or U7267 (N_7267,N_4791,N_5315);
nor U7268 (N_7268,N_5442,N_5113);
xnor U7269 (N_7269,N_4298,N_4794);
nor U7270 (N_7270,N_5300,N_5917);
and U7271 (N_7271,N_4318,N_4254);
xor U7272 (N_7272,N_5192,N_4646);
and U7273 (N_7273,N_4493,N_4169);
nor U7274 (N_7274,N_4235,N_5351);
and U7275 (N_7275,N_5361,N_5162);
or U7276 (N_7276,N_5942,N_4823);
and U7277 (N_7277,N_4609,N_4137);
xor U7278 (N_7278,N_5518,N_5738);
xnor U7279 (N_7279,N_5950,N_4191);
or U7280 (N_7280,N_4801,N_5678);
nor U7281 (N_7281,N_5391,N_4625);
nor U7282 (N_7282,N_5177,N_5703);
nand U7283 (N_7283,N_4646,N_5448);
and U7284 (N_7284,N_4927,N_4407);
or U7285 (N_7285,N_4191,N_5496);
and U7286 (N_7286,N_4653,N_4291);
nor U7287 (N_7287,N_5552,N_5841);
and U7288 (N_7288,N_5103,N_4117);
and U7289 (N_7289,N_4648,N_4354);
nand U7290 (N_7290,N_4420,N_4821);
nand U7291 (N_7291,N_4021,N_4348);
or U7292 (N_7292,N_4631,N_4195);
nor U7293 (N_7293,N_5158,N_5105);
nand U7294 (N_7294,N_5773,N_4847);
nor U7295 (N_7295,N_4948,N_4517);
or U7296 (N_7296,N_4748,N_5440);
nor U7297 (N_7297,N_4976,N_5275);
or U7298 (N_7298,N_4905,N_5685);
nor U7299 (N_7299,N_5449,N_5074);
and U7300 (N_7300,N_4906,N_5468);
and U7301 (N_7301,N_5866,N_4731);
xor U7302 (N_7302,N_5611,N_5434);
and U7303 (N_7303,N_4172,N_4553);
nor U7304 (N_7304,N_4541,N_4899);
or U7305 (N_7305,N_5204,N_5092);
and U7306 (N_7306,N_4899,N_5694);
and U7307 (N_7307,N_4120,N_5907);
nor U7308 (N_7308,N_4905,N_5756);
nor U7309 (N_7309,N_4607,N_4534);
nor U7310 (N_7310,N_4698,N_4398);
or U7311 (N_7311,N_4244,N_4774);
nand U7312 (N_7312,N_5143,N_5071);
nor U7313 (N_7313,N_5741,N_5792);
nor U7314 (N_7314,N_5067,N_5592);
and U7315 (N_7315,N_4347,N_5150);
and U7316 (N_7316,N_5864,N_4873);
xor U7317 (N_7317,N_4843,N_5759);
and U7318 (N_7318,N_5168,N_4363);
and U7319 (N_7319,N_4627,N_4852);
or U7320 (N_7320,N_4077,N_4260);
or U7321 (N_7321,N_4299,N_5772);
nor U7322 (N_7322,N_5634,N_4327);
nor U7323 (N_7323,N_5162,N_4401);
and U7324 (N_7324,N_4165,N_4711);
nand U7325 (N_7325,N_4306,N_5816);
or U7326 (N_7326,N_4875,N_4060);
nor U7327 (N_7327,N_5928,N_4475);
nor U7328 (N_7328,N_4941,N_5892);
or U7329 (N_7329,N_4296,N_4639);
nand U7330 (N_7330,N_5244,N_4949);
nor U7331 (N_7331,N_4920,N_4349);
or U7332 (N_7332,N_4963,N_4712);
nand U7333 (N_7333,N_5410,N_4013);
nor U7334 (N_7334,N_4341,N_4620);
and U7335 (N_7335,N_5658,N_5190);
or U7336 (N_7336,N_4304,N_5311);
nor U7337 (N_7337,N_4300,N_5405);
or U7338 (N_7338,N_4572,N_5532);
nand U7339 (N_7339,N_4488,N_5110);
or U7340 (N_7340,N_4107,N_5425);
and U7341 (N_7341,N_4951,N_4699);
and U7342 (N_7342,N_5610,N_5432);
nor U7343 (N_7343,N_4755,N_4165);
nor U7344 (N_7344,N_5235,N_4416);
or U7345 (N_7345,N_4132,N_5135);
and U7346 (N_7346,N_4969,N_4993);
nor U7347 (N_7347,N_5892,N_4699);
nand U7348 (N_7348,N_5845,N_5559);
or U7349 (N_7349,N_5105,N_5669);
nor U7350 (N_7350,N_5428,N_4956);
and U7351 (N_7351,N_4831,N_4050);
and U7352 (N_7352,N_4401,N_5993);
and U7353 (N_7353,N_5811,N_5210);
nand U7354 (N_7354,N_4818,N_5260);
and U7355 (N_7355,N_5876,N_4056);
nor U7356 (N_7356,N_5745,N_5279);
and U7357 (N_7357,N_5758,N_4124);
nand U7358 (N_7358,N_4187,N_4093);
nand U7359 (N_7359,N_5097,N_5348);
and U7360 (N_7360,N_4011,N_5544);
nand U7361 (N_7361,N_5071,N_5657);
xnor U7362 (N_7362,N_5908,N_5325);
and U7363 (N_7363,N_4937,N_4811);
and U7364 (N_7364,N_5413,N_4028);
nor U7365 (N_7365,N_4723,N_4748);
or U7366 (N_7366,N_4566,N_4396);
and U7367 (N_7367,N_4277,N_4551);
nor U7368 (N_7368,N_5538,N_5435);
or U7369 (N_7369,N_4792,N_5729);
and U7370 (N_7370,N_5503,N_4237);
nor U7371 (N_7371,N_5190,N_4074);
nor U7372 (N_7372,N_5019,N_4250);
and U7373 (N_7373,N_5016,N_4369);
and U7374 (N_7374,N_4835,N_4842);
nor U7375 (N_7375,N_4686,N_5192);
and U7376 (N_7376,N_4915,N_4639);
nor U7377 (N_7377,N_4535,N_4993);
nor U7378 (N_7378,N_4592,N_4379);
xor U7379 (N_7379,N_4716,N_5834);
nor U7380 (N_7380,N_4901,N_4384);
or U7381 (N_7381,N_5129,N_5668);
or U7382 (N_7382,N_4920,N_4316);
and U7383 (N_7383,N_4702,N_4535);
nor U7384 (N_7384,N_4120,N_4784);
nor U7385 (N_7385,N_5538,N_4864);
nor U7386 (N_7386,N_4956,N_5926);
and U7387 (N_7387,N_4581,N_5628);
and U7388 (N_7388,N_5286,N_5024);
nand U7389 (N_7389,N_5759,N_4522);
xnor U7390 (N_7390,N_4810,N_5917);
nand U7391 (N_7391,N_4203,N_5601);
nand U7392 (N_7392,N_4174,N_5619);
nor U7393 (N_7393,N_4284,N_5645);
nand U7394 (N_7394,N_4091,N_4055);
or U7395 (N_7395,N_5253,N_4582);
and U7396 (N_7396,N_4743,N_4548);
nor U7397 (N_7397,N_4058,N_5519);
or U7398 (N_7398,N_5720,N_5813);
nor U7399 (N_7399,N_4479,N_5338);
or U7400 (N_7400,N_5868,N_4973);
nand U7401 (N_7401,N_5194,N_4115);
nand U7402 (N_7402,N_5178,N_5319);
xnor U7403 (N_7403,N_4061,N_5396);
and U7404 (N_7404,N_4001,N_5494);
or U7405 (N_7405,N_4560,N_5838);
xor U7406 (N_7406,N_5137,N_5913);
nand U7407 (N_7407,N_4147,N_5846);
nor U7408 (N_7408,N_5027,N_4104);
or U7409 (N_7409,N_5321,N_4986);
and U7410 (N_7410,N_4582,N_5501);
nand U7411 (N_7411,N_4699,N_4413);
and U7412 (N_7412,N_5208,N_4258);
nand U7413 (N_7413,N_5673,N_4794);
and U7414 (N_7414,N_4037,N_5924);
or U7415 (N_7415,N_5667,N_4251);
or U7416 (N_7416,N_4872,N_4851);
nor U7417 (N_7417,N_4914,N_5697);
nor U7418 (N_7418,N_4513,N_4417);
nor U7419 (N_7419,N_5279,N_5049);
nor U7420 (N_7420,N_5414,N_4600);
or U7421 (N_7421,N_4444,N_4700);
nor U7422 (N_7422,N_5356,N_5303);
nand U7423 (N_7423,N_4060,N_5746);
and U7424 (N_7424,N_5140,N_5315);
nor U7425 (N_7425,N_5173,N_5736);
and U7426 (N_7426,N_5715,N_4793);
or U7427 (N_7427,N_4715,N_4318);
and U7428 (N_7428,N_5499,N_4439);
xor U7429 (N_7429,N_4894,N_4403);
xnor U7430 (N_7430,N_4611,N_5510);
or U7431 (N_7431,N_4443,N_5120);
and U7432 (N_7432,N_4641,N_4103);
xnor U7433 (N_7433,N_5561,N_5431);
or U7434 (N_7434,N_4429,N_4256);
nand U7435 (N_7435,N_4352,N_4545);
and U7436 (N_7436,N_5815,N_5464);
and U7437 (N_7437,N_4718,N_5275);
or U7438 (N_7438,N_4788,N_5217);
or U7439 (N_7439,N_4050,N_5010);
nand U7440 (N_7440,N_5381,N_5791);
and U7441 (N_7441,N_5463,N_5220);
or U7442 (N_7442,N_5849,N_4505);
nand U7443 (N_7443,N_4099,N_4495);
nand U7444 (N_7444,N_4378,N_5715);
nand U7445 (N_7445,N_4745,N_5829);
xnor U7446 (N_7446,N_5234,N_4774);
nor U7447 (N_7447,N_4516,N_4435);
or U7448 (N_7448,N_5652,N_5377);
and U7449 (N_7449,N_4044,N_5786);
or U7450 (N_7450,N_4417,N_5141);
or U7451 (N_7451,N_4246,N_5504);
nor U7452 (N_7452,N_5498,N_4512);
nand U7453 (N_7453,N_4364,N_4166);
or U7454 (N_7454,N_5382,N_5327);
or U7455 (N_7455,N_4339,N_4616);
nand U7456 (N_7456,N_5665,N_4199);
and U7457 (N_7457,N_4534,N_4780);
nand U7458 (N_7458,N_5531,N_5226);
and U7459 (N_7459,N_5279,N_5685);
or U7460 (N_7460,N_4521,N_5636);
and U7461 (N_7461,N_5394,N_4916);
nor U7462 (N_7462,N_4882,N_4857);
xor U7463 (N_7463,N_5158,N_5040);
or U7464 (N_7464,N_4217,N_5379);
nand U7465 (N_7465,N_4892,N_5135);
or U7466 (N_7466,N_5136,N_4697);
nor U7467 (N_7467,N_5264,N_4375);
nand U7468 (N_7468,N_4510,N_4902);
nor U7469 (N_7469,N_5173,N_4179);
and U7470 (N_7470,N_4824,N_4579);
or U7471 (N_7471,N_5505,N_5957);
nand U7472 (N_7472,N_4314,N_5124);
nor U7473 (N_7473,N_5656,N_4008);
or U7474 (N_7474,N_5513,N_5482);
nor U7475 (N_7475,N_5705,N_5426);
and U7476 (N_7476,N_4226,N_5952);
and U7477 (N_7477,N_4549,N_4477);
or U7478 (N_7478,N_5329,N_5455);
nand U7479 (N_7479,N_4584,N_4091);
nor U7480 (N_7480,N_4702,N_5711);
nor U7481 (N_7481,N_4128,N_5153);
nor U7482 (N_7482,N_4675,N_4791);
or U7483 (N_7483,N_5178,N_5506);
nand U7484 (N_7484,N_4038,N_4820);
or U7485 (N_7485,N_5461,N_5488);
and U7486 (N_7486,N_4962,N_5296);
nor U7487 (N_7487,N_5684,N_4295);
and U7488 (N_7488,N_4434,N_4780);
nor U7489 (N_7489,N_5406,N_4499);
xnor U7490 (N_7490,N_5669,N_5559);
or U7491 (N_7491,N_4004,N_4470);
or U7492 (N_7492,N_4617,N_4530);
nor U7493 (N_7493,N_5785,N_4522);
and U7494 (N_7494,N_4491,N_4058);
or U7495 (N_7495,N_4007,N_4845);
nor U7496 (N_7496,N_4013,N_4454);
nor U7497 (N_7497,N_5719,N_4163);
or U7498 (N_7498,N_5664,N_4695);
and U7499 (N_7499,N_4214,N_5687);
nor U7500 (N_7500,N_4712,N_4589);
nor U7501 (N_7501,N_5292,N_5508);
or U7502 (N_7502,N_4817,N_4621);
or U7503 (N_7503,N_4241,N_4829);
nand U7504 (N_7504,N_4090,N_5861);
or U7505 (N_7505,N_4788,N_5984);
and U7506 (N_7506,N_5498,N_5050);
nand U7507 (N_7507,N_4969,N_4283);
xor U7508 (N_7508,N_4508,N_4885);
or U7509 (N_7509,N_4651,N_5213);
nand U7510 (N_7510,N_4118,N_5417);
nor U7511 (N_7511,N_4215,N_5607);
and U7512 (N_7512,N_4729,N_5629);
nor U7513 (N_7513,N_4327,N_4974);
nand U7514 (N_7514,N_4119,N_5963);
and U7515 (N_7515,N_5093,N_4854);
and U7516 (N_7516,N_5894,N_5948);
nor U7517 (N_7517,N_4778,N_5863);
and U7518 (N_7518,N_5333,N_5663);
or U7519 (N_7519,N_5732,N_4247);
nand U7520 (N_7520,N_4148,N_5640);
nand U7521 (N_7521,N_4560,N_4469);
nand U7522 (N_7522,N_5413,N_4810);
xnor U7523 (N_7523,N_5211,N_5333);
nand U7524 (N_7524,N_5225,N_4276);
nor U7525 (N_7525,N_4524,N_5910);
and U7526 (N_7526,N_5272,N_5312);
nor U7527 (N_7527,N_4342,N_5664);
nor U7528 (N_7528,N_5203,N_5307);
or U7529 (N_7529,N_4759,N_4625);
and U7530 (N_7530,N_5214,N_5062);
and U7531 (N_7531,N_4885,N_5549);
nor U7532 (N_7532,N_4249,N_4531);
and U7533 (N_7533,N_5783,N_4588);
nand U7534 (N_7534,N_5001,N_5475);
and U7535 (N_7535,N_5120,N_5130);
or U7536 (N_7536,N_5413,N_4996);
and U7537 (N_7537,N_5827,N_4170);
or U7538 (N_7538,N_5262,N_5831);
nor U7539 (N_7539,N_5959,N_4097);
xnor U7540 (N_7540,N_5209,N_5954);
nor U7541 (N_7541,N_5521,N_4751);
nor U7542 (N_7542,N_5754,N_4400);
or U7543 (N_7543,N_4851,N_5909);
and U7544 (N_7544,N_4585,N_4107);
nor U7545 (N_7545,N_4919,N_5669);
nand U7546 (N_7546,N_5617,N_5496);
and U7547 (N_7547,N_4337,N_4043);
xnor U7548 (N_7548,N_4550,N_5304);
or U7549 (N_7549,N_5602,N_4533);
or U7550 (N_7550,N_4563,N_5978);
and U7551 (N_7551,N_4435,N_4682);
or U7552 (N_7552,N_4522,N_4191);
xor U7553 (N_7553,N_5096,N_5195);
nand U7554 (N_7554,N_5471,N_5335);
xor U7555 (N_7555,N_4215,N_5730);
nor U7556 (N_7556,N_5121,N_4491);
xnor U7557 (N_7557,N_5109,N_5018);
or U7558 (N_7558,N_4761,N_4567);
nand U7559 (N_7559,N_5455,N_5675);
nor U7560 (N_7560,N_4826,N_4760);
and U7561 (N_7561,N_4063,N_5085);
nand U7562 (N_7562,N_5396,N_5886);
or U7563 (N_7563,N_5105,N_5284);
nand U7564 (N_7564,N_4535,N_4762);
nor U7565 (N_7565,N_5232,N_4215);
xor U7566 (N_7566,N_4618,N_5556);
or U7567 (N_7567,N_4201,N_4810);
nor U7568 (N_7568,N_4226,N_4339);
and U7569 (N_7569,N_4735,N_5687);
nand U7570 (N_7570,N_5792,N_4450);
or U7571 (N_7571,N_4856,N_5654);
nor U7572 (N_7572,N_4751,N_5483);
nor U7573 (N_7573,N_5506,N_5961);
nor U7574 (N_7574,N_5562,N_4386);
nor U7575 (N_7575,N_4119,N_5345);
or U7576 (N_7576,N_4510,N_4797);
or U7577 (N_7577,N_5817,N_4941);
and U7578 (N_7578,N_5164,N_5560);
nor U7579 (N_7579,N_5796,N_5613);
nor U7580 (N_7580,N_4426,N_5135);
or U7581 (N_7581,N_5649,N_5847);
and U7582 (N_7582,N_5126,N_5061);
xor U7583 (N_7583,N_5347,N_4012);
xnor U7584 (N_7584,N_5306,N_5405);
or U7585 (N_7585,N_4083,N_4602);
or U7586 (N_7586,N_5161,N_4096);
and U7587 (N_7587,N_5460,N_4733);
and U7588 (N_7588,N_4450,N_4783);
xor U7589 (N_7589,N_4866,N_4130);
nand U7590 (N_7590,N_5486,N_5505);
nor U7591 (N_7591,N_4232,N_5063);
nand U7592 (N_7592,N_4024,N_4794);
nor U7593 (N_7593,N_4144,N_4756);
xnor U7594 (N_7594,N_4741,N_5017);
and U7595 (N_7595,N_5566,N_4226);
nand U7596 (N_7596,N_5520,N_5036);
nand U7597 (N_7597,N_5008,N_4942);
nand U7598 (N_7598,N_5659,N_5774);
and U7599 (N_7599,N_4232,N_5847);
xnor U7600 (N_7600,N_4415,N_5991);
nand U7601 (N_7601,N_4824,N_4175);
nor U7602 (N_7602,N_5394,N_4874);
nor U7603 (N_7603,N_5056,N_5615);
nand U7604 (N_7604,N_4785,N_4426);
or U7605 (N_7605,N_5999,N_5013);
or U7606 (N_7606,N_5221,N_5256);
nor U7607 (N_7607,N_5940,N_5146);
nand U7608 (N_7608,N_5750,N_4361);
xnor U7609 (N_7609,N_5589,N_4094);
nand U7610 (N_7610,N_4866,N_4274);
nand U7611 (N_7611,N_5906,N_5440);
nand U7612 (N_7612,N_5325,N_5995);
nor U7613 (N_7613,N_5125,N_4150);
xor U7614 (N_7614,N_5658,N_5079);
and U7615 (N_7615,N_4493,N_4785);
xor U7616 (N_7616,N_5431,N_4244);
and U7617 (N_7617,N_4166,N_5318);
xor U7618 (N_7618,N_4645,N_5523);
nand U7619 (N_7619,N_4328,N_5800);
nor U7620 (N_7620,N_5782,N_4750);
and U7621 (N_7621,N_5155,N_5267);
and U7622 (N_7622,N_4251,N_4826);
nor U7623 (N_7623,N_4746,N_5782);
and U7624 (N_7624,N_5241,N_4687);
or U7625 (N_7625,N_5321,N_5337);
nor U7626 (N_7626,N_4367,N_5063);
and U7627 (N_7627,N_4121,N_4559);
nand U7628 (N_7628,N_4091,N_4888);
and U7629 (N_7629,N_5021,N_4668);
nand U7630 (N_7630,N_4657,N_5730);
nand U7631 (N_7631,N_4587,N_5641);
nand U7632 (N_7632,N_4127,N_4811);
nor U7633 (N_7633,N_5439,N_5934);
xor U7634 (N_7634,N_5869,N_4583);
nand U7635 (N_7635,N_5689,N_5111);
nand U7636 (N_7636,N_4380,N_4162);
and U7637 (N_7637,N_5970,N_4607);
or U7638 (N_7638,N_4394,N_4110);
nor U7639 (N_7639,N_5336,N_5165);
nor U7640 (N_7640,N_5733,N_4854);
or U7641 (N_7641,N_4624,N_4815);
nor U7642 (N_7642,N_5791,N_5290);
nand U7643 (N_7643,N_4271,N_5877);
or U7644 (N_7644,N_5099,N_5614);
nand U7645 (N_7645,N_5189,N_4530);
nand U7646 (N_7646,N_5423,N_4681);
nand U7647 (N_7647,N_4062,N_5585);
and U7648 (N_7648,N_5916,N_4589);
nand U7649 (N_7649,N_5465,N_4413);
nand U7650 (N_7650,N_4834,N_4493);
and U7651 (N_7651,N_4901,N_4020);
nor U7652 (N_7652,N_5897,N_5519);
and U7653 (N_7653,N_4437,N_4058);
or U7654 (N_7654,N_5928,N_5173);
nor U7655 (N_7655,N_5736,N_5033);
or U7656 (N_7656,N_5474,N_5754);
or U7657 (N_7657,N_5649,N_4685);
xnor U7658 (N_7658,N_4763,N_4043);
nor U7659 (N_7659,N_5299,N_5609);
and U7660 (N_7660,N_4142,N_5715);
and U7661 (N_7661,N_5510,N_5398);
and U7662 (N_7662,N_5234,N_5104);
nor U7663 (N_7663,N_5209,N_5843);
or U7664 (N_7664,N_4850,N_5993);
and U7665 (N_7665,N_4378,N_5515);
or U7666 (N_7666,N_5380,N_5531);
xnor U7667 (N_7667,N_4849,N_4413);
nor U7668 (N_7668,N_5125,N_5808);
nor U7669 (N_7669,N_4762,N_5050);
nor U7670 (N_7670,N_5344,N_5897);
or U7671 (N_7671,N_5864,N_4297);
and U7672 (N_7672,N_5988,N_4797);
and U7673 (N_7673,N_5931,N_5392);
xnor U7674 (N_7674,N_4506,N_5212);
xnor U7675 (N_7675,N_4440,N_4820);
or U7676 (N_7676,N_4467,N_5142);
nor U7677 (N_7677,N_4523,N_5311);
nor U7678 (N_7678,N_4253,N_4066);
nand U7679 (N_7679,N_5541,N_4378);
and U7680 (N_7680,N_5350,N_4275);
nand U7681 (N_7681,N_5237,N_4192);
nand U7682 (N_7682,N_5831,N_5468);
nor U7683 (N_7683,N_4274,N_4225);
or U7684 (N_7684,N_5223,N_4598);
nor U7685 (N_7685,N_4700,N_5875);
nand U7686 (N_7686,N_5144,N_5586);
and U7687 (N_7687,N_5177,N_4292);
xnor U7688 (N_7688,N_4603,N_4890);
or U7689 (N_7689,N_5252,N_5504);
xnor U7690 (N_7690,N_5268,N_5306);
and U7691 (N_7691,N_4473,N_5588);
nand U7692 (N_7692,N_4201,N_4121);
or U7693 (N_7693,N_5011,N_4205);
nand U7694 (N_7694,N_4961,N_4349);
or U7695 (N_7695,N_5911,N_5550);
or U7696 (N_7696,N_4636,N_4304);
or U7697 (N_7697,N_5352,N_4526);
and U7698 (N_7698,N_4395,N_5893);
or U7699 (N_7699,N_4722,N_5788);
nand U7700 (N_7700,N_5955,N_4195);
xnor U7701 (N_7701,N_4106,N_5082);
and U7702 (N_7702,N_5656,N_4555);
nand U7703 (N_7703,N_4026,N_5369);
and U7704 (N_7704,N_5954,N_4824);
xnor U7705 (N_7705,N_4396,N_5513);
and U7706 (N_7706,N_5475,N_4693);
and U7707 (N_7707,N_5719,N_4829);
nand U7708 (N_7708,N_5006,N_5315);
xor U7709 (N_7709,N_4864,N_5806);
and U7710 (N_7710,N_5717,N_4323);
and U7711 (N_7711,N_5206,N_5344);
xor U7712 (N_7712,N_5829,N_4810);
xnor U7713 (N_7713,N_4113,N_5662);
nand U7714 (N_7714,N_5068,N_5487);
nor U7715 (N_7715,N_5920,N_5701);
nand U7716 (N_7716,N_5891,N_4325);
or U7717 (N_7717,N_5379,N_5999);
and U7718 (N_7718,N_4128,N_5596);
and U7719 (N_7719,N_5877,N_4944);
and U7720 (N_7720,N_5641,N_4430);
nor U7721 (N_7721,N_4013,N_4836);
nand U7722 (N_7722,N_4534,N_4356);
nor U7723 (N_7723,N_5662,N_5757);
or U7724 (N_7724,N_4160,N_4077);
nand U7725 (N_7725,N_5725,N_4233);
and U7726 (N_7726,N_4083,N_4513);
and U7727 (N_7727,N_4860,N_5980);
nand U7728 (N_7728,N_4278,N_4204);
xor U7729 (N_7729,N_5014,N_4452);
and U7730 (N_7730,N_4985,N_5257);
or U7731 (N_7731,N_5509,N_4410);
nand U7732 (N_7732,N_4289,N_5713);
nor U7733 (N_7733,N_5381,N_4092);
and U7734 (N_7734,N_5196,N_4518);
nor U7735 (N_7735,N_5132,N_4566);
nand U7736 (N_7736,N_5399,N_5600);
and U7737 (N_7737,N_4040,N_4222);
nand U7738 (N_7738,N_5647,N_4524);
and U7739 (N_7739,N_5603,N_4557);
nor U7740 (N_7740,N_4623,N_5741);
or U7741 (N_7741,N_4068,N_4656);
nand U7742 (N_7742,N_5842,N_5156);
or U7743 (N_7743,N_4134,N_5061);
or U7744 (N_7744,N_5597,N_5914);
and U7745 (N_7745,N_4894,N_4338);
nand U7746 (N_7746,N_4470,N_4347);
and U7747 (N_7747,N_4003,N_5800);
and U7748 (N_7748,N_5675,N_4587);
or U7749 (N_7749,N_4785,N_4068);
nand U7750 (N_7750,N_5652,N_5994);
or U7751 (N_7751,N_5238,N_5137);
or U7752 (N_7752,N_5337,N_4899);
or U7753 (N_7753,N_5263,N_4576);
nand U7754 (N_7754,N_5902,N_5680);
nor U7755 (N_7755,N_4238,N_5814);
nand U7756 (N_7756,N_5698,N_5977);
or U7757 (N_7757,N_4965,N_5142);
or U7758 (N_7758,N_4254,N_5919);
or U7759 (N_7759,N_5940,N_4725);
xnor U7760 (N_7760,N_4485,N_4825);
xnor U7761 (N_7761,N_5672,N_5440);
nor U7762 (N_7762,N_4006,N_5486);
nand U7763 (N_7763,N_4102,N_4285);
and U7764 (N_7764,N_5076,N_4704);
nor U7765 (N_7765,N_4603,N_5552);
nor U7766 (N_7766,N_5518,N_4901);
nand U7767 (N_7767,N_4511,N_4143);
or U7768 (N_7768,N_4297,N_5190);
nand U7769 (N_7769,N_4132,N_5453);
and U7770 (N_7770,N_4082,N_5892);
nor U7771 (N_7771,N_4638,N_5346);
or U7772 (N_7772,N_5512,N_4395);
nand U7773 (N_7773,N_5237,N_5852);
or U7774 (N_7774,N_4898,N_5895);
or U7775 (N_7775,N_5242,N_4630);
or U7776 (N_7776,N_4445,N_5393);
nand U7777 (N_7777,N_4832,N_5075);
and U7778 (N_7778,N_5466,N_4174);
nand U7779 (N_7779,N_4707,N_5182);
or U7780 (N_7780,N_5444,N_4846);
nor U7781 (N_7781,N_4810,N_5411);
nand U7782 (N_7782,N_4834,N_4317);
nor U7783 (N_7783,N_4513,N_4124);
and U7784 (N_7784,N_5369,N_4318);
nor U7785 (N_7785,N_5896,N_4964);
and U7786 (N_7786,N_4120,N_4468);
nand U7787 (N_7787,N_5795,N_5708);
or U7788 (N_7788,N_4051,N_5579);
and U7789 (N_7789,N_5430,N_4374);
and U7790 (N_7790,N_4528,N_5568);
nor U7791 (N_7791,N_4238,N_5918);
nor U7792 (N_7792,N_4764,N_5446);
and U7793 (N_7793,N_5967,N_4298);
or U7794 (N_7794,N_5784,N_5797);
and U7795 (N_7795,N_4629,N_4764);
nand U7796 (N_7796,N_5323,N_4832);
or U7797 (N_7797,N_5200,N_5902);
and U7798 (N_7798,N_4145,N_4681);
nor U7799 (N_7799,N_4926,N_4407);
xnor U7800 (N_7800,N_5914,N_5444);
xor U7801 (N_7801,N_5751,N_4965);
nand U7802 (N_7802,N_4152,N_5563);
or U7803 (N_7803,N_5814,N_4337);
nor U7804 (N_7804,N_4391,N_4425);
and U7805 (N_7805,N_5837,N_4810);
and U7806 (N_7806,N_5474,N_5196);
and U7807 (N_7807,N_4984,N_4695);
nor U7808 (N_7808,N_4916,N_5682);
xor U7809 (N_7809,N_4029,N_4951);
and U7810 (N_7810,N_5534,N_5722);
or U7811 (N_7811,N_5796,N_5300);
nor U7812 (N_7812,N_4094,N_5825);
nand U7813 (N_7813,N_5850,N_4722);
nor U7814 (N_7814,N_5505,N_5128);
nand U7815 (N_7815,N_4035,N_4605);
or U7816 (N_7816,N_4001,N_4107);
and U7817 (N_7817,N_4801,N_5676);
nand U7818 (N_7818,N_4764,N_5928);
nor U7819 (N_7819,N_4789,N_5063);
xnor U7820 (N_7820,N_5767,N_5464);
nor U7821 (N_7821,N_4458,N_4995);
and U7822 (N_7822,N_5346,N_5450);
nor U7823 (N_7823,N_4445,N_5636);
nand U7824 (N_7824,N_4169,N_5628);
and U7825 (N_7825,N_4068,N_5680);
or U7826 (N_7826,N_4104,N_4718);
nor U7827 (N_7827,N_5508,N_5056);
nand U7828 (N_7828,N_5827,N_5521);
and U7829 (N_7829,N_4379,N_4195);
and U7830 (N_7830,N_4990,N_5305);
nor U7831 (N_7831,N_5979,N_4864);
or U7832 (N_7832,N_5818,N_5251);
and U7833 (N_7833,N_5766,N_4201);
nand U7834 (N_7834,N_4530,N_4202);
nand U7835 (N_7835,N_5715,N_5652);
nand U7836 (N_7836,N_5818,N_4623);
nor U7837 (N_7837,N_4648,N_5273);
and U7838 (N_7838,N_4025,N_5457);
and U7839 (N_7839,N_4850,N_4963);
nor U7840 (N_7840,N_5759,N_4681);
nand U7841 (N_7841,N_4865,N_4963);
nor U7842 (N_7842,N_5843,N_5252);
nand U7843 (N_7843,N_5107,N_4613);
nand U7844 (N_7844,N_4321,N_4697);
nand U7845 (N_7845,N_4119,N_5891);
xnor U7846 (N_7846,N_5749,N_5142);
and U7847 (N_7847,N_5248,N_4819);
nor U7848 (N_7848,N_5174,N_4843);
nor U7849 (N_7849,N_4229,N_5140);
nor U7850 (N_7850,N_4711,N_5363);
nor U7851 (N_7851,N_4975,N_5822);
and U7852 (N_7852,N_4017,N_5223);
xnor U7853 (N_7853,N_5076,N_4489);
or U7854 (N_7854,N_5311,N_4489);
nor U7855 (N_7855,N_5028,N_5605);
or U7856 (N_7856,N_4094,N_5151);
nand U7857 (N_7857,N_4949,N_5429);
or U7858 (N_7858,N_4271,N_5105);
nor U7859 (N_7859,N_5337,N_5525);
and U7860 (N_7860,N_4183,N_4599);
or U7861 (N_7861,N_5795,N_5657);
and U7862 (N_7862,N_5368,N_5659);
nand U7863 (N_7863,N_4917,N_4009);
nand U7864 (N_7864,N_5242,N_5546);
nor U7865 (N_7865,N_5395,N_5878);
nand U7866 (N_7866,N_5718,N_5422);
and U7867 (N_7867,N_5966,N_5545);
nand U7868 (N_7868,N_4094,N_5894);
or U7869 (N_7869,N_5058,N_5672);
nand U7870 (N_7870,N_4831,N_4344);
xor U7871 (N_7871,N_4047,N_4460);
nor U7872 (N_7872,N_5137,N_5165);
and U7873 (N_7873,N_5317,N_4099);
nor U7874 (N_7874,N_4479,N_4128);
nand U7875 (N_7875,N_4299,N_4284);
nor U7876 (N_7876,N_4159,N_4879);
and U7877 (N_7877,N_4214,N_5717);
nor U7878 (N_7878,N_5994,N_5191);
nor U7879 (N_7879,N_5835,N_4487);
nor U7880 (N_7880,N_5857,N_5408);
nor U7881 (N_7881,N_5756,N_4862);
nor U7882 (N_7882,N_4817,N_5890);
nand U7883 (N_7883,N_5833,N_5178);
nand U7884 (N_7884,N_5512,N_4499);
nand U7885 (N_7885,N_5468,N_5764);
nor U7886 (N_7886,N_4217,N_4428);
nor U7887 (N_7887,N_5355,N_4298);
xnor U7888 (N_7888,N_4213,N_5776);
nand U7889 (N_7889,N_4382,N_5157);
nor U7890 (N_7890,N_4560,N_5987);
nor U7891 (N_7891,N_5309,N_5225);
nor U7892 (N_7892,N_5288,N_4710);
nand U7893 (N_7893,N_4262,N_5186);
nand U7894 (N_7894,N_4894,N_4250);
xnor U7895 (N_7895,N_5954,N_4281);
nor U7896 (N_7896,N_4577,N_4768);
or U7897 (N_7897,N_5978,N_5158);
and U7898 (N_7898,N_5111,N_5223);
nor U7899 (N_7899,N_4485,N_4565);
or U7900 (N_7900,N_5169,N_4173);
nor U7901 (N_7901,N_5372,N_4272);
and U7902 (N_7902,N_5241,N_5738);
or U7903 (N_7903,N_4399,N_5386);
or U7904 (N_7904,N_5964,N_5732);
xor U7905 (N_7905,N_4088,N_4305);
nor U7906 (N_7906,N_5971,N_5478);
and U7907 (N_7907,N_5496,N_5795);
nand U7908 (N_7908,N_4471,N_5763);
or U7909 (N_7909,N_4773,N_5607);
or U7910 (N_7910,N_5848,N_5403);
or U7911 (N_7911,N_5155,N_4679);
nor U7912 (N_7912,N_5993,N_4164);
or U7913 (N_7913,N_4861,N_4486);
nor U7914 (N_7914,N_5518,N_4960);
xor U7915 (N_7915,N_4811,N_4260);
and U7916 (N_7916,N_5479,N_4356);
nand U7917 (N_7917,N_5455,N_5672);
nor U7918 (N_7918,N_4409,N_5386);
and U7919 (N_7919,N_4243,N_4848);
nand U7920 (N_7920,N_4064,N_5402);
nand U7921 (N_7921,N_4507,N_4182);
nand U7922 (N_7922,N_4316,N_5184);
or U7923 (N_7923,N_4989,N_5486);
nand U7924 (N_7924,N_5686,N_5314);
and U7925 (N_7925,N_4828,N_5674);
or U7926 (N_7926,N_5732,N_4791);
nor U7927 (N_7927,N_5316,N_5028);
or U7928 (N_7928,N_5275,N_5121);
nand U7929 (N_7929,N_5879,N_5181);
nor U7930 (N_7930,N_5435,N_5068);
and U7931 (N_7931,N_4563,N_4850);
and U7932 (N_7932,N_4569,N_5964);
or U7933 (N_7933,N_5501,N_4726);
nand U7934 (N_7934,N_5644,N_5349);
and U7935 (N_7935,N_4029,N_5998);
nor U7936 (N_7936,N_5080,N_5887);
or U7937 (N_7937,N_5823,N_5310);
nor U7938 (N_7938,N_5123,N_5393);
nand U7939 (N_7939,N_5712,N_4562);
and U7940 (N_7940,N_4473,N_4861);
and U7941 (N_7941,N_4660,N_5935);
xnor U7942 (N_7942,N_5163,N_5007);
nand U7943 (N_7943,N_5475,N_4519);
or U7944 (N_7944,N_4292,N_4271);
nor U7945 (N_7945,N_5090,N_5151);
and U7946 (N_7946,N_4207,N_4297);
or U7947 (N_7947,N_5161,N_5140);
nand U7948 (N_7948,N_5044,N_4971);
nand U7949 (N_7949,N_5910,N_4045);
and U7950 (N_7950,N_4201,N_5207);
nand U7951 (N_7951,N_5027,N_4879);
and U7952 (N_7952,N_5630,N_5679);
nor U7953 (N_7953,N_4601,N_5645);
and U7954 (N_7954,N_4417,N_4180);
and U7955 (N_7955,N_4598,N_4362);
nand U7956 (N_7956,N_4421,N_5314);
nand U7957 (N_7957,N_4216,N_5539);
nand U7958 (N_7958,N_5904,N_4846);
or U7959 (N_7959,N_5780,N_5543);
nor U7960 (N_7960,N_4667,N_5294);
and U7961 (N_7961,N_5857,N_5848);
nand U7962 (N_7962,N_4171,N_4054);
nand U7963 (N_7963,N_5420,N_5144);
or U7964 (N_7964,N_5097,N_5997);
and U7965 (N_7965,N_5379,N_4015);
nor U7966 (N_7966,N_4358,N_5108);
or U7967 (N_7967,N_4946,N_5276);
nand U7968 (N_7968,N_5354,N_4642);
and U7969 (N_7969,N_5520,N_5915);
nand U7970 (N_7970,N_5124,N_4366);
or U7971 (N_7971,N_4597,N_4746);
or U7972 (N_7972,N_5344,N_4179);
or U7973 (N_7973,N_4010,N_5306);
xnor U7974 (N_7974,N_4851,N_4117);
nor U7975 (N_7975,N_4526,N_4930);
nor U7976 (N_7976,N_5416,N_4632);
and U7977 (N_7977,N_5570,N_5070);
or U7978 (N_7978,N_5349,N_4917);
and U7979 (N_7979,N_4032,N_5672);
nor U7980 (N_7980,N_4102,N_5721);
or U7981 (N_7981,N_5901,N_5293);
nand U7982 (N_7982,N_4893,N_5242);
nor U7983 (N_7983,N_5394,N_5036);
or U7984 (N_7984,N_5987,N_5719);
nand U7985 (N_7985,N_5666,N_4972);
nor U7986 (N_7986,N_4542,N_4986);
xnor U7987 (N_7987,N_4830,N_5572);
nand U7988 (N_7988,N_4979,N_4856);
nor U7989 (N_7989,N_5318,N_4081);
and U7990 (N_7990,N_5836,N_4444);
and U7991 (N_7991,N_4864,N_4985);
and U7992 (N_7992,N_4043,N_5996);
nor U7993 (N_7993,N_5144,N_5732);
nor U7994 (N_7994,N_5612,N_5399);
nand U7995 (N_7995,N_4085,N_4464);
nor U7996 (N_7996,N_5643,N_4269);
or U7997 (N_7997,N_4616,N_4081);
and U7998 (N_7998,N_4662,N_5227);
and U7999 (N_7999,N_4436,N_4881);
nand U8000 (N_8000,N_7570,N_7627);
and U8001 (N_8001,N_6638,N_7920);
nand U8002 (N_8002,N_7982,N_7315);
nand U8003 (N_8003,N_7836,N_7531);
xor U8004 (N_8004,N_6919,N_7921);
or U8005 (N_8005,N_7259,N_7950);
or U8006 (N_8006,N_6714,N_7254);
and U8007 (N_8007,N_7962,N_7853);
nand U8008 (N_8008,N_7352,N_7490);
nor U8009 (N_8009,N_6456,N_6136);
nor U8010 (N_8010,N_6414,N_7575);
or U8011 (N_8011,N_7754,N_7038);
or U8012 (N_8012,N_7759,N_6366);
or U8013 (N_8013,N_6242,N_7119);
nor U8014 (N_8014,N_7156,N_7766);
and U8015 (N_8015,N_6920,N_7456);
xnor U8016 (N_8016,N_6803,N_6047);
nand U8017 (N_8017,N_6590,N_7367);
nor U8018 (N_8018,N_7772,N_7187);
or U8019 (N_8019,N_7232,N_6856);
xnor U8020 (N_8020,N_7103,N_6142);
nand U8021 (N_8021,N_6293,N_6932);
and U8022 (N_8022,N_7319,N_7428);
nand U8023 (N_8023,N_6426,N_6143);
nand U8024 (N_8024,N_7663,N_7943);
or U8025 (N_8025,N_6380,N_7910);
and U8026 (N_8026,N_6194,N_7713);
and U8027 (N_8027,N_7897,N_7122);
nand U8028 (N_8028,N_7376,N_7878);
or U8029 (N_8029,N_6875,N_6783);
or U8030 (N_8030,N_6934,N_7970);
or U8031 (N_8031,N_7025,N_6977);
xnor U8032 (N_8032,N_7208,N_6421);
nand U8033 (N_8033,N_6168,N_6525);
nand U8034 (N_8034,N_7653,N_6359);
or U8035 (N_8035,N_6401,N_7652);
nor U8036 (N_8036,N_7662,N_6623);
or U8037 (N_8037,N_6321,N_6035);
nand U8038 (N_8038,N_6184,N_6704);
and U8039 (N_8039,N_6952,N_6526);
and U8040 (N_8040,N_7667,N_6412);
or U8041 (N_8041,N_7194,N_7072);
or U8042 (N_8042,N_7401,N_6436);
or U8043 (N_8043,N_6542,N_6280);
or U8044 (N_8044,N_7565,N_6227);
xor U8045 (N_8045,N_6652,N_7796);
xor U8046 (N_8046,N_7159,N_7391);
xor U8047 (N_8047,N_6802,N_6100);
nor U8048 (N_8048,N_6651,N_6234);
nand U8049 (N_8049,N_6330,N_7102);
or U8050 (N_8050,N_6568,N_6648);
or U8051 (N_8051,N_6267,N_7461);
nor U8052 (N_8052,N_6465,N_6998);
or U8053 (N_8053,N_7478,N_6351);
and U8054 (N_8054,N_6086,N_6643);
nor U8055 (N_8055,N_6554,N_7071);
nand U8056 (N_8056,N_6183,N_6138);
nor U8057 (N_8057,N_6809,N_6709);
nand U8058 (N_8058,N_6043,N_7705);
or U8059 (N_8059,N_7212,N_7394);
and U8060 (N_8060,N_7735,N_7483);
or U8061 (N_8061,N_6780,N_7128);
or U8062 (N_8062,N_6406,N_7585);
or U8063 (N_8063,N_6828,N_7246);
xor U8064 (N_8064,N_7034,N_7137);
or U8065 (N_8065,N_7614,N_6898);
and U8066 (N_8066,N_7683,N_7462);
xor U8067 (N_8067,N_7825,N_6499);
xor U8068 (N_8068,N_7186,N_7057);
xor U8069 (N_8069,N_7534,N_7292);
nand U8070 (N_8070,N_6451,N_6693);
nor U8071 (N_8071,N_7540,N_7473);
or U8072 (N_8072,N_6445,N_7114);
or U8073 (N_8073,N_7323,N_6153);
nand U8074 (N_8074,N_7346,N_7647);
nor U8075 (N_8075,N_6326,N_6766);
xnor U8076 (N_8076,N_7619,N_6307);
or U8077 (N_8077,N_6679,N_7835);
nor U8078 (N_8078,N_7726,N_6073);
nand U8079 (N_8079,N_6974,N_7104);
or U8080 (N_8080,N_6389,N_6983);
nand U8081 (N_8081,N_7582,N_6862);
nor U8082 (N_8082,N_6560,N_6133);
nand U8083 (N_8083,N_7769,N_7058);
nand U8084 (N_8084,N_6925,N_6762);
or U8085 (N_8085,N_6195,N_6287);
nand U8086 (N_8086,N_7499,N_7750);
xor U8087 (N_8087,N_7302,N_6441);
xor U8088 (N_8088,N_7420,N_7266);
and U8089 (N_8089,N_6782,N_6896);
or U8090 (N_8090,N_6805,N_6193);
or U8091 (N_8091,N_6923,N_6569);
and U8092 (N_8092,N_6458,N_6015);
or U8093 (N_8093,N_7996,N_7474);
or U8094 (N_8094,N_6840,N_7841);
or U8095 (N_8095,N_6763,N_7297);
or U8096 (N_8096,N_7320,N_7160);
nand U8097 (N_8097,N_6202,N_6903);
nor U8098 (N_8098,N_7279,N_7060);
xor U8099 (N_8099,N_7800,N_7642);
nand U8100 (N_8100,N_7556,N_7882);
or U8101 (N_8101,N_6595,N_6667);
xor U8102 (N_8102,N_7030,N_6883);
nand U8103 (N_8103,N_7063,N_7694);
nand U8104 (N_8104,N_6502,N_6378);
or U8105 (N_8105,N_7405,N_6570);
nor U8106 (N_8106,N_6586,N_7665);
and U8107 (N_8107,N_7555,N_6311);
nor U8108 (N_8108,N_6812,N_6355);
xor U8109 (N_8109,N_6274,N_7544);
nor U8110 (N_8110,N_6544,N_6771);
nand U8111 (N_8111,N_7550,N_7709);
nor U8112 (N_8112,N_6868,N_6636);
nand U8113 (N_8113,N_6124,N_7560);
or U8114 (N_8114,N_6180,N_6216);
nand U8115 (N_8115,N_7286,N_6446);
xnor U8116 (N_8116,N_6518,N_6395);
and U8117 (N_8117,N_6437,N_7516);
and U8118 (N_8118,N_6323,N_7202);
nand U8119 (N_8119,N_6796,N_6386);
nand U8120 (N_8120,N_7440,N_6928);
or U8121 (N_8121,N_6930,N_6946);
nor U8122 (N_8122,N_6089,N_6251);
nand U8123 (N_8123,N_7887,N_7609);
nand U8124 (N_8124,N_7724,N_6384);
and U8125 (N_8125,N_7249,N_7789);
nor U8126 (N_8126,N_6788,N_6772);
or U8127 (N_8127,N_6684,N_6506);
nand U8128 (N_8128,N_7577,N_6674);
xor U8129 (N_8129,N_7377,N_7347);
or U8130 (N_8130,N_6167,N_6931);
nand U8131 (N_8131,N_6134,N_7728);
nand U8132 (N_8132,N_6675,N_6689);
and U8133 (N_8133,N_6734,N_6831);
or U8134 (N_8134,N_6865,N_6511);
nand U8135 (N_8135,N_7902,N_6591);
or U8136 (N_8136,N_6678,N_7387);
and U8137 (N_8137,N_7118,N_6087);
nor U8138 (N_8138,N_6830,N_7427);
and U8139 (N_8139,N_6147,N_7861);
or U8140 (N_8140,N_6486,N_7725);
nand U8141 (N_8141,N_6484,N_7183);
or U8142 (N_8142,N_6564,N_7009);
or U8143 (N_8143,N_6338,N_6383);
nand U8144 (N_8144,N_7755,N_7078);
nand U8145 (N_8145,N_6580,N_6091);
nand U8146 (N_8146,N_7335,N_7032);
xnor U8147 (N_8147,N_6255,N_6320);
xor U8148 (N_8148,N_7016,N_7244);
nor U8149 (N_8149,N_6341,N_6573);
nand U8150 (N_8150,N_7200,N_6978);
and U8151 (N_8151,N_6177,N_6507);
nand U8152 (N_8152,N_7816,N_6276);
xor U8153 (N_8153,N_6706,N_6254);
nand U8154 (N_8154,N_7088,N_6157);
or U8155 (N_8155,N_7304,N_6808);
or U8156 (N_8156,N_6980,N_6645);
nor U8157 (N_8157,N_7777,N_6516);
and U8158 (N_8158,N_6697,N_6619);
nor U8159 (N_8159,N_6935,N_6661);
or U8160 (N_8160,N_6206,N_7898);
nor U8161 (N_8161,N_6863,N_6083);
nor U8162 (N_8162,N_7955,N_7937);
nor U8163 (N_8163,N_6247,N_7444);
nor U8164 (N_8164,N_7704,N_7406);
xor U8165 (N_8165,N_6936,N_7739);
nand U8166 (N_8166,N_7168,N_6474);
nand U8167 (N_8167,N_6792,N_7947);
or U8168 (N_8168,N_7164,N_6529);
or U8169 (N_8169,N_7052,N_7819);
or U8170 (N_8170,N_7171,N_7701);
nand U8171 (N_8171,N_7975,N_7133);
nor U8172 (N_8172,N_6292,N_6361);
or U8173 (N_8173,N_6747,N_7893);
or U8174 (N_8174,N_6732,N_6713);
nand U8175 (N_8175,N_7888,N_7508);
nand U8176 (N_8176,N_6243,N_7056);
nand U8177 (N_8177,N_6557,N_7365);
nor U8178 (N_8178,N_6328,N_6587);
nand U8179 (N_8179,N_6600,N_6847);
nor U8180 (N_8180,N_6742,N_6239);
nand U8181 (N_8181,N_7722,N_6550);
nor U8182 (N_8182,N_6207,N_7811);
and U8183 (N_8183,N_7929,N_7040);
nand U8184 (N_8184,N_7964,N_6531);
or U8185 (N_8185,N_7572,N_7558);
nor U8186 (N_8186,N_7120,N_7293);
nand U8187 (N_8187,N_7068,N_6765);
nand U8188 (N_8188,N_6937,N_6673);
nand U8189 (N_8189,N_7916,N_6631);
and U8190 (N_8190,N_6635,N_7966);
xor U8191 (N_8191,N_6904,N_6768);
nor U8192 (N_8192,N_6589,N_6343);
xnor U8193 (N_8193,N_7677,N_6253);
or U8194 (N_8194,N_7014,N_7820);
nor U8195 (N_8195,N_6447,N_6781);
xnor U8196 (N_8196,N_6036,N_6284);
nand U8197 (N_8197,N_7075,N_6189);
nor U8198 (N_8198,N_6052,N_7007);
and U8199 (N_8199,N_7423,N_7398);
and U8200 (N_8200,N_7933,N_6533);
nor U8201 (N_8201,N_7054,N_6565);
or U8202 (N_8202,N_7659,N_7219);
or U8203 (N_8203,N_7143,N_6941);
nor U8204 (N_8204,N_7596,N_7760);
nor U8205 (N_8205,N_6439,N_7793);
nor U8206 (N_8206,N_6873,N_7746);
or U8207 (N_8207,N_6902,N_6221);
and U8208 (N_8208,N_7889,N_6427);
or U8209 (N_8209,N_6373,N_6114);
or U8210 (N_8210,N_7859,N_6807);
xnor U8211 (N_8211,N_6773,N_6354);
and U8212 (N_8212,N_6791,N_7903);
or U8213 (N_8213,N_6039,N_6721);
and U8214 (N_8214,N_6670,N_7008);
or U8215 (N_8215,N_7011,N_6612);
and U8216 (N_8216,N_7435,N_7493);
nand U8217 (N_8217,N_6356,N_7954);
nand U8218 (N_8218,N_7633,N_6479);
or U8219 (N_8219,N_7203,N_7334);
nor U8220 (N_8220,N_7446,N_7908);
nor U8221 (N_8221,N_7877,N_7421);
nand U8222 (N_8222,N_7867,N_7096);
or U8223 (N_8223,N_7281,N_7767);
nor U8224 (N_8224,N_7115,N_7094);
nor U8225 (N_8225,N_6859,N_7250);
nand U8226 (N_8226,N_6231,N_7256);
nand U8227 (N_8227,N_7370,N_6158);
nand U8228 (N_8228,N_6972,N_6265);
and U8229 (N_8229,N_6131,N_6758);
or U8230 (N_8230,N_7076,N_6237);
or U8231 (N_8231,N_6815,N_7953);
or U8232 (N_8232,N_6115,N_6761);
or U8233 (N_8233,N_6151,N_6348);
or U8234 (N_8234,N_7576,N_7274);
nor U8235 (N_8235,N_7106,N_6261);
and U8236 (N_8236,N_6614,N_6332);
and U8237 (N_8237,N_6113,N_7031);
nand U8238 (N_8238,N_6599,N_7361);
and U8239 (N_8239,N_6085,N_6214);
xnor U8240 (N_8240,N_6279,N_7794);
xor U8241 (N_8241,N_7695,N_6470);
nor U8242 (N_8242,N_7233,N_6491);
or U8243 (N_8243,N_6744,N_7180);
nor U8244 (N_8244,N_6527,N_7419);
xnor U8245 (N_8245,N_7255,N_7239);
and U8246 (N_8246,N_6101,N_7468);
nor U8247 (N_8247,N_7991,N_6929);
and U8248 (N_8248,N_7533,N_7856);
nand U8249 (N_8249,N_6140,N_7773);
or U8250 (N_8250,N_6461,N_6749);
nor U8251 (N_8251,N_7023,N_6741);
or U8252 (N_8252,N_7395,N_6634);
or U8253 (N_8253,N_6145,N_7736);
or U8254 (N_8254,N_7494,N_7716);
and U8255 (N_8255,N_7300,N_7216);
nor U8256 (N_8256,N_6676,N_7998);
or U8257 (N_8257,N_6466,N_7326);
nand U8258 (N_8258,N_6849,N_6285);
nand U8259 (N_8259,N_6425,N_7876);
and U8260 (N_8260,N_7949,N_6508);
nand U8261 (N_8261,N_7290,N_6583);
and U8262 (N_8262,N_7961,N_6806);
or U8263 (N_8263,N_6109,N_7524);
nor U8264 (N_8264,N_6260,N_7698);
and U8265 (N_8265,N_6213,N_6695);
nand U8266 (N_8266,N_6801,N_7834);
nor U8267 (N_8267,N_7702,N_6534);
and U8268 (N_8268,N_6767,N_6894);
nor U8269 (N_8269,N_6660,N_6942);
xnor U8270 (N_8270,N_6092,N_7855);
nor U8271 (N_8271,N_7229,N_6381);
or U8272 (N_8272,N_7697,N_7042);
nor U8273 (N_8273,N_7827,N_7918);
nand U8274 (N_8274,N_6229,N_6979);
nor U8275 (N_8275,N_7209,N_6129);
nor U8276 (N_8276,N_7097,N_7004);
or U8277 (N_8277,N_7514,N_7803);
or U8278 (N_8278,N_7776,N_7214);
and U8279 (N_8279,N_7673,N_7477);
or U8280 (N_8280,N_6000,N_6141);
nor U8281 (N_8281,N_7476,N_7699);
or U8282 (N_8282,N_7337,N_7931);
nor U8283 (N_8283,N_7817,N_7756);
nor U8284 (N_8284,N_7821,N_6174);
nor U8285 (N_8285,N_6017,N_7313);
nor U8286 (N_8286,N_7938,N_7806);
nand U8287 (N_8287,N_7282,N_6752);
or U8288 (N_8288,N_7605,N_7485);
or U8289 (N_8289,N_6379,N_6751);
and U8290 (N_8290,N_6068,N_6513);
xnor U8291 (N_8291,N_7181,N_6018);
or U8292 (N_8292,N_6517,N_7712);
nor U8293 (N_8293,N_6462,N_7312);
nor U8294 (N_8294,N_7552,N_7808);
xnor U8295 (N_8295,N_7080,N_6116);
or U8296 (N_8296,N_7866,N_6798);
nand U8297 (N_8297,N_7927,N_6112);
nand U8298 (N_8298,N_6236,N_6509);
nor U8299 (N_8299,N_7854,N_7646);
or U8300 (N_8300,N_7567,N_7041);
or U8301 (N_8301,N_7362,N_7449);
nand U8302 (N_8302,N_7668,N_6249);
or U8303 (N_8303,N_6686,N_7551);
or U8304 (N_8304,N_7616,N_7113);
nand U8305 (N_8305,N_7418,N_7740);
nand U8306 (N_8306,N_6077,N_7172);
and U8307 (N_8307,N_6520,N_7610);
xnor U8308 (N_8308,N_7348,N_7590);
nand U8309 (N_8309,N_6913,N_7924);
xnor U8310 (N_8310,N_6729,N_7222);
or U8311 (N_8311,N_7385,N_6548);
or U8312 (N_8312,N_6592,N_7936);
and U8313 (N_8313,N_6905,N_6944);
or U8314 (N_8314,N_7378,N_6270);
nand U8315 (N_8315,N_6082,N_6867);
nor U8316 (N_8316,N_6764,N_6901);
nor U8317 (N_8317,N_7146,N_6754);
nor U8318 (N_8318,N_6165,N_7612);
and U8319 (N_8319,N_7457,N_6048);
nor U8320 (N_8320,N_7466,N_6879);
xnor U8321 (N_8321,N_6720,N_6376);
nand U8322 (N_8322,N_6738,N_7588);
nand U8323 (N_8323,N_7981,N_7407);
and U8324 (N_8324,N_7517,N_6030);
nor U8325 (N_8325,N_7368,N_6668);
nand U8326 (N_8326,N_7850,N_6672);
nand U8327 (N_8327,N_6387,N_7436);
and U8328 (N_8328,N_7331,N_7942);
and U8329 (N_8329,N_7069,N_7424);
nor U8330 (N_8330,N_6481,N_6662);
nand U8331 (N_8331,N_6492,N_7148);
nand U8332 (N_8332,N_6468,N_7583);
nor U8333 (N_8333,N_7770,N_6852);
nor U8334 (N_8334,N_7340,N_6199);
and U8335 (N_8335,N_6232,N_7498);
or U8336 (N_8336,N_6297,N_7752);
nand U8337 (N_8337,N_7986,N_6572);
and U8338 (N_8338,N_6318,N_6795);
and U8339 (N_8339,N_6154,N_7404);
nand U8340 (N_8340,N_6405,N_6759);
nor U8341 (N_8341,N_7879,N_7641);
nand U8342 (N_8342,N_6605,N_6006);
nor U8343 (N_8343,N_6130,N_7559);
or U8344 (N_8344,N_7545,N_7350);
or U8345 (N_8345,N_7851,N_6669);
nand U8346 (N_8346,N_7613,N_6735);
or U8347 (N_8347,N_6995,N_7205);
and U8348 (N_8348,N_7360,N_7504);
nor U8349 (N_8349,N_6857,N_7977);
or U8350 (N_8350,N_7655,N_6302);
and U8351 (N_8351,N_7357,N_7321);
nand U8352 (N_8352,N_6968,N_6870);
nor U8353 (N_8353,N_7373,N_6020);
and U8354 (N_8354,N_6659,N_7757);
nor U8355 (N_8355,N_7912,N_7375);
nand U8356 (N_8356,N_6431,N_7957);
xor U8357 (N_8357,N_6244,N_6914);
nor U8358 (N_8358,N_7564,N_6965);
and U8359 (N_8359,N_6336,N_7193);
nand U8360 (N_8360,N_7671,N_6057);
nor U8361 (N_8361,N_7992,N_7174);
xnor U8362 (N_8362,N_7003,N_6505);
nand U8363 (N_8363,N_6223,N_6454);
nor U8364 (N_8364,N_6575,N_7253);
or U8365 (N_8365,N_6219,N_6278);
and U8366 (N_8366,N_7393,N_7838);
and U8367 (N_8367,N_6753,N_6973);
nor U8368 (N_8368,N_7432,N_7000);
nor U8369 (N_8369,N_7211,N_7681);
or U8370 (N_8370,N_6460,N_7520);
nor U8371 (N_8371,N_6372,N_7204);
or U8372 (N_8372,N_6555,N_7079);
and U8373 (N_8373,N_7883,N_6305);
nor U8374 (N_8374,N_7852,N_7358);
nor U8375 (N_8375,N_6958,N_7537);
nor U8376 (N_8376,N_7651,N_7287);
or U8377 (N_8377,N_7813,N_7956);
nor U8378 (N_8378,N_6429,N_6413);
xor U8379 (N_8379,N_6956,N_7919);
nor U8380 (N_8380,N_6452,N_7270);
or U8381 (N_8381,N_7245,N_7251);
and U8382 (N_8382,N_6313,N_6072);
nand U8383 (N_8383,N_6549,N_6726);
nor U8384 (N_8384,N_7084,N_6625);
nand U8385 (N_8385,N_6122,N_6708);
and U8386 (N_8386,N_6690,N_7145);
or U8387 (N_8387,N_6897,N_6273);
or U8388 (N_8388,N_6111,N_6639);
and U8389 (N_8389,N_7688,N_6164);
xnor U8390 (N_8390,N_6010,N_7206);
nor U8391 (N_8391,N_7891,N_6211);
or U8392 (N_8392,N_6388,N_7169);
nor U8393 (N_8393,N_6546,N_7603);
or U8394 (N_8394,N_7764,N_7822);
or U8395 (N_8395,N_7422,N_6696);
or U8396 (N_8396,N_7344,N_7522);
nand U8397 (N_8397,N_6155,N_7090);
nor U8398 (N_8398,N_7322,N_6620);
and U8399 (N_8399,N_7625,N_6633);
nor U8400 (N_8400,N_6854,N_7748);
nor U8401 (N_8401,N_6711,N_6220);
or U8402 (N_8402,N_6833,N_6784);
nor U8403 (N_8403,N_7664,N_6820);
nand U8404 (N_8404,N_6295,N_6700);
nor U8405 (N_8405,N_7098,N_7536);
and U8406 (N_8406,N_6367,N_7675);
nor U8407 (N_8407,N_6810,N_7291);
and U8408 (N_8408,N_6420,N_7965);
and U8409 (N_8409,N_6576,N_6855);
or U8410 (N_8410,N_7351,N_6392);
nand U8411 (N_8411,N_7708,N_7785);
or U8412 (N_8412,N_7549,N_6882);
nand U8413 (N_8413,N_7309,N_7940);
nand U8414 (N_8414,N_7492,N_6422);
nand U8415 (N_8415,N_6892,N_6540);
or U8416 (N_8416,N_7826,N_7976);
or U8417 (N_8417,N_7615,N_7507);
nand U8418 (N_8418,N_6818,N_7349);
nand U8419 (N_8419,N_6777,N_6779);
xnor U8420 (N_8420,N_7198,N_7467);
nand U8421 (N_8421,N_6345,N_7894);
nand U8422 (N_8422,N_7587,N_7768);
nor U8423 (N_8423,N_7968,N_7718);
and U8424 (N_8424,N_7325,N_7265);
or U8425 (N_8425,N_7472,N_6423);
and U8426 (N_8426,N_7914,N_7260);
and U8427 (N_8427,N_7065,N_7338);
or U8428 (N_8428,N_6622,N_6150);
xor U8429 (N_8429,N_7283,N_7692);
or U8430 (N_8430,N_7580,N_6821);
or U8431 (N_8431,N_7445,N_7630);
nor U8432 (N_8432,N_6059,N_6182);
and U8433 (N_8433,N_6271,N_7043);
or U8434 (N_8434,N_7125,N_7412);
nand U8435 (N_8435,N_7743,N_7890);
nor U8436 (N_8436,N_6786,N_6582);
or U8437 (N_8437,N_6374,N_7660);
and U8438 (N_8438,N_7618,N_7243);
or U8439 (N_8439,N_7871,N_6347);
or U8440 (N_8440,N_6987,N_7599);
or U8441 (N_8441,N_7602,N_7454);
and U8442 (N_8442,N_7109,N_6996);
and U8443 (N_8443,N_7248,N_6362);
and U8444 (N_8444,N_6562,N_7901);
or U8445 (N_8445,N_6963,N_6515);
nand U8446 (N_8446,N_7134,N_7730);
or U8447 (N_8447,N_6483,N_7363);
and U8448 (N_8448,N_7074,N_7082);
nor U8449 (N_8449,N_6418,N_7546);
or U8450 (N_8450,N_7230,N_6075);
nand U8451 (N_8451,N_7721,N_7343);
or U8452 (N_8452,N_7299,N_6536);
nor U8453 (N_8453,N_6774,N_7684);
or U8454 (N_8454,N_7329,N_7433);
xor U8455 (N_8455,N_7926,N_6252);
nand U8456 (N_8456,N_7880,N_6149);
nand U8457 (N_8457,N_6558,N_6722);
or U8458 (N_8458,N_6495,N_7509);
nand U8459 (N_8459,N_6365,N_6262);
nand U8460 (N_8460,N_6778,N_7557);
xor U8461 (N_8461,N_7036,N_7676);
and U8462 (N_8462,N_6415,N_7276);
and U8463 (N_8463,N_6680,N_6275);
nand U8464 (N_8464,N_6248,N_7455);
xor U8465 (N_8465,N_7479,N_7220);
or U8466 (N_8466,N_7228,N_7788);
nor U8467 (N_8467,N_6246,N_7224);
or U8468 (N_8468,N_6301,N_7858);
or U8469 (N_8469,N_7941,N_7167);
nand U8470 (N_8470,N_7562,N_6841);
xor U8471 (N_8471,N_6463,N_7814);
nor U8472 (N_8472,N_7166,N_7020);
nor U8473 (N_8473,N_6547,N_7915);
nand U8474 (N_8474,N_7451,N_6393);
or U8475 (N_8475,N_7301,N_7586);
or U8476 (N_8476,N_7050,N_6698);
and U8477 (N_8477,N_6196,N_7425);
xnor U8478 (N_8478,N_7053,N_7129);
or U8479 (N_8479,N_6078,N_7284);
and U8480 (N_8480,N_6120,N_6496);
nand U8481 (N_8481,N_7341,N_6655);
nand U8482 (N_8482,N_6013,N_7584);
nand U8483 (N_8483,N_6008,N_7548);
or U8484 (N_8484,N_7707,N_6071);
or U8485 (N_8485,N_7414,N_7332);
nor U8486 (N_8486,N_6521,N_6688);
nor U8487 (N_8487,N_7028,N_7196);
nor U8488 (N_8488,N_6397,N_6061);
nand U8489 (N_8489,N_6126,N_7018);
nand U8490 (N_8490,N_7802,N_7990);
and U8491 (N_8491,N_7930,N_7872);
or U8492 (N_8492,N_7392,N_7917);
or U8493 (N_8493,N_6398,N_6402);
nand U8494 (N_8494,N_6081,N_7995);
and U8495 (N_8495,N_6309,N_6844);
nor U8496 (N_8496,N_6604,N_7272);
or U8497 (N_8497,N_6719,N_6745);
and U8498 (N_8498,N_6563,N_6291);
and U8499 (N_8499,N_6666,N_7781);
nand U8500 (N_8500,N_6200,N_6482);
nand U8501 (N_8501,N_6611,N_7581);
and U8502 (N_8502,N_6535,N_6467);
nand U8503 (N_8503,N_6848,N_6298);
xnor U8504 (N_8504,N_7223,N_7945);
or U8505 (N_8505,N_6524,N_6029);
and U8506 (N_8506,N_6475,N_7448);
nand U8507 (N_8507,N_6350,N_7875);
nor U8508 (N_8508,N_6241,N_6198);
and U8509 (N_8509,N_6245,N_6472);
nand U8510 (N_8510,N_6300,N_7142);
nand U8511 (N_8511,N_6585,N_6893);
or U8512 (N_8512,N_7775,N_7809);
nand U8513 (N_8513,N_7298,N_7989);
or U8514 (N_8514,N_6871,N_6950);
nand U8515 (N_8515,N_6340,N_6218);
nand U8516 (N_8516,N_7111,N_6663);
nand U8517 (N_8517,N_6624,N_6646);
and U8518 (N_8518,N_6478,N_6915);
nor U8519 (N_8519,N_6657,N_7807);
and U8520 (N_8520,N_6681,N_6316);
and U8521 (N_8521,N_7091,N_6408);
and U8522 (N_8522,N_6028,N_7460);
nor U8523 (N_8523,N_6926,N_6022);
nor U8524 (N_8524,N_6816,N_6579);
nor U8525 (N_8525,N_7443,N_7408);
nand U8526 (N_8526,N_7758,N_6884);
nor U8527 (N_8527,N_7062,N_7369);
nor U8528 (N_8528,N_6240,N_7197);
or U8529 (N_8529,N_7077,N_6632);
or U8530 (N_8530,N_7415,N_7027);
nor U8531 (N_8531,N_6294,N_7849);
and U8532 (N_8532,N_7573,N_7994);
or U8533 (N_8533,N_6055,N_6208);
xnor U8534 (N_8534,N_6746,N_6811);
or U8535 (N_8535,N_6128,N_6175);
xor U8536 (N_8536,N_6895,N_6717);
nor U8537 (N_8537,N_6464,N_6621);
nor U8538 (N_8538,N_7710,N_6718);
nand U8539 (N_8539,N_7939,N_7727);
and U8540 (N_8540,N_7798,N_7538);
and U8541 (N_8541,N_7999,N_6991);
and U8542 (N_8542,N_7857,N_7022);
or U8543 (N_8543,N_7459,N_6266);
nand U8544 (N_8544,N_6485,N_6961);
nand U8545 (N_8545,N_7399,N_6962);
nand U8546 (N_8546,N_6186,N_6449);
nand U8547 (N_8547,N_6501,N_6957);
and U8548 (N_8548,N_7828,N_7262);
nor U8549 (N_8549,N_7247,N_6836);
or U8550 (N_8550,N_6442,N_6916);
nand U8551 (N_8551,N_7881,N_7640);
nor U8552 (N_8552,N_7431,N_7689);
and U8553 (N_8553,N_7845,N_6982);
nand U8554 (N_8554,N_6238,N_6712);
and U8555 (N_8555,N_6891,N_7390);
nor U8556 (N_8556,N_7489,N_7691);
or U8557 (N_8557,N_6026,N_6588);
nor U8558 (N_8558,N_7486,N_6790);
or U8559 (N_8559,N_6993,N_6097);
nand U8560 (N_8560,N_6192,N_7706);
nand U8561 (N_8561,N_6396,N_6203);
and U8562 (N_8562,N_7561,N_7842);
nor U8563 (N_8563,N_6994,N_7316);
nand U8564 (N_8564,N_6337,N_6890);
and U8565 (N_8565,N_6685,N_6990);
or U8566 (N_8566,N_7190,N_7308);
nand U8567 (N_8567,N_7786,N_7830);
nor U8568 (N_8568,N_7801,N_7184);
nand U8569 (N_8569,N_6607,N_7453);
nand U8570 (N_8570,N_7591,N_6785);
and U8571 (N_8571,N_7993,N_6038);
or U8572 (N_8572,N_7201,N_6487);
nand U8573 (N_8573,N_6106,N_7086);
and U8574 (N_8574,N_7805,N_7149);
nand U8575 (N_8575,N_7130,N_7132);
nor U8576 (N_8576,N_6967,N_7521);
and U8577 (N_8577,N_7153,N_6939);
nand U8578 (N_8578,N_7574,N_6692);
xor U8579 (N_8579,N_7026,N_7978);
and U8580 (N_8580,N_7906,N_7661);
nor U8581 (N_8581,N_6179,N_6789);
nor U8582 (N_8582,N_6869,N_7001);
nor U8583 (N_8583,N_7799,N_7535);
and U8584 (N_8584,N_7899,N_6473);
xor U8585 (N_8585,N_6304,N_7934);
nor U8586 (N_8586,N_6368,N_7566);
nand U8587 (N_8587,N_7946,N_6606);
or U8588 (N_8588,N_6201,N_7123);
or U8589 (N_8589,N_7922,N_7624);
nand U8590 (N_8590,N_6574,N_7353);
or U8591 (N_8591,N_6888,N_7774);
xor U8592 (N_8592,N_7177,N_7967);
nand U8593 (N_8593,N_6834,N_6088);
nand U8594 (N_8594,N_7513,N_6108);
nand U8595 (N_8595,N_7044,N_6205);
and U8596 (N_8596,N_7355,N_6500);
or U8597 (N_8597,N_6876,N_7333);
and U8598 (N_8598,N_7024,N_6023);
or U8599 (N_8599,N_7317,N_6283);
nor U8600 (N_8600,N_7374,N_7107);
and U8601 (N_8601,N_6419,N_6776);
and U8602 (N_8602,N_6556,N_7629);
or U8603 (N_8603,N_6650,N_7532);
nand U8604 (N_8604,N_6021,N_6566);
and U8605 (N_8605,N_6212,N_6162);
or U8606 (N_8606,N_7231,N_6725);
or U8607 (N_8607,N_7873,N_7568);
or U8608 (N_8608,N_6058,N_7192);
nor U8609 (N_8609,N_6289,N_6728);
and U8610 (N_8610,N_7154,N_7310);
xor U8611 (N_8611,N_6878,N_6969);
nor U8612 (N_8612,N_6924,N_7608);
nor U8613 (N_8613,N_7089,N_6268);
nand U8614 (N_8614,N_7085,N_7737);
nand U8615 (N_8615,N_6178,N_6578);
and U8616 (N_8616,N_7403,N_6471);
or U8617 (N_8617,N_6839,N_7242);
xor U8618 (N_8618,N_7185,N_7844);
and U8619 (N_8619,N_6999,N_6596);
and U8620 (N_8620,N_6953,N_7059);
nor U8621 (N_8621,N_6497,N_7409);
xnor U8622 (N_8622,N_7429,N_6103);
nand U8623 (N_8623,N_7136,N_7210);
nand U8624 (N_8624,N_6617,N_6716);
and U8625 (N_8625,N_6949,N_7682);
nor U8626 (N_8626,N_7542,N_7696);
or U8627 (N_8627,N_6335,N_7592);
nor U8628 (N_8628,N_7563,N_6671);
nor U8629 (N_8629,N_6737,N_6594);
nand U8630 (N_8630,N_7824,N_6352);
and U8631 (N_8631,N_7496,N_7182);
or U8632 (N_8632,N_6264,N_6090);
nor U8633 (N_8633,N_7463,N_6197);
and U8634 (N_8634,N_7178,N_7617);
and U8635 (N_8635,N_6132,N_6981);
or U8636 (N_8636,N_6257,N_7339);
or U8637 (N_8637,N_7904,N_7306);
and U8638 (N_8638,N_7678,N_6817);
or U8639 (N_8639,N_7263,N_6955);
and U8640 (N_8640,N_6288,N_6185);
nor U8641 (N_8641,N_7221,N_7874);
nor U8642 (N_8642,N_7047,N_6609);
xnor U8643 (N_8643,N_7139,N_7236);
nor U8644 (N_8644,N_6874,N_6656);
nand U8645 (N_8645,N_6308,N_6156);
or U8646 (N_8646,N_6435,N_7045);
and U8647 (N_8647,N_7503,N_6031);
nand U8648 (N_8648,N_6567,N_6121);
and U8649 (N_8649,N_7241,N_6512);
and U8650 (N_8650,N_7328,N_7731);
or U8651 (N_8651,N_7162,N_7778);
and U8652 (N_8652,N_6002,N_6433);
and U8653 (N_8653,N_7234,N_7411);
and U8654 (N_8654,N_7029,N_6144);
nand U8655 (N_8655,N_7869,N_6921);
nand U8656 (N_8656,N_7359,N_6364);
nor U8657 (N_8657,N_6710,N_7997);
nand U8658 (N_8658,N_6322,N_6009);
or U8659 (N_8659,N_7037,N_7469);
or U8660 (N_8660,N_7356,N_6222);
and U8661 (N_8661,N_7973,N_6912);
xor U8662 (N_8662,N_6049,N_6209);
nor U8663 (N_8663,N_6910,N_7386);
or U8664 (N_8664,N_6084,N_6947);
or U8665 (N_8665,N_7110,N_6826);
nand U8666 (N_8666,N_7717,N_7127);
nand U8667 (N_8667,N_7554,N_7742);
nor U8668 (N_8668,N_6331,N_6135);
nor U8669 (N_8669,N_7410,N_6098);
and U8670 (N_8670,N_6074,N_7013);
or U8671 (N_8671,N_7649,N_7634);
nand U8672 (N_8672,N_6601,N_7864);
and U8673 (N_8673,N_7784,N_7987);
nor U8674 (N_8674,N_6306,N_6312);
nor U8675 (N_8675,N_7846,N_6166);
or U8676 (N_8676,N_6432,N_6004);
and U8677 (N_8677,N_7296,N_6382);
or U8678 (N_8678,N_7441,N_6045);
or U8679 (N_8679,N_6736,N_7092);
and U8680 (N_8680,N_7400,N_6523);
nand U8681 (N_8681,N_7960,N_6480);
and U8682 (N_8682,N_7847,N_6537);
nor U8683 (N_8683,N_7131,N_7318);
and U8684 (N_8684,N_6943,N_7482);
nor U8685 (N_8685,N_7620,N_6152);
and U8686 (N_8686,N_7589,N_7543);
nand U8687 (N_8687,N_6853,N_7442);
nor U8688 (N_8688,N_6377,N_7578);
and U8689 (N_8689,N_7112,N_7762);
nor U8690 (N_8690,N_7863,N_7848);
nand U8691 (N_8691,N_7458,N_7650);
xnor U8692 (N_8692,N_7658,N_7832);
nor U8693 (N_8693,N_7621,N_7765);
nand U8694 (N_8694,N_7744,N_7277);
and U8695 (N_8695,N_6705,N_7126);
nand U8696 (N_8696,N_6545,N_6864);
and U8697 (N_8697,N_7066,N_7070);
nand U8698 (N_8698,N_6846,N_6494);
and U8699 (N_8699,N_6889,N_6411);
and U8700 (N_8700,N_7579,N_7170);
nand U8701 (N_8701,N_7715,N_7389);
nand U8702 (N_8702,N_7672,N_7868);
nor U8703 (N_8703,N_6391,N_6850);
and U8704 (N_8704,N_6825,N_6315);
or U8705 (N_8705,N_7783,N_6519);
nor U8706 (N_8706,N_6014,N_7837);
nor U8707 (N_8707,N_7475,N_7021);
and U8708 (N_8708,N_6314,N_7925);
and U8709 (N_8709,N_7645,N_7980);
and U8710 (N_8710,N_7703,N_7860);
nand U8711 (N_8711,N_7175,N_7006);
nand U8712 (N_8712,N_6824,N_6756);
or U8713 (N_8713,N_6851,N_7238);
nor U8714 (N_8714,N_7215,N_7140);
nand U8715 (N_8715,N_6067,N_6760);
or U8716 (N_8716,N_7345,N_7447);
or U8717 (N_8717,N_7372,N_7285);
and U8718 (N_8718,N_6065,N_7511);
xnor U8719 (N_8719,N_7779,N_6105);
nand U8720 (N_8720,N_6358,N_6256);
and U8721 (N_8721,N_6804,N_7165);
and U8722 (N_8722,N_7720,N_6453);
xnor U8723 (N_8723,N_6699,N_7598);
and U8724 (N_8724,N_6064,N_7896);
nor U8725 (N_8725,N_7049,N_7656);
nand U8726 (N_8726,N_7763,N_6561);
nand U8727 (N_8727,N_7073,N_7152);
nand U8728 (N_8728,N_6349,N_6543);
nor U8729 (N_8729,N_6724,N_7971);
nor U8730 (N_8730,N_6258,N_7342);
nor U8731 (N_8731,N_6748,N_6842);
nor U8732 (N_8732,N_6989,N_6885);
nor U8733 (N_8733,N_6911,N_6954);
and U8734 (N_8734,N_6769,N_7268);
nor U8735 (N_8735,N_7275,N_7526);
and U8736 (N_8736,N_7885,N_6228);
and U8737 (N_8737,N_7252,N_7364);
and U8738 (N_8738,N_6339,N_7151);
and U8739 (N_8739,N_6428,N_6019);
and U8740 (N_8740,N_7865,N_6593);
and U8741 (N_8741,N_6363,N_7729);
xor U8742 (N_8742,N_7892,N_6317);
nor U8743 (N_8743,N_7280,N_6739);
nand U8744 (N_8744,N_6887,N_6430);
nand U8745 (N_8745,N_7439,N_6046);
and U8746 (N_8746,N_6522,N_6188);
nor U8747 (N_8747,N_7135,N_6938);
nor U8748 (N_8748,N_7269,N_6375);
nor U8749 (N_8749,N_7815,N_6490);
or U8750 (N_8750,N_6683,N_6093);
nand U8751 (N_8751,N_7383,N_7491);
nand U8752 (N_8752,N_7909,N_6899);
or U8753 (N_8753,N_6394,N_7379);
and U8754 (N_8754,N_7033,N_6740);
or U8755 (N_8755,N_7124,N_7095);
xor U8756 (N_8756,N_6510,N_7257);
or U8757 (N_8757,N_7771,N_6390);
nor U8758 (N_8758,N_7795,N_6615);
nor U8759 (N_8759,N_6044,N_7628);
or U8760 (N_8760,N_6603,N_6450);
nand U8761 (N_8761,N_7147,N_6076);
nand U8762 (N_8762,N_6571,N_6033);
nor U8763 (N_8763,N_7005,N_6702);
and U8764 (N_8764,N_6334,N_7745);
nor U8765 (N_8765,N_6730,N_7144);
xor U8766 (N_8766,N_7810,N_7623);
nand U8767 (N_8767,N_7900,N_7179);
nand U8768 (N_8768,N_7637,N_7430);
nor U8769 (N_8769,N_6514,N_7693);
or U8770 (N_8770,N_6770,N_7481);
nand U8771 (N_8771,N_6626,N_6723);
nor U8772 (N_8772,N_6701,N_6800);
nor U8773 (N_8773,N_6664,N_6843);
or U8774 (N_8774,N_7607,N_7010);
nand U8775 (N_8775,N_7217,N_7959);
nor U8776 (N_8776,N_7314,N_7121);
or U8777 (N_8777,N_7749,N_7638);
nor U8778 (N_8778,N_7188,N_7594);
or U8779 (N_8779,N_6658,N_7690);
and U8780 (N_8780,N_7138,N_7952);
xnor U8781 (N_8781,N_7932,N_6050);
xnor U8782 (N_8782,N_7240,N_7311);
or U8783 (N_8783,N_7500,N_7388);
nand U8784 (N_8784,N_6110,N_7117);
or U8785 (N_8785,N_6104,N_6369);
or U8786 (N_8786,N_6610,N_6933);
nand U8787 (N_8787,N_7988,N_6827);
and U8788 (N_8788,N_7714,N_7547);
nor U8789 (N_8789,N_6984,N_6455);
or U8790 (N_8790,N_6404,N_7213);
nor U8791 (N_8791,N_7985,N_6434);
nor U8792 (N_8792,N_7099,N_7751);
or U8793 (N_8793,N_6489,N_7539);
or U8794 (N_8794,N_6118,N_7923);
or U8795 (N_8795,N_7733,N_7654);
or U8796 (N_8796,N_6079,N_7515);
and U8797 (N_8797,N_7264,N_6504);
nand U8798 (N_8798,N_7812,N_7015);
nor U8799 (N_8799,N_7734,N_7913);
nor U8800 (N_8800,N_7324,N_6370);
or U8801 (N_8801,N_6613,N_6616);
or U8802 (N_8802,N_7601,N_7843);
nor U8803 (N_8803,N_6024,N_6066);
nand U8804 (N_8804,N_6799,N_6409);
nor U8805 (N_8805,N_7657,N_7969);
nand U8806 (N_8806,N_7541,N_7643);
and U8807 (N_8807,N_7413,N_6584);
nor U8808 (N_8808,N_6007,N_7862);
nor U8809 (N_8809,N_7958,N_7336);
and U8810 (N_8810,N_6860,N_6794);
nand U8811 (N_8811,N_6095,N_7261);
or U8812 (N_8812,N_6233,N_6703);
and U8813 (N_8813,N_6403,N_6823);
and U8814 (N_8814,N_6069,N_6629);
nor U8815 (N_8815,N_6272,N_7687);
nor U8816 (N_8816,N_7685,N_7141);
xor U8817 (N_8817,N_7571,N_6299);
nand U8818 (N_8818,N_7518,N_6160);
nor U8819 (N_8819,N_7396,N_7983);
or U8820 (N_8820,N_7267,N_6997);
or U8821 (N_8821,N_6225,N_7484);
and U8822 (N_8822,N_7417,N_7818);
or U8823 (N_8823,N_7506,N_6959);
nor U8824 (N_8824,N_7218,N_7679);
nand U8825 (N_8825,N_6011,N_7761);
and U8826 (N_8826,N_6707,N_7792);
nand U8827 (N_8827,N_6125,N_7648);
or U8828 (N_8828,N_6005,N_6161);
xnor U8829 (N_8829,N_7064,N_6063);
xnor U8830 (N_8830,N_6003,N_6682);
and U8831 (N_8831,N_6457,N_6027);
nor U8832 (N_8832,N_6900,N_7738);
or U8833 (N_8833,N_6360,N_7780);
nand U8834 (N_8834,N_7604,N_6385);
nor U8835 (N_8835,N_6123,N_7227);
or U8836 (N_8836,N_6169,N_6476);
nand U8837 (N_8837,N_7782,N_6559);
nor U8838 (N_8838,N_6775,N_6148);
xor U8839 (N_8839,N_6653,N_6303);
xnor U8840 (N_8840,N_6644,N_6630);
nor U8841 (N_8841,N_7093,N_7670);
nor U8842 (N_8842,N_7840,N_7487);
and U8843 (N_8843,N_7741,N_6597);
xor U8844 (N_8844,N_6040,N_7235);
and U8845 (N_8845,N_6976,N_7380);
and U8846 (N_8846,N_7116,N_6637);
and U8847 (N_8847,N_7790,N_6025);
and U8848 (N_8848,N_6880,N_7327);
xnor U8849 (N_8849,N_6966,N_7944);
nand U8850 (N_8850,N_7294,N_6641);
nor U8851 (N_8851,N_7787,N_7600);
nand U8852 (N_8852,N_6443,N_6647);
or U8853 (N_8853,N_6845,N_7700);
nor U8854 (N_8854,N_7606,N_6333);
or U8855 (N_8855,N_7416,N_7002);
nor U8856 (N_8856,N_7470,N_7051);
nor U8857 (N_8857,N_6410,N_6837);
xor U8858 (N_8858,N_7510,N_7626);
nor U8859 (N_8859,N_6060,N_6357);
and U8860 (N_8860,N_6908,N_7488);
and U8861 (N_8861,N_7450,N_7158);
xor U8862 (N_8862,N_6498,N_6056);
nor U8863 (N_8863,N_7176,N_7381);
nor U8864 (N_8864,N_6986,N_6012);
and U8865 (N_8865,N_6269,N_6835);
nand U8866 (N_8866,N_6159,N_6551);
or U8867 (N_8867,N_6743,N_7189);
nand U8868 (N_8868,N_6493,N_6204);
or U8869 (N_8869,N_7505,N_7870);
or U8870 (N_8870,N_7972,N_6787);
nand U8871 (N_8871,N_7528,N_6102);
nor U8872 (N_8872,N_6861,N_6170);
nor U8873 (N_8873,N_6037,N_6224);
xor U8874 (N_8874,N_7191,N_6530);
and U8875 (N_8875,N_6757,N_7747);
or U8876 (N_8876,N_6324,N_7195);
or U8877 (N_8877,N_7402,N_6438);
or U8878 (N_8878,N_7258,N_7907);
nor U8879 (N_8879,N_6146,N_7083);
and U8880 (N_8880,N_7501,N_6577);
nand U8881 (N_8881,N_7829,N_7530);
or U8882 (N_8882,N_7382,N_6172);
xnor U8883 (N_8883,N_6715,N_7595);
or U8884 (N_8884,N_6948,N_6096);
nor U8885 (N_8885,N_6907,N_7237);
and U8886 (N_8886,N_7948,N_6832);
nand U8887 (N_8887,N_6259,N_6424);
xor U8888 (N_8888,N_6342,N_7288);
or U8889 (N_8889,N_6539,N_6053);
nand U8890 (N_8890,N_6016,N_6750);
nand U8891 (N_8891,N_6677,N_7622);
nor U8892 (N_8892,N_6985,N_7161);
nor U8893 (N_8893,N_6094,N_6325);
nor U8894 (N_8894,N_6235,N_7048);
nand U8895 (N_8895,N_7017,N_7974);
or U8896 (N_8896,N_6813,N_7046);
and U8897 (N_8897,N_7831,N_7199);
or U8898 (N_8898,N_7081,N_6922);
nor U8899 (N_8899,N_7225,N_7886);
nand U8900 (N_8900,N_6444,N_6731);
and U8901 (N_8901,N_6327,N_7055);
nand U8902 (N_8902,N_7512,N_6642);
nand U8903 (N_8903,N_6970,N_6286);
nor U8904 (N_8904,N_7464,N_7597);
nand U8905 (N_8905,N_6872,N_6886);
and U8906 (N_8906,N_7039,N_7437);
nand U8907 (N_8907,N_7307,N_7434);
or U8908 (N_8908,N_7438,N_6866);
nand U8909 (N_8909,N_6173,N_7569);
nor U8910 (N_8910,N_7593,N_6909);
and U8911 (N_8911,N_7295,N_7100);
or U8912 (N_8912,N_6344,N_6488);
nand U8913 (N_8913,N_6217,N_6176);
and U8914 (N_8914,N_6917,N_6906);
nor U8915 (N_8915,N_7278,N_6665);
nand U8916 (N_8916,N_7105,N_6691);
and U8917 (N_8917,N_6940,N_7984);
xor U8918 (N_8918,N_7502,N_6282);
or U8919 (N_8919,N_7884,N_6459);
and U8920 (N_8920,N_6687,N_7928);
xnor U8921 (N_8921,N_7371,N_6070);
nand U8922 (N_8922,N_7631,N_6819);
or U8923 (N_8923,N_6829,N_6190);
and U8924 (N_8924,N_7644,N_6417);
nor U8925 (N_8925,N_7711,N_7905);
nand U8926 (N_8926,N_7666,N_6927);
nor U8927 (N_8927,N_6310,N_6971);
nand U8928 (N_8928,N_7305,N_6319);
or U8929 (N_8929,N_7674,N_7525);
or U8930 (N_8930,N_6992,N_6263);
xor U8931 (N_8931,N_7680,N_7173);
nor U8932 (N_8932,N_7471,N_7330);
and U8933 (N_8933,N_6127,N_6640);
xor U8934 (N_8934,N_6477,N_7271);
xor U8935 (N_8935,N_7753,N_7108);
or U8936 (N_8936,N_7804,N_6042);
nand U8937 (N_8937,N_6407,N_7495);
or U8938 (N_8938,N_6552,N_6399);
nand U8939 (N_8939,N_7833,N_6277);
and U8940 (N_8940,N_7061,N_7067);
and U8941 (N_8941,N_6532,N_7823);
nand U8942 (N_8942,N_6793,N_7087);
or U8943 (N_8943,N_6034,N_6975);
and U8944 (N_8944,N_6541,N_6416);
nor U8945 (N_8945,N_7384,N_6503);
and U8946 (N_8946,N_7669,N_6230);
or U8947 (N_8947,N_6598,N_6163);
nor U8948 (N_8948,N_7303,N_7497);
nand U8949 (N_8949,N_6797,N_7150);
and U8950 (N_8950,N_6215,N_6553);
nor U8951 (N_8951,N_6627,N_6822);
or U8952 (N_8952,N_7719,N_7529);
or U8953 (N_8953,N_7366,N_7452);
nand U8954 (N_8954,N_6226,N_7519);
nor U8955 (N_8955,N_6727,N_7951);
or U8956 (N_8956,N_7732,N_6119);
nor U8957 (N_8957,N_7157,N_7035);
and U8958 (N_8958,N_7632,N_6951);
and U8959 (N_8959,N_7354,N_6181);
nor U8960 (N_8960,N_6602,N_6187);
nand U8961 (N_8961,N_7019,N_6051);
nand U8962 (N_8962,N_6608,N_7155);
or U8963 (N_8963,N_7635,N_6041);
and U8964 (N_8964,N_6538,N_6062);
nor U8965 (N_8965,N_7273,N_7979);
xor U8966 (N_8966,N_6755,N_6448);
or U8967 (N_8967,N_6400,N_6960);
and U8968 (N_8968,N_6054,N_6107);
nor U8969 (N_8969,N_6371,N_6988);
nand U8970 (N_8970,N_6346,N_6139);
xor U8971 (N_8971,N_7839,N_7639);
nand U8972 (N_8972,N_6581,N_6171);
or U8973 (N_8973,N_6858,N_6654);
and U8974 (N_8974,N_7163,N_6099);
xnor U8975 (N_8975,N_6918,N_6353);
nand U8976 (N_8976,N_7226,N_6877);
nand U8977 (N_8977,N_6329,N_7611);
nor U8978 (N_8978,N_7963,N_6838);
nand U8979 (N_8979,N_6945,N_7723);
xnor U8980 (N_8980,N_7791,N_6694);
and U8981 (N_8981,N_6964,N_6290);
nor U8982 (N_8982,N_7686,N_7012);
and U8983 (N_8983,N_6001,N_6469);
nand U8984 (N_8984,N_6250,N_7911);
or U8985 (N_8985,N_7553,N_6137);
nor U8986 (N_8986,N_7426,N_6628);
nor U8987 (N_8987,N_7636,N_7797);
and U8988 (N_8988,N_7523,N_6649);
xor U8989 (N_8989,N_6528,N_6814);
and U8990 (N_8990,N_7480,N_7207);
and U8991 (N_8991,N_7895,N_6080);
or U8992 (N_8992,N_6881,N_6440);
and U8993 (N_8993,N_6618,N_6210);
or U8994 (N_8994,N_6296,N_6117);
nor U8995 (N_8995,N_7289,N_7465);
or U8996 (N_8996,N_7527,N_7397);
nand U8997 (N_8997,N_6191,N_7935);
nand U8998 (N_8998,N_6032,N_7101);
nand U8999 (N_8999,N_6733,N_6281);
and U9000 (N_9000,N_7574,N_6176);
or U9001 (N_9001,N_6913,N_6345);
or U9002 (N_9002,N_7069,N_7446);
and U9003 (N_9003,N_7629,N_6875);
nor U9004 (N_9004,N_7869,N_7372);
nor U9005 (N_9005,N_6209,N_7292);
or U9006 (N_9006,N_7477,N_7067);
nand U9007 (N_9007,N_6782,N_7716);
or U9008 (N_9008,N_6268,N_6105);
and U9009 (N_9009,N_7237,N_7944);
nor U9010 (N_9010,N_6758,N_6014);
nor U9011 (N_9011,N_7758,N_6287);
and U9012 (N_9012,N_6433,N_6979);
and U9013 (N_9013,N_6806,N_7895);
nor U9014 (N_9014,N_7633,N_6731);
nor U9015 (N_9015,N_7025,N_7358);
nor U9016 (N_9016,N_7187,N_6461);
xnor U9017 (N_9017,N_6819,N_7107);
and U9018 (N_9018,N_6695,N_6744);
or U9019 (N_9019,N_7721,N_6505);
nor U9020 (N_9020,N_7515,N_7792);
or U9021 (N_9021,N_7065,N_6891);
nor U9022 (N_9022,N_6387,N_7196);
or U9023 (N_9023,N_6275,N_7264);
or U9024 (N_9024,N_7013,N_6530);
nor U9025 (N_9025,N_7234,N_7843);
or U9026 (N_9026,N_7953,N_7876);
nor U9027 (N_9027,N_7111,N_7983);
nor U9028 (N_9028,N_6923,N_7760);
xnor U9029 (N_9029,N_6165,N_6948);
nor U9030 (N_9030,N_7112,N_6910);
or U9031 (N_9031,N_7699,N_7629);
or U9032 (N_9032,N_7712,N_7121);
xor U9033 (N_9033,N_7746,N_6071);
and U9034 (N_9034,N_6141,N_6378);
nor U9035 (N_9035,N_6595,N_6892);
nor U9036 (N_9036,N_6765,N_6340);
and U9037 (N_9037,N_6619,N_7840);
nand U9038 (N_9038,N_6854,N_6298);
and U9039 (N_9039,N_6541,N_7303);
nor U9040 (N_9040,N_7902,N_6979);
and U9041 (N_9041,N_7497,N_6140);
and U9042 (N_9042,N_7146,N_7317);
nand U9043 (N_9043,N_7657,N_7048);
and U9044 (N_9044,N_7774,N_7128);
xnor U9045 (N_9045,N_6723,N_7124);
nand U9046 (N_9046,N_6792,N_7683);
xor U9047 (N_9047,N_6410,N_7053);
or U9048 (N_9048,N_6846,N_7997);
xnor U9049 (N_9049,N_7140,N_6699);
or U9050 (N_9050,N_6852,N_7019);
and U9051 (N_9051,N_6216,N_6686);
or U9052 (N_9052,N_7296,N_6207);
or U9053 (N_9053,N_6153,N_6512);
nor U9054 (N_9054,N_7965,N_6515);
nor U9055 (N_9055,N_6737,N_7080);
and U9056 (N_9056,N_7603,N_6855);
and U9057 (N_9057,N_6837,N_7989);
or U9058 (N_9058,N_6597,N_6208);
xnor U9059 (N_9059,N_7751,N_6298);
or U9060 (N_9060,N_7951,N_7880);
or U9061 (N_9061,N_6926,N_7015);
and U9062 (N_9062,N_6045,N_7417);
nand U9063 (N_9063,N_6858,N_7643);
and U9064 (N_9064,N_7624,N_6957);
nand U9065 (N_9065,N_7842,N_6453);
or U9066 (N_9066,N_7714,N_7899);
and U9067 (N_9067,N_7846,N_6777);
or U9068 (N_9068,N_6586,N_7914);
or U9069 (N_9069,N_6751,N_7975);
nor U9070 (N_9070,N_6219,N_7169);
or U9071 (N_9071,N_6510,N_6972);
nand U9072 (N_9072,N_7635,N_6836);
xor U9073 (N_9073,N_7370,N_6233);
or U9074 (N_9074,N_7236,N_6496);
nor U9075 (N_9075,N_6711,N_6539);
nand U9076 (N_9076,N_7171,N_7146);
nand U9077 (N_9077,N_6566,N_6748);
nand U9078 (N_9078,N_6784,N_6603);
nor U9079 (N_9079,N_7833,N_7705);
nand U9080 (N_9080,N_6401,N_7520);
nand U9081 (N_9081,N_7602,N_6435);
nor U9082 (N_9082,N_6104,N_7733);
xnor U9083 (N_9083,N_7519,N_7922);
nor U9084 (N_9084,N_6742,N_6939);
nor U9085 (N_9085,N_6032,N_7436);
or U9086 (N_9086,N_6232,N_7750);
nand U9087 (N_9087,N_7311,N_7607);
and U9088 (N_9088,N_7719,N_7777);
nand U9089 (N_9089,N_7092,N_7743);
nor U9090 (N_9090,N_7844,N_7653);
or U9091 (N_9091,N_7567,N_6425);
nor U9092 (N_9092,N_6071,N_7425);
and U9093 (N_9093,N_6184,N_6151);
and U9094 (N_9094,N_7420,N_6609);
or U9095 (N_9095,N_7794,N_6989);
or U9096 (N_9096,N_7002,N_6780);
or U9097 (N_9097,N_6344,N_6396);
nand U9098 (N_9098,N_6428,N_7408);
nor U9099 (N_9099,N_6990,N_6213);
nor U9100 (N_9100,N_6864,N_7999);
nor U9101 (N_9101,N_6851,N_7735);
and U9102 (N_9102,N_6922,N_7603);
or U9103 (N_9103,N_6425,N_6772);
or U9104 (N_9104,N_7465,N_6962);
xnor U9105 (N_9105,N_7291,N_7697);
or U9106 (N_9106,N_7896,N_6115);
or U9107 (N_9107,N_7543,N_7352);
nand U9108 (N_9108,N_6508,N_6182);
nor U9109 (N_9109,N_6523,N_7403);
nor U9110 (N_9110,N_6145,N_7524);
and U9111 (N_9111,N_7058,N_7217);
nor U9112 (N_9112,N_6447,N_7727);
nand U9113 (N_9113,N_6511,N_6815);
xnor U9114 (N_9114,N_6077,N_7994);
nor U9115 (N_9115,N_6746,N_7848);
or U9116 (N_9116,N_6929,N_7101);
xnor U9117 (N_9117,N_7395,N_7453);
and U9118 (N_9118,N_6750,N_7944);
nand U9119 (N_9119,N_7656,N_6531);
or U9120 (N_9120,N_6177,N_7133);
nand U9121 (N_9121,N_7429,N_6952);
nor U9122 (N_9122,N_7104,N_6358);
nand U9123 (N_9123,N_7078,N_6213);
nand U9124 (N_9124,N_7834,N_6288);
xnor U9125 (N_9125,N_6841,N_7637);
or U9126 (N_9126,N_7251,N_6878);
xnor U9127 (N_9127,N_6430,N_6690);
or U9128 (N_9128,N_6675,N_7617);
nand U9129 (N_9129,N_7866,N_7587);
or U9130 (N_9130,N_6470,N_6864);
and U9131 (N_9131,N_7727,N_7450);
xor U9132 (N_9132,N_7135,N_7413);
nand U9133 (N_9133,N_7636,N_7159);
nand U9134 (N_9134,N_7615,N_6133);
nand U9135 (N_9135,N_7607,N_6821);
nand U9136 (N_9136,N_7091,N_7803);
or U9137 (N_9137,N_6301,N_7409);
nor U9138 (N_9138,N_6931,N_7325);
nor U9139 (N_9139,N_7433,N_6900);
and U9140 (N_9140,N_6289,N_6843);
nand U9141 (N_9141,N_6390,N_6710);
or U9142 (N_9142,N_7447,N_7114);
nand U9143 (N_9143,N_6040,N_6462);
xnor U9144 (N_9144,N_7431,N_6569);
and U9145 (N_9145,N_7432,N_7211);
or U9146 (N_9146,N_7395,N_7812);
nor U9147 (N_9147,N_6680,N_6302);
and U9148 (N_9148,N_6668,N_6265);
xor U9149 (N_9149,N_6677,N_7280);
nor U9150 (N_9150,N_7355,N_6817);
and U9151 (N_9151,N_6653,N_6178);
and U9152 (N_9152,N_7473,N_6587);
and U9153 (N_9153,N_7906,N_6289);
and U9154 (N_9154,N_7225,N_7793);
nand U9155 (N_9155,N_6743,N_7743);
or U9156 (N_9156,N_7227,N_6725);
and U9157 (N_9157,N_7073,N_6486);
and U9158 (N_9158,N_6246,N_7951);
and U9159 (N_9159,N_6608,N_7070);
or U9160 (N_9160,N_7260,N_7161);
nor U9161 (N_9161,N_6653,N_6535);
nand U9162 (N_9162,N_7929,N_6591);
nor U9163 (N_9163,N_7686,N_7397);
nor U9164 (N_9164,N_6926,N_6404);
nor U9165 (N_9165,N_6903,N_6710);
and U9166 (N_9166,N_7121,N_7352);
or U9167 (N_9167,N_7062,N_6910);
nor U9168 (N_9168,N_6029,N_6439);
nor U9169 (N_9169,N_7059,N_7959);
nor U9170 (N_9170,N_6543,N_6819);
xnor U9171 (N_9171,N_6619,N_6565);
or U9172 (N_9172,N_6751,N_6011);
and U9173 (N_9173,N_7508,N_7486);
or U9174 (N_9174,N_6330,N_6631);
nand U9175 (N_9175,N_6017,N_6435);
nor U9176 (N_9176,N_6322,N_7941);
and U9177 (N_9177,N_6675,N_6203);
nand U9178 (N_9178,N_7612,N_7436);
or U9179 (N_9179,N_6185,N_7245);
xnor U9180 (N_9180,N_7164,N_7120);
nand U9181 (N_9181,N_7831,N_6991);
nor U9182 (N_9182,N_6729,N_6418);
or U9183 (N_9183,N_6617,N_6930);
nand U9184 (N_9184,N_6539,N_6513);
or U9185 (N_9185,N_7533,N_7507);
nand U9186 (N_9186,N_6414,N_6223);
xor U9187 (N_9187,N_7573,N_7983);
or U9188 (N_9188,N_6262,N_6279);
nor U9189 (N_9189,N_6500,N_7592);
and U9190 (N_9190,N_6353,N_6859);
nor U9191 (N_9191,N_6686,N_6005);
and U9192 (N_9192,N_6958,N_6656);
and U9193 (N_9193,N_6986,N_6499);
nand U9194 (N_9194,N_6720,N_7451);
nor U9195 (N_9195,N_6800,N_7607);
nor U9196 (N_9196,N_6071,N_7352);
nand U9197 (N_9197,N_6020,N_6545);
or U9198 (N_9198,N_7610,N_6518);
and U9199 (N_9199,N_6104,N_6862);
xnor U9200 (N_9200,N_7043,N_7159);
nand U9201 (N_9201,N_6938,N_6088);
nor U9202 (N_9202,N_7199,N_6303);
or U9203 (N_9203,N_6938,N_6845);
nand U9204 (N_9204,N_6291,N_7597);
and U9205 (N_9205,N_7430,N_7503);
nand U9206 (N_9206,N_6671,N_6876);
or U9207 (N_9207,N_7394,N_6713);
and U9208 (N_9208,N_6658,N_7417);
and U9209 (N_9209,N_7666,N_7074);
xnor U9210 (N_9210,N_7894,N_6295);
nand U9211 (N_9211,N_7411,N_7394);
nor U9212 (N_9212,N_6431,N_6453);
or U9213 (N_9213,N_6230,N_7274);
and U9214 (N_9214,N_6569,N_6786);
xnor U9215 (N_9215,N_7804,N_6895);
xor U9216 (N_9216,N_7521,N_6869);
nor U9217 (N_9217,N_6616,N_6378);
or U9218 (N_9218,N_6564,N_7901);
nor U9219 (N_9219,N_6018,N_6356);
xor U9220 (N_9220,N_6255,N_6576);
or U9221 (N_9221,N_7347,N_6142);
nand U9222 (N_9222,N_6609,N_7938);
and U9223 (N_9223,N_7894,N_6633);
xor U9224 (N_9224,N_7602,N_7041);
or U9225 (N_9225,N_6684,N_7656);
nor U9226 (N_9226,N_7001,N_6179);
nand U9227 (N_9227,N_6955,N_7229);
xnor U9228 (N_9228,N_6714,N_7844);
xnor U9229 (N_9229,N_7345,N_6278);
nand U9230 (N_9230,N_6099,N_6097);
and U9231 (N_9231,N_6674,N_7190);
or U9232 (N_9232,N_6691,N_7221);
and U9233 (N_9233,N_7797,N_7058);
and U9234 (N_9234,N_7056,N_6666);
and U9235 (N_9235,N_7463,N_6792);
nand U9236 (N_9236,N_7287,N_6946);
nand U9237 (N_9237,N_7517,N_6677);
and U9238 (N_9238,N_6089,N_6683);
nor U9239 (N_9239,N_7467,N_7580);
nand U9240 (N_9240,N_7299,N_6272);
or U9241 (N_9241,N_7129,N_6796);
or U9242 (N_9242,N_7475,N_6414);
nor U9243 (N_9243,N_7603,N_7368);
nor U9244 (N_9244,N_7414,N_6891);
nor U9245 (N_9245,N_6027,N_6902);
and U9246 (N_9246,N_7940,N_6475);
and U9247 (N_9247,N_6941,N_6293);
xnor U9248 (N_9248,N_7133,N_7088);
nor U9249 (N_9249,N_6276,N_7349);
and U9250 (N_9250,N_6504,N_6175);
nor U9251 (N_9251,N_7204,N_7185);
nor U9252 (N_9252,N_7720,N_7559);
or U9253 (N_9253,N_6033,N_7994);
nand U9254 (N_9254,N_7386,N_7736);
nor U9255 (N_9255,N_7318,N_6981);
nor U9256 (N_9256,N_6125,N_6522);
nor U9257 (N_9257,N_6223,N_6507);
nor U9258 (N_9258,N_6876,N_6446);
xor U9259 (N_9259,N_6734,N_7319);
nand U9260 (N_9260,N_6263,N_6858);
nand U9261 (N_9261,N_6843,N_6620);
or U9262 (N_9262,N_7298,N_7848);
nand U9263 (N_9263,N_6784,N_6885);
nor U9264 (N_9264,N_6007,N_7048);
and U9265 (N_9265,N_7612,N_7666);
or U9266 (N_9266,N_7722,N_7593);
nor U9267 (N_9267,N_7928,N_6721);
or U9268 (N_9268,N_6950,N_6084);
or U9269 (N_9269,N_7214,N_6451);
nand U9270 (N_9270,N_7943,N_7678);
nand U9271 (N_9271,N_6619,N_7337);
nand U9272 (N_9272,N_6460,N_7967);
nand U9273 (N_9273,N_7951,N_6381);
nand U9274 (N_9274,N_6672,N_6504);
nor U9275 (N_9275,N_7899,N_6259);
nand U9276 (N_9276,N_6207,N_7137);
and U9277 (N_9277,N_7775,N_6776);
or U9278 (N_9278,N_6158,N_6298);
nor U9279 (N_9279,N_7204,N_6839);
and U9280 (N_9280,N_7409,N_6569);
nor U9281 (N_9281,N_7055,N_6383);
or U9282 (N_9282,N_7554,N_6813);
nand U9283 (N_9283,N_7039,N_6787);
or U9284 (N_9284,N_6447,N_7133);
or U9285 (N_9285,N_6336,N_6803);
xnor U9286 (N_9286,N_6120,N_6184);
xor U9287 (N_9287,N_7365,N_7796);
nor U9288 (N_9288,N_7331,N_7949);
or U9289 (N_9289,N_6501,N_6024);
or U9290 (N_9290,N_6734,N_7428);
nor U9291 (N_9291,N_6837,N_7051);
and U9292 (N_9292,N_6244,N_7180);
xnor U9293 (N_9293,N_6433,N_6699);
nor U9294 (N_9294,N_7744,N_6286);
and U9295 (N_9295,N_7267,N_6499);
nor U9296 (N_9296,N_7522,N_6690);
nor U9297 (N_9297,N_6462,N_6461);
and U9298 (N_9298,N_7237,N_7396);
nand U9299 (N_9299,N_7758,N_6375);
and U9300 (N_9300,N_7183,N_6617);
nor U9301 (N_9301,N_7056,N_7480);
nand U9302 (N_9302,N_7784,N_7369);
or U9303 (N_9303,N_7125,N_7957);
nand U9304 (N_9304,N_7491,N_6127);
or U9305 (N_9305,N_6100,N_7339);
nor U9306 (N_9306,N_7762,N_6131);
nor U9307 (N_9307,N_7693,N_7287);
and U9308 (N_9308,N_7612,N_6120);
or U9309 (N_9309,N_7173,N_7773);
or U9310 (N_9310,N_6418,N_7426);
nor U9311 (N_9311,N_6049,N_7218);
or U9312 (N_9312,N_7877,N_7664);
nor U9313 (N_9313,N_7466,N_6352);
nor U9314 (N_9314,N_6096,N_7328);
or U9315 (N_9315,N_6867,N_6996);
xnor U9316 (N_9316,N_7931,N_6132);
or U9317 (N_9317,N_6377,N_7034);
nor U9318 (N_9318,N_7243,N_6858);
and U9319 (N_9319,N_7429,N_7015);
nand U9320 (N_9320,N_6316,N_6296);
nand U9321 (N_9321,N_7512,N_7719);
nand U9322 (N_9322,N_6216,N_7921);
and U9323 (N_9323,N_7837,N_6605);
xnor U9324 (N_9324,N_6412,N_6406);
nand U9325 (N_9325,N_7280,N_7983);
xor U9326 (N_9326,N_7443,N_7005);
and U9327 (N_9327,N_6652,N_7094);
nand U9328 (N_9328,N_6447,N_7635);
nand U9329 (N_9329,N_7088,N_6238);
nor U9330 (N_9330,N_6737,N_7660);
nand U9331 (N_9331,N_6497,N_7270);
nor U9332 (N_9332,N_6933,N_6463);
or U9333 (N_9333,N_6106,N_6107);
nand U9334 (N_9334,N_7892,N_7138);
and U9335 (N_9335,N_7907,N_6497);
nor U9336 (N_9336,N_6635,N_7512);
nor U9337 (N_9337,N_7134,N_6995);
nor U9338 (N_9338,N_7258,N_6476);
and U9339 (N_9339,N_6704,N_6540);
xnor U9340 (N_9340,N_6150,N_7546);
or U9341 (N_9341,N_6071,N_7574);
nor U9342 (N_9342,N_6354,N_6754);
nor U9343 (N_9343,N_6365,N_7035);
nor U9344 (N_9344,N_7279,N_7611);
nor U9345 (N_9345,N_7702,N_7467);
and U9346 (N_9346,N_7192,N_6601);
or U9347 (N_9347,N_7239,N_7455);
and U9348 (N_9348,N_7755,N_7045);
and U9349 (N_9349,N_6145,N_7583);
and U9350 (N_9350,N_6273,N_7499);
or U9351 (N_9351,N_7867,N_7108);
nor U9352 (N_9352,N_6342,N_7674);
xor U9353 (N_9353,N_6276,N_7773);
and U9354 (N_9354,N_6418,N_7652);
or U9355 (N_9355,N_7395,N_6351);
xnor U9356 (N_9356,N_6198,N_6266);
xor U9357 (N_9357,N_6682,N_6785);
nand U9358 (N_9358,N_6453,N_7002);
nor U9359 (N_9359,N_7984,N_7332);
nand U9360 (N_9360,N_6386,N_6720);
or U9361 (N_9361,N_6239,N_7798);
and U9362 (N_9362,N_6717,N_6627);
nand U9363 (N_9363,N_6439,N_7534);
nor U9364 (N_9364,N_7573,N_6908);
nand U9365 (N_9365,N_6737,N_6147);
nand U9366 (N_9366,N_6182,N_7983);
and U9367 (N_9367,N_6693,N_7115);
and U9368 (N_9368,N_6646,N_7222);
or U9369 (N_9369,N_6019,N_7771);
nand U9370 (N_9370,N_7655,N_7966);
xnor U9371 (N_9371,N_6658,N_6207);
and U9372 (N_9372,N_6337,N_6184);
nor U9373 (N_9373,N_6010,N_6082);
nand U9374 (N_9374,N_7323,N_6902);
xnor U9375 (N_9375,N_7363,N_6470);
nand U9376 (N_9376,N_6455,N_6063);
and U9377 (N_9377,N_7119,N_6189);
nor U9378 (N_9378,N_6228,N_6757);
and U9379 (N_9379,N_6942,N_6972);
and U9380 (N_9380,N_7930,N_6132);
and U9381 (N_9381,N_6348,N_6606);
nand U9382 (N_9382,N_7134,N_6160);
nor U9383 (N_9383,N_6893,N_7690);
nor U9384 (N_9384,N_7228,N_6444);
nand U9385 (N_9385,N_7602,N_7031);
nand U9386 (N_9386,N_7402,N_6721);
nor U9387 (N_9387,N_7413,N_7459);
and U9388 (N_9388,N_7717,N_6649);
nand U9389 (N_9389,N_6791,N_7232);
and U9390 (N_9390,N_7844,N_7286);
and U9391 (N_9391,N_6970,N_7938);
and U9392 (N_9392,N_6746,N_6273);
xor U9393 (N_9393,N_7063,N_6665);
nand U9394 (N_9394,N_7228,N_6916);
and U9395 (N_9395,N_6925,N_7387);
or U9396 (N_9396,N_6290,N_6669);
xnor U9397 (N_9397,N_6245,N_6034);
and U9398 (N_9398,N_7140,N_7653);
or U9399 (N_9399,N_7610,N_7583);
or U9400 (N_9400,N_7231,N_6494);
and U9401 (N_9401,N_7717,N_6221);
nand U9402 (N_9402,N_6987,N_7496);
nor U9403 (N_9403,N_7181,N_6816);
and U9404 (N_9404,N_7252,N_6074);
nand U9405 (N_9405,N_7188,N_7206);
nor U9406 (N_9406,N_7707,N_6629);
xor U9407 (N_9407,N_6062,N_7341);
nor U9408 (N_9408,N_7937,N_7077);
and U9409 (N_9409,N_6017,N_7484);
or U9410 (N_9410,N_7306,N_7868);
and U9411 (N_9411,N_6408,N_7194);
and U9412 (N_9412,N_6816,N_7874);
xnor U9413 (N_9413,N_6190,N_6212);
or U9414 (N_9414,N_6880,N_7198);
nor U9415 (N_9415,N_7827,N_7240);
or U9416 (N_9416,N_6015,N_6122);
nand U9417 (N_9417,N_7432,N_6178);
or U9418 (N_9418,N_7968,N_6249);
nand U9419 (N_9419,N_6369,N_7751);
nor U9420 (N_9420,N_7801,N_6627);
and U9421 (N_9421,N_7592,N_6578);
nor U9422 (N_9422,N_7235,N_7389);
or U9423 (N_9423,N_6678,N_7995);
nand U9424 (N_9424,N_6151,N_7585);
nand U9425 (N_9425,N_6858,N_6840);
xnor U9426 (N_9426,N_6442,N_6914);
or U9427 (N_9427,N_6298,N_6558);
nand U9428 (N_9428,N_6923,N_6774);
nand U9429 (N_9429,N_7404,N_7903);
xnor U9430 (N_9430,N_7799,N_7472);
nor U9431 (N_9431,N_7116,N_7180);
xnor U9432 (N_9432,N_7627,N_6632);
or U9433 (N_9433,N_7352,N_6249);
nand U9434 (N_9434,N_6892,N_7354);
nand U9435 (N_9435,N_6136,N_7765);
or U9436 (N_9436,N_7167,N_7250);
and U9437 (N_9437,N_7538,N_7197);
nand U9438 (N_9438,N_6600,N_6197);
and U9439 (N_9439,N_6277,N_7136);
nor U9440 (N_9440,N_6867,N_7517);
xor U9441 (N_9441,N_7150,N_7817);
and U9442 (N_9442,N_6039,N_7077);
or U9443 (N_9443,N_6421,N_7318);
nand U9444 (N_9444,N_6313,N_6648);
nor U9445 (N_9445,N_7881,N_6234);
xor U9446 (N_9446,N_7958,N_6116);
or U9447 (N_9447,N_6540,N_7602);
nand U9448 (N_9448,N_6894,N_6857);
nand U9449 (N_9449,N_6769,N_6342);
and U9450 (N_9450,N_6707,N_7854);
nor U9451 (N_9451,N_7442,N_7097);
nand U9452 (N_9452,N_7879,N_7593);
or U9453 (N_9453,N_6904,N_7054);
nor U9454 (N_9454,N_6878,N_7370);
nand U9455 (N_9455,N_7811,N_7889);
nor U9456 (N_9456,N_7126,N_7445);
nand U9457 (N_9457,N_7719,N_6505);
and U9458 (N_9458,N_6910,N_6468);
nor U9459 (N_9459,N_6338,N_6514);
or U9460 (N_9460,N_6092,N_6136);
or U9461 (N_9461,N_6389,N_6518);
or U9462 (N_9462,N_7540,N_6017);
nor U9463 (N_9463,N_7761,N_7887);
nor U9464 (N_9464,N_6548,N_7955);
nor U9465 (N_9465,N_7841,N_7599);
and U9466 (N_9466,N_7484,N_6531);
nor U9467 (N_9467,N_6577,N_7526);
or U9468 (N_9468,N_6493,N_6438);
nor U9469 (N_9469,N_6624,N_7506);
nor U9470 (N_9470,N_7709,N_7773);
or U9471 (N_9471,N_6436,N_7121);
or U9472 (N_9472,N_7263,N_7867);
nand U9473 (N_9473,N_7587,N_7597);
nor U9474 (N_9474,N_7111,N_6245);
or U9475 (N_9475,N_7237,N_6204);
nor U9476 (N_9476,N_7504,N_7305);
or U9477 (N_9477,N_6502,N_6294);
nor U9478 (N_9478,N_7517,N_6651);
nor U9479 (N_9479,N_7437,N_6252);
or U9480 (N_9480,N_6331,N_7237);
or U9481 (N_9481,N_7773,N_6656);
xor U9482 (N_9482,N_7557,N_6634);
xor U9483 (N_9483,N_7488,N_6071);
nand U9484 (N_9484,N_7493,N_7577);
xor U9485 (N_9485,N_6235,N_6310);
or U9486 (N_9486,N_7356,N_7017);
and U9487 (N_9487,N_7119,N_6773);
nor U9488 (N_9488,N_6276,N_6671);
and U9489 (N_9489,N_7837,N_7622);
and U9490 (N_9490,N_7849,N_7778);
and U9491 (N_9491,N_7529,N_6873);
nor U9492 (N_9492,N_7888,N_6755);
nor U9493 (N_9493,N_7930,N_7358);
xnor U9494 (N_9494,N_6274,N_7839);
xor U9495 (N_9495,N_7515,N_7444);
or U9496 (N_9496,N_7001,N_6460);
and U9497 (N_9497,N_6041,N_6097);
xnor U9498 (N_9498,N_6997,N_6286);
nor U9499 (N_9499,N_7052,N_6307);
and U9500 (N_9500,N_7482,N_7859);
nand U9501 (N_9501,N_6281,N_6228);
or U9502 (N_9502,N_6682,N_7096);
and U9503 (N_9503,N_6224,N_6864);
nand U9504 (N_9504,N_7532,N_6302);
nand U9505 (N_9505,N_6405,N_6917);
and U9506 (N_9506,N_6506,N_7196);
and U9507 (N_9507,N_7543,N_7728);
or U9508 (N_9508,N_7308,N_7894);
and U9509 (N_9509,N_7035,N_7896);
nor U9510 (N_9510,N_6916,N_6324);
xnor U9511 (N_9511,N_7806,N_6096);
and U9512 (N_9512,N_6423,N_6669);
and U9513 (N_9513,N_7721,N_7337);
or U9514 (N_9514,N_6769,N_6357);
nand U9515 (N_9515,N_6683,N_7221);
or U9516 (N_9516,N_7832,N_7510);
nand U9517 (N_9517,N_6550,N_7243);
nand U9518 (N_9518,N_7541,N_6452);
and U9519 (N_9519,N_7882,N_6448);
and U9520 (N_9520,N_7227,N_6914);
and U9521 (N_9521,N_6240,N_6401);
nand U9522 (N_9522,N_6832,N_6850);
and U9523 (N_9523,N_7830,N_7896);
or U9524 (N_9524,N_7279,N_6327);
or U9525 (N_9525,N_6859,N_6684);
or U9526 (N_9526,N_7685,N_6943);
and U9527 (N_9527,N_6203,N_7837);
and U9528 (N_9528,N_7089,N_6094);
nor U9529 (N_9529,N_6887,N_6626);
xnor U9530 (N_9530,N_7329,N_7644);
nand U9531 (N_9531,N_6972,N_7901);
or U9532 (N_9532,N_7901,N_7506);
or U9533 (N_9533,N_6437,N_6338);
and U9534 (N_9534,N_7588,N_7166);
nand U9535 (N_9535,N_7279,N_7119);
and U9536 (N_9536,N_6755,N_7156);
nand U9537 (N_9537,N_6398,N_7461);
nor U9538 (N_9538,N_6666,N_7621);
and U9539 (N_9539,N_6063,N_6907);
nand U9540 (N_9540,N_7856,N_6505);
nand U9541 (N_9541,N_6195,N_6759);
xnor U9542 (N_9542,N_6422,N_6650);
nor U9543 (N_9543,N_7501,N_7460);
xnor U9544 (N_9544,N_6055,N_6715);
nand U9545 (N_9545,N_7347,N_6321);
nand U9546 (N_9546,N_6138,N_6857);
nor U9547 (N_9547,N_7991,N_6535);
and U9548 (N_9548,N_7872,N_6717);
xnor U9549 (N_9549,N_6604,N_7379);
and U9550 (N_9550,N_7601,N_6960);
or U9551 (N_9551,N_7558,N_6859);
or U9552 (N_9552,N_6373,N_7898);
nand U9553 (N_9553,N_6752,N_7641);
and U9554 (N_9554,N_6736,N_7571);
or U9555 (N_9555,N_6907,N_7118);
nor U9556 (N_9556,N_6904,N_6017);
nand U9557 (N_9557,N_7164,N_7081);
and U9558 (N_9558,N_7680,N_6184);
and U9559 (N_9559,N_7163,N_6839);
and U9560 (N_9560,N_7129,N_7576);
and U9561 (N_9561,N_6645,N_7044);
and U9562 (N_9562,N_6522,N_6017);
or U9563 (N_9563,N_6707,N_6720);
nor U9564 (N_9564,N_6761,N_6984);
and U9565 (N_9565,N_7931,N_7358);
and U9566 (N_9566,N_6208,N_6847);
or U9567 (N_9567,N_6934,N_7914);
or U9568 (N_9568,N_7852,N_6659);
xnor U9569 (N_9569,N_6586,N_6631);
or U9570 (N_9570,N_7257,N_6293);
nand U9571 (N_9571,N_6459,N_6787);
nor U9572 (N_9572,N_6787,N_7424);
nand U9573 (N_9573,N_7635,N_7122);
xor U9574 (N_9574,N_7066,N_7489);
xnor U9575 (N_9575,N_6947,N_6249);
and U9576 (N_9576,N_6331,N_6600);
nor U9577 (N_9577,N_6240,N_6222);
nand U9578 (N_9578,N_7737,N_6090);
or U9579 (N_9579,N_7942,N_7459);
and U9580 (N_9580,N_7644,N_6298);
xnor U9581 (N_9581,N_6868,N_7797);
nand U9582 (N_9582,N_7591,N_7028);
nor U9583 (N_9583,N_6416,N_6845);
and U9584 (N_9584,N_7327,N_7464);
and U9585 (N_9585,N_6936,N_6110);
nor U9586 (N_9586,N_7007,N_6510);
or U9587 (N_9587,N_6386,N_6580);
and U9588 (N_9588,N_7414,N_7949);
nor U9589 (N_9589,N_6309,N_6480);
or U9590 (N_9590,N_6102,N_6710);
nand U9591 (N_9591,N_7139,N_6110);
nor U9592 (N_9592,N_6838,N_7066);
or U9593 (N_9593,N_7995,N_6876);
or U9594 (N_9594,N_7891,N_7500);
nand U9595 (N_9595,N_6946,N_6702);
and U9596 (N_9596,N_6839,N_6892);
nor U9597 (N_9597,N_7774,N_7670);
and U9598 (N_9598,N_7659,N_7305);
nor U9599 (N_9599,N_7279,N_7232);
nor U9600 (N_9600,N_7834,N_6844);
xnor U9601 (N_9601,N_7991,N_6434);
nor U9602 (N_9602,N_6895,N_7165);
or U9603 (N_9603,N_7593,N_7607);
nand U9604 (N_9604,N_6053,N_6232);
or U9605 (N_9605,N_6024,N_7769);
or U9606 (N_9606,N_6584,N_6468);
nor U9607 (N_9607,N_6702,N_7857);
nor U9608 (N_9608,N_7161,N_6382);
or U9609 (N_9609,N_7977,N_7347);
or U9610 (N_9610,N_7249,N_6647);
xnor U9611 (N_9611,N_7089,N_6460);
nand U9612 (N_9612,N_7273,N_7300);
and U9613 (N_9613,N_6866,N_6741);
or U9614 (N_9614,N_7104,N_7371);
and U9615 (N_9615,N_7952,N_7544);
xor U9616 (N_9616,N_6291,N_6721);
nand U9617 (N_9617,N_7880,N_6276);
or U9618 (N_9618,N_6008,N_7545);
or U9619 (N_9619,N_6199,N_6983);
or U9620 (N_9620,N_7973,N_7219);
nand U9621 (N_9621,N_7450,N_7849);
nand U9622 (N_9622,N_6499,N_6664);
and U9623 (N_9623,N_7390,N_6660);
nor U9624 (N_9624,N_6027,N_7447);
and U9625 (N_9625,N_7502,N_7493);
nand U9626 (N_9626,N_7870,N_7368);
nand U9627 (N_9627,N_6212,N_6247);
and U9628 (N_9628,N_6241,N_7877);
and U9629 (N_9629,N_7068,N_7104);
nor U9630 (N_9630,N_6289,N_6920);
or U9631 (N_9631,N_6598,N_6520);
nand U9632 (N_9632,N_6018,N_6608);
xnor U9633 (N_9633,N_6582,N_6634);
nor U9634 (N_9634,N_6302,N_7483);
or U9635 (N_9635,N_7604,N_7395);
or U9636 (N_9636,N_7558,N_7763);
nand U9637 (N_9637,N_7458,N_7291);
nand U9638 (N_9638,N_6874,N_7598);
and U9639 (N_9639,N_7566,N_7476);
nand U9640 (N_9640,N_6303,N_7807);
or U9641 (N_9641,N_7889,N_7425);
nand U9642 (N_9642,N_6552,N_7147);
or U9643 (N_9643,N_6366,N_7090);
nor U9644 (N_9644,N_6836,N_6400);
nor U9645 (N_9645,N_6127,N_6450);
xnor U9646 (N_9646,N_7764,N_7994);
or U9647 (N_9647,N_6833,N_7719);
xor U9648 (N_9648,N_7954,N_7161);
and U9649 (N_9649,N_7332,N_7166);
nand U9650 (N_9650,N_7796,N_6782);
and U9651 (N_9651,N_6401,N_7435);
nor U9652 (N_9652,N_7208,N_7363);
and U9653 (N_9653,N_6660,N_6631);
nor U9654 (N_9654,N_6417,N_7047);
nand U9655 (N_9655,N_7972,N_6805);
nand U9656 (N_9656,N_6461,N_6560);
nand U9657 (N_9657,N_7530,N_7939);
or U9658 (N_9658,N_6105,N_6188);
nor U9659 (N_9659,N_7528,N_7399);
nor U9660 (N_9660,N_7449,N_7691);
or U9661 (N_9661,N_6476,N_6605);
or U9662 (N_9662,N_6955,N_7697);
nand U9663 (N_9663,N_7031,N_6952);
nand U9664 (N_9664,N_6000,N_7142);
nor U9665 (N_9665,N_7786,N_7194);
nand U9666 (N_9666,N_7761,N_6803);
or U9667 (N_9667,N_7820,N_6771);
nor U9668 (N_9668,N_6952,N_6957);
or U9669 (N_9669,N_7655,N_6372);
or U9670 (N_9670,N_7352,N_7249);
nor U9671 (N_9671,N_6009,N_6187);
xnor U9672 (N_9672,N_7844,N_6677);
or U9673 (N_9673,N_6751,N_6230);
or U9674 (N_9674,N_6603,N_7447);
nor U9675 (N_9675,N_6954,N_7325);
nor U9676 (N_9676,N_7847,N_7991);
and U9677 (N_9677,N_6878,N_7337);
nor U9678 (N_9678,N_7179,N_6830);
nand U9679 (N_9679,N_7509,N_6665);
nor U9680 (N_9680,N_7637,N_6677);
and U9681 (N_9681,N_7627,N_7032);
nand U9682 (N_9682,N_6832,N_7135);
nor U9683 (N_9683,N_7942,N_7811);
nand U9684 (N_9684,N_7518,N_7934);
xnor U9685 (N_9685,N_6368,N_6362);
xor U9686 (N_9686,N_6498,N_6678);
and U9687 (N_9687,N_7219,N_6810);
or U9688 (N_9688,N_7504,N_7085);
and U9689 (N_9689,N_7501,N_6044);
nand U9690 (N_9690,N_6633,N_6600);
or U9691 (N_9691,N_7238,N_7600);
nand U9692 (N_9692,N_7348,N_7300);
xor U9693 (N_9693,N_7908,N_7847);
xnor U9694 (N_9694,N_7398,N_7464);
and U9695 (N_9695,N_6558,N_6037);
nor U9696 (N_9696,N_6325,N_7669);
and U9697 (N_9697,N_7754,N_6197);
nor U9698 (N_9698,N_7900,N_7915);
and U9699 (N_9699,N_6441,N_6030);
or U9700 (N_9700,N_7242,N_7118);
xor U9701 (N_9701,N_6785,N_6087);
or U9702 (N_9702,N_6894,N_6570);
xor U9703 (N_9703,N_7885,N_7849);
and U9704 (N_9704,N_6274,N_6165);
nand U9705 (N_9705,N_6625,N_6095);
and U9706 (N_9706,N_6909,N_7246);
and U9707 (N_9707,N_7678,N_6295);
nand U9708 (N_9708,N_7889,N_6407);
nor U9709 (N_9709,N_7081,N_7510);
nor U9710 (N_9710,N_7320,N_7053);
or U9711 (N_9711,N_6075,N_7798);
nand U9712 (N_9712,N_7863,N_6827);
or U9713 (N_9713,N_6568,N_6315);
nand U9714 (N_9714,N_6961,N_6387);
nor U9715 (N_9715,N_6915,N_6356);
or U9716 (N_9716,N_7431,N_7786);
nand U9717 (N_9717,N_6034,N_7283);
or U9718 (N_9718,N_6705,N_7859);
nor U9719 (N_9719,N_7030,N_7644);
xor U9720 (N_9720,N_6108,N_7216);
or U9721 (N_9721,N_6701,N_7372);
and U9722 (N_9722,N_6375,N_6939);
and U9723 (N_9723,N_7942,N_6013);
or U9724 (N_9724,N_7904,N_7843);
nand U9725 (N_9725,N_7966,N_7185);
nand U9726 (N_9726,N_7305,N_7184);
or U9727 (N_9727,N_7593,N_7006);
nand U9728 (N_9728,N_7983,N_7810);
nor U9729 (N_9729,N_7046,N_6665);
and U9730 (N_9730,N_6757,N_6701);
or U9731 (N_9731,N_6097,N_6456);
nand U9732 (N_9732,N_6866,N_6789);
and U9733 (N_9733,N_6923,N_6790);
and U9734 (N_9734,N_6262,N_6315);
and U9735 (N_9735,N_7044,N_7115);
or U9736 (N_9736,N_7990,N_7370);
or U9737 (N_9737,N_7182,N_7273);
or U9738 (N_9738,N_6578,N_7942);
and U9739 (N_9739,N_6537,N_6129);
and U9740 (N_9740,N_7703,N_6953);
or U9741 (N_9741,N_7222,N_6766);
nand U9742 (N_9742,N_6210,N_7817);
or U9743 (N_9743,N_6006,N_6417);
or U9744 (N_9744,N_7023,N_7255);
or U9745 (N_9745,N_6876,N_6329);
nand U9746 (N_9746,N_7388,N_6503);
and U9747 (N_9747,N_7614,N_7827);
and U9748 (N_9748,N_6163,N_7439);
and U9749 (N_9749,N_7692,N_7710);
and U9750 (N_9750,N_7139,N_7816);
nor U9751 (N_9751,N_7174,N_7257);
nor U9752 (N_9752,N_7987,N_7996);
and U9753 (N_9753,N_7231,N_7610);
nor U9754 (N_9754,N_6988,N_6841);
and U9755 (N_9755,N_7584,N_7248);
nand U9756 (N_9756,N_7427,N_7112);
nor U9757 (N_9757,N_6808,N_6464);
nor U9758 (N_9758,N_7193,N_6601);
nand U9759 (N_9759,N_7138,N_6470);
nor U9760 (N_9760,N_7984,N_7190);
nand U9761 (N_9761,N_7744,N_7794);
xnor U9762 (N_9762,N_6939,N_6357);
nor U9763 (N_9763,N_7803,N_7558);
or U9764 (N_9764,N_6476,N_7982);
nor U9765 (N_9765,N_7179,N_6345);
nand U9766 (N_9766,N_6882,N_7483);
nor U9767 (N_9767,N_6259,N_6344);
or U9768 (N_9768,N_7960,N_7785);
or U9769 (N_9769,N_7871,N_7301);
nor U9770 (N_9770,N_6786,N_7499);
or U9771 (N_9771,N_7560,N_7858);
nand U9772 (N_9772,N_7372,N_7711);
nand U9773 (N_9773,N_7533,N_6346);
or U9774 (N_9774,N_6193,N_6569);
or U9775 (N_9775,N_7760,N_7955);
or U9776 (N_9776,N_7705,N_7195);
or U9777 (N_9777,N_6318,N_6341);
and U9778 (N_9778,N_6891,N_6752);
nand U9779 (N_9779,N_7336,N_7063);
nor U9780 (N_9780,N_6813,N_6465);
nor U9781 (N_9781,N_7075,N_7243);
and U9782 (N_9782,N_6318,N_6924);
xor U9783 (N_9783,N_7761,N_6771);
xnor U9784 (N_9784,N_7445,N_7167);
and U9785 (N_9785,N_6933,N_6443);
nor U9786 (N_9786,N_7132,N_6206);
xnor U9787 (N_9787,N_6856,N_7824);
nand U9788 (N_9788,N_7419,N_6258);
xnor U9789 (N_9789,N_6910,N_6554);
nor U9790 (N_9790,N_6501,N_6456);
nor U9791 (N_9791,N_6614,N_6216);
xnor U9792 (N_9792,N_6994,N_6868);
xor U9793 (N_9793,N_6958,N_6020);
xor U9794 (N_9794,N_6888,N_6951);
nor U9795 (N_9795,N_7695,N_7951);
and U9796 (N_9796,N_6353,N_6236);
nor U9797 (N_9797,N_7217,N_6897);
and U9798 (N_9798,N_7719,N_6781);
and U9799 (N_9799,N_7955,N_6052);
nand U9800 (N_9800,N_6247,N_6906);
nor U9801 (N_9801,N_6467,N_6089);
nand U9802 (N_9802,N_6616,N_7365);
xnor U9803 (N_9803,N_6713,N_7171);
nor U9804 (N_9804,N_7858,N_7696);
nand U9805 (N_9805,N_6585,N_6313);
nand U9806 (N_9806,N_7624,N_7733);
xnor U9807 (N_9807,N_6060,N_6526);
xor U9808 (N_9808,N_6601,N_6798);
and U9809 (N_9809,N_7566,N_6126);
nand U9810 (N_9810,N_6733,N_7517);
nor U9811 (N_9811,N_7004,N_6731);
or U9812 (N_9812,N_6735,N_6390);
or U9813 (N_9813,N_7620,N_6943);
and U9814 (N_9814,N_6899,N_6069);
or U9815 (N_9815,N_6006,N_6085);
nand U9816 (N_9816,N_6123,N_7920);
or U9817 (N_9817,N_6586,N_7442);
and U9818 (N_9818,N_7927,N_6384);
nand U9819 (N_9819,N_7316,N_6777);
xnor U9820 (N_9820,N_7652,N_6559);
and U9821 (N_9821,N_6377,N_7909);
nor U9822 (N_9822,N_7713,N_7541);
nand U9823 (N_9823,N_7333,N_7978);
and U9824 (N_9824,N_7712,N_6503);
and U9825 (N_9825,N_6063,N_6296);
nor U9826 (N_9826,N_7163,N_7635);
or U9827 (N_9827,N_7383,N_6372);
nor U9828 (N_9828,N_7740,N_7323);
or U9829 (N_9829,N_7374,N_7437);
nand U9830 (N_9830,N_6469,N_6175);
xnor U9831 (N_9831,N_7753,N_7297);
nor U9832 (N_9832,N_6032,N_7620);
or U9833 (N_9833,N_7844,N_7003);
or U9834 (N_9834,N_6338,N_6002);
nor U9835 (N_9835,N_7115,N_6612);
or U9836 (N_9836,N_7593,N_6258);
nor U9837 (N_9837,N_6372,N_6391);
nand U9838 (N_9838,N_7681,N_6957);
nand U9839 (N_9839,N_6483,N_6890);
and U9840 (N_9840,N_7677,N_7025);
or U9841 (N_9841,N_7266,N_6097);
nand U9842 (N_9842,N_6949,N_6248);
nand U9843 (N_9843,N_7461,N_6707);
and U9844 (N_9844,N_7455,N_7587);
or U9845 (N_9845,N_6398,N_6462);
nor U9846 (N_9846,N_6139,N_7819);
nor U9847 (N_9847,N_6691,N_7972);
and U9848 (N_9848,N_7226,N_6051);
or U9849 (N_9849,N_6355,N_7704);
nand U9850 (N_9850,N_6321,N_7301);
nand U9851 (N_9851,N_6704,N_6386);
nor U9852 (N_9852,N_7938,N_6011);
xor U9853 (N_9853,N_7218,N_6649);
nor U9854 (N_9854,N_7847,N_6606);
nand U9855 (N_9855,N_6796,N_7375);
or U9856 (N_9856,N_7097,N_6649);
nand U9857 (N_9857,N_6728,N_7237);
nor U9858 (N_9858,N_7834,N_7356);
and U9859 (N_9859,N_7266,N_6483);
or U9860 (N_9860,N_7087,N_6367);
nand U9861 (N_9861,N_7062,N_6187);
nand U9862 (N_9862,N_6774,N_6570);
nor U9863 (N_9863,N_7100,N_7164);
and U9864 (N_9864,N_7467,N_6705);
and U9865 (N_9865,N_6980,N_7411);
nor U9866 (N_9866,N_6014,N_6245);
or U9867 (N_9867,N_6425,N_6205);
xor U9868 (N_9868,N_7198,N_6057);
nand U9869 (N_9869,N_7170,N_7952);
nor U9870 (N_9870,N_7187,N_7224);
and U9871 (N_9871,N_7307,N_7090);
and U9872 (N_9872,N_6846,N_6680);
and U9873 (N_9873,N_6433,N_7329);
nand U9874 (N_9874,N_6250,N_6796);
nor U9875 (N_9875,N_6261,N_7407);
and U9876 (N_9876,N_6858,N_6980);
nand U9877 (N_9877,N_6628,N_6031);
or U9878 (N_9878,N_6732,N_6051);
nor U9879 (N_9879,N_6732,N_7146);
nor U9880 (N_9880,N_7776,N_6940);
nand U9881 (N_9881,N_7664,N_7505);
xor U9882 (N_9882,N_6130,N_7785);
or U9883 (N_9883,N_7471,N_6319);
nor U9884 (N_9884,N_6004,N_6964);
nand U9885 (N_9885,N_7063,N_6920);
nand U9886 (N_9886,N_6152,N_6003);
or U9887 (N_9887,N_6275,N_7244);
xnor U9888 (N_9888,N_7614,N_6214);
or U9889 (N_9889,N_6610,N_6505);
and U9890 (N_9890,N_7239,N_7131);
and U9891 (N_9891,N_7318,N_7327);
or U9892 (N_9892,N_7767,N_7433);
nand U9893 (N_9893,N_7732,N_7707);
nor U9894 (N_9894,N_7532,N_7423);
or U9895 (N_9895,N_6295,N_6779);
and U9896 (N_9896,N_7278,N_6270);
nor U9897 (N_9897,N_6043,N_6010);
nor U9898 (N_9898,N_7533,N_6996);
and U9899 (N_9899,N_6950,N_6636);
nor U9900 (N_9900,N_6562,N_6958);
nand U9901 (N_9901,N_6369,N_6848);
or U9902 (N_9902,N_6370,N_7590);
and U9903 (N_9903,N_7680,N_7051);
and U9904 (N_9904,N_6309,N_6584);
nor U9905 (N_9905,N_7761,N_7652);
nand U9906 (N_9906,N_7951,N_6153);
nand U9907 (N_9907,N_6024,N_6917);
nor U9908 (N_9908,N_7712,N_6311);
and U9909 (N_9909,N_6278,N_7032);
or U9910 (N_9910,N_7890,N_7770);
or U9911 (N_9911,N_6621,N_6393);
and U9912 (N_9912,N_6609,N_7289);
or U9913 (N_9913,N_7294,N_6908);
or U9914 (N_9914,N_7234,N_7995);
and U9915 (N_9915,N_6312,N_7374);
nand U9916 (N_9916,N_6228,N_7771);
and U9917 (N_9917,N_7301,N_6843);
nor U9918 (N_9918,N_7763,N_7014);
or U9919 (N_9919,N_6322,N_6814);
and U9920 (N_9920,N_7037,N_6434);
or U9921 (N_9921,N_7775,N_7634);
and U9922 (N_9922,N_7930,N_6033);
or U9923 (N_9923,N_7605,N_7081);
and U9924 (N_9924,N_7795,N_6073);
or U9925 (N_9925,N_7892,N_6573);
and U9926 (N_9926,N_7314,N_7573);
nand U9927 (N_9927,N_6959,N_7378);
nor U9928 (N_9928,N_6566,N_6747);
nor U9929 (N_9929,N_6106,N_7512);
nor U9930 (N_9930,N_6621,N_7047);
nand U9931 (N_9931,N_7361,N_7454);
nand U9932 (N_9932,N_6109,N_6032);
and U9933 (N_9933,N_7622,N_6211);
xor U9934 (N_9934,N_7010,N_6829);
and U9935 (N_9935,N_6293,N_6415);
nand U9936 (N_9936,N_7293,N_6024);
and U9937 (N_9937,N_7247,N_7477);
xor U9938 (N_9938,N_6647,N_7379);
nand U9939 (N_9939,N_7592,N_6352);
nor U9940 (N_9940,N_7844,N_7193);
or U9941 (N_9941,N_7645,N_6806);
nor U9942 (N_9942,N_6618,N_6718);
xnor U9943 (N_9943,N_6728,N_6943);
xnor U9944 (N_9944,N_7473,N_6352);
and U9945 (N_9945,N_6180,N_7472);
or U9946 (N_9946,N_6386,N_7074);
or U9947 (N_9947,N_6275,N_7994);
or U9948 (N_9948,N_7481,N_6008);
or U9949 (N_9949,N_7397,N_6357);
nand U9950 (N_9950,N_6726,N_6430);
nand U9951 (N_9951,N_7931,N_7977);
nor U9952 (N_9952,N_6883,N_7975);
or U9953 (N_9953,N_7499,N_6873);
or U9954 (N_9954,N_7269,N_7984);
or U9955 (N_9955,N_7901,N_7566);
and U9956 (N_9956,N_6865,N_7643);
nor U9957 (N_9957,N_7405,N_6574);
nand U9958 (N_9958,N_6328,N_6062);
or U9959 (N_9959,N_7311,N_7769);
or U9960 (N_9960,N_7206,N_6800);
or U9961 (N_9961,N_7526,N_6638);
or U9962 (N_9962,N_6381,N_7970);
nor U9963 (N_9963,N_6594,N_6882);
and U9964 (N_9964,N_7583,N_7913);
or U9965 (N_9965,N_7975,N_6278);
nand U9966 (N_9966,N_7552,N_6627);
nor U9967 (N_9967,N_7032,N_7943);
nand U9968 (N_9968,N_6304,N_6112);
or U9969 (N_9969,N_7430,N_7626);
nand U9970 (N_9970,N_6686,N_6513);
nor U9971 (N_9971,N_7157,N_7423);
nor U9972 (N_9972,N_7517,N_6844);
and U9973 (N_9973,N_7172,N_6109);
and U9974 (N_9974,N_7817,N_7686);
or U9975 (N_9975,N_7471,N_7129);
xor U9976 (N_9976,N_7555,N_6932);
nor U9977 (N_9977,N_7654,N_7860);
and U9978 (N_9978,N_6985,N_6237);
nand U9979 (N_9979,N_6828,N_6505);
and U9980 (N_9980,N_7189,N_6551);
or U9981 (N_9981,N_6218,N_6445);
nor U9982 (N_9982,N_6076,N_6422);
and U9983 (N_9983,N_7315,N_7217);
or U9984 (N_9984,N_7367,N_7975);
nor U9985 (N_9985,N_7469,N_6182);
nand U9986 (N_9986,N_6568,N_7840);
nor U9987 (N_9987,N_7785,N_6849);
and U9988 (N_9988,N_6293,N_6565);
nand U9989 (N_9989,N_7884,N_6159);
nand U9990 (N_9990,N_7502,N_6509);
nor U9991 (N_9991,N_6317,N_7791);
xnor U9992 (N_9992,N_6053,N_6604);
nor U9993 (N_9993,N_7821,N_7645);
nor U9994 (N_9994,N_6415,N_7174);
nor U9995 (N_9995,N_7360,N_7451);
nor U9996 (N_9996,N_7180,N_6720);
nand U9997 (N_9997,N_6010,N_7073);
or U9998 (N_9998,N_7504,N_6429);
nor U9999 (N_9999,N_7170,N_6183);
or U10000 (N_10000,N_8282,N_8658);
and U10001 (N_10001,N_9127,N_8443);
and U10002 (N_10002,N_9066,N_9864);
nor U10003 (N_10003,N_9419,N_9297);
nor U10004 (N_10004,N_8362,N_8932);
and U10005 (N_10005,N_8575,N_9711);
xnor U10006 (N_10006,N_8463,N_8855);
or U10007 (N_10007,N_8270,N_8579);
or U10008 (N_10008,N_8035,N_9984);
or U10009 (N_10009,N_8147,N_9214);
and U10010 (N_10010,N_8217,N_9936);
and U10011 (N_10011,N_9304,N_8605);
or U10012 (N_10012,N_8833,N_9045);
and U10013 (N_10013,N_8054,N_9008);
nor U10014 (N_10014,N_9628,N_9540);
nand U10015 (N_10015,N_8484,N_9097);
and U10016 (N_10016,N_8345,N_8310);
or U10017 (N_10017,N_9988,N_9291);
or U10018 (N_10018,N_8713,N_9973);
xor U10019 (N_10019,N_8535,N_9273);
or U10020 (N_10020,N_8966,N_9779);
or U10021 (N_10021,N_8827,N_9530);
nor U10022 (N_10022,N_9844,N_8051);
and U10023 (N_10023,N_8913,N_9911);
and U10024 (N_10024,N_8512,N_8832);
or U10025 (N_10025,N_9560,N_8329);
xnor U10026 (N_10026,N_8903,N_8444);
nor U10027 (N_10027,N_9772,N_9661);
or U10028 (N_10028,N_8016,N_8255);
nand U10029 (N_10029,N_8729,N_8702);
nand U10030 (N_10030,N_8047,N_9733);
nor U10031 (N_10031,N_9789,N_9978);
nor U10032 (N_10032,N_9437,N_9506);
nor U10033 (N_10033,N_9270,N_8079);
and U10034 (N_10034,N_8243,N_9263);
and U10035 (N_10035,N_8754,N_9591);
or U10036 (N_10036,N_8887,N_8701);
and U10037 (N_10037,N_9333,N_8026);
nand U10038 (N_10038,N_9735,N_8465);
and U10039 (N_10039,N_9011,N_9755);
and U10040 (N_10040,N_9104,N_9309);
and U10041 (N_10041,N_8870,N_9310);
and U10042 (N_10042,N_9116,N_8140);
or U10043 (N_10043,N_9326,N_8339);
and U10044 (N_10044,N_9536,N_9373);
nand U10045 (N_10045,N_8170,N_9537);
and U10046 (N_10046,N_9525,N_9856);
nand U10047 (N_10047,N_9528,N_9181);
nor U10048 (N_10048,N_9646,N_9036);
and U10049 (N_10049,N_9023,N_9826);
nand U10050 (N_10050,N_8541,N_9126);
or U10051 (N_10051,N_8802,N_9169);
or U10052 (N_10052,N_9059,N_9794);
nor U10053 (N_10053,N_8543,N_8820);
nand U10054 (N_10054,N_8759,N_9015);
nand U10055 (N_10055,N_9171,N_8335);
or U10056 (N_10056,N_8417,N_8772);
or U10057 (N_10057,N_8354,N_9717);
and U10058 (N_10058,N_9738,N_9925);
or U10059 (N_10059,N_9369,N_8184);
and U10060 (N_10060,N_9824,N_8319);
and U10061 (N_10061,N_9545,N_8994);
and U10062 (N_10062,N_8317,N_9742);
nand U10063 (N_10063,N_8737,N_9344);
nor U10064 (N_10064,N_9150,N_9423);
xnor U10065 (N_10065,N_8782,N_9072);
nor U10066 (N_10066,N_9922,N_9107);
xor U10067 (N_10067,N_8192,N_9960);
xnor U10068 (N_10068,N_9586,N_8076);
nand U10069 (N_10069,N_8404,N_8916);
and U10070 (N_10070,N_9793,N_9024);
nand U10071 (N_10071,N_9800,N_8379);
or U10072 (N_10072,N_9714,N_8059);
or U10073 (N_10073,N_9474,N_8005);
or U10074 (N_10074,N_8272,N_8922);
and U10075 (N_10075,N_8756,N_8485);
nor U10076 (N_10076,N_8876,N_8518);
and U10077 (N_10077,N_8371,N_9436);
nor U10078 (N_10078,N_9145,N_8235);
or U10079 (N_10079,N_9180,N_9165);
and U10080 (N_10080,N_8623,N_9211);
or U10081 (N_10081,N_8072,N_8933);
or U10082 (N_10082,N_8636,N_9820);
nor U10083 (N_10083,N_9421,N_8914);
nor U10084 (N_10084,N_8284,N_8992);
xor U10085 (N_10085,N_8571,N_8186);
or U10086 (N_10086,N_8608,N_8323);
nor U10087 (N_10087,N_9534,N_8407);
or U10088 (N_10088,N_9523,N_8018);
nand U10089 (N_10089,N_8945,N_9642);
nand U10090 (N_10090,N_8818,N_8098);
and U10091 (N_10091,N_9161,N_9699);
nand U10092 (N_10092,N_9814,N_8591);
nand U10093 (N_10093,N_8908,N_9961);
or U10094 (N_10094,N_8764,N_8346);
xnor U10095 (N_10095,N_8784,N_9640);
xnor U10096 (N_10096,N_9515,N_8169);
and U10097 (N_10097,N_8561,N_9902);
nor U10098 (N_10098,N_9042,N_8293);
or U10099 (N_10099,N_9977,N_8618);
and U10100 (N_10100,N_9808,N_8011);
and U10101 (N_10101,N_8088,N_8995);
nand U10102 (N_10102,N_8934,N_9645);
xor U10103 (N_10103,N_9890,N_8332);
or U10104 (N_10104,N_8686,N_9802);
nand U10105 (N_10105,N_8368,N_8682);
and U10106 (N_10106,N_8227,N_9604);
or U10107 (N_10107,N_9092,N_9593);
nor U10108 (N_10108,N_8146,N_9601);
or U10109 (N_10109,N_9972,N_9550);
nand U10110 (N_10110,N_8927,N_8071);
nor U10111 (N_10111,N_8373,N_9394);
nor U10112 (N_10112,N_9328,N_8711);
or U10113 (N_10113,N_8931,N_8479);
nand U10114 (N_10114,N_8514,N_8889);
xnor U10115 (N_10115,N_9607,N_8178);
and U10116 (N_10116,N_9160,N_8999);
nand U10117 (N_10117,N_9576,N_8464);
xnor U10118 (N_10118,N_8476,N_8955);
nand U10119 (N_10119,N_9153,N_8313);
nor U10120 (N_10120,N_9086,N_9941);
xnor U10121 (N_10121,N_8730,N_9602);
or U10122 (N_10122,N_8250,N_9582);
and U10123 (N_10123,N_9842,N_8722);
nand U10124 (N_10124,N_8988,N_9775);
and U10125 (N_10125,N_8228,N_9098);
nand U10126 (N_10126,N_8638,N_9233);
and U10127 (N_10127,N_9431,N_8321);
and U10128 (N_10128,N_8288,N_9823);
xnor U10129 (N_10129,N_9848,N_8924);
and U10130 (N_10130,N_9201,N_8568);
or U10131 (N_10131,N_9608,N_8100);
and U10132 (N_10132,N_9222,N_8232);
or U10133 (N_10133,N_8734,N_9644);
xnor U10134 (N_10134,N_8306,N_9004);
or U10135 (N_10135,N_9937,N_8322);
and U10136 (N_10136,N_8418,N_8635);
nand U10137 (N_10137,N_9198,N_9447);
nor U10138 (N_10138,N_9449,N_8705);
and U10139 (N_10139,N_9473,N_9278);
and U10140 (N_10140,N_9833,N_9010);
and U10141 (N_10141,N_9346,N_8849);
and U10142 (N_10142,N_8482,N_8625);
and U10143 (N_10143,N_8207,N_8644);
xnor U10144 (N_10144,N_8126,N_8634);
nor U10145 (N_10145,N_9438,N_9991);
or U10146 (N_10146,N_9874,N_9505);
or U10147 (N_10147,N_9479,N_9368);
nor U10148 (N_10148,N_9957,N_9355);
nand U10149 (N_10149,N_9187,N_9627);
nand U10150 (N_10150,N_8537,N_8359);
nand U10151 (N_10151,N_8841,N_8829);
or U10152 (N_10152,N_8566,N_9684);
xnor U10153 (N_10153,N_9425,N_9228);
xor U10154 (N_10154,N_9568,N_9021);
and U10155 (N_10155,N_9279,N_9354);
nand U10156 (N_10156,N_8249,N_9812);
or U10157 (N_10157,N_8172,N_8360);
nor U10158 (N_10158,N_9511,N_8891);
nor U10159 (N_10159,N_9791,N_9889);
or U10160 (N_10160,N_9347,N_8540);
and U10161 (N_10161,N_8167,N_8271);
nand U10162 (N_10162,N_8956,N_8381);
xor U10163 (N_10163,N_9685,N_9884);
nand U10164 (N_10164,N_9167,N_8452);
and U10165 (N_10165,N_9641,N_8470);
or U10166 (N_10166,N_8196,N_9632);
nor U10167 (N_10167,N_8923,N_8388);
nor U10168 (N_10168,N_8168,N_9725);
and U10169 (N_10169,N_9598,N_8180);
nand U10170 (N_10170,N_9217,N_8811);
or U10171 (N_10171,N_9485,N_8599);
and U10172 (N_10172,N_8794,N_8307);
and U10173 (N_10173,N_9965,N_8967);
nor U10174 (N_10174,N_8584,N_8337);
and U10175 (N_10175,N_8646,N_8156);
or U10176 (N_10176,N_8344,N_9865);
or U10177 (N_10177,N_9231,N_9442);
nand U10178 (N_10178,N_9037,N_9189);
and U10179 (N_10179,N_9331,N_9185);
nor U10180 (N_10180,N_8781,N_9134);
or U10181 (N_10181,N_8691,N_9982);
and U10182 (N_10182,N_9781,N_9096);
or U10183 (N_10183,N_8879,N_8052);
and U10184 (N_10184,N_9953,N_8256);
or U10185 (N_10185,N_8130,N_9048);
or U10186 (N_10186,N_8036,N_8695);
or U10187 (N_10187,N_8174,N_8403);
nand U10188 (N_10188,N_8108,N_8218);
xor U10189 (N_10189,N_9335,N_8901);
and U10190 (N_10190,N_9558,N_9410);
and U10191 (N_10191,N_9910,N_8002);
xor U10192 (N_10192,N_8336,N_9840);
and U10193 (N_10193,N_8708,N_9541);
and U10194 (N_10194,N_9516,N_8939);
nand U10195 (N_10195,N_9241,N_9778);
or U10196 (N_10196,N_9559,N_8395);
nor U10197 (N_10197,N_9188,N_9696);
nor U10198 (N_10198,N_9337,N_9843);
nor U10199 (N_10199,N_8019,N_9477);
and U10200 (N_10200,N_9302,N_8300);
or U10201 (N_10201,N_8869,N_8659);
and U10202 (N_10202,N_9799,N_9056);
nor U10203 (N_10203,N_8183,N_9796);
nand U10204 (N_10204,N_9868,N_9664);
and U10205 (N_10205,N_9486,N_9689);
nand U10206 (N_10206,N_8245,N_9702);
nor U10207 (N_10207,N_9080,N_9359);
or U10208 (N_10208,N_9895,N_9782);
or U10209 (N_10209,N_9091,N_8439);
or U10210 (N_10210,N_9260,N_8238);
xnor U10211 (N_10211,N_8075,N_8921);
and U10212 (N_10212,N_8765,N_9353);
nor U10213 (N_10213,N_9698,N_8063);
or U10214 (N_10214,N_8806,N_9815);
or U10215 (N_10215,N_9009,N_8983);
and U10216 (N_10216,N_8220,N_8893);
and U10217 (N_10217,N_8555,N_9268);
nor U10218 (N_10218,N_9434,N_8954);
nand U10219 (N_10219,N_8763,N_9102);
nor U10220 (N_10220,N_8134,N_9517);
and U10221 (N_10221,N_8986,N_8214);
xor U10222 (N_10222,N_9115,N_9716);
nand U10223 (N_10223,N_9117,N_9583);
or U10224 (N_10224,N_8340,N_9636);
nor U10225 (N_10225,N_9544,N_8799);
and U10226 (N_10226,N_9365,N_8166);
and U10227 (N_10227,N_8865,N_9863);
nand U10228 (N_10228,N_8997,N_9964);
and U10229 (N_10229,N_9599,N_9146);
nor U10230 (N_10230,N_9592,N_9514);
or U10231 (N_10231,N_9934,N_8269);
or U10232 (N_10232,N_8456,N_9543);
nand U10233 (N_10233,N_9352,N_8853);
nor U10234 (N_10234,N_8836,N_9396);
xnor U10235 (N_10235,N_8024,N_9459);
nand U10236 (N_10236,N_8621,N_8008);
and U10237 (N_10237,N_8960,N_9235);
and U10238 (N_10238,N_9557,N_9663);
or U10239 (N_10239,N_9497,N_8803);
nor U10240 (N_10240,N_9881,N_8970);
nor U10241 (N_10241,N_8428,N_9053);
and U10242 (N_10242,N_9247,N_8926);
xnor U10243 (N_10243,N_9886,N_8478);
or U10244 (N_10244,N_9805,N_8355);
xor U10245 (N_10245,N_8867,N_9518);
nand U10246 (N_10246,N_9708,N_8352);
nand U10247 (N_10247,N_9921,N_8067);
nor U10248 (N_10248,N_8102,N_9413);
and U10249 (N_10249,N_9500,N_8048);
or U10250 (N_10250,N_9345,N_9949);
and U10251 (N_10251,N_9891,N_8607);
nand U10252 (N_10252,N_9736,N_8033);
nand U10253 (N_10253,N_9305,N_8420);
nor U10254 (N_10254,N_9513,N_9367);
or U10255 (N_10255,N_8442,N_8065);
nor U10256 (N_10256,N_8560,N_9058);
and U10257 (N_10257,N_9963,N_8538);
nor U10258 (N_10258,N_9016,N_8424);
and U10259 (N_10259,N_9580,N_8055);
and U10260 (N_10260,N_9729,N_8953);
nand U10261 (N_10261,N_8502,N_8043);
and U10262 (N_10262,N_8259,N_8610);
nand U10263 (N_10263,N_9786,N_8374);
and U10264 (N_10264,N_8370,N_8828);
and U10265 (N_10265,N_9424,N_9759);
nand U10266 (N_10266,N_8461,N_9932);
xor U10267 (N_10267,N_9931,N_9503);
nor U10268 (N_10268,N_9596,N_8978);
and U10269 (N_10269,N_9967,N_8287);
nor U10270 (N_10270,N_9920,N_9283);
nand U10271 (N_10271,N_8438,N_9139);
nand U10272 (N_10272,N_9626,N_9147);
and U10273 (N_10273,N_9435,N_9594);
nand U10274 (N_10274,N_8408,N_9197);
and U10275 (N_10275,N_8350,N_8455);
xnor U10276 (N_10276,N_8117,N_8351);
and U10277 (N_10277,N_8712,N_9252);
nor U10278 (N_10278,N_9014,N_8624);
or U10279 (N_10279,N_8637,N_9770);
nor U10280 (N_10280,N_9039,N_9205);
and U10281 (N_10281,N_8261,N_8044);
nand U10282 (N_10282,N_8440,N_9081);
or U10283 (N_10283,N_8520,N_9028);
or U10284 (N_10284,N_9792,N_8738);
xnor U10285 (N_10285,N_8750,N_8657);
and U10286 (N_10286,N_8603,N_9184);
or U10287 (N_10287,N_9451,N_8380);
nor U10288 (N_10288,N_8703,N_9532);
nor U10289 (N_10289,N_9285,N_9194);
and U10290 (N_10290,N_9570,N_8755);
or U10291 (N_10291,N_9099,N_9510);
or U10292 (N_10292,N_8390,N_9851);
xor U10293 (N_10293,N_8819,N_8679);
nor U10294 (N_10294,N_8205,N_9569);
and U10295 (N_10295,N_8690,N_8837);
nor U10296 (N_10296,N_8640,N_9658);
and U10297 (N_10297,N_8328,N_8675);
and U10298 (N_10298,N_9624,N_8357);
or U10299 (N_10299,N_8006,N_9401);
nand U10300 (N_10300,N_9682,N_8961);
nand U10301 (N_10301,N_8057,N_8678);
nor U10302 (N_10302,N_9867,N_8431);
nor U10303 (N_10303,N_8771,N_9549);
nand U10304 (N_10304,N_9392,N_8137);
nand U10305 (N_10305,N_9670,N_9261);
nor U10306 (N_10306,N_8399,N_8155);
nor U10307 (N_10307,N_8116,N_9740);
and U10308 (N_10308,N_9075,N_9494);
and U10309 (N_10309,N_8551,N_8487);
nor U10310 (N_10310,N_9001,N_9384);
or U10311 (N_10311,N_8330,N_8215);
or U10312 (N_10312,N_8533,N_8124);
or U10313 (N_10313,N_9588,N_8376);
or U10314 (N_10314,N_8495,N_9718);
nand U10315 (N_10315,N_8101,N_8132);
nand U10316 (N_10316,N_8861,N_9176);
or U10317 (N_10317,N_8414,N_8548);
nor U10318 (N_10318,N_9484,N_8740);
xnor U10319 (N_10319,N_9721,N_9264);
or U10320 (N_10320,N_8706,N_9332);
nor U10321 (N_10321,N_8058,N_9258);
nor U10322 (N_10322,N_8257,N_8735);
nor U10323 (N_10323,N_9149,N_8549);
nor U10324 (N_10324,N_9512,N_9981);
nand U10325 (N_10325,N_8546,N_8292);
and U10326 (N_10326,N_9177,N_8663);
and U10327 (N_10327,N_8299,N_8696);
and U10328 (N_10328,N_9956,N_9199);
or U10329 (N_10329,N_9723,N_8987);
and U10330 (N_10330,N_9120,N_9831);
and U10331 (N_10331,N_8219,N_8433);
and U10332 (N_10332,N_9356,N_8023);
or U10333 (N_10333,N_9630,N_8662);
xor U10334 (N_10334,N_8038,N_9440);
nand U10335 (N_10335,N_8494,N_8015);
or U10336 (N_10336,N_9019,N_9930);
nand U10337 (N_10337,N_9478,N_8831);
and U10338 (N_10338,N_8613,N_9662);
and U10339 (N_10339,N_9143,N_8990);
or U10340 (N_10340,N_8466,N_9554);
and U10341 (N_10341,N_8894,N_8092);
nor U10342 (N_10342,N_8974,N_9676);
and U10343 (N_10343,N_9521,N_9565);
nand U10344 (N_10344,N_9130,N_8904);
or U10345 (N_10345,N_9025,N_9316);
or U10346 (N_10346,N_8628,N_9142);
or U10347 (N_10347,N_8776,N_9818);
and U10348 (N_10348,N_9940,N_9206);
nor U10349 (N_10349,N_9371,N_9595);
or U10350 (N_10350,N_8073,N_9763);
and U10351 (N_10351,N_8162,N_9952);
xor U10352 (N_10352,N_8587,N_9675);
nand U10353 (N_10353,N_9342,N_9915);
nor U10354 (N_10354,N_8509,N_8716);
or U10355 (N_10355,N_8886,N_9387);
nand U10356 (N_10356,N_9219,N_8815);
nand U10357 (N_10357,N_9374,N_8731);
nand U10358 (N_10358,N_9509,N_8206);
nand U10359 (N_10359,N_8211,N_9329);
or U10360 (N_10360,N_8212,N_9695);
nor U10361 (N_10361,N_9154,N_8040);
nand U10362 (N_10362,N_9128,N_9106);
nor U10363 (N_10363,N_9005,N_9271);
or U10364 (N_10364,N_8991,N_9667);
nor U10365 (N_10365,N_8632,N_9912);
and U10366 (N_10366,N_9055,N_8112);
or U10367 (N_10367,N_9462,N_9531);
nand U10368 (N_10368,N_9340,N_9221);
or U10369 (N_10369,N_8203,N_8860);
nand U10370 (N_10370,N_9993,N_9680);
or U10371 (N_10371,N_8389,N_9012);
nor U10372 (N_10372,N_9606,N_8979);
or U10373 (N_10373,N_9616,N_8745);
and U10374 (N_10374,N_8209,N_8748);
nor U10375 (N_10375,N_8077,N_8539);
nand U10376 (N_10376,N_9766,N_9958);
nand U10377 (N_10377,N_9614,N_9454);
nand U10378 (N_10378,N_9597,N_9315);
xor U10379 (N_10379,N_9909,N_8157);
and U10380 (N_10380,N_8700,N_9460);
and U10381 (N_10381,N_9090,N_8268);
xor U10382 (N_10382,N_8797,N_8830);
or U10383 (N_10383,N_9888,N_8226);
nor U10384 (N_10384,N_9100,N_8736);
and U10385 (N_10385,N_9827,N_8435);
nor U10386 (N_10386,N_8042,N_9089);
nor U10387 (N_10387,N_9686,N_9880);
nor U10388 (N_10388,N_9311,N_9338);
and U10389 (N_10389,N_8789,N_9215);
or U10390 (N_10390,N_8198,N_9649);
nor U10391 (N_10391,N_9681,N_8937);
nor U10392 (N_10392,N_8925,N_9444);
or U10393 (N_10393,N_9555,N_9566);
nand U10394 (N_10394,N_8767,N_8145);
nand U10395 (N_10395,N_9955,N_9151);
nand U10396 (N_10396,N_9162,N_9746);
or U10397 (N_10397,N_8111,N_8800);
nand U10398 (N_10398,N_8273,N_9136);
and U10399 (N_10399,N_9507,N_9320);
or U10400 (N_10400,N_9455,N_8519);
and U10401 (N_10401,N_9672,N_9467);
and U10402 (N_10402,N_9807,N_8508);
nor U10403 (N_10403,N_9905,N_8809);
nand U10404 (N_10404,N_8030,N_9109);
or U10405 (N_10405,N_9208,N_9829);
nand U10406 (N_10406,N_9051,N_8483);
or U10407 (N_10407,N_8324,N_8325);
nor U10408 (N_10408,N_9919,N_9140);
nor U10409 (N_10409,N_9852,N_9527);
or U10410 (N_10410,N_9893,N_9861);
and U10411 (N_10411,N_8899,N_8128);
nand U10412 (N_10412,N_8153,N_9892);
xnor U10413 (N_10413,N_9069,N_9765);
nor U10414 (N_10414,N_9105,N_8798);
or U10415 (N_10415,N_9617,N_9994);
or U10416 (N_10416,N_9414,N_8872);
and U10417 (N_10417,N_9622,N_8594);
nor U10418 (N_10418,N_8918,N_9780);
and U10419 (N_10419,N_8884,N_9704);
and U10420 (N_10420,N_9432,N_8338);
and U10421 (N_10421,N_8779,N_9050);
nand U10422 (N_10422,N_8447,N_8910);
nor U10423 (N_10423,N_8046,N_8411);
nand U10424 (N_10424,N_8471,N_9108);
or U10425 (N_10425,N_9519,N_9853);
nor U10426 (N_10426,N_8917,N_8505);
and U10427 (N_10427,N_8761,N_9398);
nand U10428 (N_10428,N_8823,N_9966);
or U10429 (N_10429,N_9006,N_8254);
and U10430 (N_10430,N_8796,N_8720);
and U10431 (N_10431,N_8064,N_8240);
or U10432 (N_10432,N_9286,N_8847);
nor U10433 (N_10433,N_9041,N_8410);
and U10434 (N_10434,N_9192,N_9299);
and U10435 (N_10435,N_9971,N_9490);
or U10436 (N_10436,N_8320,N_9694);
or U10437 (N_10437,N_8105,N_9539);
nand U10438 (N_10438,N_9655,N_8118);
nor U10439 (N_10439,N_9357,N_9574);
nor U10440 (N_10440,N_8813,N_9618);
nand U10441 (N_10441,N_8825,N_8187);
xnor U10442 (N_10442,N_9846,N_9903);
nand U10443 (N_10443,N_8687,N_8786);
nor U10444 (N_10444,N_8427,N_9870);
xnor U10445 (N_10445,N_8326,N_9872);
xnor U10446 (N_10446,N_9251,N_8526);
xor U10447 (N_10447,N_8515,N_8941);
and U10448 (N_10448,N_9253,N_8681);
nor U10449 (N_10449,N_9730,N_9634);
or U10450 (N_10450,N_8291,N_8387);
nand U10451 (N_10451,N_8888,N_8839);
nor U10452 (N_10452,N_8199,N_8586);
nor U10453 (N_10453,N_8697,N_8302);
and U10454 (N_10454,N_8525,N_8715);
nand U10455 (N_10455,N_8467,N_9111);
and U10456 (N_10456,N_8554,N_8161);
nor U10457 (N_10457,N_8106,N_9897);
and U10458 (N_10458,N_8375,N_9813);
xor U10459 (N_10459,N_9378,N_8182);
or U10460 (N_10460,N_8001,N_9237);
nand U10461 (N_10461,N_9313,N_8597);
or U10462 (N_10462,N_8666,N_8493);
and U10463 (N_10463,N_8630,N_8915);
nand U10464 (N_10464,N_9375,N_8457);
or U10465 (N_10465,N_9416,N_9838);
and U10466 (N_10466,N_9489,N_9976);
nor U10467 (N_10467,N_9970,N_8429);
nand U10468 (N_10468,N_8139,N_8980);
or U10469 (N_10469,N_8074,N_8083);
and U10470 (N_10470,N_9450,N_8179);
and U10471 (N_10471,N_8757,N_9619);
nand U10472 (N_10472,N_9244,N_9488);
or U10473 (N_10473,N_8513,N_9204);
or U10474 (N_10474,N_9364,N_9213);
nor U10475 (N_10475,N_8563,N_8692);
nand U10476 (N_10476,N_8749,N_9227);
nand U10477 (N_10477,N_9361,N_9481);
nor U10478 (N_10478,N_9998,N_8557);
nand U10479 (N_10479,N_9088,N_8532);
and U10480 (N_10480,N_9700,N_9179);
nand U10481 (N_10481,N_8286,N_8262);
nand U10482 (N_10482,N_9790,N_9491);
nand U10483 (N_10483,N_8843,N_9929);
nand U10484 (N_10484,N_9475,N_9216);
nor U10485 (N_10485,N_9280,N_8685);
or U10486 (N_10486,N_9629,N_9064);
or U10487 (N_10487,N_8280,N_9281);
nor U10488 (N_10488,N_8208,N_9330);
or U10489 (N_10489,N_8593,N_8905);
nor U10490 (N_10490,N_8396,N_9164);
nand U10491 (N_10491,N_8601,N_8726);
nor U10492 (N_10492,N_8400,N_8585);
nand U10493 (N_10493,N_8896,N_9393);
nor U10494 (N_10494,N_9262,N_9722);
nand U10495 (N_10495,N_9715,N_8349);
and U10496 (N_10496,N_8553,N_9633);
nor U10497 (N_10497,N_9638,N_8564);
nor U10498 (N_10498,N_8998,N_9529);
or U10499 (N_10499,N_9385,N_8171);
and U10500 (N_10500,N_8394,N_8565);
or U10501 (N_10501,N_9047,N_9307);
nor U10502 (N_10502,N_9229,N_8160);
or U10503 (N_10503,N_9987,N_8501);
nand U10504 (N_10504,N_9110,N_9660);
nand U10505 (N_10505,N_9869,N_9719);
nor U10506 (N_10506,N_8405,N_8234);
nor U10507 (N_10507,N_8303,N_8148);
and U10508 (N_10508,N_8906,N_9428);
nand U10509 (N_10509,N_9654,N_9399);
nor U10510 (N_10510,N_9526,N_8516);
or U10511 (N_10511,N_8615,N_8912);
nand U10512 (N_10512,N_8305,N_8787);
nor U10513 (N_10513,N_9017,N_8489);
or U10514 (N_10514,N_8274,N_8239);
and U10515 (N_10515,N_8119,N_9034);
xnor U10516 (N_10516,N_8928,N_8972);
or U10517 (N_10517,N_8804,N_9882);
nand U10518 (N_10518,N_8817,N_8545);
nand U10519 (N_10519,N_8096,N_9621);
nor U10520 (N_10520,N_8430,N_9938);
nand U10521 (N_10521,N_8885,N_8045);
and U10522 (N_10522,N_8616,N_9697);
nand U10523 (N_10523,N_9402,N_9057);
xor U10524 (N_10524,N_9168,N_8604);
nor U10525 (N_10525,N_8406,N_8397);
nand U10526 (N_10526,N_8462,N_9567);
and U10527 (N_10527,N_8027,N_8542);
nor U10528 (N_10528,N_8423,N_9170);
nand U10529 (N_10529,N_8622,N_9470);
nand U10530 (N_10530,N_8009,N_8450);
and U10531 (N_10531,N_9175,N_8698);
nor U10532 (N_10532,N_9657,N_8684);
nand U10533 (N_10533,N_8107,N_8242);
nand U10534 (N_10534,N_9849,N_9504);
nand U10535 (N_10535,N_9832,N_9022);
nor U10536 (N_10536,N_8957,N_8871);
or U10537 (N_10537,N_8263,N_8936);
and U10538 (N_10538,N_9535,N_9182);
nand U10539 (N_10539,N_9209,N_8947);
and U10540 (N_10540,N_9860,N_8898);
nor U10541 (N_10541,N_9040,N_8216);
or U10542 (N_10542,N_8458,N_9339);
nor U10543 (N_10543,N_9785,N_8230);
nor U10544 (N_10544,N_9665,N_8385);
and U10545 (N_10545,N_9809,N_8308);
or U10546 (N_10546,N_9997,N_9743);
and U10547 (N_10547,N_8358,N_8993);
and U10548 (N_10548,N_8649,N_8530);
nor U10549 (N_10549,N_9635,N_9383);
xor U10550 (N_10550,N_8958,N_8244);
nor U10551 (N_10551,N_9277,N_8699);
nand U10552 (N_10552,N_8012,N_8660);
or U10553 (N_10553,N_8095,N_9095);
and U10554 (N_10554,N_9835,N_8747);
and U10555 (N_10555,N_8151,N_9391);
or U10556 (N_10556,N_8093,N_8582);
nor U10557 (N_10557,N_9033,N_8386);
nand U10558 (N_10558,N_9589,N_8655);
or U10559 (N_10559,N_8053,N_9300);
and U10560 (N_10560,N_9433,N_9321);
and U10561 (N_10561,N_9085,N_9254);
nand U10562 (N_10562,N_9020,N_8296);
nor U10563 (N_10563,N_9144,N_8060);
and U10564 (N_10564,N_9751,N_8612);
nor U10565 (N_10565,N_8577,N_9979);
nand U10566 (N_10566,N_8084,N_9713);
nand U10567 (N_10567,N_8890,N_9980);
nand U10568 (N_10568,N_9927,N_8946);
or U10569 (N_10569,N_8143,N_9113);
nor U10570 (N_10570,N_8141,N_8719);
or U10571 (N_10571,N_9408,N_9821);
nor U10572 (N_10572,N_9112,N_8835);
or U10573 (N_10573,N_8807,N_8266);
or U10574 (N_10574,N_8866,N_8710);
and U10575 (N_10575,N_8356,N_9054);
nor U10576 (N_10576,N_9266,N_9990);
nor U10577 (N_10577,N_8552,N_9312);
and U10578 (N_10578,N_8741,N_9389);
nand U10579 (N_10579,N_9220,N_9575);
xnor U10580 (N_10580,N_9819,N_9508);
or U10581 (N_10581,N_9426,N_9173);
nand U10582 (N_10582,N_8277,N_8619);
and U10583 (N_10583,N_9464,N_8940);
or U10584 (N_10584,N_8733,N_9084);
and U10585 (N_10585,N_9876,N_8857);
nand U10586 (N_10586,N_8531,N_9752);
nor U10587 (N_10587,N_9031,N_9155);
nand U10588 (N_10588,N_9533,N_9292);
nor U10589 (N_10589,N_8892,N_8334);
nand U10590 (N_10590,N_9078,N_8480);
or U10591 (N_10591,N_8529,N_9584);
nand U10592 (N_10592,N_9226,N_9087);
nand U10593 (N_10593,N_9293,N_9230);
and U10594 (N_10594,N_8774,N_9637);
and U10595 (N_10595,N_9841,N_9679);
nand U10596 (N_10596,N_8129,N_8311);
or U10597 (N_10597,N_8078,N_9928);
nand U10598 (N_10598,N_8600,N_9707);
nor U10599 (N_10599,N_9974,N_9400);
nor U10600 (N_10600,N_8070,N_9129);
nand U10601 (N_10601,N_8845,N_8851);
and U10602 (N_10602,N_8981,N_8041);
and U10603 (N_10603,N_9773,N_9653);
or U10604 (N_10604,N_8780,N_9850);
and U10605 (N_10605,N_8241,N_9666);
nor U10606 (N_10606,N_9724,N_8295);
nor U10607 (N_10607,N_8838,N_9314);
or U10608 (N_10608,N_8309,N_8446);
and U10609 (N_10609,N_9585,N_9551);
nand U10610 (N_10610,N_8365,N_9857);
and U10611 (N_10611,N_8080,N_8775);
nor U10612 (N_10612,N_8810,N_8175);
xor U10613 (N_10613,N_8445,N_9873);
and U10614 (N_10614,N_8343,N_8004);
or U10615 (N_10615,N_9951,N_9327);
and U10616 (N_10616,N_9196,N_9687);
nand U10617 (N_10617,N_9319,N_9122);
nand U10618 (N_10618,N_9933,N_9372);
nor U10619 (N_10619,N_8347,N_8181);
nand U10620 (N_10620,N_9712,N_8583);
xor U10621 (N_10621,N_9659,N_9858);
and U10622 (N_10622,N_9225,N_9250);
and U10623 (N_10623,N_9784,N_9032);
nor U10624 (N_10624,N_8377,N_8975);
xor U10625 (N_10625,N_8363,N_9376);
nand U10626 (N_10626,N_9547,N_8739);
nand U10627 (N_10627,N_8275,N_9581);
nand U10628 (N_10628,N_8788,N_8877);
and U10629 (N_10629,N_9082,N_8652);
or U10630 (N_10630,N_8842,N_8276);
and U10631 (N_10631,N_8620,N_8665);
nand U10632 (N_10632,N_8562,N_9000);
nand U10633 (N_10633,N_8645,N_8822);
nor U10634 (N_10634,N_8880,N_9900);
nor U10635 (N_10635,N_9427,N_8589);
nand U10636 (N_10636,N_8578,N_9896);
and U10637 (N_10637,N_9769,N_9124);
nand U10638 (N_10638,N_9077,N_8943);
and U10639 (N_10639,N_9690,N_8651);
or U10640 (N_10640,N_8826,N_8989);
nand U10641 (N_10641,N_9959,N_8669);
nor U10642 (N_10642,N_8523,N_9062);
nor U10643 (N_10643,N_9883,N_8982);
nand U10644 (N_10644,N_8844,N_8413);
nor U10645 (N_10645,N_8475,N_8769);
xnor U10646 (N_10646,N_8361,N_8881);
or U10647 (N_10647,N_9210,N_9801);
nand U10648 (N_10648,N_9381,N_9183);
nand U10649 (N_10649,N_8856,N_8671);
or U10650 (N_10650,N_9701,N_9986);
and U10651 (N_10651,N_8976,N_9296);
nand U10652 (N_10652,N_8911,N_8793);
nor U10653 (N_10653,N_9243,N_8223);
nand U10654 (N_10654,N_8846,N_9070);
and U10655 (N_10655,N_9323,N_8233);
xnor U10656 (N_10656,N_8673,N_9224);
or U10657 (N_10657,N_8210,N_9542);
nor U10658 (N_10658,N_8590,N_9317);
nand U10659 (N_10659,N_8082,N_9797);
nor U10660 (N_10660,N_8304,N_9678);
and U10661 (N_10661,N_8294,N_9068);
or U10662 (N_10662,N_9457,N_8617);
nor U10663 (N_10663,N_8109,N_9693);
nand U10664 (N_10664,N_8068,N_9125);
and U10665 (N_10665,N_8672,N_8588);
or U10666 (N_10666,N_8197,N_9406);
or U10667 (N_10667,N_8732,N_9904);
and U10668 (N_10668,N_9612,N_8721);
xor U10669 (N_10669,N_9771,N_9018);
nor U10670 (N_10670,N_8907,N_9671);
or U10671 (N_10671,N_9071,N_8674);
and U10672 (N_10672,N_8746,N_8034);
and U10673 (N_10673,N_8816,N_8177);
and U10674 (N_10674,N_9174,N_8963);
nand U10675 (N_10675,N_9272,N_8195);
xnor U10676 (N_10676,N_9343,N_8087);
xnor U10677 (N_10677,N_9962,N_9992);
xnor U10678 (N_10678,N_8185,N_8372);
nor U10679 (N_10679,N_8527,N_8790);
nor U10680 (N_10680,N_8099,N_9476);
nor U10681 (N_10681,N_9610,N_8676);
and U10682 (N_10682,N_8609,N_8840);
and U10683 (N_10683,N_9445,N_8144);
and U10684 (N_10684,N_8661,N_8965);
nand U10685 (N_10685,N_9318,N_9246);
xnor U10686 (N_10686,N_9388,N_9674);
and U10687 (N_10687,N_8188,N_8425);
and U10688 (N_10688,N_8298,N_9573);
nor U10689 (N_10689,N_9668,N_9380);
xnor U10690 (N_10690,N_8289,N_9157);
or U10691 (N_10691,N_8265,N_9855);
nor U10692 (N_10692,N_9728,N_9223);
or U10693 (N_10693,N_8778,N_8247);
nand U10694 (N_10694,N_9191,N_8944);
or U10695 (N_10695,N_9745,N_9178);
nor U10696 (N_10696,N_9207,N_8252);
or U10697 (N_10697,N_8222,N_9727);
nor U10698 (N_10698,N_8570,N_8598);
nand U10699 (N_10699,N_9487,N_9358);
nand U10700 (N_10700,N_8364,N_8473);
and U10701 (N_10701,N_9063,N_8654);
xor U10702 (N_10702,N_8110,N_9968);
nor U10703 (N_10703,N_9276,N_9412);
and U10704 (N_10704,N_9609,N_8481);
and U10705 (N_10705,N_9935,N_8688);
and U10706 (N_10706,N_8258,N_8007);
nor U10707 (N_10707,N_9044,N_8426);
and U10708 (N_10708,N_8333,N_8031);
nor U10709 (N_10709,N_8486,N_9322);
or U10710 (N_10710,N_9924,N_8760);
and U10711 (N_10711,N_9720,N_8868);
and U10712 (N_10712,N_8558,N_8163);
and U10713 (N_10713,N_9325,N_9603);
and U10714 (N_10714,N_8003,N_8854);
nand U10715 (N_10715,N_8049,N_8454);
and U10716 (N_10716,N_9744,N_8728);
and U10717 (N_10717,N_8801,N_9362);
nand U10718 (N_10718,N_8014,N_9411);
xor U10719 (N_10719,N_8113,N_9395);
nand U10720 (N_10720,N_8556,N_8814);
nand U10721 (N_10721,N_9232,N_8032);
and U10722 (N_10722,N_9615,N_9926);
nand U10723 (N_10723,N_9907,N_9236);
and U10724 (N_10724,N_8951,N_8919);
and U10725 (N_10725,N_8316,N_8882);
or U10726 (N_10726,N_8534,N_8419);
and U10727 (N_10727,N_9275,N_8902);
or U10728 (N_10728,N_9788,N_8094);
nand U10729 (N_10729,N_9822,N_9248);
nor U10730 (N_10730,N_9762,N_9803);
and U10731 (N_10731,N_8176,N_8878);
nand U10732 (N_10732,N_8398,N_9159);
and U10733 (N_10733,N_8191,N_9705);
nor U10734 (N_10734,N_9652,N_8142);
nand U10735 (N_10735,N_8704,N_9121);
nand U10736 (N_10736,N_9692,N_9954);
xor U10737 (N_10737,N_9828,N_8572);
or U10738 (N_10738,N_8547,N_8777);
or U10739 (N_10739,N_9710,N_9439);
and U10740 (N_10740,N_8920,N_8342);
and U10741 (N_10741,N_8000,N_9847);
xnor U10742 (N_10742,N_9571,N_8808);
nor U10743 (N_10743,N_8091,N_9669);
or U10744 (N_10744,N_8490,N_8504);
nand U10745 (N_10745,N_9749,N_9639);
nand U10746 (N_10746,N_9578,N_8401);
or U10747 (N_10747,N_9245,N_8574);
and U10748 (N_10748,N_9899,N_8753);
nor U10749 (N_10749,N_9734,N_8752);
and U10750 (N_10750,N_9563,N_8125);
xnor U10751 (N_10751,N_9906,N_9046);
nand U10752 (N_10752,N_9469,N_8567);
or U10753 (N_10753,N_8792,N_9677);
or U10754 (N_10754,N_8069,N_9158);
or U10755 (N_10755,N_8517,N_9825);
or U10756 (N_10756,N_8341,N_9334);
or U10757 (N_10757,N_9947,N_9397);
nand U10758 (N_10758,N_9553,N_9648);
nor U10759 (N_10759,N_9572,N_9520);
or U10760 (N_10760,N_9163,N_8236);
nor U10761 (N_10761,N_9753,N_9195);
nand U10762 (N_10762,N_9417,N_8850);
nand U10763 (N_10763,N_8602,N_8948);
nor U10764 (N_10764,N_9409,N_9295);
nand U10765 (N_10765,N_8959,N_8511);
or U10766 (N_10766,N_9811,N_8498);
nand U10767 (N_10767,N_9495,N_8670);
nor U10768 (N_10768,N_8279,N_9943);
or U10769 (N_10769,N_9152,N_8725);
nor U10770 (N_10770,N_8441,N_8020);
nand U10771 (N_10771,N_9234,N_9837);
nand U10772 (N_10772,N_8497,N_8500);
nand U10773 (N_10773,N_8121,N_9502);
nor U10774 (N_10774,N_8611,N_8492);
or U10775 (N_10775,N_9002,N_8971);
or U10776 (N_10776,N_9901,N_8131);
nor U10777 (N_10777,N_9186,N_9308);
nand U10778 (N_10778,N_8650,N_9739);
nand U10779 (N_10779,N_8221,N_9871);
nor U10780 (N_10780,N_9029,N_9975);
and U10781 (N_10781,N_9776,N_9732);
and U10782 (N_10782,N_8536,N_8596);
nor U10783 (N_10783,N_9141,N_9461);
nor U10784 (N_10784,N_9377,N_8935);
or U10785 (N_10785,N_9350,N_9468);
and U10786 (N_10786,N_8648,N_9123);
nor U10787 (N_10787,N_9590,N_8929);
or U10788 (N_10788,N_9118,N_8639);
and U10789 (N_10789,N_9631,N_8022);
nand U10790 (N_10790,N_8283,N_8576);
or U10791 (N_10791,N_9463,N_8528);
or U10792 (N_10792,N_9026,N_9498);
xnor U10793 (N_10793,N_9370,N_9360);
nor U10794 (N_10794,N_8950,N_9303);
and U10795 (N_10795,N_8938,N_9239);
nand U10796 (N_10796,N_9767,N_9492);
or U10797 (N_10797,N_8874,N_8061);
and U10798 (N_10798,N_8062,N_8524);
nand U10799 (N_10799,N_8474,N_8290);
nor U10800 (N_10800,N_9131,N_9448);
or U10801 (N_10801,N_9212,N_8089);
and U10802 (N_10802,N_8821,N_9166);
and U10803 (N_10803,N_8237,N_8862);
or U10804 (N_10804,N_9561,N_9076);
nor U10805 (N_10805,N_9190,N_9748);
and U10806 (N_10806,N_9452,N_9382);
and U10807 (N_10807,N_9913,N_9939);
nor U10808 (N_10808,N_8367,N_8246);
nor U10809 (N_10809,N_9038,N_8202);
xor U10810 (N_10810,N_8056,N_8090);
nand U10811 (N_10811,N_9289,N_8985);
nor U10812 (N_10812,N_9989,N_9148);
nand U10813 (N_10813,N_9810,N_9562);
nor U10814 (N_10814,N_9499,N_8707);
and U10815 (N_10815,N_9651,N_8984);
and U10816 (N_10816,N_9379,N_9203);
and U10817 (N_10817,N_8848,N_9049);
and U10818 (N_10818,N_9859,N_8154);
and U10819 (N_10819,N_9298,N_8795);
or U10820 (N_10820,N_9341,N_8477);
and U10821 (N_10821,N_8066,N_8173);
nand U10822 (N_10822,N_8680,N_9731);
and U10823 (N_10823,N_9079,N_9996);
or U10824 (N_10824,N_8248,N_8434);
or U10825 (N_10825,N_9946,N_9948);
or U10826 (N_10826,N_9403,N_9119);
nor U10827 (N_10827,N_9898,N_8559);
and U10828 (N_10828,N_8521,N_9404);
nor U10829 (N_10829,N_8996,N_9845);
nand U10830 (N_10830,N_9917,N_8973);
and U10831 (N_10831,N_8165,N_8135);
nor U10832 (N_10832,N_8496,N_8942);
or U10833 (N_10833,N_8114,N_8768);
nand U10834 (N_10834,N_9061,N_8264);
and U10835 (N_10835,N_9349,N_9067);
xor U10836 (N_10836,N_9783,N_8460);
or U10837 (N_10837,N_8653,N_8949);
nor U10838 (N_10838,N_8312,N_9757);
or U10839 (N_10839,N_9923,N_9862);
and U10840 (N_10840,N_8488,N_9950);
nor U10841 (N_10841,N_9747,N_9456);
xnor U10842 (N_10842,N_9866,N_9726);
nor U10843 (N_10843,N_8327,N_8204);
nand U10844 (N_10844,N_9761,N_9620);
nor U10845 (N_10845,N_8421,N_8085);
xor U10846 (N_10846,N_9027,N_8858);
nand U10847 (N_10847,N_8422,N_8873);
nand U10848 (N_10848,N_8863,N_9035);
and U10849 (N_10849,N_8717,N_9703);
and U10850 (N_10850,N_8812,N_8724);
and U10851 (N_10851,N_9706,N_8123);
nor U10852 (N_10852,N_8614,N_9249);
or U10853 (N_10853,N_8499,N_9493);
xnor U10854 (N_10854,N_8503,N_9650);
nor U10855 (N_10855,N_8201,N_9114);
nor U10856 (N_10856,N_9673,N_8152);
nand U10857 (N_10857,N_8253,N_8969);
xor U10858 (N_10858,N_8522,N_8366);
or U10859 (N_10859,N_8159,N_8580);
nand U10860 (N_10860,N_8081,N_9052);
and U10861 (N_10861,N_9834,N_8251);
xnor U10862 (N_10862,N_9577,N_8968);
nor U10863 (N_10863,N_8727,N_8150);
or U10864 (N_10864,N_9750,N_9587);
nand U10865 (N_10865,N_9875,N_8766);
nand U10866 (N_10866,N_8595,N_8633);
nor U10867 (N_10867,N_9945,N_8581);
nor U10868 (N_10868,N_9482,N_9816);
or U10869 (N_10869,N_9787,N_8694);
and U10870 (N_10870,N_9501,N_9471);
and U10871 (N_10871,N_9324,N_9999);
or U10872 (N_10872,N_8791,N_8369);
nand U10873 (N_10873,N_8573,N_9546);
and U10874 (N_10874,N_9287,N_8050);
nor U10875 (N_10875,N_9798,N_9430);
nor U10876 (N_10876,N_8449,N_8267);
nor U10877 (N_10877,N_8834,N_8491);
nor U10878 (N_10878,N_8895,N_8550);
nor U10879 (N_10879,N_9193,N_8864);
and U10880 (N_10880,N_9415,N_8977);
or U10881 (N_10881,N_9453,N_8627);
nor U10882 (N_10882,N_9133,N_8436);
and U10883 (N_10883,N_9101,N_8930);
and U10884 (N_10884,N_8409,N_8021);
xnor U10885 (N_10885,N_9760,N_9496);
or U10886 (N_10886,N_8744,N_8507);
nor U10887 (N_10887,N_9007,N_9579);
nand U10888 (N_10888,N_9683,N_9282);
nor U10889 (N_10889,N_8626,N_9944);
or U10890 (N_10890,N_9552,N_9242);
and U10891 (N_10891,N_8158,N_8416);
nand U10892 (N_10892,N_8393,N_9709);
nand U10893 (N_10893,N_9556,N_9267);
nand U10894 (N_10894,N_9443,N_8013);
nor U10895 (N_10895,N_8824,N_9691);
nand U10896 (N_10896,N_8037,N_9483);
xor U10897 (N_10897,N_9284,N_8301);
nor U10898 (N_10898,N_9255,N_8149);
nor U10899 (N_10899,N_9774,N_8689);
or U10900 (N_10900,N_8805,N_8472);
and U10901 (N_10901,N_9132,N_9887);
nor U10902 (N_10902,N_9103,N_9741);
and U10903 (N_10903,N_9839,N_9446);
nor U10904 (N_10904,N_8200,N_9564);
and U10905 (N_10905,N_9093,N_8909);
and U10906 (N_10906,N_8224,N_9135);
nor U10907 (N_10907,N_9065,N_8193);
or U10908 (N_10908,N_8086,N_9854);
nor U10909 (N_10909,N_8641,N_9754);
nand U10910 (N_10910,N_9777,N_9985);
and U10911 (N_10911,N_9465,N_8642);
nor U10912 (N_10912,N_8773,N_9240);
and U10913 (N_10913,N_9172,N_9257);
nor U10914 (N_10914,N_9420,N_8415);
and U10915 (N_10915,N_8285,N_8133);
and U10916 (N_10916,N_9877,N_8751);
nor U10917 (N_10917,N_9138,N_8097);
or U10918 (N_10918,N_9914,N_8631);
and U10919 (N_10919,N_8103,N_9073);
nand U10920 (N_10920,N_9407,N_8213);
nor U10921 (N_10921,N_9405,N_8353);
and U10922 (N_10922,N_9600,N_9879);
or U10923 (N_10923,N_8451,N_8468);
or U10924 (N_10924,N_9094,N_9647);
or U10925 (N_10925,N_8010,N_8297);
and U10926 (N_10926,N_9480,N_8709);
or U10927 (N_10927,N_8647,N_8225);
nand U10928 (N_10928,N_9060,N_8331);
and U10929 (N_10929,N_8318,N_8315);
nor U10930 (N_10930,N_9137,N_9656);
and U10931 (N_10931,N_8592,N_8028);
and U10932 (N_10932,N_9238,N_9200);
nand U10933 (N_10933,N_8391,N_9942);
nor U10934 (N_10934,N_9804,N_9030);
and U10935 (N_10935,N_9625,N_9202);
or U10936 (N_10936,N_8164,N_8392);
xor U10937 (N_10937,N_8278,N_8025);
xnor U10938 (N_10938,N_8785,N_9301);
or U10939 (N_10939,N_9548,N_8378);
and U10940 (N_10940,N_8718,N_8384);
nand U10941 (N_10941,N_8770,N_8883);
or U10942 (N_10942,N_8510,N_8859);
nand U10943 (N_10943,N_9969,N_9737);
xor U10944 (N_10944,N_8606,N_8138);
xnor U10945 (N_10945,N_9363,N_8852);
or U10946 (N_10946,N_8120,N_9538);
nor U10947 (N_10947,N_8656,N_8743);
and U10948 (N_10948,N_8783,N_9768);
and U10949 (N_10949,N_8412,N_9806);
nand U10950 (N_10950,N_9083,N_9013);
nor U10951 (N_10951,N_8952,N_8758);
or U10952 (N_10952,N_8348,N_8762);
nor U10953 (N_10953,N_8693,N_9524);
nand U10954 (N_10954,N_9830,N_8189);
nand U10955 (N_10955,N_9306,N_8039);
and U10956 (N_10956,N_9623,N_8629);
and U10957 (N_10957,N_8643,N_8104);
nor U10958 (N_10958,N_9878,N_8402);
and U10959 (N_10959,N_9074,N_8714);
xnor U10960 (N_10960,N_8667,N_9218);
or U10961 (N_10961,N_8437,N_9795);
nand U10962 (N_10962,N_9472,N_9003);
nor U10963 (N_10963,N_9894,N_8569);
nand U10964 (N_10964,N_9764,N_8017);
nand U10965 (N_10965,N_8194,N_8127);
nand U10966 (N_10966,N_9269,N_8962);
or U10967 (N_10967,N_8723,N_9918);
nand U10968 (N_10968,N_8115,N_8448);
nor U10969 (N_10969,N_9043,N_8136);
and U10970 (N_10970,N_8029,N_9265);
nand U10971 (N_10971,N_9995,N_9611);
and U10972 (N_10972,N_8453,N_9756);
or U10973 (N_10973,N_9908,N_9885);
nor U10974 (N_10974,N_9522,N_9916);
nand U10975 (N_10975,N_9458,N_9429);
nand U10976 (N_10976,N_9836,N_8229);
or U10977 (N_10977,N_9366,N_9688);
nor U10978 (N_10978,N_8382,N_8260);
nor U10979 (N_10979,N_9256,N_9390);
nand U10980 (N_10980,N_8383,N_9386);
or U10981 (N_10981,N_9605,N_9348);
nor U10982 (N_10982,N_9156,N_9288);
and U10983 (N_10983,N_9336,N_8122);
and U10984 (N_10984,N_8683,N_8742);
nand U10985 (N_10985,N_9418,N_8469);
xor U10986 (N_10986,N_9294,N_8875);
or U10987 (N_10987,N_9441,N_9613);
nor U10988 (N_10988,N_9259,N_9466);
and U10989 (N_10989,N_9422,N_8506);
and U10990 (N_10990,N_8964,N_8900);
nand U10991 (N_10991,N_9290,N_8668);
nand U10992 (N_10992,N_8314,N_8281);
or U10993 (N_10993,N_9817,N_8231);
nor U10994 (N_10994,N_9983,N_8677);
or U10995 (N_10995,N_8897,N_8190);
nor U10996 (N_10996,N_9351,N_8432);
or U10997 (N_10997,N_8459,N_8544);
and U10998 (N_10998,N_9274,N_8664);
nor U10999 (N_10999,N_9758,N_9643);
and U11000 (N_11000,N_9700,N_9048);
or U11001 (N_11001,N_8056,N_8075);
or U11002 (N_11002,N_8333,N_9147);
and U11003 (N_11003,N_9076,N_9700);
nor U11004 (N_11004,N_8751,N_9752);
nand U11005 (N_11005,N_9507,N_8881);
nor U11006 (N_11006,N_8223,N_9036);
or U11007 (N_11007,N_9860,N_9322);
or U11008 (N_11008,N_9391,N_8352);
nor U11009 (N_11009,N_8754,N_8876);
and U11010 (N_11010,N_8498,N_8932);
nand U11011 (N_11011,N_8122,N_9219);
or U11012 (N_11012,N_9702,N_8012);
nor U11013 (N_11013,N_9027,N_9433);
nand U11014 (N_11014,N_9929,N_8013);
nor U11015 (N_11015,N_9830,N_9893);
or U11016 (N_11016,N_8326,N_9355);
or U11017 (N_11017,N_8063,N_8740);
and U11018 (N_11018,N_8497,N_8999);
and U11019 (N_11019,N_9791,N_9803);
nand U11020 (N_11020,N_9163,N_9931);
and U11021 (N_11021,N_8124,N_9881);
nand U11022 (N_11022,N_8747,N_9839);
and U11023 (N_11023,N_8524,N_9220);
nor U11024 (N_11024,N_9936,N_9803);
nor U11025 (N_11025,N_9874,N_9840);
xor U11026 (N_11026,N_9148,N_9283);
nor U11027 (N_11027,N_8835,N_9324);
and U11028 (N_11028,N_8948,N_8376);
nand U11029 (N_11029,N_9981,N_9966);
xor U11030 (N_11030,N_9239,N_9436);
nor U11031 (N_11031,N_8272,N_9860);
and U11032 (N_11032,N_8586,N_9417);
and U11033 (N_11033,N_9944,N_9240);
nor U11034 (N_11034,N_8396,N_9523);
nor U11035 (N_11035,N_8034,N_9112);
xnor U11036 (N_11036,N_8241,N_8293);
nand U11037 (N_11037,N_8660,N_9108);
or U11038 (N_11038,N_9734,N_8089);
and U11039 (N_11039,N_9774,N_9429);
nand U11040 (N_11040,N_9395,N_9470);
and U11041 (N_11041,N_8390,N_8443);
and U11042 (N_11042,N_8373,N_9441);
or U11043 (N_11043,N_9960,N_9959);
nor U11044 (N_11044,N_8878,N_9329);
nor U11045 (N_11045,N_9775,N_8639);
nor U11046 (N_11046,N_8648,N_8934);
nor U11047 (N_11047,N_9046,N_9803);
and U11048 (N_11048,N_9678,N_8275);
or U11049 (N_11049,N_8506,N_8155);
nor U11050 (N_11050,N_8575,N_9105);
nor U11051 (N_11051,N_8039,N_9390);
and U11052 (N_11052,N_9240,N_8289);
nand U11053 (N_11053,N_8075,N_8116);
or U11054 (N_11054,N_8378,N_9118);
or U11055 (N_11055,N_8856,N_9223);
nand U11056 (N_11056,N_8404,N_8577);
or U11057 (N_11057,N_9759,N_8368);
or U11058 (N_11058,N_9465,N_9046);
xnor U11059 (N_11059,N_9154,N_9550);
nand U11060 (N_11060,N_9913,N_9821);
nor U11061 (N_11061,N_8708,N_8309);
and U11062 (N_11062,N_9661,N_8362);
and U11063 (N_11063,N_8034,N_9532);
nand U11064 (N_11064,N_8219,N_9154);
and U11065 (N_11065,N_9225,N_8001);
and U11066 (N_11066,N_9356,N_9937);
nor U11067 (N_11067,N_8507,N_9929);
and U11068 (N_11068,N_9439,N_8633);
or U11069 (N_11069,N_8513,N_8094);
nand U11070 (N_11070,N_8046,N_9554);
or U11071 (N_11071,N_8901,N_9063);
and U11072 (N_11072,N_8159,N_9302);
or U11073 (N_11073,N_9255,N_8409);
or U11074 (N_11074,N_9180,N_9216);
and U11075 (N_11075,N_9489,N_9723);
or U11076 (N_11076,N_9491,N_8918);
nor U11077 (N_11077,N_8080,N_9804);
or U11078 (N_11078,N_8200,N_9773);
nor U11079 (N_11079,N_8038,N_8029);
nor U11080 (N_11080,N_9262,N_9047);
nand U11081 (N_11081,N_9917,N_8373);
or U11082 (N_11082,N_9250,N_9027);
and U11083 (N_11083,N_8204,N_9097);
nand U11084 (N_11084,N_9587,N_9675);
xnor U11085 (N_11085,N_9878,N_9269);
nor U11086 (N_11086,N_8945,N_9875);
nand U11087 (N_11087,N_9069,N_8142);
nor U11088 (N_11088,N_8505,N_9400);
nand U11089 (N_11089,N_9273,N_9931);
or U11090 (N_11090,N_9958,N_8998);
nor U11091 (N_11091,N_9739,N_8884);
nor U11092 (N_11092,N_8951,N_9003);
nand U11093 (N_11093,N_8093,N_9352);
and U11094 (N_11094,N_9810,N_9732);
or U11095 (N_11095,N_9779,N_9081);
or U11096 (N_11096,N_8008,N_9179);
or U11097 (N_11097,N_9820,N_9111);
and U11098 (N_11098,N_9809,N_9188);
xnor U11099 (N_11099,N_8560,N_9668);
xnor U11100 (N_11100,N_9686,N_9742);
or U11101 (N_11101,N_9370,N_9069);
and U11102 (N_11102,N_9330,N_8037);
or U11103 (N_11103,N_9624,N_8195);
xnor U11104 (N_11104,N_8848,N_8980);
and U11105 (N_11105,N_9813,N_8728);
nand U11106 (N_11106,N_8348,N_8345);
nor U11107 (N_11107,N_9796,N_9694);
and U11108 (N_11108,N_8429,N_9379);
nand U11109 (N_11109,N_8740,N_9959);
and U11110 (N_11110,N_9400,N_8787);
or U11111 (N_11111,N_9264,N_9200);
xor U11112 (N_11112,N_9435,N_9734);
and U11113 (N_11113,N_8480,N_8075);
xor U11114 (N_11114,N_9378,N_8087);
and U11115 (N_11115,N_8365,N_8277);
nor U11116 (N_11116,N_8251,N_8768);
nand U11117 (N_11117,N_9614,N_8588);
xor U11118 (N_11118,N_9001,N_9896);
or U11119 (N_11119,N_9260,N_8703);
nand U11120 (N_11120,N_8344,N_9651);
nand U11121 (N_11121,N_9297,N_9204);
and U11122 (N_11122,N_9804,N_8111);
or U11123 (N_11123,N_8228,N_9875);
nor U11124 (N_11124,N_9004,N_8254);
nor U11125 (N_11125,N_8168,N_8740);
nand U11126 (N_11126,N_9797,N_8394);
nand U11127 (N_11127,N_8354,N_8864);
nor U11128 (N_11128,N_8536,N_9320);
or U11129 (N_11129,N_8812,N_9065);
nor U11130 (N_11130,N_8329,N_9734);
nand U11131 (N_11131,N_8918,N_9542);
or U11132 (N_11132,N_9198,N_9230);
nor U11133 (N_11133,N_9585,N_8571);
and U11134 (N_11134,N_9708,N_9098);
nand U11135 (N_11135,N_9298,N_8398);
and U11136 (N_11136,N_9882,N_9401);
nor U11137 (N_11137,N_9018,N_9727);
xor U11138 (N_11138,N_8625,N_8368);
nor U11139 (N_11139,N_9377,N_9967);
nand U11140 (N_11140,N_9230,N_9141);
xnor U11141 (N_11141,N_8865,N_8550);
nand U11142 (N_11142,N_8031,N_9954);
and U11143 (N_11143,N_9772,N_8438);
and U11144 (N_11144,N_8142,N_8479);
nor U11145 (N_11145,N_9529,N_8182);
and U11146 (N_11146,N_8818,N_8572);
and U11147 (N_11147,N_8391,N_8240);
xnor U11148 (N_11148,N_9612,N_9772);
xnor U11149 (N_11149,N_8415,N_9722);
nand U11150 (N_11150,N_9896,N_9446);
nand U11151 (N_11151,N_9261,N_8818);
or U11152 (N_11152,N_9826,N_9013);
nor U11153 (N_11153,N_9475,N_9418);
nand U11154 (N_11154,N_9016,N_9351);
and U11155 (N_11155,N_9286,N_9562);
or U11156 (N_11156,N_9306,N_9810);
xor U11157 (N_11157,N_8689,N_9263);
nand U11158 (N_11158,N_9941,N_8792);
nand U11159 (N_11159,N_8623,N_8211);
nand U11160 (N_11160,N_9831,N_8027);
or U11161 (N_11161,N_9185,N_9755);
nor U11162 (N_11162,N_8514,N_9593);
nor U11163 (N_11163,N_8976,N_9942);
and U11164 (N_11164,N_8852,N_8162);
nor U11165 (N_11165,N_8239,N_9026);
and U11166 (N_11166,N_9583,N_9219);
nor U11167 (N_11167,N_8852,N_9313);
nand U11168 (N_11168,N_8448,N_9370);
and U11169 (N_11169,N_8943,N_8669);
and U11170 (N_11170,N_8739,N_9912);
or U11171 (N_11171,N_9147,N_9637);
and U11172 (N_11172,N_8784,N_8366);
xor U11173 (N_11173,N_8369,N_8946);
and U11174 (N_11174,N_9735,N_9053);
xnor U11175 (N_11175,N_9552,N_9187);
and U11176 (N_11176,N_8202,N_8756);
nor U11177 (N_11177,N_8612,N_9905);
and U11178 (N_11178,N_9270,N_8314);
or U11179 (N_11179,N_8556,N_9481);
and U11180 (N_11180,N_8148,N_9539);
nand U11181 (N_11181,N_9146,N_8060);
or U11182 (N_11182,N_8701,N_8939);
or U11183 (N_11183,N_8172,N_9921);
nand U11184 (N_11184,N_9117,N_9643);
nor U11185 (N_11185,N_9149,N_9652);
xnor U11186 (N_11186,N_8981,N_8128);
or U11187 (N_11187,N_8607,N_9918);
nand U11188 (N_11188,N_8089,N_8092);
nand U11189 (N_11189,N_8531,N_9596);
nand U11190 (N_11190,N_9807,N_8024);
xor U11191 (N_11191,N_8174,N_9733);
nor U11192 (N_11192,N_9393,N_9236);
nor U11193 (N_11193,N_8254,N_8491);
and U11194 (N_11194,N_9960,N_9408);
and U11195 (N_11195,N_9555,N_9352);
nor U11196 (N_11196,N_9232,N_8027);
nor U11197 (N_11197,N_9327,N_8025);
nand U11198 (N_11198,N_9553,N_9717);
or U11199 (N_11199,N_9794,N_9186);
nor U11200 (N_11200,N_8647,N_8323);
and U11201 (N_11201,N_8318,N_8823);
nand U11202 (N_11202,N_9522,N_9691);
or U11203 (N_11203,N_9890,N_9111);
and U11204 (N_11204,N_9612,N_8733);
and U11205 (N_11205,N_9811,N_9568);
nor U11206 (N_11206,N_8806,N_8148);
nand U11207 (N_11207,N_8947,N_9795);
and U11208 (N_11208,N_8035,N_9032);
nor U11209 (N_11209,N_8436,N_9600);
nor U11210 (N_11210,N_8628,N_9145);
xor U11211 (N_11211,N_8101,N_9184);
nand U11212 (N_11212,N_8897,N_9476);
or U11213 (N_11213,N_9256,N_9430);
nor U11214 (N_11214,N_9998,N_8205);
xnor U11215 (N_11215,N_9653,N_8317);
nor U11216 (N_11216,N_8551,N_9236);
nand U11217 (N_11217,N_8827,N_9836);
or U11218 (N_11218,N_8116,N_8944);
nor U11219 (N_11219,N_8289,N_9145);
nor U11220 (N_11220,N_9734,N_8623);
or U11221 (N_11221,N_8426,N_8451);
or U11222 (N_11222,N_8902,N_8145);
nand U11223 (N_11223,N_9764,N_9716);
or U11224 (N_11224,N_8270,N_9869);
or U11225 (N_11225,N_9409,N_9825);
and U11226 (N_11226,N_8405,N_9226);
or U11227 (N_11227,N_9099,N_8533);
nor U11228 (N_11228,N_9509,N_9212);
nor U11229 (N_11229,N_9900,N_8076);
nor U11230 (N_11230,N_8917,N_9959);
or U11231 (N_11231,N_8817,N_8872);
or U11232 (N_11232,N_8398,N_8903);
nor U11233 (N_11233,N_9375,N_8592);
or U11234 (N_11234,N_8031,N_8418);
xor U11235 (N_11235,N_8717,N_9745);
or U11236 (N_11236,N_9554,N_8874);
and U11237 (N_11237,N_8773,N_9034);
and U11238 (N_11238,N_8835,N_9598);
or U11239 (N_11239,N_9732,N_8082);
and U11240 (N_11240,N_9604,N_9844);
nand U11241 (N_11241,N_9834,N_9254);
xnor U11242 (N_11242,N_9822,N_9771);
nor U11243 (N_11243,N_9623,N_8237);
and U11244 (N_11244,N_8849,N_8154);
and U11245 (N_11245,N_8082,N_8552);
or U11246 (N_11246,N_9178,N_9758);
or U11247 (N_11247,N_8729,N_8559);
or U11248 (N_11248,N_8189,N_8338);
and U11249 (N_11249,N_9504,N_9181);
and U11250 (N_11250,N_9521,N_8985);
and U11251 (N_11251,N_8236,N_8216);
nand U11252 (N_11252,N_9029,N_8384);
xnor U11253 (N_11253,N_9431,N_8271);
nor U11254 (N_11254,N_9291,N_9977);
and U11255 (N_11255,N_9046,N_8825);
nor U11256 (N_11256,N_8099,N_8301);
xnor U11257 (N_11257,N_8131,N_9466);
or U11258 (N_11258,N_9006,N_9693);
and U11259 (N_11259,N_8290,N_9048);
nor U11260 (N_11260,N_9930,N_8791);
nor U11261 (N_11261,N_8585,N_8800);
nand U11262 (N_11262,N_8278,N_8606);
xnor U11263 (N_11263,N_8086,N_8348);
nor U11264 (N_11264,N_8890,N_8613);
xor U11265 (N_11265,N_8171,N_9457);
nand U11266 (N_11266,N_9809,N_9299);
nand U11267 (N_11267,N_8059,N_8634);
or U11268 (N_11268,N_9892,N_9896);
nor U11269 (N_11269,N_9299,N_8113);
nor U11270 (N_11270,N_9260,N_9441);
or U11271 (N_11271,N_9427,N_9069);
or U11272 (N_11272,N_8540,N_8484);
nand U11273 (N_11273,N_9720,N_9174);
and U11274 (N_11274,N_8542,N_8368);
nand U11275 (N_11275,N_9869,N_8419);
xor U11276 (N_11276,N_8288,N_8525);
nand U11277 (N_11277,N_8054,N_8203);
and U11278 (N_11278,N_8169,N_9794);
nand U11279 (N_11279,N_8287,N_8849);
and U11280 (N_11280,N_8500,N_9657);
and U11281 (N_11281,N_8502,N_9712);
or U11282 (N_11282,N_9662,N_9471);
or U11283 (N_11283,N_9647,N_8795);
and U11284 (N_11284,N_8678,N_9917);
nand U11285 (N_11285,N_9543,N_9681);
nand U11286 (N_11286,N_8912,N_8516);
or U11287 (N_11287,N_8077,N_9361);
nand U11288 (N_11288,N_8257,N_8642);
or U11289 (N_11289,N_8367,N_9855);
xor U11290 (N_11290,N_9035,N_8766);
or U11291 (N_11291,N_8411,N_8242);
and U11292 (N_11292,N_9295,N_9697);
or U11293 (N_11293,N_9963,N_9644);
nand U11294 (N_11294,N_9505,N_8790);
nand U11295 (N_11295,N_8956,N_9199);
nand U11296 (N_11296,N_8567,N_8874);
xnor U11297 (N_11297,N_9472,N_8904);
nor U11298 (N_11298,N_9992,N_9730);
nand U11299 (N_11299,N_8373,N_8309);
or U11300 (N_11300,N_8111,N_9566);
nor U11301 (N_11301,N_8303,N_9797);
nand U11302 (N_11302,N_8883,N_8476);
nor U11303 (N_11303,N_8834,N_8975);
or U11304 (N_11304,N_9888,N_8642);
nand U11305 (N_11305,N_8850,N_8325);
nor U11306 (N_11306,N_8051,N_9254);
or U11307 (N_11307,N_9874,N_8111);
nand U11308 (N_11308,N_9411,N_9744);
nor U11309 (N_11309,N_8614,N_9955);
nor U11310 (N_11310,N_8352,N_9820);
or U11311 (N_11311,N_8809,N_8713);
or U11312 (N_11312,N_8965,N_9320);
nand U11313 (N_11313,N_8348,N_9084);
or U11314 (N_11314,N_9821,N_9783);
nor U11315 (N_11315,N_9357,N_9142);
nand U11316 (N_11316,N_8714,N_8022);
nand U11317 (N_11317,N_9027,N_8679);
nor U11318 (N_11318,N_9423,N_9178);
or U11319 (N_11319,N_9012,N_9909);
nor U11320 (N_11320,N_9636,N_8859);
nand U11321 (N_11321,N_8945,N_9499);
and U11322 (N_11322,N_9214,N_8601);
xnor U11323 (N_11323,N_9940,N_9804);
xnor U11324 (N_11324,N_8781,N_9356);
and U11325 (N_11325,N_9776,N_9200);
nor U11326 (N_11326,N_8803,N_8726);
nor U11327 (N_11327,N_9414,N_9042);
or U11328 (N_11328,N_8002,N_9149);
or U11329 (N_11329,N_9777,N_9460);
xor U11330 (N_11330,N_8029,N_9626);
xor U11331 (N_11331,N_8544,N_9808);
xnor U11332 (N_11332,N_8051,N_9314);
and U11333 (N_11333,N_9070,N_9991);
or U11334 (N_11334,N_9675,N_9288);
nand U11335 (N_11335,N_9227,N_8830);
xor U11336 (N_11336,N_9794,N_9957);
and U11337 (N_11337,N_8491,N_9736);
nor U11338 (N_11338,N_9666,N_8933);
xnor U11339 (N_11339,N_8230,N_8802);
and U11340 (N_11340,N_9869,N_8163);
or U11341 (N_11341,N_8899,N_9513);
nor U11342 (N_11342,N_8754,N_8263);
xnor U11343 (N_11343,N_9593,N_8484);
and U11344 (N_11344,N_9307,N_9691);
nor U11345 (N_11345,N_8391,N_8460);
xor U11346 (N_11346,N_9120,N_8163);
or U11347 (N_11347,N_9017,N_9052);
and U11348 (N_11348,N_9013,N_8113);
nand U11349 (N_11349,N_8260,N_9700);
xor U11350 (N_11350,N_8648,N_8207);
nand U11351 (N_11351,N_9287,N_9963);
nor U11352 (N_11352,N_8838,N_9967);
or U11353 (N_11353,N_8399,N_9398);
and U11354 (N_11354,N_9914,N_9591);
nand U11355 (N_11355,N_8336,N_8034);
or U11356 (N_11356,N_9669,N_9985);
or U11357 (N_11357,N_8645,N_8477);
nand U11358 (N_11358,N_8791,N_9271);
or U11359 (N_11359,N_8119,N_9661);
nor U11360 (N_11360,N_8180,N_9048);
and U11361 (N_11361,N_9910,N_9995);
or U11362 (N_11362,N_9467,N_8061);
nand U11363 (N_11363,N_8632,N_9199);
and U11364 (N_11364,N_9816,N_9871);
or U11365 (N_11365,N_9995,N_9006);
nand U11366 (N_11366,N_9249,N_9051);
nor U11367 (N_11367,N_9229,N_8378);
and U11368 (N_11368,N_8702,N_8464);
nand U11369 (N_11369,N_8347,N_8189);
nand U11370 (N_11370,N_9483,N_9925);
nor U11371 (N_11371,N_9749,N_9631);
nor U11372 (N_11372,N_8590,N_8678);
xor U11373 (N_11373,N_9046,N_9779);
and U11374 (N_11374,N_8278,N_9804);
nor U11375 (N_11375,N_8198,N_8339);
or U11376 (N_11376,N_9966,N_9843);
and U11377 (N_11377,N_9664,N_9475);
nand U11378 (N_11378,N_9114,N_9869);
or U11379 (N_11379,N_9210,N_8959);
xor U11380 (N_11380,N_8587,N_8602);
nor U11381 (N_11381,N_9775,N_9334);
nor U11382 (N_11382,N_9501,N_9635);
and U11383 (N_11383,N_8952,N_8155);
nor U11384 (N_11384,N_9612,N_9236);
nor U11385 (N_11385,N_9174,N_8586);
and U11386 (N_11386,N_8149,N_9226);
nand U11387 (N_11387,N_9484,N_8848);
or U11388 (N_11388,N_9326,N_9933);
nor U11389 (N_11389,N_8228,N_9818);
nor U11390 (N_11390,N_8542,N_9710);
xor U11391 (N_11391,N_8673,N_8537);
nand U11392 (N_11392,N_8668,N_9602);
and U11393 (N_11393,N_8354,N_8942);
nand U11394 (N_11394,N_9941,N_8842);
nor U11395 (N_11395,N_8691,N_9858);
nor U11396 (N_11396,N_8798,N_9925);
nor U11397 (N_11397,N_8615,N_9783);
nand U11398 (N_11398,N_8090,N_9229);
nand U11399 (N_11399,N_8507,N_9212);
nand U11400 (N_11400,N_9489,N_9928);
and U11401 (N_11401,N_9189,N_9597);
and U11402 (N_11402,N_8179,N_9826);
and U11403 (N_11403,N_9189,N_8899);
or U11404 (N_11404,N_8856,N_9136);
nand U11405 (N_11405,N_9561,N_9187);
nor U11406 (N_11406,N_9830,N_8524);
nand U11407 (N_11407,N_9204,N_8074);
xnor U11408 (N_11408,N_8951,N_8482);
and U11409 (N_11409,N_9102,N_8631);
nand U11410 (N_11410,N_8966,N_9195);
nand U11411 (N_11411,N_9306,N_9572);
xor U11412 (N_11412,N_9086,N_8727);
nor U11413 (N_11413,N_9096,N_8026);
and U11414 (N_11414,N_8495,N_9487);
nand U11415 (N_11415,N_9954,N_9119);
or U11416 (N_11416,N_9097,N_8781);
nand U11417 (N_11417,N_9333,N_9045);
and U11418 (N_11418,N_8291,N_8180);
and U11419 (N_11419,N_8540,N_8343);
nor U11420 (N_11420,N_8999,N_8883);
and U11421 (N_11421,N_8281,N_8106);
xor U11422 (N_11422,N_9881,N_9173);
and U11423 (N_11423,N_8198,N_9271);
nand U11424 (N_11424,N_9505,N_9253);
or U11425 (N_11425,N_9256,N_9285);
nand U11426 (N_11426,N_9766,N_9105);
nor U11427 (N_11427,N_8795,N_9928);
or U11428 (N_11428,N_8547,N_9057);
or U11429 (N_11429,N_9870,N_9383);
xor U11430 (N_11430,N_9129,N_9310);
or U11431 (N_11431,N_9633,N_9350);
or U11432 (N_11432,N_9720,N_8841);
nand U11433 (N_11433,N_9523,N_9761);
nand U11434 (N_11434,N_8830,N_8250);
and U11435 (N_11435,N_8605,N_9462);
nor U11436 (N_11436,N_8717,N_9099);
nand U11437 (N_11437,N_9760,N_9721);
and U11438 (N_11438,N_8304,N_8604);
or U11439 (N_11439,N_8329,N_9286);
and U11440 (N_11440,N_8447,N_9117);
and U11441 (N_11441,N_8921,N_8927);
xnor U11442 (N_11442,N_8980,N_9771);
or U11443 (N_11443,N_9624,N_9874);
xor U11444 (N_11444,N_9733,N_9902);
or U11445 (N_11445,N_8095,N_8462);
nor U11446 (N_11446,N_8306,N_9811);
or U11447 (N_11447,N_8918,N_9722);
nand U11448 (N_11448,N_9207,N_8049);
nand U11449 (N_11449,N_8244,N_8007);
xnor U11450 (N_11450,N_9714,N_9694);
and U11451 (N_11451,N_9985,N_9272);
nand U11452 (N_11452,N_8837,N_8728);
or U11453 (N_11453,N_9370,N_8807);
nand U11454 (N_11454,N_8937,N_9234);
or U11455 (N_11455,N_8252,N_8387);
and U11456 (N_11456,N_9906,N_8898);
and U11457 (N_11457,N_8047,N_8182);
nand U11458 (N_11458,N_8279,N_9365);
nand U11459 (N_11459,N_8673,N_9777);
xnor U11460 (N_11460,N_8438,N_8518);
nand U11461 (N_11461,N_9235,N_9605);
nand U11462 (N_11462,N_9628,N_9282);
nor U11463 (N_11463,N_8161,N_8333);
or U11464 (N_11464,N_9207,N_9700);
nand U11465 (N_11465,N_8288,N_8260);
and U11466 (N_11466,N_8300,N_9882);
or U11467 (N_11467,N_9095,N_8588);
nand U11468 (N_11468,N_9341,N_9749);
or U11469 (N_11469,N_8854,N_8094);
and U11470 (N_11470,N_8300,N_8195);
nor U11471 (N_11471,N_8104,N_9019);
nor U11472 (N_11472,N_9541,N_8055);
or U11473 (N_11473,N_9970,N_8667);
or U11474 (N_11474,N_9509,N_9424);
nand U11475 (N_11475,N_8865,N_9530);
and U11476 (N_11476,N_8749,N_9013);
xnor U11477 (N_11477,N_9603,N_9323);
nor U11478 (N_11478,N_9320,N_9609);
nor U11479 (N_11479,N_9996,N_8646);
and U11480 (N_11480,N_8356,N_9294);
xor U11481 (N_11481,N_8395,N_8146);
and U11482 (N_11482,N_8735,N_9638);
and U11483 (N_11483,N_8895,N_9415);
and U11484 (N_11484,N_9683,N_9314);
or U11485 (N_11485,N_9407,N_8288);
nand U11486 (N_11486,N_8113,N_8111);
nand U11487 (N_11487,N_8428,N_9253);
or U11488 (N_11488,N_9924,N_8236);
or U11489 (N_11489,N_8029,N_9395);
or U11490 (N_11490,N_9747,N_9818);
and U11491 (N_11491,N_8563,N_9345);
xnor U11492 (N_11492,N_9056,N_9279);
and U11493 (N_11493,N_9276,N_8506);
and U11494 (N_11494,N_8632,N_8493);
or U11495 (N_11495,N_9844,N_9382);
nor U11496 (N_11496,N_8424,N_8941);
nor U11497 (N_11497,N_8944,N_8169);
nor U11498 (N_11498,N_8155,N_9551);
and U11499 (N_11499,N_9616,N_9597);
xor U11500 (N_11500,N_9450,N_8481);
nor U11501 (N_11501,N_8871,N_8750);
or U11502 (N_11502,N_8950,N_9721);
nand U11503 (N_11503,N_9726,N_8842);
or U11504 (N_11504,N_9106,N_8983);
nor U11505 (N_11505,N_8491,N_8720);
nand U11506 (N_11506,N_9592,N_8831);
or U11507 (N_11507,N_9686,N_8881);
nor U11508 (N_11508,N_8713,N_9694);
or U11509 (N_11509,N_8969,N_9075);
nor U11510 (N_11510,N_8402,N_8438);
and U11511 (N_11511,N_8540,N_9353);
nand U11512 (N_11512,N_9777,N_8951);
nor U11513 (N_11513,N_8043,N_9335);
or U11514 (N_11514,N_8781,N_8805);
nand U11515 (N_11515,N_8151,N_9090);
and U11516 (N_11516,N_8932,N_8364);
and U11517 (N_11517,N_8256,N_8794);
nand U11518 (N_11518,N_9126,N_9001);
or U11519 (N_11519,N_8747,N_8750);
and U11520 (N_11520,N_8948,N_9223);
and U11521 (N_11521,N_8148,N_9285);
nand U11522 (N_11522,N_8764,N_9189);
or U11523 (N_11523,N_9176,N_9760);
and U11524 (N_11524,N_8741,N_8641);
xnor U11525 (N_11525,N_9326,N_8483);
or U11526 (N_11526,N_8939,N_9339);
and U11527 (N_11527,N_8668,N_9829);
nand U11528 (N_11528,N_8849,N_8834);
nand U11529 (N_11529,N_9069,N_8021);
and U11530 (N_11530,N_8072,N_8448);
or U11531 (N_11531,N_9357,N_8296);
nand U11532 (N_11532,N_9270,N_8412);
and U11533 (N_11533,N_8438,N_9517);
or U11534 (N_11534,N_9992,N_9784);
nand U11535 (N_11535,N_9289,N_8980);
nor U11536 (N_11536,N_8255,N_9937);
nand U11537 (N_11537,N_9335,N_9978);
nand U11538 (N_11538,N_8392,N_8838);
nand U11539 (N_11539,N_9717,N_8658);
nand U11540 (N_11540,N_9764,N_8676);
or U11541 (N_11541,N_9905,N_9417);
nor U11542 (N_11542,N_8236,N_8048);
nand U11543 (N_11543,N_8294,N_9754);
and U11544 (N_11544,N_8335,N_9748);
nand U11545 (N_11545,N_8058,N_8755);
or U11546 (N_11546,N_9048,N_9675);
nand U11547 (N_11547,N_8993,N_8760);
nand U11548 (N_11548,N_8567,N_8956);
nor U11549 (N_11549,N_9282,N_8299);
nand U11550 (N_11550,N_9275,N_9253);
nand U11551 (N_11551,N_8072,N_9418);
and U11552 (N_11552,N_8454,N_9938);
or U11553 (N_11553,N_8228,N_8167);
nand U11554 (N_11554,N_9845,N_8671);
or U11555 (N_11555,N_9321,N_8657);
xor U11556 (N_11556,N_9950,N_8875);
or U11557 (N_11557,N_9152,N_9285);
nor U11558 (N_11558,N_9569,N_8311);
nor U11559 (N_11559,N_8707,N_8317);
and U11560 (N_11560,N_9430,N_8038);
and U11561 (N_11561,N_8301,N_9347);
xnor U11562 (N_11562,N_8324,N_8796);
or U11563 (N_11563,N_9378,N_9899);
or U11564 (N_11564,N_9932,N_8018);
nand U11565 (N_11565,N_9365,N_8974);
and U11566 (N_11566,N_9450,N_9207);
or U11567 (N_11567,N_9193,N_8889);
nand U11568 (N_11568,N_9049,N_8729);
nor U11569 (N_11569,N_8917,N_9629);
xor U11570 (N_11570,N_9177,N_9811);
nor U11571 (N_11571,N_8807,N_8431);
or U11572 (N_11572,N_9138,N_8096);
and U11573 (N_11573,N_8367,N_9086);
nor U11574 (N_11574,N_8591,N_9147);
nor U11575 (N_11575,N_9166,N_9377);
xnor U11576 (N_11576,N_9275,N_9583);
or U11577 (N_11577,N_8929,N_9387);
or U11578 (N_11578,N_9794,N_9971);
nor U11579 (N_11579,N_9100,N_8366);
xnor U11580 (N_11580,N_8237,N_9125);
or U11581 (N_11581,N_8725,N_9360);
xnor U11582 (N_11582,N_8523,N_8473);
nor U11583 (N_11583,N_8735,N_9826);
or U11584 (N_11584,N_9236,N_9373);
and U11585 (N_11585,N_9680,N_8702);
xnor U11586 (N_11586,N_9366,N_9449);
and U11587 (N_11587,N_8605,N_9759);
nand U11588 (N_11588,N_8295,N_8895);
nor U11589 (N_11589,N_8701,N_9306);
or U11590 (N_11590,N_8114,N_9712);
nor U11591 (N_11591,N_9173,N_9877);
and U11592 (N_11592,N_8501,N_9124);
nand U11593 (N_11593,N_9908,N_8918);
and U11594 (N_11594,N_8530,N_9312);
xor U11595 (N_11595,N_9524,N_9515);
or U11596 (N_11596,N_8395,N_8967);
or U11597 (N_11597,N_9466,N_8422);
nand U11598 (N_11598,N_8735,N_9298);
and U11599 (N_11599,N_8205,N_8073);
or U11600 (N_11600,N_9351,N_9935);
nor U11601 (N_11601,N_9704,N_8899);
nor U11602 (N_11602,N_8376,N_8523);
or U11603 (N_11603,N_9870,N_9232);
or U11604 (N_11604,N_9096,N_8527);
or U11605 (N_11605,N_9517,N_8552);
nand U11606 (N_11606,N_8393,N_8042);
nand U11607 (N_11607,N_8475,N_8968);
nand U11608 (N_11608,N_8923,N_8253);
nor U11609 (N_11609,N_8454,N_9514);
nand U11610 (N_11610,N_9766,N_8527);
and U11611 (N_11611,N_8159,N_9146);
nand U11612 (N_11612,N_8843,N_8621);
and U11613 (N_11613,N_9746,N_8974);
or U11614 (N_11614,N_9636,N_8944);
nand U11615 (N_11615,N_8702,N_9388);
nand U11616 (N_11616,N_8303,N_9238);
nor U11617 (N_11617,N_9025,N_8417);
nand U11618 (N_11618,N_8329,N_8052);
nand U11619 (N_11619,N_8788,N_8583);
nand U11620 (N_11620,N_8523,N_9309);
or U11621 (N_11621,N_9153,N_8921);
nor U11622 (N_11622,N_9258,N_8921);
and U11623 (N_11623,N_8870,N_9655);
nand U11624 (N_11624,N_8868,N_8692);
nand U11625 (N_11625,N_8374,N_8114);
and U11626 (N_11626,N_9783,N_8405);
nand U11627 (N_11627,N_8680,N_8852);
or U11628 (N_11628,N_8681,N_9305);
and U11629 (N_11629,N_9739,N_8651);
nand U11630 (N_11630,N_8070,N_8214);
or U11631 (N_11631,N_9364,N_8827);
and U11632 (N_11632,N_8512,N_8936);
nor U11633 (N_11633,N_9550,N_8309);
nor U11634 (N_11634,N_8692,N_8344);
and U11635 (N_11635,N_8774,N_9249);
nand U11636 (N_11636,N_8893,N_9307);
or U11637 (N_11637,N_8623,N_9313);
and U11638 (N_11638,N_9168,N_9770);
xor U11639 (N_11639,N_9585,N_8216);
nand U11640 (N_11640,N_8095,N_8425);
nor U11641 (N_11641,N_8878,N_9383);
nor U11642 (N_11642,N_8364,N_9614);
xnor U11643 (N_11643,N_9123,N_8140);
nor U11644 (N_11644,N_8495,N_8270);
nor U11645 (N_11645,N_8242,N_9536);
and U11646 (N_11646,N_8719,N_8805);
and U11647 (N_11647,N_9133,N_8403);
nand U11648 (N_11648,N_8112,N_8563);
or U11649 (N_11649,N_9959,N_8741);
xor U11650 (N_11650,N_8870,N_8928);
nand U11651 (N_11651,N_8861,N_9624);
nor U11652 (N_11652,N_9853,N_9348);
nand U11653 (N_11653,N_9906,N_8199);
xnor U11654 (N_11654,N_8680,N_8079);
and U11655 (N_11655,N_8038,N_8146);
or U11656 (N_11656,N_9447,N_9493);
nand U11657 (N_11657,N_9355,N_9321);
nor U11658 (N_11658,N_9304,N_8391);
xor U11659 (N_11659,N_9724,N_9140);
or U11660 (N_11660,N_8684,N_8087);
or U11661 (N_11661,N_8562,N_8641);
nand U11662 (N_11662,N_8410,N_9857);
nand U11663 (N_11663,N_8181,N_9148);
xor U11664 (N_11664,N_9544,N_9318);
nor U11665 (N_11665,N_9633,N_8881);
or U11666 (N_11666,N_8490,N_9387);
nand U11667 (N_11667,N_8452,N_9537);
or U11668 (N_11668,N_8382,N_9035);
and U11669 (N_11669,N_9732,N_8944);
and U11670 (N_11670,N_8245,N_9709);
and U11671 (N_11671,N_8154,N_8086);
or U11672 (N_11672,N_9016,N_9318);
and U11673 (N_11673,N_9011,N_8408);
nor U11674 (N_11674,N_8526,N_9896);
nand U11675 (N_11675,N_9123,N_9792);
and U11676 (N_11676,N_8850,N_9494);
nor U11677 (N_11677,N_9809,N_9016);
or U11678 (N_11678,N_9696,N_8711);
and U11679 (N_11679,N_8307,N_9868);
xor U11680 (N_11680,N_9885,N_9014);
nand U11681 (N_11681,N_9287,N_8459);
or U11682 (N_11682,N_8211,N_9157);
or U11683 (N_11683,N_8394,N_8951);
nand U11684 (N_11684,N_8758,N_8267);
or U11685 (N_11685,N_9373,N_9250);
nand U11686 (N_11686,N_9943,N_9972);
nor U11687 (N_11687,N_8738,N_8162);
or U11688 (N_11688,N_9298,N_8088);
and U11689 (N_11689,N_9213,N_9431);
xnor U11690 (N_11690,N_9363,N_8934);
or U11691 (N_11691,N_9540,N_8329);
nor U11692 (N_11692,N_8845,N_8850);
nand U11693 (N_11693,N_8190,N_8433);
and U11694 (N_11694,N_8129,N_8070);
and U11695 (N_11695,N_9219,N_9068);
nand U11696 (N_11696,N_9891,N_8975);
xor U11697 (N_11697,N_9636,N_9659);
or U11698 (N_11698,N_8078,N_9198);
nand U11699 (N_11699,N_8344,N_8637);
nor U11700 (N_11700,N_9918,N_9277);
and U11701 (N_11701,N_8949,N_8382);
nand U11702 (N_11702,N_9983,N_8558);
or U11703 (N_11703,N_8339,N_9178);
and U11704 (N_11704,N_8160,N_8803);
nand U11705 (N_11705,N_8348,N_8493);
xnor U11706 (N_11706,N_9313,N_8774);
and U11707 (N_11707,N_8635,N_9831);
and U11708 (N_11708,N_9518,N_8099);
nor U11709 (N_11709,N_9275,N_8773);
and U11710 (N_11710,N_8748,N_8047);
nor U11711 (N_11711,N_9532,N_9143);
or U11712 (N_11712,N_9314,N_9341);
or U11713 (N_11713,N_9433,N_9954);
xor U11714 (N_11714,N_9770,N_9265);
and U11715 (N_11715,N_9174,N_8909);
and U11716 (N_11716,N_9122,N_8517);
and U11717 (N_11717,N_8875,N_8834);
or U11718 (N_11718,N_8664,N_8972);
xor U11719 (N_11719,N_8527,N_8163);
or U11720 (N_11720,N_9560,N_9337);
xnor U11721 (N_11721,N_8869,N_8671);
or U11722 (N_11722,N_8224,N_9275);
nand U11723 (N_11723,N_8652,N_8637);
or U11724 (N_11724,N_9096,N_9700);
and U11725 (N_11725,N_9320,N_8275);
nor U11726 (N_11726,N_9576,N_9582);
nand U11727 (N_11727,N_9872,N_8187);
or U11728 (N_11728,N_9973,N_9594);
nand U11729 (N_11729,N_8034,N_8151);
and U11730 (N_11730,N_9553,N_8875);
xnor U11731 (N_11731,N_9537,N_8853);
or U11732 (N_11732,N_8405,N_8784);
or U11733 (N_11733,N_8180,N_9614);
nand U11734 (N_11734,N_9304,N_9989);
and U11735 (N_11735,N_8304,N_8044);
nor U11736 (N_11736,N_9749,N_9009);
nor U11737 (N_11737,N_9991,N_8468);
and U11738 (N_11738,N_8277,N_9850);
and U11739 (N_11739,N_9684,N_8559);
and U11740 (N_11740,N_9078,N_9020);
and U11741 (N_11741,N_9382,N_8019);
nor U11742 (N_11742,N_8905,N_9240);
or U11743 (N_11743,N_8558,N_8370);
or U11744 (N_11744,N_9109,N_8625);
and U11745 (N_11745,N_9298,N_9200);
or U11746 (N_11746,N_8939,N_8004);
nand U11747 (N_11747,N_9682,N_8926);
or U11748 (N_11748,N_8604,N_8635);
nand U11749 (N_11749,N_8036,N_9386);
or U11750 (N_11750,N_8876,N_8555);
and U11751 (N_11751,N_8561,N_8402);
and U11752 (N_11752,N_8994,N_8549);
and U11753 (N_11753,N_8539,N_8800);
nand U11754 (N_11754,N_9631,N_9127);
and U11755 (N_11755,N_8721,N_8467);
or U11756 (N_11756,N_9060,N_8603);
nor U11757 (N_11757,N_9980,N_9304);
nand U11758 (N_11758,N_9366,N_8443);
nor U11759 (N_11759,N_9902,N_9668);
or U11760 (N_11760,N_8184,N_8692);
xor U11761 (N_11761,N_8001,N_9407);
nor U11762 (N_11762,N_8730,N_9995);
or U11763 (N_11763,N_9249,N_8161);
or U11764 (N_11764,N_9053,N_9031);
xnor U11765 (N_11765,N_9057,N_9479);
nand U11766 (N_11766,N_8833,N_9866);
nand U11767 (N_11767,N_9450,N_9819);
nor U11768 (N_11768,N_9463,N_8762);
nor U11769 (N_11769,N_8643,N_8213);
or U11770 (N_11770,N_8222,N_9576);
or U11771 (N_11771,N_9671,N_8633);
xor U11772 (N_11772,N_9194,N_9919);
nand U11773 (N_11773,N_8696,N_9749);
xor U11774 (N_11774,N_9346,N_9053);
nand U11775 (N_11775,N_9356,N_8464);
nor U11776 (N_11776,N_8875,N_8214);
xor U11777 (N_11777,N_8298,N_9583);
nand U11778 (N_11778,N_9416,N_8880);
or U11779 (N_11779,N_9143,N_8300);
or U11780 (N_11780,N_8348,N_9642);
or U11781 (N_11781,N_9096,N_8879);
xnor U11782 (N_11782,N_8120,N_8054);
xor U11783 (N_11783,N_8373,N_8792);
or U11784 (N_11784,N_8206,N_8545);
nor U11785 (N_11785,N_9865,N_9228);
or U11786 (N_11786,N_9138,N_8108);
nor U11787 (N_11787,N_9722,N_8865);
nor U11788 (N_11788,N_8399,N_9358);
nand U11789 (N_11789,N_9119,N_8070);
and U11790 (N_11790,N_9344,N_9679);
and U11791 (N_11791,N_8930,N_9531);
nor U11792 (N_11792,N_9863,N_9548);
or U11793 (N_11793,N_9842,N_8899);
and U11794 (N_11794,N_8284,N_8927);
nand U11795 (N_11795,N_9407,N_8957);
xor U11796 (N_11796,N_9387,N_8134);
and U11797 (N_11797,N_9628,N_9967);
nor U11798 (N_11798,N_8534,N_8376);
or U11799 (N_11799,N_8996,N_9631);
and U11800 (N_11800,N_9202,N_8609);
nor U11801 (N_11801,N_9693,N_9044);
nand U11802 (N_11802,N_8931,N_8868);
nor U11803 (N_11803,N_8576,N_9083);
nand U11804 (N_11804,N_9744,N_9791);
or U11805 (N_11805,N_9101,N_8990);
or U11806 (N_11806,N_9614,N_9577);
xor U11807 (N_11807,N_9882,N_8873);
nor U11808 (N_11808,N_8807,N_8706);
nor U11809 (N_11809,N_9531,N_8606);
and U11810 (N_11810,N_8095,N_8342);
nor U11811 (N_11811,N_9127,N_8829);
xnor U11812 (N_11812,N_9318,N_8478);
nor U11813 (N_11813,N_8794,N_8780);
or U11814 (N_11814,N_8536,N_8692);
or U11815 (N_11815,N_8218,N_8121);
or U11816 (N_11816,N_9109,N_8149);
and U11817 (N_11817,N_9238,N_8283);
nor U11818 (N_11818,N_8457,N_8402);
nand U11819 (N_11819,N_9840,N_9314);
nand U11820 (N_11820,N_9528,N_9534);
and U11821 (N_11821,N_8727,N_9053);
nor U11822 (N_11822,N_9293,N_9713);
or U11823 (N_11823,N_8026,N_9971);
nand U11824 (N_11824,N_8722,N_8382);
and U11825 (N_11825,N_8049,N_8104);
and U11826 (N_11826,N_9772,N_9574);
or U11827 (N_11827,N_8287,N_9149);
nand U11828 (N_11828,N_9433,N_9155);
nor U11829 (N_11829,N_9065,N_9932);
and U11830 (N_11830,N_9854,N_9621);
nor U11831 (N_11831,N_8087,N_9084);
nand U11832 (N_11832,N_9485,N_8654);
and U11833 (N_11833,N_8018,N_8327);
nor U11834 (N_11834,N_8570,N_9403);
nand U11835 (N_11835,N_8392,N_9011);
or U11836 (N_11836,N_8642,N_8597);
nand U11837 (N_11837,N_8893,N_9366);
and U11838 (N_11838,N_8443,N_8393);
or U11839 (N_11839,N_8232,N_9577);
and U11840 (N_11840,N_8262,N_9358);
nor U11841 (N_11841,N_9045,N_8859);
and U11842 (N_11842,N_8601,N_9130);
and U11843 (N_11843,N_9003,N_9230);
xnor U11844 (N_11844,N_8878,N_8167);
and U11845 (N_11845,N_9755,N_8114);
nand U11846 (N_11846,N_8628,N_8728);
xor U11847 (N_11847,N_9276,N_8465);
or U11848 (N_11848,N_8489,N_9130);
nor U11849 (N_11849,N_9380,N_9924);
and U11850 (N_11850,N_8079,N_8420);
or U11851 (N_11851,N_9324,N_9098);
nor U11852 (N_11852,N_9126,N_9314);
or U11853 (N_11853,N_9540,N_8041);
nand U11854 (N_11854,N_9256,N_8140);
xnor U11855 (N_11855,N_9119,N_9686);
nand U11856 (N_11856,N_9671,N_9281);
nor U11857 (N_11857,N_9961,N_9980);
nand U11858 (N_11858,N_9156,N_9517);
nand U11859 (N_11859,N_8558,N_9636);
nor U11860 (N_11860,N_8630,N_9091);
nor U11861 (N_11861,N_8025,N_9359);
or U11862 (N_11862,N_8927,N_9842);
nor U11863 (N_11863,N_8657,N_9524);
nand U11864 (N_11864,N_8890,N_8004);
xor U11865 (N_11865,N_8265,N_8952);
and U11866 (N_11866,N_8531,N_9329);
nor U11867 (N_11867,N_8946,N_9592);
nand U11868 (N_11868,N_9103,N_9495);
nor U11869 (N_11869,N_9144,N_9210);
or U11870 (N_11870,N_9977,N_9898);
or U11871 (N_11871,N_8804,N_9755);
nor U11872 (N_11872,N_8660,N_9194);
nor U11873 (N_11873,N_8253,N_9274);
xor U11874 (N_11874,N_8261,N_8200);
and U11875 (N_11875,N_9533,N_9823);
nor U11876 (N_11876,N_8453,N_8202);
nor U11877 (N_11877,N_8695,N_8051);
and U11878 (N_11878,N_9928,N_9652);
nor U11879 (N_11879,N_8241,N_9226);
nand U11880 (N_11880,N_9818,N_8232);
nand U11881 (N_11881,N_9530,N_8021);
and U11882 (N_11882,N_8510,N_8333);
or U11883 (N_11883,N_9313,N_8607);
nand U11884 (N_11884,N_9742,N_8410);
nor U11885 (N_11885,N_8218,N_8528);
xnor U11886 (N_11886,N_9864,N_9105);
nor U11887 (N_11887,N_8020,N_9483);
or U11888 (N_11888,N_8780,N_8316);
and U11889 (N_11889,N_8891,N_9383);
nor U11890 (N_11890,N_9272,N_9337);
xor U11891 (N_11891,N_9374,N_8245);
nor U11892 (N_11892,N_9798,N_8817);
nor U11893 (N_11893,N_8500,N_8830);
nand U11894 (N_11894,N_8470,N_9255);
or U11895 (N_11895,N_8060,N_9661);
nor U11896 (N_11896,N_9759,N_8981);
and U11897 (N_11897,N_8603,N_9205);
nand U11898 (N_11898,N_8575,N_9138);
nor U11899 (N_11899,N_9300,N_8162);
xor U11900 (N_11900,N_9668,N_8374);
or U11901 (N_11901,N_8871,N_9716);
and U11902 (N_11902,N_9360,N_9381);
nor U11903 (N_11903,N_8997,N_9804);
or U11904 (N_11904,N_9269,N_8421);
and U11905 (N_11905,N_8557,N_9604);
nor U11906 (N_11906,N_9011,N_8965);
nor U11907 (N_11907,N_9662,N_8220);
and U11908 (N_11908,N_8590,N_8193);
or U11909 (N_11909,N_9350,N_8593);
and U11910 (N_11910,N_8694,N_8036);
nor U11911 (N_11911,N_9666,N_9110);
nand U11912 (N_11912,N_9488,N_8071);
xor U11913 (N_11913,N_9922,N_8505);
xnor U11914 (N_11914,N_8829,N_8831);
or U11915 (N_11915,N_8256,N_8407);
or U11916 (N_11916,N_9876,N_8919);
nor U11917 (N_11917,N_9149,N_8614);
nand U11918 (N_11918,N_8344,N_8295);
and U11919 (N_11919,N_9316,N_8129);
nand U11920 (N_11920,N_9182,N_9271);
xnor U11921 (N_11921,N_9262,N_9214);
nand U11922 (N_11922,N_8338,N_8020);
or U11923 (N_11923,N_9948,N_8952);
nor U11924 (N_11924,N_9151,N_9084);
nor U11925 (N_11925,N_8366,N_8305);
nand U11926 (N_11926,N_8412,N_8773);
nand U11927 (N_11927,N_9395,N_9269);
nor U11928 (N_11928,N_9604,N_9423);
or U11929 (N_11929,N_9781,N_9851);
or U11930 (N_11930,N_9410,N_8497);
nand U11931 (N_11931,N_8986,N_8552);
and U11932 (N_11932,N_9409,N_9404);
xor U11933 (N_11933,N_9087,N_9722);
and U11934 (N_11934,N_9331,N_9292);
nor U11935 (N_11935,N_9143,N_8020);
and U11936 (N_11936,N_9859,N_9960);
nand U11937 (N_11937,N_8640,N_9612);
xor U11938 (N_11938,N_8236,N_8259);
xor U11939 (N_11939,N_9551,N_8972);
and U11940 (N_11940,N_8570,N_8892);
and U11941 (N_11941,N_8975,N_8395);
nand U11942 (N_11942,N_9046,N_8868);
nand U11943 (N_11943,N_9116,N_9471);
nand U11944 (N_11944,N_9774,N_8026);
xnor U11945 (N_11945,N_9415,N_8180);
and U11946 (N_11946,N_8141,N_9309);
nand U11947 (N_11947,N_8506,N_9945);
nand U11948 (N_11948,N_8513,N_8522);
and U11949 (N_11949,N_9586,N_8675);
nand U11950 (N_11950,N_9528,N_8195);
and U11951 (N_11951,N_9719,N_8585);
xnor U11952 (N_11952,N_8006,N_8046);
or U11953 (N_11953,N_9946,N_8235);
or U11954 (N_11954,N_8924,N_9407);
or U11955 (N_11955,N_9053,N_8608);
and U11956 (N_11956,N_8535,N_8376);
nand U11957 (N_11957,N_9078,N_8821);
and U11958 (N_11958,N_8775,N_9792);
nand U11959 (N_11959,N_9809,N_9000);
nand U11960 (N_11960,N_9554,N_9359);
nor U11961 (N_11961,N_8300,N_9059);
and U11962 (N_11962,N_9581,N_8005);
or U11963 (N_11963,N_9423,N_8542);
or U11964 (N_11964,N_8088,N_8148);
and U11965 (N_11965,N_8513,N_9095);
and U11966 (N_11966,N_8288,N_8981);
xnor U11967 (N_11967,N_8071,N_9232);
xor U11968 (N_11968,N_8853,N_9509);
nand U11969 (N_11969,N_9077,N_8124);
or U11970 (N_11970,N_9012,N_8400);
and U11971 (N_11971,N_8268,N_9298);
nand U11972 (N_11972,N_9965,N_9146);
or U11973 (N_11973,N_8389,N_9049);
and U11974 (N_11974,N_9554,N_9597);
nor U11975 (N_11975,N_9630,N_8231);
nand U11976 (N_11976,N_8514,N_9475);
xnor U11977 (N_11977,N_8890,N_8907);
nand U11978 (N_11978,N_9138,N_8467);
nor U11979 (N_11979,N_8036,N_9738);
nor U11980 (N_11980,N_9581,N_8536);
nor U11981 (N_11981,N_8568,N_9347);
or U11982 (N_11982,N_8699,N_9762);
nand U11983 (N_11983,N_8701,N_8863);
nand U11984 (N_11984,N_9909,N_9393);
nand U11985 (N_11985,N_9588,N_9488);
xor U11986 (N_11986,N_9873,N_8433);
nor U11987 (N_11987,N_8500,N_8898);
and U11988 (N_11988,N_8840,N_9399);
and U11989 (N_11989,N_9188,N_8577);
nor U11990 (N_11990,N_9190,N_9870);
or U11991 (N_11991,N_8000,N_9605);
nor U11992 (N_11992,N_8321,N_8171);
nor U11993 (N_11993,N_9852,N_8604);
and U11994 (N_11994,N_9562,N_9374);
nand U11995 (N_11995,N_8947,N_9406);
nand U11996 (N_11996,N_8432,N_9118);
nand U11997 (N_11997,N_8356,N_8939);
and U11998 (N_11998,N_8770,N_9903);
nor U11999 (N_11999,N_9186,N_8738);
nand U12000 (N_12000,N_11635,N_11332);
or U12001 (N_12001,N_11414,N_11543);
or U12002 (N_12002,N_10301,N_10058);
and U12003 (N_12003,N_11567,N_10647);
and U12004 (N_12004,N_11004,N_10595);
nand U12005 (N_12005,N_11303,N_11812);
or U12006 (N_12006,N_10959,N_11961);
and U12007 (N_12007,N_11940,N_11459);
xnor U12008 (N_12008,N_10599,N_10442);
nor U12009 (N_12009,N_10687,N_11150);
nand U12010 (N_12010,N_10001,N_10960);
and U12011 (N_12011,N_11458,N_10129);
nor U12012 (N_12012,N_11252,N_11148);
nor U12013 (N_12013,N_10234,N_10265);
nor U12014 (N_12014,N_11813,N_11796);
or U12015 (N_12015,N_11662,N_11279);
nand U12016 (N_12016,N_11088,N_10643);
nand U12017 (N_12017,N_11649,N_10889);
nand U12018 (N_12018,N_11080,N_11198);
or U12019 (N_12019,N_10856,N_10166);
xnor U12020 (N_12020,N_10774,N_10768);
and U12021 (N_12021,N_10310,N_11733);
nand U12022 (N_12022,N_10814,N_11029);
nand U12023 (N_12023,N_10440,N_10082);
nand U12024 (N_12024,N_11299,N_10458);
and U12025 (N_12025,N_11062,N_11228);
nand U12026 (N_12026,N_10655,N_11162);
or U12027 (N_12027,N_11885,N_10360);
or U12028 (N_12028,N_10588,N_11192);
and U12029 (N_12029,N_10878,N_11443);
or U12030 (N_12030,N_10165,N_11850);
nor U12031 (N_12031,N_11405,N_10463);
and U12032 (N_12032,N_10982,N_10771);
or U12033 (N_12033,N_11871,N_11486);
nand U12034 (N_12034,N_11310,N_11103);
nand U12035 (N_12035,N_10282,N_10696);
nand U12036 (N_12036,N_11160,N_11351);
nor U12037 (N_12037,N_11355,N_11383);
and U12038 (N_12038,N_11102,N_10339);
or U12039 (N_12039,N_11138,N_10587);
nand U12040 (N_12040,N_11311,N_10292);
and U12041 (N_12041,N_11046,N_10886);
nor U12042 (N_12042,N_10117,N_11845);
or U12043 (N_12043,N_11322,N_10908);
xnor U12044 (N_12044,N_11260,N_10324);
nand U12045 (N_12045,N_11586,N_11691);
nand U12046 (N_12046,N_11523,N_10349);
nor U12047 (N_12047,N_11875,N_11125);
and U12048 (N_12048,N_10710,N_11978);
nand U12049 (N_12049,N_11516,N_10744);
nand U12050 (N_12050,N_11061,N_11240);
and U12051 (N_12051,N_11638,N_11435);
and U12052 (N_12052,N_11952,N_10183);
nor U12053 (N_12053,N_10152,N_10773);
nor U12054 (N_12054,N_10704,N_10722);
or U12055 (N_12055,N_10944,N_10898);
and U12056 (N_12056,N_10873,N_11873);
and U12057 (N_12057,N_10356,N_11413);
nand U12058 (N_12058,N_11899,N_10943);
nor U12059 (N_12059,N_10323,N_11792);
or U12060 (N_12060,N_11320,N_11382);
and U12061 (N_12061,N_11597,N_10306);
nand U12062 (N_12062,N_11384,N_11715);
nand U12063 (N_12063,N_10991,N_10961);
and U12064 (N_12064,N_10009,N_10930);
nand U12065 (N_12065,N_11257,N_11087);
and U12066 (N_12066,N_11831,N_10688);
or U12067 (N_12067,N_11718,N_10615);
or U12068 (N_12068,N_11177,N_10691);
nor U12069 (N_12069,N_11713,N_10321);
or U12070 (N_12070,N_11506,N_10302);
and U12071 (N_12071,N_11137,N_10093);
and U12072 (N_12072,N_11761,N_11654);
and U12073 (N_12073,N_11579,N_10596);
and U12074 (N_12074,N_10716,N_11447);
or U12075 (N_12075,N_10462,N_11729);
nand U12076 (N_12076,N_11937,N_10000);
and U12077 (N_12077,N_11637,N_11653);
or U12078 (N_12078,N_11736,N_11000);
or U12079 (N_12079,N_10749,N_10346);
and U12080 (N_12080,N_11782,N_10160);
or U12081 (N_12081,N_11737,N_10954);
nor U12082 (N_12082,N_10392,N_10550);
and U12083 (N_12083,N_10019,N_11318);
nor U12084 (N_12084,N_11633,N_11731);
nand U12085 (N_12085,N_10181,N_11787);
and U12086 (N_12086,N_10482,N_11795);
and U12087 (N_12087,N_10988,N_11902);
nand U12088 (N_12088,N_11949,N_10167);
nand U12089 (N_12089,N_11955,N_11356);
and U12090 (N_12090,N_11181,N_11780);
or U12091 (N_12091,N_10351,N_10464);
or U12092 (N_12092,N_10205,N_11412);
or U12093 (N_12093,N_10876,N_10924);
xnor U12094 (N_12094,N_10371,N_10103);
nand U12095 (N_12095,N_10445,N_10934);
xnor U12096 (N_12096,N_10592,N_11193);
and U12097 (N_12097,N_10147,N_10638);
nand U12098 (N_12098,N_11645,N_11839);
nand U12099 (N_12099,N_11109,N_11953);
nand U12100 (N_12100,N_11107,N_10359);
nor U12101 (N_12101,N_11624,N_11998);
or U12102 (N_12102,N_11706,N_10729);
nand U12103 (N_12103,N_11188,N_11604);
or U12104 (N_12104,N_11034,N_10362);
nand U12105 (N_12105,N_11403,N_10622);
nand U12106 (N_12106,N_10724,N_10702);
nand U12107 (N_12107,N_10753,N_11212);
nor U12108 (N_12108,N_10497,N_10833);
or U12109 (N_12109,N_11379,N_10134);
xnor U12110 (N_12110,N_11788,N_11755);
xor U12111 (N_12111,N_11520,N_11956);
nand U12112 (N_12112,N_10335,N_10607);
or U12113 (N_12113,N_10380,N_10646);
or U12114 (N_12114,N_10740,N_11686);
or U12115 (N_12115,N_11475,N_10893);
xor U12116 (N_12116,N_11225,N_11124);
or U12117 (N_12117,N_10941,N_10437);
and U12118 (N_12118,N_11540,N_10678);
nand U12119 (N_12119,N_11933,N_10970);
nand U12120 (N_12120,N_11941,N_10350);
or U12121 (N_12121,N_11560,N_10764);
nand U12122 (N_12122,N_11600,N_11099);
nand U12123 (N_12123,N_10614,N_11595);
or U12124 (N_12124,N_10085,N_10798);
xnor U12125 (N_12125,N_11400,N_11993);
or U12126 (N_12126,N_11183,N_10769);
or U12127 (N_12127,N_10329,N_11176);
or U12128 (N_12128,N_10683,N_11853);
or U12129 (N_12129,N_10668,N_10423);
nor U12130 (N_12130,N_11263,N_10849);
xnor U12131 (N_12131,N_10322,N_10491);
nor U12132 (N_12132,N_11246,N_11019);
or U12133 (N_12133,N_11868,N_11292);
or U12134 (N_12134,N_10487,N_10541);
xnor U12135 (N_12135,N_11497,N_10062);
nor U12136 (N_12136,N_10429,N_10582);
nor U12137 (N_12137,N_11305,N_10973);
nor U12138 (N_12138,N_10826,N_10176);
nor U12139 (N_12139,N_10490,N_10718);
nand U12140 (N_12140,N_11465,N_10011);
nand U12141 (N_12141,N_10372,N_11507);
nand U12142 (N_12142,N_11696,N_11574);
xor U12143 (N_12143,N_10572,N_11483);
nand U12144 (N_12144,N_10695,N_11077);
and U12145 (N_12145,N_10274,N_10252);
and U12146 (N_12146,N_11849,N_11455);
or U12147 (N_12147,N_10531,N_10231);
or U12148 (N_12148,N_11499,N_11295);
or U12149 (N_12149,N_11298,N_11337);
nand U12150 (N_12150,N_10444,N_11023);
xor U12151 (N_12151,N_10186,N_11513);
nor U12152 (N_12152,N_11865,N_11419);
or U12153 (N_12153,N_10338,N_10028);
xor U12154 (N_12154,N_11463,N_11683);
nor U12155 (N_12155,N_11282,N_10828);
xor U12156 (N_12156,N_11829,N_10778);
or U12157 (N_12157,N_11655,N_10340);
xor U12158 (N_12158,N_11496,N_11220);
nor U12159 (N_12159,N_10585,N_10032);
nor U12160 (N_12160,N_10225,N_10963);
or U12161 (N_12161,N_11530,N_10745);
xor U12162 (N_12162,N_11362,N_11682);
nand U12163 (N_12163,N_11128,N_11766);
and U12164 (N_12164,N_11428,N_11048);
and U12165 (N_12165,N_10672,N_10211);
nand U12166 (N_12166,N_11927,N_11963);
and U12167 (N_12167,N_10577,N_10249);
and U12168 (N_12168,N_10698,N_10259);
nand U12169 (N_12169,N_11376,N_10616);
nand U12170 (N_12170,N_11461,N_10027);
xnor U12171 (N_12171,N_10971,N_10962);
and U12172 (N_12172,N_11477,N_10258);
and U12173 (N_12173,N_11620,N_11083);
nor U12174 (N_12174,N_11009,N_10715);
nand U12175 (N_12175,N_11036,N_10883);
or U12176 (N_12176,N_10575,N_11489);
xnor U12177 (N_12177,N_10840,N_11559);
nor U12178 (N_12178,N_10369,N_10850);
or U12179 (N_12179,N_10039,N_10297);
or U12180 (N_12180,N_11734,N_10169);
nand U12181 (N_12181,N_11521,N_11857);
and U12182 (N_12182,N_11281,N_11482);
nor U12183 (N_12183,N_10996,N_10594);
nor U12184 (N_12184,N_11484,N_10467);
nand U12185 (N_12185,N_10403,N_11485);
nand U12186 (N_12186,N_11585,N_11067);
xnor U12187 (N_12187,N_11283,N_10818);
or U12188 (N_12188,N_11056,N_11328);
or U12189 (N_12189,N_11154,N_10885);
or U12190 (N_12190,N_11182,N_10476);
and U12191 (N_12191,N_10692,N_10061);
nor U12192 (N_12192,N_11721,N_10547);
xnor U12193 (N_12193,N_10314,N_11702);
or U12194 (N_12194,N_11646,N_11794);
and U12195 (N_12195,N_10847,N_10975);
nor U12196 (N_12196,N_10786,N_11254);
nor U12197 (N_12197,N_10517,N_11970);
xnor U12198 (N_12198,N_11456,N_10382);
nand U12199 (N_12199,N_11074,N_11313);
nor U12200 (N_12200,N_10053,N_10125);
nor U12201 (N_12201,N_10221,N_10964);
nand U12202 (N_12202,N_11648,N_11016);
xnor U12203 (N_12203,N_11991,N_10071);
nor U12204 (N_12204,N_11110,N_11290);
and U12205 (N_12205,N_11338,N_10098);
nor U12206 (N_12206,N_11271,N_11209);
and U12207 (N_12207,N_10556,N_10526);
nand U12208 (N_12208,N_11757,N_11844);
or U12209 (N_12209,N_10378,N_10939);
or U12210 (N_12210,N_11820,N_10427);
nand U12211 (N_12211,N_10420,N_10373);
nand U12212 (N_12212,N_10277,N_11660);
nor U12213 (N_12213,N_10727,N_11418);
nand U12214 (N_12214,N_11752,N_11753);
or U12215 (N_12215,N_10570,N_10313);
and U12216 (N_12216,N_10393,N_10389);
or U12217 (N_12217,N_10925,N_10581);
nor U12218 (N_12218,N_10843,N_10483);
nor U12219 (N_12219,N_10999,N_10037);
nand U12220 (N_12220,N_10888,N_11877);
nand U12221 (N_12221,N_11641,N_10024);
nand U12222 (N_12222,N_11134,N_11402);
nand U12223 (N_12223,N_11404,N_10240);
nand U12224 (N_12224,N_10750,N_11642);
or U12225 (N_12225,N_11221,N_10366);
nand U12226 (N_12226,N_11444,N_10627);
nand U12227 (N_12227,N_10534,N_10938);
xor U12228 (N_12228,N_11663,N_10477);
or U12229 (N_12229,N_10025,N_10521);
nand U12230 (N_12230,N_10198,N_10290);
or U12231 (N_12231,N_11568,N_10838);
or U12232 (N_12232,N_10417,N_10560);
and U12233 (N_12233,N_11503,N_10611);
nand U12234 (N_12234,N_11407,N_10045);
and U12235 (N_12235,N_10918,N_11913);
nor U12236 (N_12236,N_10679,N_11315);
nand U12237 (N_12237,N_10185,N_10140);
or U12238 (N_12238,N_11719,N_10008);
xnor U12239 (N_12239,N_10800,N_10164);
nor U12240 (N_12240,N_11480,N_10034);
xnor U12241 (N_12241,N_10119,N_11621);
nand U12242 (N_12242,N_11126,N_11202);
xor U12243 (N_12243,N_11002,N_11255);
xor U12244 (N_12244,N_11408,N_10714);
or U12245 (N_12245,N_10603,N_10319);
xnor U12246 (N_12246,N_11769,N_11129);
and U12247 (N_12247,N_11081,N_10502);
and U12248 (N_12248,N_11098,N_10227);
nand U12249 (N_12249,N_11808,N_11416);
or U12250 (N_12250,N_11607,N_11467);
xnor U12251 (N_12251,N_11005,N_10620);
and U12252 (N_12252,N_10731,N_11608);
nand U12253 (N_12253,N_10904,N_10839);
or U12254 (N_12254,N_11058,N_11592);
or U12255 (N_12255,N_11665,N_11601);
and U12256 (N_12256,N_11415,N_10177);
nor U12257 (N_12257,N_10107,N_11306);
nand U12258 (N_12258,N_11533,N_11388);
nand U12259 (N_12259,N_10105,N_10866);
xnor U12260 (N_12260,N_11051,N_10633);
or U12261 (N_12261,N_10114,N_11743);
nand U12262 (N_12262,N_11816,N_11569);
xor U12263 (N_12263,N_11399,N_10080);
nor U12264 (N_12264,N_11393,N_11578);
nor U12265 (N_12265,N_11307,N_10789);
and U12266 (N_12266,N_10228,N_10469);
xor U12267 (N_12267,N_10161,N_10757);
nand U12268 (N_12268,N_11909,N_11916);
nor U12269 (N_12269,N_11040,N_10990);
or U12270 (N_12270,N_11884,N_10005);
and U12271 (N_12271,N_10783,N_11008);
nand U12272 (N_12272,N_11492,N_10253);
and U12273 (N_12273,N_10549,N_10909);
nand U12274 (N_12274,N_11449,N_11116);
xnor U12275 (N_12275,N_11013,N_11161);
nand U12276 (N_12276,N_11754,N_11422);
nor U12277 (N_12277,N_10222,N_11558);
nor U12278 (N_12278,N_11500,N_11363);
nand U12279 (N_12279,N_10414,N_10052);
or U12280 (N_12280,N_10293,N_11928);
nand U12281 (N_12281,N_10174,N_11823);
or U12282 (N_12282,N_11872,N_11587);
or U12283 (N_12283,N_11911,N_11050);
nor U12284 (N_12284,N_10554,N_11498);
or U12285 (N_12285,N_11717,N_11020);
and U12286 (N_12286,N_10387,N_11106);
and U12287 (N_12287,N_11840,N_11535);
and U12288 (N_12288,N_10072,N_10515);
xor U12289 (N_12289,N_11759,N_11078);
nor U12290 (N_12290,N_10184,N_11745);
or U12291 (N_12291,N_11417,N_10618);
nor U12292 (N_12292,N_11326,N_10056);
nand U12293 (N_12293,N_10398,N_11440);
nand U12294 (N_12294,N_11060,N_11992);
and U12295 (N_12295,N_11291,N_11350);
and U12296 (N_12296,N_11697,N_11681);
nand U12297 (N_12297,N_11554,N_10929);
or U12298 (N_12298,N_11312,N_11488);
or U12299 (N_12299,N_10984,N_11280);
and U12300 (N_12300,N_10004,N_10266);
nor U12301 (N_12301,N_10626,N_11028);
nor U12302 (N_12302,N_11610,N_11052);
nand U12303 (N_12303,N_11760,N_11802);
nor U12304 (N_12304,N_11541,N_11709);
nand U12305 (N_12305,N_11335,N_11617);
or U12306 (N_12306,N_10223,N_11187);
or U12307 (N_12307,N_10247,N_10969);
nand U12308 (N_12308,N_11975,N_11155);
nand U12309 (N_12309,N_10533,N_10065);
nor U12310 (N_12310,N_11195,N_10717);
xor U12311 (N_12311,N_11847,N_11158);
nor U12312 (N_12312,N_11385,N_11175);
or U12313 (N_12313,N_10712,N_11333);
or U12314 (N_12314,N_11324,N_11895);
or U12315 (N_12315,N_11256,N_11864);
nor U12316 (N_12316,N_10370,N_11748);
nor U12317 (N_12317,N_10583,N_10891);
and U12318 (N_12318,N_10995,N_11448);
and U12319 (N_12319,N_11344,N_11490);
nor U12320 (N_12320,N_11861,N_10263);
nand U12321 (N_12321,N_11190,N_11366);
nand U12322 (N_12322,N_11272,N_10586);
and U12323 (N_12323,N_10180,N_10645);
and U12324 (N_12324,N_10667,N_11830);
nor U12325 (N_12325,N_10513,N_11836);
nor U12326 (N_12326,N_10628,N_10431);
and U12327 (N_12327,N_11108,N_11210);
nor U12328 (N_12328,N_10481,N_10078);
or U12329 (N_12329,N_11528,N_11226);
xor U12330 (N_12330,N_10153,N_11776);
nand U12331 (N_12331,N_10419,N_10248);
nor U12332 (N_12332,N_10112,N_11241);
nand U12333 (N_12333,N_11264,N_10881);
or U12334 (N_12334,N_11122,N_10545);
or U12335 (N_12335,N_10751,N_11623);
and U12336 (N_12336,N_11781,N_11445);
nand U12337 (N_12337,N_11677,N_10279);
or U12338 (N_12338,N_11544,N_10077);
and U12339 (N_12339,N_11636,N_10780);
nand U12340 (N_12340,N_11906,N_11304);
nand U12341 (N_12341,N_11340,N_11097);
or U12342 (N_12342,N_10475,N_10430);
and U12343 (N_12343,N_11694,N_10830);
nand U12344 (N_12344,N_10998,N_11401);
nor U12345 (N_12345,N_11920,N_10374);
nand U12346 (N_12346,N_10311,N_10391);
nand U12347 (N_12347,N_10874,N_10242);
nor U12348 (N_12348,N_10709,N_11901);
or U12349 (N_12349,N_11708,N_11369);
or U12350 (N_12350,N_11468,N_10837);
nand U12351 (N_12351,N_11804,N_11247);
and U12352 (N_12352,N_10538,N_10073);
nand U12353 (N_12353,N_11505,N_11863);
or U12354 (N_12354,N_11710,N_10877);
xnor U12355 (N_12355,N_11855,N_10262);
nor U12356 (N_12356,N_11025,N_10662);
nand U12357 (N_12357,N_10660,N_10199);
xnor U12358 (N_12358,N_11777,N_11742);
and U12359 (N_12359,N_10489,N_11724);
nand U12360 (N_12360,N_10523,N_10665);
or U12361 (N_12361,N_11015,N_10608);
xor U12362 (N_12362,N_10926,N_10516);
or U12363 (N_12363,N_10746,N_10428);
and U12364 (N_12364,N_10997,N_10207);
nor U12365 (N_12365,N_11151,N_10871);
xor U12366 (N_12366,N_11049,N_11908);
nand U12367 (N_12367,N_10418,N_10224);
or U12368 (N_12368,N_11072,N_11185);
nand U12369 (N_12369,N_10743,N_10699);
nor U12370 (N_12370,N_11093,N_10612);
and U12371 (N_12371,N_11529,N_11590);
nand U12372 (N_12372,N_10162,N_11073);
nor U12373 (N_12373,N_11631,N_11512);
or U12374 (N_12374,N_10530,N_10742);
nand U12375 (N_12375,N_10289,N_11003);
nor U12376 (N_12376,N_10194,N_10215);
or U12377 (N_12377,N_10634,N_11818);
nand U12378 (N_12378,N_11197,N_11156);
nand U12379 (N_12379,N_10551,N_10286);
nor U12380 (N_12380,N_11047,N_11771);
nor U12381 (N_12381,N_10357,N_10284);
or U12382 (N_12382,N_11939,N_11935);
nand U12383 (N_12383,N_11573,N_11976);
nor U12384 (N_12384,N_11171,N_10685);
nand U12385 (N_12385,N_11999,N_11464);
nand U12386 (N_12386,N_10561,N_10193);
and U12387 (N_12387,N_11852,N_11958);
or U12388 (N_12388,N_11426,N_10233);
nor U12389 (N_12389,N_10546,N_11206);
or U12390 (N_12390,N_11789,N_11689);
nor U12391 (N_12391,N_11286,N_10609);
and U12392 (N_12392,N_11564,N_11972);
nand U12393 (N_12393,N_10684,N_10763);
nor U12394 (N_12394,N_10735,N_10096);
nor U12395 (N_12395,N_11945,N_11518);
nor U12396 (N_12396,N_10213,N_10844);
and U12397 (N_12397,N_11472,N_11325);
or U12398 (N_12398,N_10777,N_11778);
or U12399 (N_12399,N_11300,N_11673);
and U12400 (N_12400,N_11599,N_11994);
or U12401 (N_12401,N_11764,N_10950);
and U12402 (N_12402,N_11091,N_10197);
or U12403 (N_12403,N_11679,N_10086);
nand U12404 (N_12404,N_11826,N_10042);
or U12405 (N_12405,N_11259,N_11234);
xor U12406 (N_12406,N_10203,N_10807);
or U12407 (N_12407,N_11450,N_10725);
nor U12408 (N_12408,N_10132,N_10355);
xnor U12409 (N_12409,N_10070,N_10048);
nor U12410 (N_12410,N_10456,N_11065);
and U12411 (N_12411,N_11897,N_11526);
or U12412 (N_12412,N_10486,N_10157);
and U12413 (N_12413,N_10738,N_11647);
or U12414 (N_12414,N_10536,N_10793);
or U12415 (N_12415,N_10661,N_10424);
nor U12416 (N_12416,N_10432,N_10590);
nor U12417 (N_12417,N_10565,N_11168);
nor U12418 (N_12418,N_10148,N_11127);
or U12419 (N_12419,N_11085,N_11959);
nand U12420 (N_12420,N_10641,N_11285);
and U12421 (N_12421,N_11772,N_10122);
nand U12422 (N_12422,N_10495,N_10189);
or U12423 (N_12423,N_10190,N_11374);
and U12424 (N_12424,N_11997,N_11938);
nor U12425 (N_12425,N_10178,N_11071);
nand U12426 (N_12426,N_11879,N_10064);
nor U12427 (N_12427,N_10041,N_11314);
nor U12428 (N_12428,N_11105,N_11545);
nand U12429 (N_12429,N_11876,N_11453);
and U12430 (N_12430,N_11981,N_10260);
and U12431 (N_12431,N_10455,N_11261);
and U12432 (N_12432,N_10848,N_10368);
nor U12433 (N_12433,N_11044,N_10525);
nor U12434 (N_12434,N_10511,N_11725);
and U12435 (N_12435,N_11980,N_10133);
nor U12436 (N_12436,N_11606,N_11577);
or U12437 (N_12437,N_10472,N_11410);
nand U12438 (N_12438,N_10204,N_10361);
and U12439 (N_12439,N_11075,N_10580);
and U12440 (N_12440,N_11960,N_10170);
xor U12441 (N_12441,N_10448,N_10613);
nand U12442 (N_12442,N_11053,N_10674);
nand U12443 (N_12443,N_11924,N_10461);
or U12444 (N_12444,N_11200,N_11907);
or U12445 (N_12445,N_10083,N_10326);
or U12446 (N_12446,N_10473,N_10325);
or U12447 (N_12447,N_11208,N_10602);
nand U12448 (N_12448,N_11842,N_10425);
nand U12449 (N_12449,N_10723,N_10468);
xnor U12450 (N_12450,N_11973,N_11966);
and U12451 (N_12451,N_11353,N_11035);
or U12452 (N_12452,N_10300,N_10060);
nor U12453 (N_12453,N_11705,N_10294);
nor U12454 (N_12454,N_10690,N_10200);
and U12455 (N_12455,N_11249,N_10689);
and U12456 (N_12456,N_11224,N_11294);
xor U12457 (N_12457,N_10268,N_10415);
nor U12458 (N_12458,N_11532,N_11473);
and U12459 (N_12459,N_10334,N_10928);
nand U12460 (N_12460,N_10981,N_11843);
nor U12461 (N_12461,N_11141,N_10956);
nor U12462 (N_12462,N_11707,N_11786);
nand U12463 (N_12463,N_10673,N_10968);
or U12464 (N_12464,N_10238,N_10318);
nand U12465 (N_12465,N_10498,N_11323);
or U12466 (N_12466,N_10573,N_10841);
nor U12467 (N_12467,N_10488,N_11644);
xnor U12468 (N_12468,N_11701,N_10344);
and U12469 (N_12469,N_10509,N_10038);
and U12470 (N_12470,N_11793,N_11390);
nor U12471 (N_12471,N_11481,N_10452);
nand U12472 (N_12472,N_11238,N_11007);
nand U12473 (N_12473,N_10030,N_10254);
nand U12474 (N_12474,N_11667,N_10353);
nor U12475 (N_12475,N_10663,N_10752);
xor U12476 (N_12476,N_10721,N_10816);
and U12477 (N_12477,N_10985,N_11552);
nor U12478 (N_12478,N_11951,N_10701);
or U12479 (N_12479,N_11570,N_10316);
or U12480 (N_12480,N_11359,N_10868);
nor U12481 (N_12481,N_10192,N_10946);
or U12482 (N_12482,N_11178,N_10022);
and U12483 (N_12483,N_10955,N_11767);
and U12484 (N_12484,N_10821,N_11121);
nor U12485 (N_12485,N_10031,N_10273);
nand U12486 (N_12486,N_10074,N_11522);
nand U12487 (N_12487,N_10621,N_10097);
nor U12488 (N_12488,N_11368,N_10872);
nand U12489 (N_12489,N_11639,N_10739);
and U12490 (N_12490,N_10343,N_10682);
nor U12491 (N_12491,N_11203,N_11880);
nor U12492 (N_12492,N_10307,N_11735);
and U12493 (N_12493,N_11846,N_10214);
and U12494 (N_12494,N_10953,N_10906);
or U12495 (N_12495,N_10046,N_10851);
or U12496 (N_12496,N_11095,N_10212);
nand U12497 (N_12497,N_10896,N_11184);
nand U12498 (N_12498,N_10861,N_11117);
xor U12499 (N_12499,N_10173,N_10532);
nand U12500 (N_12500,N_11113,N_10466);
and U12501 (N_12501,N_11274,N_11656);
and U12502 (N_12502,N_11354,N_10345);
xnor U12503 (N_12503,N_11429,N_11824);
or U12504 (N_12504,N_10719,N_11803);
nor U12505 (N_12505,N_10501,N_11216);
and U12506 (N_12506,N_11634,N_10557);
nor U12507 (N_12507,N_10797,N_10457);
and U12508 (N_12508,N_10449,N_11012);
or U12509 (N_12509,N_11801,N_11278);
and U12510 (N_12510,N_11277,N_10182);
xnor U12511 (N_12511,N_10095,N_10923);
and U12512 (N_12512,N_11730,N_11273);
nor U12513 (N_12513,N_10365,N_11431);
nor U12514 (N_12514,N_10519,N_10348);
xor U12515 (N_12515,N_10412,N_11179);
nand U12516 (N_12516,N_11425,N_10755);
or U12517 (N_12517,N_11236,N_10974);
and U12518 (N_12518,N_10694,N_11205);
or U12519 (N_12519,N_11017,N_10298);
nand U12520 (N_12520,N_10075,N_10782);
and U12521 (N_12521,N_10591,N_11515);
nand U12522 (N_12522,N_11828,N_10044);
nor U12523 (N_12523,N_10766,N_10548);
or U12524 (N_12524,N_10823,N_10210);
nor U12525 (N_12525,N_11508,N_11131);
nand U12526 (N_12526,N_10255,N_10949);
or U12527 (N_12527,N_10528,N_11346);
or U12528 (N_12528,N_11301,N_10539);
nand U12529 (N_12529,N_11014,N_11947);
or U12530 (N_12530,N_10813,N_11140);
nand U12531 (N_12531,N_10865,N_11191);
nand U12532 (N_12532,N_11946,N_10651);
and U12533 (N_12533,N_10680,N_11149);
nand U12534 (N_12534,N_10900,N_11476);
nor U12535 (N_12535,N_11827,N_10853);
or U12536 (N_12536,N_11343,N_11043);
nor U12537 (N_12537,N_10822,N_10994);
and U12538 (N_12538,N_11438,N_11276);
or U12539 (N_12539,N_10804,N_11239);
and U12540 (N_12540,N_11917,N_11229);
nand U12541 (N_12541,N_10106,N_11309);
nand U12542 (N_12542,N_11874,N_10283);
nor U12543 (N_12543,N_10862,N_10859);
nand U12544 (N_12544,N_11632,N_11805);
nor U12545 (N_12545,N_11001,N_11094);
and U12546 (N_12546,N_11248,N_10894);
and U12547 (N_12547,N_11266,N_11575);
nand U12548 (N_12548,N_11762,N_11882);
nor U12549 (N_12549,N_10503,N_11517);
nand U12550 (N_12550,N_11809,N_11245);
nand U12551 (N_12551,N_11214,N_10337);
and U12552 (N_12552,N_11237,N_10013);
and U12553 (N_12553,N_11687,N_10905);
or U12554 (N_12554,N_11851,N_10506);
or U12555 (N_12555,N_10332,N_11547);
and U12556 (N_12556,N_11348,N_10016);
nor U12557 (N_12557,N_11217,N_10836);
nand U12558 (N_12558,N_11092,N_10902);
nor U12559 (N_12559,N_11658,N_11302);
xnor U12560 (N_12560,N_10809,N_11948);
or U12561 (N_12561,N_10705,N_11684);
nor U12562 (N_12562,N_10825,N_11974);
nor U12563 (N_12563,N_11627,N_11123);
and U12564 (N_12564,N_11815,N_11437);
nand U12565 (N_12565,N_10675,N_11242);
or U12566 (N_12566,N_10584,N_11167);
and U12567 (N_12567,N_10664,N_11493);
nor U12568 (N_12568,N_10377,N_10512);
nand U12569 (N_12569,N_11364,N_11726);
nand U12570 (N_12570,N_11358,N_10220);
and U12571 (N_12571,N_11614,N_10295);
nor U12572 (N_12572,N_11166,N_11045);
or U12573 (N_12573,N_11563,N_10381);
nor U12574 (N_12574,N_11082,N_11537);
nand U12575 (N_12575,N_11651,N_11548);
nand U12576 (N_12576,N_11785,N_10251);
and U12577 (N_12577,N_10629,N_11330);
nor U12578 (N_12578,N_10067,N_11096);
and U12579 (N_12579,N_11576,N_10492);
nand U12580 (N_12580,N_10935,N_10094);
or U12581 (N_12581,N_11929,N_11603);
or U12582 (N_12582,N_11389,N_11704);
nor U12583 (N_12583,N_11319,N_10239);
nor U12584 (N_12584,N_11919,N_10385);
and U12585 (N_12585,N_10921,N_10728);
nand U12586 (N_12586,N_11965,N_10230);
and U12587 (N_12587,N_10658,N_11250);
nand U12588 (N_12588,N_11538,N_11006);
or U12589 (N_12589,N_10748,N_10737);
and U12590 (N_12590,N_11571,N_10315);
or U12591 (N_12591,N_11284,N_11170);
nor U12592 (N_12592,N_11531,N_10088);
and U12593 (N_12593,N_10010,N_11732);
nand U12594 (N_12594,N_10406,N_11923);
and U12595 (N_12595,N_10330,N_11930);
or U12596 (N_12596,N_10784,N_11918);
nor U12597 (N_12597,N_10676,N_10305);
xor U12598 (N_12598,N_10388,N_10051);
or U12599 (N_12599,N_10101,N_11784);
xnor U12600 (N_12600,N_10500,N_11591);
nand U12601 (N_12601,N_10781,N_10146);
nand U12602 (N_12602,N_10931,N_11987);
xnor U12603 (N_12603,N_11194,N_10331);
nor U12604 (N_12604,N_11527,N_11728);
nand U12605 (N_12605,N_10972,N_10741);
nand U12606 (N_12606,N_11666,N_11146);
nand U12607 (N_12607,N_11659,N_11434);
and U12608 (N_12608,N_10845,N_10624);
nor U12609 (N_12609,N_11347,N_10732);
nor U12610 (N_12610,N_10540,N_10912);
or U12611 (N_12611,N_10226,N_10130);
nor U12612 (N_12612,N_10099,N_11822);
xor U12613 (N_12613,N_11112,N_11561);
xnor U12614 (N_12614,N_10439,N_10299);
nor U12615 (N_12615,N_10630,N_10747);
nand U12616 (N_12616,N_10202,N_11881);
or U12617 (N_12617,N_10907,N_10035);
or U12618 (N_12618,N_11891,N_10120);
nor U12619 (N_12619,N_10693,N_10504);
nor U12620 (N_12620,N_10867,N_10272);
nand U12621 (N_12621,N_10109,N_11222);
nand U12622 (N_12622,N_10707,N_10657);
nor U12623 (N_12623,N_10216,N_11611);
nand U12624 (N_12624,N_10168,N_11834);
xnor U12625 (N_12625,N_11268,N_10358);
nand U12626 (N_12626,N_11367,N_11903);
and U12627 (N_12627,N_10312,N_11157);
and U12628 (N_12628,N_11756,N_11751);
nand U12629 (N_12629,N_10375,N_11964);
or U12630 (N_12630,N_11186,N_10188);
nor U12631 (N_12631,N_11700,N_11765);
and U12632 (N_12632,N_11396,N_11668);
nand U12633 (N_12633,N_10454,N_10659);
nand U12634 (N_12634,N_11460,N_10810);
nand U12635 (N_12635,N_10328,N_11670);
nand U12636 (N_12636,N_11063,N_11619);
or U12637 (N_12637,N_11996,N_11605);
and U12638 (N_12638,N_11233,N_11427);
or U12639 (N_12639,N_10895,N_10196);
nand U12640 (N_12640,N_11406,N_10141);
xor U12641 (N_12641,N_11598,N_10040);
and U12642 (N_12642,N_10537,N_11807);
nor U12643 (N_12643,N_10631,N_10155);
nor U12644 (N_12644,N_10520,N_11452);
or U12645 (N_12645,N_11550,N_11365);
xor U12646 (N_12646,N_11165,N_10806);
or U12647 (N_12647,N_10159,N_10320);
and U12648 (N_12648,N_11750,N_11511);
nor U12649 (N_12649,N_10887,N_10394);
and U12650 (N_12650,N_10812,N_10597);
or U12651 (N_12651,N_11153,N_11136);
and U12652 (N_12652,N_11423,N_10564);
xnor U12653 (N_12653,N_11491,N_11287);
nand U12654 (N_12654,N_10124,N_10451);
nand U12655 (N_12655,N_11076,N_10790);
nand U12656 (N_12656,N_11038,N_10447);
nor U12657 (N_12657,N_11041,N_10474);
xor U12658 (N_12658,N_11712,N_11010);
or U12659 (N_12659,N_11478,N_11594);
or U12660 (N_12660,N_11409,N_10574);
nand U12661 (N_12661,N_10671,N_11381);
and U12662 (N_12662,N_11565,N_10054);
or U12663 (N_12663,N_11230,N_11693);
and U12664 (N_12664,N_10794,N_10736);
and U12665 (N_12665,N_11716,N_11172);
nand U12666 (N_12666,N_11817,N_11269);
nor U12667 (N_12667,N_10553,N_10945);
nand U12668 (N_12668,N_10017,N_10171);
and U12669 (N_12669,N_11580,N_10136);
and U12670 (N_12670,N_11196,N_11386);
nor U12671 (N_12671,N_11339,N_11669);
xor U12672 (N_12672,N_11596,N_11797);
xnor U12673 (N_12673,N_11479,N_10855);
xor U12674 (N_12674,N_11211,N_11678);
or U12675 (N_12675,N_11352,N_10787);
and U12676 (N_12676,N_10832,N_10617);
nor U12677 (N_12677,N_11714,N_11265);
nand U12678 (N_12678,N_10020,N_11556);
or U12679 (N_12679,N_10858,N_10820);
and U12680 (N_12680,N_10275,N_11838);
nor U12681 (N_12681,N_10527,N_11744);
nor U12682 (N_12682,N_10649,N_11144);
and U12683 (N_12683,N_11139,N_11922);
or U12684 (N_12684,N_11914,N_10879);
or U12685 (N_12685,N_10123,N_10232);
and U12686 (N_12686,N_11119,N_11775);
and U12687 (N_12687,N_10811,N_11747);
nor U12688 (N_12688,N_11692,N_10076);
nand U12689 (N_12689,N_10091,N_11799);
or U12690 (N_12690,N_10759,N_10568);
nand U12691 (N_12691,N_10108,N_10558);
and U12692 (N_12692,N_10518,N_11031);
and U12693 (N_12693,N_10625,N_10354);
nor U12694 (N_12694,N_10917,N_10113);
nand U12695 (N_12695,N_11749,N_10708);
and U12696 (N_12696,N_10681,N_11451);
nand U12697 (N_12697,N_10494,N_11504);
and U12698 (N_12698,N_10229,N_10480);
and U12699 (N_12699,N_10669,N_11814);
nor U12700 (N_12700,N_11039,N_10110);
nand U12701 (N_12701,N_10453,N_10104);
and U12702 (N_12702,N_11219,N_10347);
and U12703 (N_12703,N_11982,N_11557);
xnor U12704 (N_12704,N_10007,N_11883);
and U12705 (N_12705,N_10264,N_10992);
nand U12706 (N_12706,N_10666,N_10656);
or U12707 (N_12707,N_11251,N_11536);
nor U12708 (N_12708,N_10796,N_10333);
and U12709 (N_12709,N_10434,N_10433);
nor U12710 (N_12710,N_10158,N_11159);
xnor U12711 (N_12711,N_11534,N_10966);
and U12712 (N_12712,N_10236,N_11936);
nor U12713 (N_12713,N_11524,N_10143);
and U12714 (N_12714,N_10271,N_10670);
xnor U12715 (N_12715,N_10402,N_11069);
nor U12716 (N_12716,N_11609,N_11433);
nand U12717 (N_12717,N_10765,N_10951);
and U12718 (N_12718,N_11421,N_10014);
nor U12719 (N_12719,N_10281,N_11630);
nor U12720 (N_12720,N_10979,N_11723);
or U12721 (N_12721,N_11866,N_10916);
and U12722 (N_12722,N_10640,N_10172);
xnor U12723 (N_12723,N_10713,N_11147);
nand U12724 (N_12724,N_10965,N_10336);
nor U12725 (N_12725,N_11057,N_11079);
nor U12726 (N_12726,N_10899,N_10278);
or U12727 (N_12727,N_11086,N_10542);
and U12728 (N_12728,N_11501,N_10697);
and U12729 (N_12729,N_10986,N_10897);
or U12730 (N_12730,N_10601,N_10217);
xor U12731 (N_12731,N_11616,N_10700);
and U12732 (N_12732,N_11841,N_10600);
or U12733 (N_12733,N_10341,N_10049);
and U12734 (N_12734,N_11664,N_10084);
or U12735 (N_12735,N_11204,N_10829);
or U12736 (N_12736,N_11055,N_11672);
and U12737 (N_12737,N_11819,N_10396);
xnor U12738 (N_12738,N_10036,N_11430);
nand U12739 (N_12739,N_11698,N_11296);
or U12740 (N_12740,N_11471,N_11164);
nand U12741 (N_12741,N_10026,N_10919);
and U12742 (N_12742,N_10775,N_10287);
nor U12743 (N_12743,N_11904,N_10405);
nand U12744 (N_12744,N_10579,N_10711);
nand U12745 (N_12745,N_10989,N_11551);
or U12746 (N_12746,N_11675,N_11925);
nand U12747 (N_12747,N_11525,N_10860);
and U12748 (N_12748,N_10063,N_11114);
xnor U12749 (N_12749,N_10012,N_11699);
nand U12750 (N_12750,N_10642,N_10792);
and U12751 (N_12751,N_11345,N_10276);
or U12752 (N_12752,N_11495,N_11207);
or U12753 (N_12753,N_11032,N_10126);
nor U12754 (N_12754,N_10441,N_11773);
nor U12755 (N_12755,N_10269,N_10443);
and U12756 (N_12756,N_11258,N_10383);
nor U12757 (N_12757,N_11424,N_11011);
nand U12758 (N_12758,N_11018,N_11546);
and U12759 (N_12759,N_11469,N_10983);
nand U12760 (N_12760,N_10023,N_11549);
xor U12761 (N_12761,N_10604,N_10246);
and U12762 (N_12762,N_11342,N_10066);
nand U12763 (N_12763,N_11395,N_11432);
and U12764 (N_12764,N_10720,N_11059);
nor U12765 (N_12765,N_10936,N_10852);
nand U12766 (N_12766,N_10654,N_10208);
nand U12767 (N_12767,N_11582,N_10589);
or U12768 (N_12768,N_11090,N_10884);
nand U12769 (N_12769,N_10195,N_11612);
and U12770 (N_12770,N_11954,N_11143);
nand U12771 (N_12771,N_10535,N_11100);
and U12772 (N_12772,N_10762,N_10241);
or U12773 (N_12773,N_10976,N_11810);
nand U12774 (N_12774,N_10937,N_10047);
nor U12775 (N_12775,N_10121,N_11889);
nor U12776 (N_12776,N_10308,N_10015);
nor U12777 (N_12777,N_10397,N_11502);
nand U12778 (N_12778,N_11373,N_10364);
nor U12779 (N_12779,N_10754,N_10808);
nor U12780 (N_12780,N_11218,N_10115);
and U12781 (N_12781,N_11640,N_10139);
and U12782 (N_12782,N_11988,N_11317);
or U12783 (N_12783,N_11995,N_10846);
nand U12784 (N_12784,N_11253,N_10914);
nor U12785 (N_12785,N_10057,N_10235);
and U12786 (N_12786,N_10772,N_10401);
or U12787 (N_12787,N_10733,N_11174);
nor U12788 (N_12788,N_10977,N_10317);
and U12789 (N_12789,N_10291,N_10243);
and U12790 (N_12790,N_11133,N_10206);
and U12791 (N_12791,N_10734,N_10245);
nor U12792 (N_12792,N_10635,N_10090);
and U12793 (N_12793,N_11971,N_11542);
or U12794 (N_12794,N_11628,N_11811);
or U12795 (N_12795,N_11783,N_11539);
and U12796 (N_12796,N_10598,N_10352);
or U12797 (N_12797,N_11232,N_11790);
and U12798 (N_12798,N_10218,N_10559);
xnor U12799 (N_12799,N_11163,N_11243);
xor U12800 (N_12800,N_11027,N_10791);
nand U12801 (N_12801,N_11262,N_11893);
and U12802 (N_12802,N_10639,N_10957);
and U12803 (N_12803,N_10450,N_10018);
nor U12804 (N_12804,N_10824,N_11943);
nor U12805 (N_12805,N_10390,N_11297);
and U12806 (N_12806,N_10257,N_11293);
and U12807 (N_12807,N_11584,N_10776);
nor U12808 (N_12808,N_11308,N_10510);
or U12809 (N_12809,N_11026,N_10478);
or U12810 (N_12810,N_11888,N_11878);
and U12811 (N_12811,N_10522,N_10363);
nor U12812 (N_12812,N_10404,N_11037);
nand U12813 (N_12813,N_11329,N_11680);
nand U12814 (N_12814,N_10288,N_11375);
and U12815 (N_12815,N_10857,N_11967);
and U12816 (N_12816,N_11727,N_10619);
or U12817 (N_12817,N_10801,N_10623);
nand U12818 (N_12818,N_11397,N_10163);
xnor U12819 (N_12819,N_10552,N_11487);
nand U12820 (N_12820,N_11135,N_11779);
nand U12821 (N_12821,N_11213,N_10758);
nor U12822 (N_12822,N_11349,N_10788);
or U12823 (N_12823,N_10496,N_11562);
or U12824 (N_12824,N_11470,N_10842);
nand U12825 (N_12825,N_11370,N_11357);
or U12826 (N_12826,N_11334,N_10785);
nand U12827 (N_12827,N_11394,N_11791);
and U12828 (N_12828,N_10920,N_11267);
or U12829 (N_12829,N_11856,N_10942);
or U12830 (N_12830,N_10493,N_11391);
and U12831 (N_12831,N_11270,N_11890);
nand U12832 (N_12832,N_11905,N_11854);
xnor U12833 (N_12833,N_10436,N_10484);
xnor U12834 (N_12834,N_10149,N_10150);
xnor U12835 (N_12835,N_10304,N_11886);
nand U12836 (N_12836,N_10578,N_11739);
or U12837 (N_12837,N_10327,N_10915);
and U12838 (N_12838,N_11380,N_11921);
nand U12839 (N_12839,N_10485,N_11862);
and U12840 (N_12840,N_10002,N_11860);
nand U12841 (N_12841,N_11084,N_10191);
or U12842 (N_12842,N_10869,N_10726);
or U12843 (N_12843,N_11774,N_11439);
nand U12844 (N_12844,N_11626,N_11833);
and U12845 (N_12845,N_10802,N_10819);
or U12846 (N_12846,N_11835,N_10081);
and U12847 (N_12847,N_10100,N_11054);
nand U12848 (N_12848,N_10151,N_11189);
nor U12849 (N_12849,N_11602,N_11387);
nor U12850 (N_12850,N_10116,N_11869);
nor U12851 (N_12851,N_10187,N_10703);
nor U12852 (N_12852,N_10069,N_11130);
nand U12853 (N_12853,N_11070,N_10952);
nor U12854 (N_12854,N_10761,N_11798);
nor U12855 (N_12855,N_11657,N_11064);
nand U12856 (N_12856,N_11572,N_11336);
and U12857 (N_12857,N_11378,N_11089);
or U12858 (N_12858,N_11510,N_11068);
nor U12859 (N_12859,N_10465,N_10342);
or U12860 (N_12860,N_10256,N_10460);
and U12861 (N_12861,N_10947,N_11615);
nand U12862 (N_12862,N_11618,N_10543);
nor U12863 (N_12863,N_11622,N_10416);
and U12864 (N_12864,N_11392,N_10201);
nand U12865 (N_12865,N_10958,N_11625);
and U12866 (N_12866,N_10779,N_10050);
nand U12867 (N_12867,N_10499,N_11985);
and U12868 (N_12868,N_11589,N_11821);
and U12869 (N_12869,N_11235,N_11514);
nand U12870 (N_12870,N_10831,N_11519);
xnor U12871 (N_12871,N_11227,N_11685);
or U12872 (N_12872,N_11142,N_11152);
or U12873 (N_12873,N_10803,N_10379);
nor U12874 (N_12874,N_11173,N_10505);
nand U12875 (N_12875,N_11912,N_11674);
nor U12876 (N_12876,N_11915,N_11553);
or U12877 (N_12877,N_11832,N_11962);
nand U12878 (N_12878,N_11661,N_10993);
nand U12879 (N_12879,N_10137,N_11867);
and U12880 (N_12880,N_10079,N_10760);
and U12881 (N_12881,N_11145,N_10903);
or U12882 (N_12882,N_10399,N_10479);
nor U12883 (N_12883,N_10237,N_11371);
nand U12884 (N_12884,N_10544,N_10834);
xnor U12885 (N_12885,N_10296,N_11671);
and U12886 (N_12886,N_11361,N_11738);
or U12887 (N_12887,N_10285,N_10507);
nor U12888 (N_12888,N_10118,N_10142);
nor U12889 (N_12889,N_11442,N_11806);
or U12890 (N_12890,N_11593,N_11870);
nand U12891 (N_12891,N_11990,N_10870);
and U12892 (N_12892,N_11741,N_10901);
nand U12893 (N_12893,N_11474,N_11033);
and U12894 (N_12894,N_11643,N_10605);
and U12895 (N_12895,N_10756,N_11720);
xnor U12896 (N_12896,N_11969,N_11042);
nor U12897 (N_12897,N_11932,N_10089);
and U12898 (N_12898,N_11931,N_11588);
or U12899 (N_12899,N_10111,N_10524);
nand U12900 (N_12900,N_10395,N_11377);
nand U12901 (N_12901,N_10767,N_11825);
nor U12902 (N_12902,N_11566,N_11984);
nor U12903 (N_12903,N_11411,N_11223);
nor U12904 (N_12904,N_10880,N_10987);
nand U12905 (N_12905,N_10529,N_10135);
nand U12906 (N_12906,N_10219,N_10384);
or U12907 (N_12907,N_11494,N_11215);
nand U12908 (N_12908,N_10179,N_11331);
nor U12909 (N_12909,N_10932,N_11466);
xor U12910 (N_12910,N_11859,N_10864);
and U12911 (N_12911,N_10006,N_10890);
nand U12912 (N_12912,N_11118,N_11509);
or U12913 (N_12913,N_10127,N_11115);
nor U12914 (N_12914,N_10576,N_11968);
and U12915 (N_12915,N_11398,N_10250);
xor U12916 (N_12916,N_10566,N_11986);
nor U12917 (N_12917,N_11934,N_10459);
nand U12918 (N_12918,N_11120,N_11244);
nand U12919 (N_12919,N_11944,N_11066);
nor U12920 (N_12920,N_10569,N_10400);
xnor U12921 (N_12921,N_11703,N_11711);
and U12922 (N_12922,N_10706,N_11768);
nor U12923 (N_12923,N_11360,N_10087);
nand U12924 (N_12924,N_11650,N_11770);
nand U12925 (N_12925,N_11180,N_10309);
nor U12926 (N_12926,N_10770,N_10410);
and U12927 (N_12927,N_10817,N_10827);
nand U12928 (N_12928,N_10911,N_10102);
xor U12929 (N_12929,N_10606,N_10055);
and U12930 (N_12930,N_11341,N_11275);
nor U12931 (N_12931,N_11989,N_11629);
or U12932 (N_12932,N_10980,N_11690);
or U12933 (N_12933,N_10209,N_10933);
xnor U12934 (N_12934,N_10411,N_10156);
nor U12935 (N_12935,N_10567,N_10653);
xor U12936 (N_12936,N_10940,N_10677);
nor U12937 (N_12937,N_10854,N_11457);
nand U12938 (N_12938,N_10863,N_10805);
and U12939 (N_12939,N_10562,N_11581);
xnor U12940 (N_12940,N_10003,N_10068);
nand U12941 (N_12941,N_10636,N_10409);
xor U12942 (N_12942,N_10422,N_11892);
or U12943 (N_12943,N_11169,N_10927);
nand U12944 (N_12944,N_10730,N_11024);
nand U12945 (N_12945,N_10978,N_10029);
or U12946 (N_12946,N_10244,N_11316);
nor U12947 (N_12947,N_10421,N_11454);
xnor U12948 (N_12948,N_10144,N_11896);
or U12949 (N_12949,N_11201,N_10795);
nor U12950 (N_12950,N_10948,N_10922);
nand U12951 (N_12951,N_11436,N_10967);
or U12952 (N_12952,N_11555,N_11800);
nand U12953 (N_12953,N_10875,N_11910);
nand U12954 (N_12954,N_11942,N_11695);
nand U12955 (N_12955,N_11132,N_10571);
nand U12956 (N_12956,N_10413,N_10386);
xnor U12957 (N_12957,N_11022,N_10913);
nor U12958 (N_12958,N_10021,N_11652);
nor U12959 (N_12959,N_10138,N_10407);
nor U12960 (N_12960,N_11030,N_11746);
and U12961 (N_12961,N_10892,N_11111);
or U12962 (N_12962,N_11289,N_10261);
or U12963 (N_12963,N_11372,N_11446);
or U12964 (N_12964,N_10471,N_11983);
nor U12965 (N_12965,N_10438,N_11887);
nor U12966 (N_12966,N_10910,N_11288);
or U12967 (N_12967,N_10267,N_11722);
and U12968 (N_12968,N_11979,N_11900);
and U12969 (N_12969,N_11613,N_10175);
and U12970 (N_12970,N_10815,N_10593);
and U12971 (N_12971,N_11950,N_11327);
and U12972 (N_12972,N_10154,N_10644);
and U12973 (N_12973,N_11688,N_10446);
nand U12974 (N_12974,N_11583,N_11894);
nor U12975 (N_12975,N_10367,N_10408);
nor U12976 (N_12976,N_10435,N_10882);
nand U12977 (N_12977,N_10280,N_11101);
nor U12978 (N_12978,N_11758,N_10470);
nand U12979 (N_12979,N_11858,N_10059);
and U12980 (N_12980,N_10835,N_10508);
nor U12981 (N_12981,N_10555,N_10303);
nor U12982 (N_12982,N_10145,N_10648);
nor U12983 (N_12983,N_11104,N_10128);
nor U12984 (N_12984,N_11837,N_10650);
nand U12985 (N_12985,N_11462,N_10686);
or U12986 (N_12986,N_11898,N_10652);
or U12987 (N_12987,N_10426,N_10799);
nor U12988 (N_12988,N_10270,N_10514);
and U12989 (N_12989,N_11021,N_10376);
nor U12990 (N_12990,N_11977,N_10610);
or U12991 (N_12991,N_10632,N_10043);
nor U12992 (N_12992,N_11763,N_11199);
nand U12993 (N_12993,N_11321,N_11848);
xnor U12994 (N_12994,N_11926,N_10092);
and U12995 (N_12995,N_10131,N_11231);
and U12996 (N_12996,N_10563,N_10637);
nor U12997 (N_12997,N_11420,N_10033);
nor U12998 (N_12998,N_11740,N_11676);
nor U12999 (N_12999,N_11441,N_11957);
or U13000 (N_13000,N_10940,N_10759);
nand U13001 (N_13001,N_11063,N_10704);
nand U13002 (N_13002,N_11742,N_10533);
or U13003 (N_13003,N_11344,N_11595);
nand U13004 (N_13004,N_10221,N_10684);
xnor U13005 (N_13005,N_10893,N_10839);
or U13006 (N_13006,N_10977,N_10478);
nand U13007 (N_13007,N_11101,N_10774);
and U13008 (N_13008,N_11145,N_11792);
nand U13009 (N_13009,N_11573,N_11643);
nor U13010 (N_13010,N_10847,N_11797);
nand U13011 (N_13011,N_11459,N_10354);
xnor U13012 (N_13012,N_11886,N_11161);
and U13013 (N_13013,N_11562,N_11626);
or U13014 (N_13014,N_10694,N_10179);
nor U13015 (N_13015,N_11312,N_11266);
nor U13016 (N_13016,N_10279,N_11034);
xnor U13017 (N_13017,N_11425,N_10169);
nand U13018 (N_13018,N_11410,N_11102);
or U13019 (N_13019,N_11405,N_10860);
and U13020 (N_13020,N_11417,N_11089);
or U13021 (N_13021,N_11519,N_10327);
and U13022 (N_13022,N_10202,N_11978);
xor U13023 (N_13023,N_11470,N_11649);
xnor U13024 (N_13024,N_10641,N_10579);
nand U13025 (N_13025,N_11639,N_10417);
nand U13026 (N_13026,N_11107,N_11076);
or U13027 (N_13027,N_11700,N_11222);
xnor U13028 (N_13028,N_10026,N_11426);
or U13029 (N_13029,N_10436,N_11428);
xnor U13030 (N_13030,N_11352,N_11833);
and U13031 (N_13031,N_10286,N_10429);
or U13032 (N_13032,N_11749,N_11780);
and U13033 (N_13033,N_10546,N_10134);
nand U13034 (N_13034,N_10333,N_10870);
xnor U13035 (N_13035,N_11131,N_11620);
nor U13036 (N_13036,N_11485,N_10374);
nor U13037 (N_13037,N_11991,N_10379);
nand U13038 (N_13038,N_10670,N_10032);
and U13039 (N_13039,N_10722,N_10222);
and U13040 (N_13040,N_11226,N_10806);
nor U13041 (N_13041,N_11304,N_10074);
nand U13042 (N_13042,N_10573,N_10112);
xor U13043 (N_13043,N_11284,N_11556);
or U13044 (N_13044,N_11937,N_10788);
or U13045 (N_13045,N_10682,N_11635);
nor U13046 (N_13046,N_10754,N_10220);
nor U13047 (N_13047,N_10018,N_11693);
nor U13048 (N_13048,N_11077,N_10645);
nand U13049 (N_13049,N_11419,N_10135);
nand U13050 (N_13050,N_11696,N_10970);
nand U13051 (N_13051,N_11844,N_11386);
or U13052 (N_13052,N_10365,N_10983);
nand U13053 (N_13053,N_10249,N_11325);
or U13054 (N_13054,N_10400,N_10211);
xnor U13055 (N_13055,N_10772,N_11547);
nand U13056 (N_13056,N_10441,N_11843);
or U13057 (N_13057,N_11965,N_10724);
nand U13058 (N_13058,N_11562,N_11409);
nand U13059 (N_13059,N_11488,N_10618);
nand U13060 (N_13060,N_10321,N_11953);
nand U13061 (N_13061,N_11467,N_11543);
nand U13062 (N_13062,N_10187,N_10131);
or U13063 (N_13063,N_10130,N_10989);
xor U13064 (N_13064,N_10352,N_10398);
nor U13065 (N_13065,N_10962,N_10264);
and U13066 (N_13066,N_10328,N_11048);
and U13067 (N_13067,N_10933,N_10653);
xor U13068 (N_13068,N_11179,N_10966);
or U13069 (N_13069,N_10242,N_10657);
and U13070 (N_13070,N_10360,N_10848);
and U13071 (N_13071,N_10832,N_11083);
nor U13072 (N_13072,N_11966,N_10924);
xor U13073 (N_13073,N_11747,N_10419);
or U13074 (N_13074,N_11755,N_11754);
xnor U13075 (N_13075,N_10991,N_10981);
nor U13076 (N_13076,N_11020,N_10586);
xor U13077 (N_13077,N_10675,N_10371);
nor U13078 (N_13078,N_10637,N_11232);
nor U13079 (N_13079,N_11091,N_11000);
or U13080 (N_13080,N_11734,N_10457);
nor U13081 (N_13081,N_11827,N_11122);
nor U13082 (N_13082,N_10374,N_11392);
nor U13083 (N_13083,N_11129,N_11348);
or U13084 (N_13084,N_11327,N_11286);
nor U13085 (N_13085,N_10922,N_11928);
or U13086 (N_13086,N_11373,N_10162);
nor U13087 (N_13087,N_10300,N_10422);
nand U13088 (N_13088,N_10908,N_11077);
and U13089 (N_13089,N_11110,N_10270);
nor U13090 (N_13090,N_10885,N_10956);
nand U13091 (N_13091,N_10847,N_10591);
or U13092 (N_13092,N_10399,N_10298);
or U13093 (N_13093,N_11459,N_10735);
nand U13094 (N_13094,N_11178,N_10108);
xor U13095 (N_13095,N_10432,N_10351);
or U13096 (N_13096,N_11543,N_10369);
or U13097 (N_13097,N_10428,N_10801);
or U13098 (N_13098,N_11187,N_10632);
and U13099 (N_13099,N_10412,N_10205);
nor U13100 (N_13100,N_11527,N_10579);
or U13101 (N_13101,N_10056,N_11464);
or U13102 (N_13102,N_11766,N_11251);
and U13103 (N_13103,N_10157,N_10799);
and U13104 (N_13104,N_10715,N_10035);
nand U13105 (N_13105,N_11071,N_10242);
nand U13106 (N_13106,N_11677,N_10953);
nand U13107 (N_13107,N_10382,N_10591);
and U13108 (N_13108,N_11656,N_10192);
nor U13109 (N_13109,N_11017,N_11012);
and U13110 (N_13110,N_10787,N_10713);
xor U13111 (N_13111,N_10768,N_10237);
or U13112 (N_13112,N_10841,N_11427);
nor U13113 (N_13113,N_10788,N_10772);
nand U13114 (N_13114,N_11440,N_11223);
nand U13115 (N_13115,N_10853,N_10585);
and U13116 (N_13116,N_10933,N_10407);
nor U13117 (N_13117,N_10828,N_10251);
nor U13118 (N_13118,N_11589,N_11159);
and U13119 (N_13119,N_11212,N_10587);
or U13120 (N_13120,N_10935,N_10991);
nand U13121 (N_13121,N_11530,N_11861);
or U13122 (N_13122,N_10931,N_10959);
and U13123 (N_13123,N_10081,N_10910);
or U13124 (N_13124,N_11035,N_11888);
nor U13125 (N_13125,N_10612,N_11910);
xnor U13126 (N_13126,N_11788,N_10588);
nor U13127 (N_13127,N_11577,N_11728);
nand U13128 (N_13128,N_11343,N_11200);
nor U13129 (N_13129,N_10849,N_10680);
nor U13130 (N_13130,N_11374,N_11289);
and U13131 (N_13131,N_11694,N_10377);
or U13132 (N_13132,N_10259,N_10800);
nand U13133 (N_13133,N_11700,N_11760);
nand U13134 (N_13134,N_11161,N_10236);
nand U13135 (N_13135,N_10881,N_11969);
nor U13136 (N_13136,N_10102,N_11535);
or U13137 (N_13137,N_10263,N_10268);
and U13138 (N_13138,N_10514,N_11479);
and U13139 (N_13139,N_10172,N_10230);
or U13140 (N_13140,N_11208,N_10253);
or U13141 (N_13141,N_11363,N_11099);
or U13142 (N_13142,N_11841,N_10859);
nand U13143 (N_13143,N_10292,N_10382);
nor U13144 (N_13144,N_11923,N_11935);
or U13145 (N_13145,N_11555,N_10058);
nand U13146 (N_13146,N_11520,N_11408);
and U13147 (N_13147,N_11654,N_11841);
and U13148 (N_13148,N_11541,N_11851);
and U13149 (N_13149,N_11364,N_10407);
nand U13150 (N_13150,N_10031,N_10577);
nor U13151 (N_13151,N_10326,N_10864);
or U13152 (N_13152,N_10709,N_11974);
and U13153 (N_13153,N_10279,N_10501);
and U13154 (N_13154,N_11562,N_11997);
nor U13155 (N_13155,N_10811,N_11703);
nor U13156 (N_13156,N_11145,N_11863);
and U13157 (N_13157,N_10797,N_10491);
nand U13158 (N_13158,N_11804,N_11416);
or U13159 (N_13159,N_10791,N_10192);
and U13160 (N_13160,N_11519,N_10906);
or U13161 (N_13161,N_11204,N_11894);
and U13162 (N_13162,N_11179,N_10899);
nor U13163 (N_13163,N_11873,N_10221);
or U13164 (N_13164,N_10450,N_11157);
nand U13165 (N_13165,N_11734,N_10077);
nor U13166 (N_13166,N_11067,N_10039);
xnor U13167 (N_13167,N_11520,N_10305);
nor U13168 (N_13168,N_10220,N_11556);
or U13169 (N_13169,N_10459,N_10256);
nor U13170 (N_13170,N_10723,N_11622);
or U13171 (N_13171,N_10841,N_11225);
nor U13172 (N_13172,N_11981,N_11419);
or U13173 (N_13173,N_11038,N_11495);
and U13174 (N_13174,N_10060,N_11108);
and U13175 (N_13175,N_11204,N_10199);
nor U13176 (N_13176,N_11581,N_10560);
nand U13177 (N_13177,N_10886,N_11966);
nor U13178 (N_13178,N_10598,N_10914);
nor U13179 (N_13179,N_11995,N_11542);
and U13180 (N_13180,N_11626,N_11950);
nand U13181 (N_13181,N_11582,N_11047);
or U13182 (N_13182,N_10853,N_11210);
and U13183 (N_13183,N_11264,N_11694);
xnor U13184 (N_13184,N_11951,N_10042);
or U13185 (N_13185,N_10715,N_10738);
nand U13186 (N_13186,N_10408,N_11985);
and U13187 (N_13187,N_11668,N_11845);
and U13188 (N_13188,N_11693,N_10922);
nor U13189 (N_13189,N_10112,N_11035);
and U13190 (N_13190,N_10805,N_11664);
nand U13191 (N_13191,N_10209,N_11022);
nor U13192 (N_13192,N_10642,N_11278);
or U13193 (N_13193,N_11711,N_11563);
nor U13194 (N_13194,N_10272,N_11808);
or U13195 (N_13195,N_11327,N_10595);
nand U13196 (N_13196,N_10713,N_10166);
or U13197 (N_13197,N_11263,N_10772);
nor U13198 (N_13198,N_11336,N_10496);
and U13199 (N_13199,N_10214,N_11870);
nor U13200 (N_13200,N_11096,N_10093);
nor U13201 (N_13201,N_10507,N_10192);
nand U13202 (N_13202,N_10597,N_10350);
nor U13203 (N_13203,N_10113,N_11625);
nor U13204 (N_13204,N_11078,N_11388);
and U13205 (N_13205,N_10709,N_10650);
xnor U13206 (N_13206,N_10585,N_10961);
and U13207 (N_13207,N_11699,N_11561);
and U13208 (N_13208,N_11976,N_10911);
and U13209 (N_13209,N_11096,N_10183);
nand U13210 (N_13210,N_10010,N_10393);
and U13211 (N_13211,N_10454,N_10971);
and U13212 (N_13212,N_11972,N_10486);
xnor U13213 (N_13213,N_11167,N_10142);
nor U13214 (N_13214,N_10890,N_10796);
nand U13215 (N_13215,N_11290,N_10775);
nand U13216 (N_13216,N_10728,N_11806);
nor U13217 (N_13217,N_10649,N_11586);
xor U13218 (N_13218,N_11295,N_10789);
xor U13219 (N_13219,N_11881,N_10370);
and U13220 (N_13220,N_10173,N_11633);
or U13221 (N_13221,N_10156,N_11213);
and U13222 (N_13222,N_11848,N_11454);
nor U13223 (N_13223,N_10561,N_10789);
nand U13224 (N_13224,N_11503,N_11883);
and U13225 (N_13225,N_11334,N_11786);
or U13226 (N_13226,N_11828,N_10642);
or U13227 (N_13227,N_10616,N_11571);
xor U13228 (N_13228,N_10037,N_11496);
nand U13229 (N_13229,N_11030,N_10459);
nand U13230 (N_13230,N_11461,N_11796);
and U13231 (N_13231,N_10471,N_10672);
nand U13232 (N_13232,N_10720,N_10657);
nor U13233 (N_13233,N_10664,N_10817);
or U13234 (N_13234,N_11941,N_11259);
xor U13235 (N_13235,N_11442,N_10647);
or U13236 (N_13236,N_11706,N_10483);
nand U13237 (N_13237,N_11269,N_11200);
or U13238 (N_13238,N_10196,N_10136);
and U13239 (N_13239,N_10609,N_11896);
nor U13240 (N_13240,N_10503,N_11717);
or U13241 (N_13241,N_10277,N_10702);
nor U13242 (N_13242,N_11900,N_10790);
nand U13243 (N_13243,N_11094,N_11627);
nor U13244 (N_13244,N_11573,N_11722);
or U13245 (N_13245,N_11326,N_11024);
and U13246 (N_13246,N_10702,N_11252);
or U13247 (N_13247,N_11378,N_10212);
or U13248 (N_13248,N_11817,N_10011);
nand U13249 (N_13249,N_11822,N_10629);
nand U13250 (N_13250,N_10298,N_10960);
and U13251 (N_13251,N_11029,N_10502);
nor U13252 (N_13252,N_11653,N_11373);
nand U13253 (N_13253,N_11079,N_11751);
nor U13254 (N_13254,N_10840,N_10081);
and U13255 (N_13255,N_10379,N_11084);
or U13256 (N_13256,N_10027,N_11129);
or U13257 (N_13257,N_11116,N_11843);
nand U13258 (N_13258,N_11746,N_10965);
and U13259 (N_13259,N_10116,N_11715);
and U13260 (N_13260,N_11695,N_11662);
nand U13261 (N_13261,N_11811,N_11731);
nor U13262 (N_13262,N_10669,N_10794);
and U13263 (N_13263,N_11701,N_11932);
and U13264 (N_13264,N_10447,N_10154);
nand U13265 (N_13265,N_10632,N_10976);
and U13266 (N_13266,N_10182,N_10924);
and U13267 (N_13267,N_10567,N_11303);
and U13268 (N_13268,N_10180,N_11522);
and U13269 (N_13269,N_10338,N_10248);
nor U13270 (N_13270,N_10250,N_10477);
and U13271 (N_13271,N_11373,N_11167);
nand U13272 (N_13272,N_11126,N_10850);
nand U13273 (N_13273,N_11718,N_11629);
and U13274 (N_13274,N_10913,N_11506);
nand U13275 (N_13275,N_11074,N_10491);
or U13276 (N_13276,N_11159,N_10990);
nand U13277 (N_13277,N_10376,N_11932);
nand U13278 (N_13278,N_11148,N_10537);
or U13279 (N_13279,N_10420,N_11031);
nand U13280 (N_13280,N_11427,N_10677);
and U13281 (N_13281,N_10783,N_10002);
xor U13282 (N_13282,N_10073,N_10068);
nor U13283 (N_13283,N_11313,N_10011);
nor U13284 (N_13284,N_11221,N_10094);
nand U13285 (N_13285,N_10503,N_11939);
or U13286 (N_13286,N_11702,N_10096);
and U13287 (N_13287,N_11042,N_11769);
nand U13288 (N_13288,N_10921,N_10599);
nand U13289 (N_13289,N_11361,N_11008);
and U13290 (N_13290,N_10644,N_10672);
nand U13291 (N_13291,N_11776,N_10087);
nor U13292 (N_13292,N_11996,N_11100);
nor U13293 (N_13293,N_10291,N_10858);
nor U13294 (N_13294,N_10005,N_10449);
nand U13295 (N_13295,N_11617,N_11709);
xnor U13296 (N_13296,N_10671,N_11656);
nand U13297 (N_13297,N_11829,N_10549);
or U13298 (N_13298,N_10318,N_10535);
and U13299 (N_13299,N_11561,N_11600);
and U13300 (N_13300,N_11994,N_11825);
and U13301 (N_13301,N_10566,N_10270);
and U13302 (N_13302,N_10258,N_10315);
or U13303 (N_13303,N_10726,N_10834);
nand U13304 (N_13304,N_10702,N_11626);
and U13305 (N_13305,N_11397,N_11304);
nor U13306 (N_13306,N_10123,N_11464);
or U13307 (N_13307,N_10053,N_11193);
nand U13308 (N_13308,N_11716,N_10881);
and U13309 (N_13309,N_11545,N_11796);
or U13310 (N_13310,N_11142,N_11995);
or U13311 (N_13311,N_11199,N_11271);
nand U13312 (N_13312,N_11739,N_11516);
nor U13313 (N_13313,N_10873,N_11810);
nor U13314 (N_13314,N_11097,N_10508);
nand U13315 (N_13315,N_11170,N_10262);
or U13316 (N_13316,N_10838,N_11727);
or U13317 (N_13317,N_11837,N_11589);
and U13318 (N_13318,N_11450,N_10952);
nand U13319 (N_13319,N_10325,N_10364);
or U13320 (N_13320,N_11767,N_11420);
or U13321 (N_13321,N_10010,N_11487);
nand U13322 (N_13322,N_10606,N_10936);
or U13323 (N_13323,N_11434,N_11167);
xor U13324 (N_13324,N_10864,N_11170);
nand U13325 (N_13325,N_11858,N_11149);
nand U13326 (N_13326,N_11224,N_11689);
or U13327 (N_13327,N_11579,N_10735);
nand U13328 (N_13328,N_10636,N_10847);
or U13329 (N_13329,N_10692,N_10280);
and U13330 (N_13330,N_10806,N_11748);
and U13331 (N_13331,N_10215,N_11480);
xor U13332 (N_13332,N_11989,N_11917);
nand U13333 (N_13333,N_10355,N_11039);
nor U13334 (N_13334,N_11357,N_10581);
or U13335 (N_13335,N_10727,N_11423);
and U13336 (N_13336,N_11153,N_11699);
nand U13337 (N_13337,N_11706,N_10848);
and U13338 (N_13338,N_11249,N_11673);
nand U13339 (N_13339,N_11760,N_10631);
xnor U13340 (N_13340,N_10867,N_10310);
nor U13341 (N_13341,N_10357,N_11578);
nand U13342 (N_13342,N_11972,N_11147);
xor U13343 (N_13343,N_11090,N_11054);
nand U13344 (N_13344,N_11023,N_10618);
and U13345 (N_13345,N_10201,N_10839);
and U13346 (N_13346,N_10290,N_11557);
or U13347 (N_13347,N_10189,N_10006);
nor U13348 (N_13348,N_10324,N_11505);
nor U13349 (N_13349,N_10216,N_11259);
and U13350 (N_13350,N_10128,N_11698);
nor U13351 (N_13351,N_11061,N_11342);
nor U13352 (N_13352,N_11818,N_11750);
nor U13353 (N_13353,N_11446,N_10233);
xor U13354 (N_13354,N_10371,N_11237);
or U13355 (N_13355,N_10436,N_10113);
nand U13356 (N_13356,N_11720,N_11676);
or U13357 (N_13357,N_10490,N_11859);
nor U13358 (N_13358,N_11058,N_10495);
or U13359 (N_13359,N_11978,N_10950);
nor U13360 (N_13360,N_11002,N_11006);
or U13361 (N_13361,N_10638,N_11448);
and U13362 (N_13362,N_11579,N_10700);
and U13363 (N_13363,N_10686,N_11281);
nand U13364 (N_13364,N_11342,N_11293);
nand U13365 (N_13365,N_10572,N_10180);
nor U13366 (N_13366,N_11327,N_11410);
nor U13367 (N_13367,N_10183,N_11701);
or U13368 (N_13368,N_11445,N_10571);
and U13369 (N_13369,N_11461,N_11010);
nor U13370 (N_13370,N_10712,N_10094);
nand U13371 (N_13371,N_10947,N_11587);
and U13372 (N_13372,N_10641,N_10552);
or U13373 (N_13373,N_11485,N_10565);
or U13374 (N_13374,N_10893,N_11311);
or U13375 (N_13375,N_10737,N_11827);
or U13376 (N_13376,N_10087,N_10146);
nand U13377 (N_13377,N_10869,N_10360);
nor U13378 (N_13378,N_11359,N_10803);
nand U13379 (N_13379,N_11601,N_11525);
nor U13380 (N_13380,N_11218,N_10747);
nor U13381 (N_13381,N_10835,N_10375);
and U13382 (N_13382,N_10280,N_11911);
nand U13383 (N_13383,N_11375,N_10727);
nand U13384 (N_13384,N_11233,N_11487);
and U13385 (N_13385,N_10811,N_11827);
nor U13386 (N_13386,N_10880,N_10518);
and U13387 (N_13387,N_10847,N_11356);
nand U13388 (N_13388,N_10053,N_11933);
or U13389 (N_13389,N_11656,N_11345);
or U13390 (N_13390,N_11559,N_11902);
xnor U13391 (N_13391,N_10769,N_11020);
nor U13392 (N_13392,N_11843,N_10354);
and U13393 (N_13393,N_11847,N_10454);
nand U13394 (N_13394,N_10256,N_11763);
nor U13395 (N_13395,N_11462,N_10014);
and U13396 (N_13396,N_10481,N_11612);
nor U13397 (N_13397,N_11482,N_11740);
or U13398 (N_13398,N_11837,N_11081);
or U13399 (N_13399,N_11356,N_10312);
and U13400 (N_13400,N_11639,N_10089);
nand U13401 (N_13401,N_11965,N_11314);
nand U13402 (N_13402,N_11910,N_10631);
and U13403 (N_13403,N_11487,N_10676);
and U13404 (N_13404,N_11869,N_10755);
and U13405 (N_13405,N_10225,N_11746);
and U13406 (N_13406,N_10910,N_10101);
nor U13407 (N_13407,N_11667,N_10954);
and U13408 (N_13408,N_10100,N_11882);
xor U13409 (N_13409,N_10649,N_10492);
and U13410 (N_13410,N_10842,N_11959);
xnor U13411 (N_13411,N_10505,N_10814);
and U13412 (N_13412,N_11812,N_11144);
nand U13413 (N_13413,N_10986,N_11184);
and U13414 (N_13414,N_10157,N_11745);
nand U13415 (N_13415,N_10609,N_10435);
nand U13416 (N_13416,N_10311,N_10493);
nor U13417 (N_13417,N_11049,N_10534);
or U13418 (N_13418,N_11378,N_10613);
nand U13419 (N_13419,N_10206,N_10330);
or U13420 (N_13420,N_11603,N_11828);
xor U13421 (N_13421,N_11172,N_10575);
or U13422 (N_13422,N_10437,N_11937);
or U13423 (N_13423,N_11065,N_10726);
nand U13424 (N_13424,N_10185,N_11701);
nand U13425 (N_13425,N_10285,N_10887);
nor U13426 (N_13426,N_11901,N_11012);
xor U13427 (N_13427,N_10673,N_11680);
nor U13428 (N_13428,N_11108,N_10290);
nor U13429 (N_13429,N_10022,N_10100);
nor U13430 (N_13430,N_10780,N_10135);
and U13431 (N_13431,N_11369,N_10199);
xnor U13432 (N_13432,N_10517,N_10085);
nor U13433 (N_13433,N_11758,N_11777);
nor U13434 (N_13434,N_10135,N_10705);
or U13435 (N_13435,N_11376,N_10633);
nor U13436 (N_13436,N_11111,N_11866);
or U13437 (N_13437,N_11623,N_11542);
and U13438 (N_13438,N_11757,N_10948);
nand U13439 (N_13439,N_10804,N_11375);
nor U13440 (N_13440,N_10497,N_11167);
nand U13441 (N_13441,N_10835,N_11116);
nand U13442 (N_13442,N_11580,N_11529);
xor U13443 (N_13443,N_10704,N_11641);
nor U13444 (N_13444,N_10869,N_11954);
nor U13445 (N_13445,N_11762,N_10635);
and U13446 (N_13446,N_10461,N_10531);
nand U13447 (N_13447,N_10900,N_11928);
and U13448 (N_13448,N_10940,N_10562);
and U13449 (N_13449,N_11920,N_11294);
nand U13450 (N_13450,N_10236,N_11628);
nor U13451 (N_13451,N_10303,N_10095);
and U13452 (N_13452,N_11082,N_10360);
nand U13453 (N_13453,N_11489,N_10661);
nor U13454 (N_13454,N_11271,N_10454);
nor U13455 (N_13455,N_11633,N_10473);
and U13456 (N_13456,N_10036,N_10886);
xor U13457 (N_13457,N_10472,N_11449);
nand U13458 (N_13458,N_11873,N_10526);
or U13459 (N_13459,N_10414,N_10378);
nand U13460 (N_13460,N_11808,N_11551);
nand U13461 (N_13461,N_10033,N_11303);
and U13462 (N_13462,N_10090,N_11830);
nand U13463 (N_13463,N_11659,N_11765);
nor U13464 (N_13464,N_11033,N_11526);
and U13465 (N_13465,N_11884,N_11128);
nor U13466 (N_13466,N_10904,N_11105);
nor U13467 (N_13467,N_11270,N_10008);
and U13468 (N_13468,N_10407,N_11895);
nand U13469 (N_13469,N_10578,N_10730);
nor U13470 (N_13470,N_11869,N_10018);
nand U13471 (N_13471,N_11431,N_10032);
nor U13472 (N_13472,N_11772,N_11266);
and U13473 (N_13473,N_10958,N_11501);
nand U13474 (N_13474,N_11883,N_11021);
nor U13475 (N_13475,N_10566,N_10482);
nor U13476 (N_13476,N_10209,N_11060);
and U13477 (N_13477,N_11915,N_11325);
xor U13478 (N_13478,N_11905,N_10465);
nor U13479 (N_13479,N_10665,N_10068);
xnor U13480 (N_13480,N_11722,N_11656);
nor U13481 (N_13481,N_11444,N_10535);
and U13482 (N_13482,N_10879,N_10130);
and U13483 (N_13483,N_10027,N_10768);
or U13484 (N_13484,N_10562,N_10049);
nand U13485 (N_13485,N_11434,N_11822);
xor U13486 (N_13486,N_11535,N_10387);
or U13487 (N_13487,N_10510,N_10396);
nand U13488 (N_13488,N_10288,N_10734);
nand U13489 (N_13489,N_10430,N_11735);
or U13490 (N_13490,N_11592,N_11602);
or U13491 (N_13491,N_11969,N_10028);
xor U13492 (N_13492,N_10104,N_10007);
or U13493 (N_13493,N_10847,N_11032);
xnor U13494 (N_13494,N_11572,N_10159);
or U13495 (N_13495,N_11665,N_11330);
and U13496 (N_13496,N_10308,N_11166);
nor U13497 (N_13497,N_10397,N_11634);
and U13498 (N_13498,N_10478,N_11555);
and U13499 (N_13499,N_10819,N_11367);
and U13500 (N_13500,N_11690,N_11131);
or U13501 (N_13501,N_10944,N_10424);
nor U13502 (N_13502,N_10370,N_10692);
nor U13503 (N_13503,N_10998,N_10069);
or U13504 (N_13504,N_10383,N_10598);
nand U13505 (N_13505,N_11186,N_11870);
or U13506 (N_13506,N_10774,N_11912);
nand U13507 (N_13507,N_11817,N_11023);
and U13508 (N_13508,N_10469,N_10915);
nand U13509 (N_13509,N_10694,N_11078);
nor U13510 (N_13510,N_11624,N_10415);
or U13511 (N_13511,N_11138,N_11269);
and U13512 (N_13512,N_10553,N_11504);
nor U13513 (N_13513,N_10579,N_10520);
or U13514 (N_13514,N_11448,N_10051);
xor U13515 (N_13515,N_10914,N_10862);
xor U13516 (N_13516,N_10173,N_11103);
nand U13517 (N_13517,N_11985,N_10368);
and U13518 (N_13518,N_11628,N_10301);
and U13519 (N_13519,N_11020,N_11763);
xor U13520 (N_13520,N_11893,N_11986);
and U13521 (N_13521,N_10491,N_10973);
nand U13522 (N_13522,N_10048,N_10414);
xnor U13523 (N_13523,N_10527,N_10711);
nand U13524 (N_13524,N_11996,N_10563);
xor U13525 (N_13525,N_10107,N_10888);
nand U13526 (N_13526,N_11077,N_10089);
nand U13527 (N_13527,N_11969,N_10642);
nor U13528 (N_13528,N_11672,N_11133);
and U13529 (N_13529,N_11639,N_10363);
nand U13530 (N_13530,N_11821,N_11128);
nand U13531 (N_13531,N_10258,N_10127);
nor U13532 (N_13532,N_11758,N_10386);
or U13533 (N_13533,N_11531,N_11737);
or U13534 (N_13534,N_11260,N_10226);
and U13535 (N_13535,N_11315,N_10842);
or U13536 (N_13536,N_10320,N_10840);
nand U13537 (N_13537,N_10969,N_11848);
nor U13538 (N_13538,N_11280,N_10704);
nor U13539 (N_13539,N_10483,N_11906);
and U13540 (N_13540,N_11044,N_11216);
or U13541 (N_13541,N_10713,N_11770);
nand U13542 (N_13542,N_11536,N_11633);
or U13543 (N_13543,N_10869,N_11630);
xor U13544 (N_13544,N_10690,N_10299);
xnor U13545 (N_13545,N_10297,N_11791);
nor U13546 (N_13546,N_10171,N_10901);
nand U13547 (N_13547,N_11298,N_10539);
or U13548 (N_13548,N_11658,N_10056);
and U13549 (N_13549,N_10042,N_11918);
xor U13550 (N_13550,N_10921,N_11060);
xnor U13551 (N_13551,N_10733,N_11743);
nand U13552 (N_13552,N_10485,N_10292);
nand U13553 (N_13553,N_10280,N_11414);
or U13554 (N_13554,N_11272,N_11138);
and U13555 (N_13555,N_11447,N_11656);
nor U13556 (N_13556,N_11130,N_11294);
and U13557 (N_13557,N_10643,N_10467);
nor U13558 (N_13558,N_11501,N_11937);
nand U13559 (N_13559,N_10243,N_10385);
or U13560 (N_13560,N_11491,N_11288);
or U13561 (N_13561,N_10421,N_11000);
nor U13562 (N_13562,N_10277,N_11759);
nor U13563 (N_13563,N_11766,N_11579);
and U13564 (N_13564,N_11060,N_10732);
and U13565 (N_13565,N_10562,N_11473);
nor U13566 (N_13566,N_10107,N_10334);
or U13567 (N_13567,N_10304,N_10083);
or U13568 (N_13568,N_11611,N_11552);
and U13569 (N_13569,N_11822,N_11112);
or U13570 (N_13570,N_11831,N_11352);
and U13571 (N_13571,N_10756,N_10289);
and U13572 (N_13572,N_10472,N_11683);
and U13573 (N_13573,N_10973,N_11414);
nand U13574 (N_13574,N_11945,N_11745);
nand U13575 (N_13575,N_10813,N_10210);
and U13576 (N_13576,N_10807,N_11118);
xor U13577 (N_13577,N_10354,N_11598);
nor U13578 (N_13578,N_10447,N_11186);
nand U13579 (N_13579,N_10877,N_10637);
and U13580 (N_13580,N_11298,N_10510);
or U13581 (N_13581,N_10168,N_10384);
nor U13582 (N_13582,N_11728,N_11448);
and U13583 (N_13583,N_10744,N_10704);
and U13584 (N_13584,N_10618,N_10698);
and U13585 (N_13585,N_11217,N_11073);
xor U13586 (N_13586,N_10057,N_11025);
or U13587 (N_13587,N_10976,N_11883);
nand U13588 (N_13588,N_11121,N_10615);
and U13589 (N_13589,N_11132,N_10714);
nand U13590 (N_13590,N_11133,N_11948);
nand U13591 (N_13591,N_10980,N_11277);
xor U13592 (N_13592,N_10264,N_11632);
and U13593 (N_13593,N_11391,N_10664);
and U13594 (N_13594,N_10512,N_10408);
xor U13595 (N_13595,N_10289,N_10497);
nand U13596 (N_13596,N_11305,N_11920);
nand U13597 (N_13597,N_10137,N_10566);
and U13598 (N_13598,N_11435,N_10492);
or U13599 (N_13599,N_11324,N_10247);
or U13600 (N_13600,N_11132,N_11877);
or U13601 (N_13601,N_10087,N_11057);
nand U13602 (N_13602,N_10610,N_11197);
or U13603 (N_13603,N_11384,N_11234);
and U13604 (N_13604,N_11153,N_10795);
nor U13605 (N_13605,N_10207,N_10130);
nand U13606 (N_13606,N_10383,N_10667);
and U13607 (N_13607,N_11346,N_11335);
or U13608 (N_13608,N_11357,N_10642);
or U13609 (N_13609,N_10224,N_11328);
or U13610 (N_13610,N_10020,N_11853);
or U13611 (N_13611,N_11778,N_11439);
nor U13612 (N_13612,N_10205,N_10636);
nor U13613 (N_13613,N_10687,N_11704);
and U13614 (N_13614,N_11291,N_11331);
and U13615 (N_13615,N_10898,N_10929);
nor U13616 (N_13616,N_10499,N_10489);
and U13617 (N_13617,N_11614,N_11191);
nor U13618 (N_13618,N_11578,N_10700);
and U13619 (N_13619,N_10819,N_11398);
nor U13620 (N_13620,N_11938,N_11904);
or U13621 (N_13621,N_10186,N_10111);
nand U13622 (N_13622,N_11452,N_10996);
nor U13623 (N_13623,N_11411,N_10109);
nor U13624 (N_13624,N_10967,N_11944);
nand U13625 (N_13625,N_10294,N_10956);
nor U13626 (N_13626,N_10934,N_10984);
nand U13627 (N_13627,N_11278,N_10050);
nand U13628 (N_13628,N_10149,N_11918);
or U13629 (N_13629,N_10848,N_10718);
nor U13630 (N_13630,N_11486,N_10743);
nor U13631 (N_13631,N_11467,N_10282);
nor U13632 (N_13632,N_11235,N_11816);
nand U13633 (N_13633,N_11416,N_11301);
or U13634 (N_13634,N_10553,N_11048);
and U13635 (N_13635,N_10111,N_10353);
and U13636 (N_13636,N_11431,N_11704);
or U13637 (N_13637,N_11874,N_11262);
or U13638 (N_13638,N_11380,N_10334);
and U13639 (N_13639,N_10128,N_10581);
nand U13640 (N_13640,N_11419,N_10782);
or U13641 (N_13641,N_11731,N_11369);
or U13642 (N_13642,N_11897,N_11246);
nand U13643 (N_13643,N_10110,N_11448);
nor U13644 (N_13644,N_11569,N_11589);
or U13645 (N_13645,N_11477,N_10406);
nand U13646 (N_13646,N_10427,N_10410);
nor U13647 (N_13647,N_11129,N_11189);
and U13648 (N_13648,N_10610,N_11029);
or U13649 (N_13649,N_10402,N_10349);
or U13650 (N_13650,N_10657,N_11914);
nand U13651 (N_13651,N_11907,N_11984);
nor U13652 (N_13652,N_11109,N_10333);
or U13653 (N_13653,N_10726,N_11825);
nor U13654 (N_13654,N_11355,N_10062);
or U13655 (N_13655,N_11613,N_10370);
and U13656 (N_13656,N_11243,N_11762);
or U13657 (N_13657,N_10645,N_11593);
xor U13658 (N_13658,N_10574,N_10784);
and U13659 (N_13659,N_11714,N_11223);
or U13660 (N_13660,N_10176,N_11182);
nand U13661 (N_13661,N_11620,N_11190);
and U13662 (N_13662,N_10333,N_10763);
nor U13663 (N_13663,N_10130,N_10463);
and U13664 (N_13664,N_10689,N_11991);
or U13665 (N_13665,N_11068,N_11642);
nor U13666 (N_13666,N_11560,N_11098);
nor U13667 (N_13667,N_10033,N_11080);
and U13668 (N_13668,N_10552,N_11548);
and U13669 (N_13669,N_11270,N_11077);
nand U13670 (N_13670,N_10861,N_10488);
nor U13671 (N_13671,N_11008,N_11562);
or U13672 (N_13672,N_11113,N_10211);
xnor U13673 (N_13673,N_11194,N_10596);
or U13674 (N_13674,N_11006,N_11490);
or U13675 (N_13675,N_11076,N_10091);
or U13676 (N_13676,N_11666,N_11316);
or U13677 (N_13677,N_11267,N_10490);
nor U13678 (N_13678,N_10932,N_11900);
and U13679 (N_13679,N_10024,N_10537);
and U13680 (N_13680,N_11548,N_11498);
nor U13681 (N_13681,N_10633,N_11463);
nand U13682 (N_13682,N_10885,N_11230);
and U13683 (N_13683,N_10130,N_10271);
nand U13684 (N_13684,N_10814,N_11774);
nor U13685 (N_13685,N_10564,N_11600);
nor U13686 (N_13686,N_10884,N_10144);
nor U13687 (N_13687,N_11992,N_10762);
or U13688 (N_13688,N_11884,N_11364);
xor U13689 (N_13689,N_10468,N_11811);
xor U13690 (N_13690,N_11331,N_11316);
nor U13691 (N_13691,N_11327,N_11688);
or U13692 (N_13692,N_10498,N_10940);
and U13693 (N_13693,N_10850,N_11940);
nand U13694 (N_13694,N_10154,N_11401);
and U13695 (N_13695,N_11176,N_11699);
and U13696 (N_13696,N_11585,N_11935);
nor U13697 (N_13697,N_11281,N_10115);
and U13698 (N_13698,N_10518,N_10834);
nor U13699 (N_13699,N_11470,N_10373);
and U13700 (N_13700,N_11155,N_10751);
nor U13701 (N_13701,N_10195,N_10118);
nand U13702 (N_13702,N_10632,N_11888);
or U13703 (N_13703,N_10872,N_10006);
and U13704 (N_13704,N_11584,N_10423);
or U13705 (N_13705,N_10179,N_11123);
or U13706 (N_13706,N_11531,N_10096);
nor U13707 (N_13707,N_11001,N_10228);
and U13708 (N_13708,N_10486,N_11445);
nor U13709 (N_13709,N_11770,N_11243);
or U13710 (N_13710,N_10681,N_10608);
nand U13711 (N_13711,N_11407,N_11907);
and U13712 (N_13712,N_11615,N_11767);
and U13713 (N_13713,N_11651,N_10163);
xor U13714 (N_13714,N_10858,N_11985);
or U13715 (N_13715,N_10401,N_10897);
or U13716 (N_13716,N_11597,N_10141);
xnor U13717 (N_13717,N_11972,N_11317);
xnor U13718 (N_13718,N_10938,N_11062);
xor U13719 (N_13719,N_11045,N_11312);
nor U13720 (N_13720,N_10446,N_11342);
nand U13721 (N_13721,N_11238,N_10432);
or U13722 (N_13722,N_11452,N_11859);
xor U13723 (N_13723,N_10614,N_11491);
and U13724 (N_13724,N_11212,N_10134);
and U13725 (N_13725,N_11375,N_11146);
or U13726 (N_13726,N_10428,N_10560);
nand U13727 (N_13727,N_10350,N_10719);
nor U13728 (N_13728,N_10939,N_11490);
and U13729 (N_13729,N_10440,N_10742);
nand U13730 (N_13730,N_11266,N_10274);
nor U13731 (N_13731,N_11490,N_11821);
or U13732 (N_13732,N_11569,N_10550);
nand U13733 (N_13733,N_11442,N_11904);
and U13734 (N_13734,N_10012,N_10366);
xnor U13735 (N_13735,N_10170,N_11528);
nor U13736 (N_13736,N_10874,N_11964);
or U13737 (N_13737,N_11856,N_11297);
nor U13738 (N_13738,N_10567,N_11581);
xor U13739 (N_13739,N_11608,N_11189);
nor U13740 (N_13740,N_11201,N_11345);
nand U13741 (N_13741,N_10388,N_10987);
nor U13742 (N_13742,N_11921,N_11357);
or U13743 (N_13743,N_10780,N_11781);
nor U13744 (N_13744,N_10569,N_10262);
xor U13745 (N_13745,N_10442,N_11019);
nor U13746 (N_13746,N_10165,N_11045);
nor U13747 (N_13747,N_10229,N_11526);
and U13748 (N_13748,N_11688,N_11965);
or U13749 (N_13749,N_10286,N_10914);
and U13750 (N_13750,N_11285,N_10777);
xnor U13751 (N_13751,N_11357,N_11416);
or U13752 (N_13752,N_10933,N_11356);
nand U13753 (N_13753,N_10966,N_10843);
xnor U13754 (N_13754,N_11015,N_11896);
nor U13755 (N_13755,N_11834,N_10726);
nand U13756 (N_13756,N_11790,N_11477);
nor U13757 (N_13757,N_11402,N_11578);
or U13758 (N_13758,N_11069,N_11523);
or U13759 (N_13759,N_10291,N_10708);
nand U13760 (N_13760,N_11337,N_11633);
and U13761 (N_13761,N_11246,N_11789);
and U13762 (N_13762,N_10509,N_11856);
or U13763 (N_13763,N_11695,N_11008);
nor U13764 (N_13764,N_10033,N_10175);
or U13765 (N_13765,N_11639,N_11901);
nor U13766 (N_13766,N_11595,N_11437);
and U13767 (N_13767,N_11904,N_11079);
xnor U13768 (N_13768,N_10380,N_11712);
xnor U13769 (N_13769,N_11836,N_11960);
xor U13770 (N_13770,N_11954,N_10608);
xnor U13771 (N_13771,N_11742,N_11374);
nor U13772 (N_13772,N_10402,N_11000);
and U13773 (N_13773,N_10751,N_11729);
nor U13774 (N_13774,N_11054,N_10457);
nor U13775 (N_13775,N_10100,N_10341);
and U13776 (N_13776,N_11451,N_10194);
or U13777 (N_13777,N_11238,N_11798);
nor U13778 (N_13778,N_11724,N_11854);
nor U13779 (N_13779,N_11517,N_11691);
nand U13780 (N_13780,N_10136,N_11723);
nand U13781 (N_13781,N_11253,N_10648);
nor U13782 (N_13782,N_11912,N_11871);
nand U13783 (N_13783,N_11083,N_11916);
nor U13784 (N_13784,N_10446,N_10897);
nor U13785 (N_13785,N_11498,N_11098);
and U13786 (N_13786,N_10801,N_11594);
nand U13787 (N_13787,N_10104,N_10153);
and U13788 (N_13788,N_10744,N_11577);
xor U13789 (N_13789,N_10334,N_11330);
and U13790 (N_13790,N_11468,N_11802);
nand U13791 (N_13791,N_10031,N_11958);
and U13792 (N_13792,N_10419,N_10708);
nor U13793 (N_13793,N_10118,N_11389);
and U13794 (N_13794,N_11012,N_10777);
nand U13795 (N_13795,N_10171,N_11889);
xnor U13796 (N_13796,N_11748,N_11647);
and U13797 (N_13797,N_11624,N_11009);
and U13798 (N_13798,N_11972,N_10907);
and U13799 (N_13799,N_11297,N_11410);
nand U13800 (N_13800,N_11017,N_11343);
and U13801 (N_13801,N_10077,N_11377);
or U13802 (N_13802,N_11681,N_11425);
nand U13803 (N_13803,N_11409,N_10634);
and U13804 (N_13804,N_10678,N_11100);
nor U13805 (N_13805,N_11744,N_11134);
or U13806 (N_13806,N_10584,N_11031);
and U13807 (N_13807,N_11311,N_10695);
or U13808 (N_13808,N_10676,N_11783);
nor U13809 (N_13809,N_11336,N_11884);
or U13810 (N_13810,N_11044,N_11696);
or U13811 (N_13811,N_10610,N_11779);
or U13812 (N_13812,N_10657,N_11116);
nand U13813 (N_13813,N_10195,N_10162);
nand U13814 (N_13814,N_11372,N_10211);
xnor U13815 (N_13815,N_10793,N_11991);
nand U13816 (N_13816,N_11538,N_10332);
or U13817 (N_13817,N_10163,N_10459);
xnor U13818 (N_13818,N_11424,N_10555);
and U13819 (N_13819,N_10014,N_11223);
and U13820 (N_13820,N_10838,N_10579);
nor U13821 (N_13821,N_10934,N_11785);
or U13822 (N_13822,N_11680,N_11006);
nor U13823 (N_13823,N_10758,N_10902);
nor U13824 (N_13824,N_10000,N_11203);
and U13825 (N_13825,N_10626,N_11483);
nand U13826 (N_13826,N_11467,N_11131);
and U13827 (N_13827,N_11458,N_11592);
nor U13828 (N_13828,N_11904,N_11145);
nor U13829 (N_13829,N_10543,N_10406);
xnor U13830 (N_13830,N_11422,N_11263);
xor U13831 (N_13831,N_10378,N_11767);
or U13832 (N_13832,N_11766,N_10329);
nand U13833 (N_13833,N_11220,N_11473);
xnor U13834 (N_13834,N_10027,N_10274);
or U13835 (N_13835,N_10731,N_11545);
nor U13836 (N_13836,N_10102,N_11296);
nand U13837 (N_13837,N_11204,N_11535);
nor U13838 (N_13838,N_11691,N_11573);
nand U13839 (N_13839,N_10109,N_11066);
or U13840 (N_13840,N_10758,N_11654);
nor U13841 (N_13841,N_10612,N_11438);
nor U13842 (N_13842,N_10647,N_11662);
or U13843 (N_13843,N_10576,N_11708);
xor U13844 (N_13844,N_11202,N_10870);
nor U13845 (N_13845,N_11945,N_10182);
nand U13846 (N_13846,N_10917,N_11659);
nand U13847 (N_13847,N_11825,N_11819);
or U13848 (N_13848,N_11789,N_11279);
nor U13849 (N_13849,N_10253,N_11672);
or U13850 (N_13850,N_10238,N_11857);
and U13851 (N_13851,N_11175,N_11446);
xnor U13852 (N_13852,N_10453,N_11557);
nor U13853 (N_13853,N_10020,N_10416);
or U13854 (N_13854,N_11820,N_11618);
and U13855 (N_13855,N_11714,N_11957);
nor U13856 (N_13856,N_11018,N_10081);
nand U13857 (N_13857,N_11719,N_11449);
or U13858 (N_13858,N_11256,N_10839);
xnor U13859 (N_13859,N_11594,N_11034);
and U13860 (N_13860,N_10467,N_11468);
and U13861 (N_13861,N_10808,N_10387);
xnor U13862 (N_13862,N_10168,N_10545);
nor U13863 (N_13863,N_10058,N_10331);
nand U13864 (N_13864,N_10360,N_10489);
nand U13865 (N_13865,N_11944,N_10328);
and U13866 (N_13866,N_11080,N_11384);
nand U13867 (N_13867,N_10117,N_11105);
and U13868 (N_13868,N_11276,N_10322);
nand U13869 (N_13869,N_11602,N_11320);
nor U13870 (N_13870,N_10379,N_10920);
or U13871 (N_13871,N_11321,N_10647);
nand U13872 (N_13872,N_11303,N_11895);
or U13873 (N_13873,N_10422,N_11484);
nand U13874 (N_13874,N_10480,N_11044);
xor U13875 (N_13875,N_10630,N_11483);
nand U13876 (N_13876,N_11172,N_10400);
nand U13877 (N_13877,N_10248,N_11792);
xnor U13878 (N_13878,N_11897,N_10116);
nand U13879 (N_13879,N_10443,N_11978);
or U13880 (N_13880,N_10271,N_11239);
or U13881 (N_13881,N_10831,N_11750);
nor U13882 (N_13882,N_11534,N_10808);
nand U13883 (N_13883,N_10313,N_10567);
or U13884 (N_13884,N_10688,N_11371);
nor U13885 (N_13885,N_11461,N_11752);
or U13886 (N_13886,N_10923,N_10561);
and U13887 (N_13887,N_10101,N_10981);
nor U13888 (N_13888,N_10273,N_10270);
nor U13889 (N_13889,N_11104,N_10221);
or U13890 (N_13890,N_10384,N_10694);
nand U13891 (N_13891,N_11653,N_11668);
nor U13892 (N_13892,N_10533,N_11672);
nor U13893 (N_13893,N_10806,N_10211);
nor U13894 (N_13894,N_11706,N_10248);
nand U13895 (N_13895,N_10736,N_11282);
or U13896 (N_13896,N_10671,N_11492);
or U13897 (N_13897,N_11529,N_10292);
or U13898 (N_13898,N_10945,N_11988);
nor U13899 (N_13899,N_10996,N_11829);
nor U13900 (N_13900,N_10230,N_11182);
nor U13901 (N_13901,N_10009,N_10589);
nor U13902 (N_13902,N_10906,N_10220);
nand U13903 (N_13903,N_10045,N_11688);
xor U13904 (N_13904,N_11601,N_11548);
or U13905 (N_13905,N_11817,N_10780);
nand U13906 (N_13906,N_11415,N_11930);
nor U13907 (N_13907,N_11381,N_10906);
or U13908 (N_13908,N_11931,N_11745);
nand U13909 (N_13909,N_10715,N_10366);
or U13910 (N_13910,N_10595,N_11482);
and U13911 (N_13911,N_10092,N_11267);
or U13912 (N_13912,N_10526,N_10323);
nand U13913 (N_13913,N_11563,N_10711);
xor U13914 (N_13914,N_10909,N_11619);
or U13915 (N_13915,N_10658,N_10253);
or U13916 (N_13916,N_11197,N_10344);
and U13917 (N_13917,N_11210,N_11592);
and U13918 (N_13918,N_10180,N_11854);
or U13919 (N_13919,N_10432,N_11493);
nor U13920 (N_13920,N_10483,N_11673);
xor U13921 (N_13921,N_10530,N_11136);
xor U13922 (N_13922,N_10976,N_10595);
and U13923 (N_13923,N_11408,N_10135);
or U13924 (N_13924,N_10906,N_11147);
nor U13925 (N_13925,N_11795,N_11934);
and U13926 (N_13926,N_10685,N_10524);
xor U13927 (N_13927,N_11625,N_10676);
nand U13928 (N_13928,N_10971,N_10587);
nor U13929 (N_13929,N_10460,N_10570);
or U13930 (N_13930,N_10027,N_10278);
xnor U13931 (N_13931,N_10181,N_11496);
or U13932 (N_13932,N_11414,N_11766);
nor U13933 (N_13933,N_10723,N_11477);
xnor U13934 (N_13934,N_10726,N_11581);
xor U13935 (N_13935,N_11217,N_11744);
nor U13936 (N_13936,N_10257,N_11201);
and U13937 (N_13937,N_11980,N_10450);
nor U13938 (N_13938,N_10802,N_11679);
and U13939 (N_13939,N_10252,N_11199);
or U13940 (N_13940,N_11479,N_10255);
or U13941 (N_13941,N_11032,N_10588);
nor U13942 (N_13942,N_10852,N_10629);
and U13943 (N_13943,N_11190,N_10461);
xor U13944 (N_13944,N_10855,N_10872);
or U13945 (N_13945,N_10270,N_11782);
nor U13946 (N_13946,N_11043,N_10994);
xnor U13947 (N_13947,N_10459,N_11294);
nor U13948 (N_13948,N_10405,N_11326);
nor U13949 (N_13949,N_10801,N_11506);
nor U13950 (N_13950,N_10857,N_11381);
and U13951 (N_13951,N_10563,N_10079);
and U13952 (N_13952,N_10920,N_11185);
and U13953 (N_13953,N_10147,N_10377);
or U13954 (N_13954,N_11454,N_10612);
nor U13955 (N_13955,N_11385,N_10676);
nand U13956 (N_13956,N_10409,N_11688);
nor U13957 (N_13957,N_10164,N_11317);
and U13958 (N_13958,N_10059,N_10549);
nor U13959 (N_13959,N_11636,N_10860);
nor U13960 (N_13960,N_10915,N_10015);
nand U13961 (N_13961,N_11752,N_11508);
and U13962 (N_13962,N_11777,N_10511);
nor U13963 (N_13963,N_11872,N_10084);
and U13964 (N_13964,N_10736,N_10028);
or U13965 (N_13965,N_10008,N_11859);
nand U13966 (N_13966,N_10895,N_10642);
nand U13967 (N_13967,N_11069,N_11426);
nor U13968 (N_13968,N_10810,N_11866);
and U13969 (N_13969,N_10053,N_10690);
or U13970 (N_13970,N_10054,N_11868);
nand U13971 (N_13971,N_10521,N_10977);
and U13972 (N_13972,N_11687,N_10747);
or U13973 (N_13973,N_11422,N_11467);
nand U13974 (N_13974,N_10768,N_11732);
or U13975 (N_13975,N_10707,N_10215);
nor U13976 (N_13976,N_10604,N_10502);
and U13977 (N_13977,N_10912,N_11798);
or U13978 (N_13978,N_10113,N_10795);
or U13979 (N_13979,N_11911,N_11262);
nor U13980 (N_13980,N_10561,N_11349);
nand U13981 (N_13981,N_10648,N_11557);
xor U13982 (N_13982,N_11509,N_10997);
xor U13983 (N_13983,N_11677,N_10984);
nor U13984 (N_13984,N_10913,N_11589);
and U13985 (N_13985,N_11776,N_11608);
xor U13986 (N_13986,N_10951,N_11942);
xor U13987 (N_13987,N_10468,N_10814);
xor U13988 (N_13988,N_10872,N_10669);
or U13989 (N_13989,N_10157,N_10260);
nor U13990 (N_13990,N_11956,N_10761);
nor U13991 (N_13991,N_10565,N_10225);
or U13992 (N_13992,N_11847,N_10322);
nand U13993 (N_13993,N_10760,N_11208);
and U13994 (N_13994,N_11697,N_11800);
or U13995 (N_13995,N_10683,N_11966);
or U13996 (N_13996,N_11314,N_10715);
or U13997 (N_13997,N_11294,N_11029);
and U13998 (N_13998,N_11695,N_10252);
and U13999 (N_13999,N_10608,N_10044);
nand U14000 (N_14000,N_13094,N_12515);
nor U14001 (N_14001,N_13255,N_12681);
nor U14002 (N_14002,N_13970,N_12524);
and U14003 (N_14003,N_12690,N_12677);
and U14004 (N_14004,N_12935,N_12883);
nand U14005 (N_14005,N_13782,N_12821);
nand U14006 (N_14006,N_12854,N_12492);
nor U14007 (N_14007,N_13979,N_13186);
xnor U14008 (N_14008,N_13381,N_12746);
and U14009 (N_14009,N_12792,N_12428);
xnor U14010 (N_14010,N_12111,N_13329);
or U14011 (N_14011,N_13508,N_12068);
nand U14012 (N_14012,N_12061,N_13232);
nor U14013 (N_14013,N_13993,N_12268);
and U14014 (N_14014,N_13967,N_12998);
and U14015 (N_14015,N_12537,N_13715);
or U14016 (N_14016,N_12619,N_12432);
or U14017 (N_14017,N_12645,N_13128);
or U14018 (N_14018,N_13224,N_13441);
nor U14019 (N_14019,N_13348,N_12714);
nor U14020 (N_14020,N_13866,N_12699);
and U14021 (N_14021,N_12323,N_13501);
or U14022 (N_14022,N_12433,N_13101);
nand U14023 (N_14023,N_13641,N_12596);
nand U14024 (N_14024,N_12188,N_13990);
or U14025 (N_14025,N_12761,N_12072);
nor U14026 (N_14026,N_13603,N_13959);
nand U14027 (N_14027,N_12488,N_12707);
or U14028 (N_14028,N_13520,N_12523);
and U14029 (N_14029,N_13007,N_12048);
or U14030 (N_14030,N_12158,N_12413);
nand U14031 (N_14031,N_12888,N_12083);
and U14032 (N_14032,N_12280,N_12286);
and U14033 (N_14033,N_13669,N_13947);
nor U14034 (N_14034,N_12261,N_13153);
nand U14035 (N_14035,N_13732,N_13734);
xor U14036 (N_14036,N_12972,N_13108);
and U14037 (N_14037,N_13871,N_13429);
and U14038 (N_14038,N_12832,N_12922);
nand U14039 (N_14039,N_12153,N_12607);
or U14040 (N_14040,N_13697,N_13614);
and U14041 (N_14041,N_12529,N_13221);
nand U14042 (N_14042,N_13371,N_13756);
or U14043 (N_14043,N_12456,N_13623);
or U14044 (N_14044,N_12866,N_12422);
nor U14045 (N_14045,N_12304,N_13066);
or U14046 (N_14046,N_13801,N_13189);
nand U14047 (N_14047,N_13927,N_12363);
xnor U14048 (N_14048,N_12631,N_12013);
or U14049 (N_14049,N_12467,N_12656);
or U14050 (N_14050,N_13410,N_12267);
or U14051 (N_14051,N_13594,N_12225);
nor U14052 (N_14052,N_12450,N_13804);
and U14053 (N_14053,N_13021,N_13686);
or U14054 (N_14054,N_12169,N_13719);
or U14055 (N_14055,N_13576,N_13952);
and U14056 (N_14056,N_13735,N_13122);
nand U14057 (N_14057,N_12898,N_12787);
and U14058 (N_14058,N_12655,N_12613);
and U14059 (N_14059,N_13730,N_13575);
nand U14060 (N_14060,N_13018,N_12771);
or U14061 (N_14061,N_12041,N_13542);
nor U14062 (N_14062,N_13815,N_13290);
nor U14063 (N_14063,N_13605,N_12675);
nand U14064 (N_14064,N_12844,N_12958);
or U14065 (N_14065,N_13176,N_13105);
nand U14066 (N_14066,N_13031,N_12510);
nor U14067 (N_14067,N_13848,N_12591);
xnor U14068 (N_14068,N_13945,N_12824);
xor U14069 (N_14069,N_13426,N_13858);
and U14070 (N_14070,N_13088,N_13302);
nor U14071 (N_14071,N_13338,N_13402);
and U14072 (N_14072,N_12633,N_13138);
nand U14073 (N_14073,N_13654,N_13928);
nor U14074 (N_14074,N_12617,N_12109);
nand U14075 (N_14075,N_13244,N_13786);
nor U14076 (N_14076,N_13687,N_13359);
and U14077 (N_14077,N_13968,N_12600);
and U14078 (N_14078,N_12748,N_12058);
nand U14079 (N_14079,N_12717,N_13091);
and U14080 (N_14080,N_13891,N_13171);
nor U14081 (N_14081,N_13494,N_12978);
or U14082 (N_14082,N_13530,N_13937);
nand U14083 (N_14083,N_13659,N_12604);
nand U14084 (N_14084,N_12130,N_13152);
and U14085 (N_14085,N_12031,N_12870);
and U14086 (N_14086,N_13405,N_13033);
nor U14087 (N_14087,N_12352,N_12419);
nor U14088 (N_14088,N_13689,N_12984);
or U14089 (N_14089,N_12723,N_12299);
and U14090 (N_14090,N_12751,N_13898);
or U14091 (N_14091,N_13397,N_12789);
and U14092 (N_14092,N_13477,N_13643);
nand U14093 (N_14093,N_13379,N_12330);
and U14094 (N_14094,N_12506,N_12000);
nor U14095 (N_14095,N_13438,N_13214);
nor U14096 (N_14096,N_13001,N_12414);
and U14097 (N_14097,N_13401,N_13292);
and U14098 (N_14098,N_13330,N_12634);
nand U14099 (N_14099,N_13295,N_12378);
or U14100 (N_14100,N_12444,N_12765);
and U14101 (N_14101,N_13747,N_13087);
and U14102 (N_14102,N_12121,N_13580);
or U14103 (N_14103,N_13256,N_12140);
xor U14104 (N_14104,N_12118,N_12172);
nand U14105 (N_14105,N_13878,N_12811);
and U14106 (N_14106,N_13874,N_13781);
nor U14107 (N_14107,N_12548,N_13608);
nor U14108 (N_14108,N_13535,N_13618);
and U14109 (N_14109,N_12520,N_13591);
nand U14110 (N_14110,N_13099,N_12359);
and U14111 (N_14111,N_12451,N_13588);
nor U14112 (N_14112,N_13355,N_13067);
or U14113 (N_14113,N_13427,N_12021);
and U14114 (N_14114,N_13272,N_13439);
and U14115 (N_14115,N_12369,N_13294);
or U14116 (N_14116,N_12217,N_13276);
or U14117 (N_14117,N_12229,N_12740);
or U14118 (N_14118,N_12878,N_12370);
or U14119 (N_14119,N_13082,N_12266);
nor U14120 (N_14120,N_13070,N_12547);
and U14121 (N_14121,N_12598,N_12705);
and U14122 (N_14122,N_12875,N_13777);
or U14123 (N_14123,N_13203,N_13502);
xnor U14124 (N_14124,N_13519,N_13054);
or U14125 (N_14125,N_13469,N_12987);
nand U14126 (N_14126,N_12610,N_12429);
xnor U14127 (N_14127,N_12231,N_13653);
and U14128 (N_14128,N_13773,N_12522);
and U14129 (N_14129,N_13022,N_12084);
or U14130 (N_14130,N_13289,N_12621);
and U14131 (N_14131,N_12049,N_13319);
nor U14132 (N_14132,N_13870,N_13960);
and U14133 (N_14133,N_13935,N_13922);
or U14134 (N_14134,N_12500,N_12016);
or U14135 (N_14135,N_13629,N_12802);
nand U14136 (N_14136,N_12496,N_12385);
nand U14137 (N_14137,N_12806,N_13452);
nand U14138 (N_14138,N_13504,N_12373);
nand U14139 (N_14139,N_13146,N_13123);
nand U14140 (N_14140,N_13262,N_12503);
xnor U14141 (N_14141,N_12146,N_12336);
or U14142 (N_14142,N_12839,N_13399);
or U14143 (N_14143,N_13482,N_12417);
and U14144 (N_14144,N_12137,N_13717);
nor U14145 (N_14145,N_12601,N_12653);
nor U14146 (N_14146,N_13060,N_13005);
xor U14147 (N_14147,N_12788,N_13322);
xor U14148 (N_14148,N_13911,N_12930);
and U14149 (N_14149,N_12669,N_12890);
xnor U14150 (N_14150,N_13881,N_12278);
xnor U14151 (N_14151,N_12850,N_12238);
or U14152 (N_14152,N_12774,N_12840);
or U14153 (N_14153,N_13627,N_13073);
nor U14154 (N_14154,N_12973,N_12003);
and U14155 (N_14155,N_13674,N_12145);
or U14156 (N_14156,N_12443,N_12697);
and U14157 (N_14157,N_12934,N_13671);
or U14158 (N_14158,N_13305,N_13523);
nand U14159 (N_14159,N_12693,N_12906);
or U14160 (N_14160,N_12994,N_12480);
nand U14161 (N_14161,N_12779,N_12818);
nand U14162 (N_14162,N_13062,N_13778);
nand U14163 (N_14163,N_13155,N_13896);
or U14164 (N_14164,N_12571,N_12383);
or U14165 (N_14165,N_12493,N_12351);
nor U14166 (N_14166,N_12482,N_12262);
or U14167 (N_14167,N_12104,N_12425);
nor U14168 (N_14168,N_12290,N_13611);
or U14169 (N_14169,N_13989,N_13373);
nor U14170 (N_14170,N_13071,N_12614);
nand U14171 (N_14171,N_13190,N_12531);
nand U14172 (N_14172,N_12347,N_12661);
xor U14173 (N_14173,N_13846,N_12495);
and U14174 (N_14174,N_12962,N_13318);
or U14175 (N_14175,N_13484,N_12243);
xnor U14176 (N_14176,N_12168,N_13829);
and U14177 (N_14177,N_12464,N_13303);
or U14178 (N_14178,N_13585,N_13586);
or U14179 (N_14179,N_12241,N_13098);
and U14180 (N_14180,N_13841,N_13115);
or U14181 (N_14181,N_13182,N_12739);
and U14182 (N_14182,N_13393,N_13263);
and U14183 (N_14183,N_13584,N_12042);
and U14184 (N_14184,N_12170,N_13178);
and U14185 (N_14185,N_12702,N_13995);
nand U14186 (N_14186,N_12341,N_12557);
nor U14187 (N_14187,N_13370,N_13795);
nor U14188 (N_14188,N_13750,N_13454);
nand U14189 (N_14189,N_12585,N_12305);
nor U14190 (N_14190,N_12222,N_13316);
nor U14191 (N_14191,N_13187,N_12986);
nor U14192 (N_14192,N_13195,N_13383);
nor U14193 (N_14193,N_12708,N_13474);
or U14194 (N_14194,N_12486,N_12476);
nand U14195 (N_14195,N_12391,N_13038);
nor U14196 (N_14196,N_12009,N_13710);
and U14197 (N_14197,N_12459,N_12865);
nor U14198 (N_14198,N_12030,N_13562);
nor U14199 (N_14199,N_13248,N_13518);
nand U14200 (N_14200,N_12975,N_13754);
nand U14201 (N_14201,N_13549,N_12289);
nor U14202 (N_14202,N_13577,N_12452);
nor U14203 (N_14203,N_13156,N_12579);
nor U14204 (N_14204,N_13388,N_12043);
or U14205 (N_14205,N_12673,N_13720);
and U14206 (N_14206,N_12635,N_13568);
and U14207 (N_14207,N_13226,N_12512);
nand U14208 (N_14208,N_13826,N_13113);
nor U14209 (N_14209,N_13444,N_12320);
nor U14210 (N_14210,N_13844,N_13657);
xor U14211 (N_14211,N_13579,N_13705);
and U14212 (N_14212,N_13432,N_13948);
nor U14213 (N_14213,N_12773,N_12107);
nor U14214 (N_14214,N_13737,N_13034);
or U14215 (N_14215,N_13408,N_13544);
xnor U14216 (N_14216,N_12680,N_12144);
nand U14217 (N_14217,N_12593,N_13764);
nand U14218 (N_14218,N_13078,N_13800);
and U14219 (N_14219,N_12536,N_13956);
and U14220 (N_14220,N_12210,N_12535);
or U14221 (N_14221,N_12882,N_13837);
or U14222 (N_14222,N_13802,N_13278);
xnor U14223 (N_14223,N_12827,N_12331);
and U14224 (N_14224,N_13218,N_12244);
and U14225 (N_14225,N_13499,N_13570);
nor U14226 (N_14226,N_13599,N_13298);
xor U14227 (N_14227,N_12295,N_12204);
and U14228 (N_14228,N_13957,N_13711);
nand U14229 (N_14229,N_12113,N_12662);
nor U14230 (N_14230,N_12993,N_12442);
nand U14231 (N_14231,N_13017,N_12559);
and U14232 (N_14232,N_13539,N_12402);
or U14233 (N_14233,N_12270,N_13930);
nor U14234 (N_14234,N_12542,N_12195);
xor U14235 (N_14235,N_12284,N_13035);
or U14236 (N_14236,N_12939,N_13617);
nor U14237 (N_14237,N_12475,N_13722);
or U14238 (N_14238,N_13739,N_12649);
nand U14239 (N_14239,N_12793,N_12065);
nand U14240 (N_14240,N_13158,N_13661);
and U14241 (N_14241,N_12110,N_13363);
and U14242 (N_14242,N_12149,N_13974);
xor U14243 (N_14243,N_13548,N_13210);
nand U14244 (N_14244,N_13762,N_12213);
nand U14245 (N_14245,N_13423,N_13431);
or U14246 (N_14246,N_13842,N_12623);
xnor U14247 (N_14247,N_13966,N_13776);
nor U14248 (N_14248,N_13695,N_12810);
xnor U14249 (N_14249,N_12497,N_13273);
xor U14250 (N_14250,N_12720,N_12660);
nor U14251 (N_14251,N_13490,N_12778);
nand U14252 (N_14252,N_13709,N_13307);
nor U14253 (N_14253,N_12205,N_12164);
nor U14254 (N_14254,N_13904,N_13699);
nand U14255 (N_14255,N_12874,N_12264);
nand U14256 (N_14256,N_12037,N_12160);
nand U14257 (N_14257,N_12240,N_13811);
nand U14258 (N_14258,N_12434,N_13486);
nor U14259 (N_14259,N_12325,N_12219);
and U14260 (N_14260,N_13257,N_13693);
nor U14261 (N_14261,N_12063,N_12629);
xor U14262 (N_14262,N_12365,N_12499);
or U14263 (N_14263,N_13933,N_13978);
nand U14264 (N_14264,N_12277,N_13511);
and U14265 (N_14265,N_12212,N_12872);
nor U14266 (N_14266,N_12200,N_12927);
nor U14267 (N_14267,N_13600,N_13415);
or U14268 (N_14268,N_12981,N_12027);
xor U14269 (N_14269,N_12823,N_13185);
or U14270 (N_14270,N_13932,N_13984);
or U14271 (N_14271,N_12904,N_13425);
nand U14272 (N_14272,N_12155,N_13336);
and U14273 (N_14273,N_13134,N_13803);
and U14274 (N_14274,N_13524,N_12586);
nor U14275 (N_14275,N_13421,N_13026);
xnor U14276 (N_14276,N_13745,N_12375);
xnor U14277 (N_14277,N_12609,N_13680);
nand U14278 (N_14278,N_12952,N_13822);
nor U14279 (N_14279,N_12296,N_13647);
or U14280 (N_14280,N_13707,N_12867);
and U14281 (N_14281,N_12902,N_12310);
or U14282 (N_14282,N_12969,N_12999);
nand U14283 (N_14283,N_13788,N_13704);
xnor U14284 (N_14284,N_12989,N_13516);
nor U14285 (N_14285,N_13166,N_13321);
nand U14286 (N_14286,N_12471,N_12851);
nand U14287 (N_14287,N_13172,N_12166);
or U14288 (N_14288,N_13250,N_12887);
xor U14289 (N_14289,N_12173,N_13840);
or U14290 (N_14290,N_13596,N_12763);
or U14291 (N_14291,N_13996,N_13897);
nor U14292 (N_14292,N_12424,N_13817);
and U14293 (N_14293,N_12466,N_13767);
or U14294 (N_14294,N_12950,N_12570);
nor U14295 (N_14295,N_13268,N_13827);
xnor U14296 (N_14296,N_13943,N_12057);
nand U14297 (N_14297,N_13857,N_12961);
nor U14298 (N_14298,N_13451,N_13412);
nand U14299 (N_14299,N_13768,N_13326);
or U14300 (N_14300,N_12576,N_12514);
and U14301 (N_14301,N_12259,N_13170);
or U14302 (N_14302,N_13147,N_13604);
nand U14303 (N_14303,N_13275,N_13664);
or U14304 (N_14304,N_12676,N_12314);
and U14305 (N_14305,N_13616,N_12915);
nor U14306 (N_14306,N_12033,N_12519);
and U14307 (N_14307,N_12148,N_13914);
nor U14308 (N_14308,N_12594,N_12005);
nor U14309 (N_14309,N_13666,N_13880);
nor U14310 (N_14310,N_13708,N_13053);
nand U14311 (N_14311,N_12606,N_12291);
nor U14312 (N_14312,N_13798,N_12807);
xor U14313 (N_14313,N_12316,N_12885);
nand U14314 (N_14314,N_12179,N_12122);
or U14315 (N_14315,N_13650,N_13656);
xnor U14316 (N_14316,N_12124,N_12324);
nand U14317 (N_14317,N_12136,N_13306);
or U14318 (N_14318,N_12154,N_13912);
and U14319 (N_14319,N_13744,N_13567);
nand U14320 (N_14320,N_12618,N_12349);
or U14321 (N_14321,N_12128,N_12097);
nor U14322 (N_14322,N_13240,N_13890);
and U14323 (N_14323,N_13217,N_12843);
nor U14324 (N_14324,N_13267,N_12937);
nand U14325 (N_14325,N_13908,N_13994);
nand U14326 (N_14326,N_13304,N_12599);
nand U14327 (N_14327,N_12929,N_13673);
xnor U14328 (N_14328,N_13068,N_12620);
nor U14329 (N_14329,N_13222,N_12230);
xnor U14330 (N_14330,N_12592,N_12207);
and U14331 (N_14331,N_13249,N_12731);
or U14332 (N_14332,N_12393,N_13929);
or U14333 (N_14333,N_12448,N_12340);
nand U14334 (N_14334,N_12400,N_12625);
nor U14335 (N_14335,N_13497,N_12199);
and U14336 (N_14336,N_13774,N_12218);
nand U14337 (N_14337,N_12756,N_12275);
nor U14338 (N_14338,N_12157,N_13339);
and U14339 (N_14339,N_13903,N_13847);
and U14340 (N_14340,N_12518,N_12006);
and U14341 (N_14341,N_13029,N_13097);
and U14342 (N_14342,N_13814,N_13785);
nor U14343 (N_14343,N_13824,N_13713);
or U14344 (N_14344,N_13706,N_12208);
xnor U14345 (N_14345,N_13049,N_13300);
or U14346 (N_14346,N_12710,N_13938);
and U14347 (N_14347,N_12931,N_12394);
or U14348 (N_14348,N_12193,N_13748);
nor U14349 (N_14349,N_12098,N_12627);
nor U14350 (N_14350,N_13965,N_13864);
and U14351 (N_14351,N_13135,N_13149);
xor U14352 (N_14352,N_12064,N_13377);
or U14353 (N_14353,N_12736,N_12747);
xor U14354 (N_14354,N_13503,N_12783);
or U14355 (N_14355,N_12300,N_13942);
xor U14356 (N_14356,N_12611,N_12313);
nand U14357 (N_14357,N_13521,N_12265);
and U14358 (N_14358,N_12010,N_12501);
or U14359 (N_14359,N_13213,N_13834);
and U14360 (N_14360,N_13064,N_12786);
nand U14361 (N_14361,N_13331,N_12076);
and U14362 (N_14362,N_12232,N_13312);
nand U14363 (N_14363,N_12504,N_12439);
nand U14364 (N_14364,N_13601,N_12580);
nor U14365 (N_14365,N_13905,N_13512);
or U14366 (N_14366,N_13724,N_12988);
nand U14367 (N_14367,N_13681,N_12901);
or U14368 (N_14368,N_13351,N_13875);
and U14369 (N_14369,N_13116,N_13685);
nor U14370 (N_14370,N_12868,N_12508);
nand U14371 (N_14371,N_13980,N_12017);
nand U14372 (N_14372,N_12597,N_12541);
or U14373 (N_14373,N_12381,N_13853);
nor U14374 (N_14374,N_12943,N_13074);
or U14375 (N_14375,N_12663,N_12859);
nand U14376 (N_14376,N_12423,N_12722);
nor U14377 (N_14377,N_13635,N_12582);
and U14378 (N_14378,N_13004,N_12877);
xnor U14379 (N_14379,N_13201,N_12054);
and U14380 (N_14380,N_12185,N_13760);
or U14381 (N_14381,N_12298,N_13027);
nand U14382 (N_14382,N_13725,N_13495);
and U14383 (N_14383,N_12646,N_12552);
and U14384 (N_14384,N_13587,N_13254);
xnor U14385 (N_14385,N_12741,N_12389);
xor U14386 (N_14386,N_12980,N_13437);
and U14387 (N_14387,N_12913,N_13531);
and U14388 (N_14388,N_13310,N_12632);
or U14389 (N_14389,N_12180,N_13416);
nor U14390 (N_14390,N_12940,N_12420);
or U14391 (N_14391,N_12431,N_13016);
nand U14392 (N_14392,N_13525,N_13683);
and U14393 (N_14393,N_12735,N_13944);
and U14394 (N_14394,N_12835,N_12641);
and U14395 (N_14395,N_12970,N_13471);
nand U14396 (N_14396,N_13237,N_12554);
or U14397 (N_14397,N_13385,N_12762);
and U14398 (N_14398,N_13610,N_13492);
nor U14399 (N_14399,N_13564,N_12654);
nand U14400 (N_14400,N_12382,N_12134);
nand U14401 (N_14401,N_12979,N_13335);
or U14402 (N_14402,N_12791,N_12116);
xor U14403 (N_14403,N_12814,N_12317);
xor U14404 (N_14404,N_12358,N_12990);
nor U14405 (N_14405,N_13882,N_13270);
or U14406 (N_14406,N_12647,N_12752);
nand U14407 (N_14407,N_13340,N_12689);
and U14408 (N_14408,N_13063,N_13574);
nand U14409 (N_14409,N_12344,N_13380);
nor U14410 (N_14410,N_12896,N_12454);
nor U14411 (N_14411,N_13085,N_12672);
and U14412 (N_14412,N_12530,N_13046);
xor U14413 (N_14413,N_13095,N_12734);
nand U14414 (N_14414,N_13855,N_13859);
nor U14415 (N_14415,N_12678,N_13793);
and U14416 (N_14416,N_12540,N_13867);
nor U14417 (N_14417,N_12051,N_12228);
and U14418 (N_14418,N_13736,N_13281);
nand U14419 (N_14419,N_12666,N_13327);
nor U14420 (N_14420,N_12318,N_13631);
and U14421 (N_14421,N_12477,N_12440);
and U14422 (N_14422,N_13663,N_13924);
or U14423 (N_14423,N_13626,N_12131);
and U14424 (N_14424,N_13301,N_12837);
nand U14425 (N_14425,N_12976,N_13821);
nand U14426 (N_14426,N_13649,N_12366);
or U14427 (N_14427,N_13532,N_13433);
or U14428 (N_14428,N_13332,N_12725);
and U14429 (N_14429,N_12384,N_12355);
or U14430 (N_14430,N_13110,N_12630);
and U14431 (N_14431,N_12465,N_13833);
nor U14432 (N_14432,N_13805,N_13458);
and U14433 (N_14433,N_13375,N_12838);
and U14434 (N_14434,N_13806,N_12463);
and U14435 (N_14435,N_12665,N_12447);
or U14436 (N_14436,N_12936,N_12095);
or U14437 (N_14437,N_13131,N_13258);
nor U14438 (N_14438,N_12982,N_12664);
or U14439 (N_14439,N_13537,N_13220);
nor U14440 (N_14440,N_12545,N_12768);
nor U14441 (N_14441,N_13212,N_13569);
nand U14442 (N_14442,N_13396,N_12018);
and U14443 (N_14443,N_12801,N_13856);
nor U14444 (N_14444,N_12511,N_13140);
and U14445 (N_14445,N_13488,N_13252);
xor U14446 (N_14446,N_12086,N_13025);
nor U14447 (N_14447,N_12667,N_12652);
nor U14448 (N_14448,N_13287,N_12082);
and U14449 (N_14449,N_13354,N_13015);
or U14450 (N_14450,N_12825,N_12997);
or U14451 (N_14451,N_12159,N_12679);
nand U14452 (N_14452,N_12845,N_12099);
nand U14453 (N_14453,N_13753,N_13797);
and U14454 (N_14454,N_12028,N_13161);
nand U14455 (N_14455,N_12588,N_13002);
nand U14456 (N_14456,N_13790,N_13314);
nand U14457 (N_14457,N_13992,N_12817);
and U14458 (N_14458,N_12093,N_12002);
nor U14459 (N_14459,N_12053,N_13463);
xnor U14460 (N_14460,N_13769,N_12303);
nor U14461 (N_14461,N_13571,N_12651);
and U14462 (N_14462,N_12047,N_12812);
xnor U14463 (N_14463,N_13360,N_12388);
nor U14464 (N_14464,N_12178,N_12957);
and U14465 (N_14465,N_12045,N_12658);
and U14466 (N_14466,N_13117,N_13173);
nor U14467 (N_14467,N_12026,N_12880);
nand U14468 (N_14468,N_13645,N_12372);
or U14469 (N_14469,N_13986,N_12800);
nand U14470 (N_14470,N_12932,N_13137);
and U14471 (N_14471,N_13919,N_12189);
nor U14472 (N_14472,N_12052,N_12250);
nand U14473 (N_14473,N_13527,N_13288);
xnor U14474 (N_14474,N_13142,N_12615);
nor U14475 (N_14475,N_12345,N_12856);
nor U14476 (N_14476,N_12184,N_13997);
nand U14477 (N_14477,N_12516,N_12775);
nor U14478 (N_14478,N_13475,N_13386);
and U14479 (N_14479,N_13677,N_13264);
xnor U14480 (N_14480,N_12112,N_12427);
nand U14481 (N_14481,N_13296,N_12462);
xnor U14482 (N_14482,N_12505,N_12386);
nor U14483 (N_14483,N_12356,N_12836);
and U14484 (N_14484,N_12377,N_12133);
nand U14485 (N_14485,N_12293,N_13164);
or U14486 (N_14486,N_13496,N_12556);
or U14487 (N_14487,N_13976,N_12067);
xnor U14488 (N_14488,N_13350,N_13077);
nand U14489 (N_14489,N_12410,N_12435);
nand U14490 (N_14490,N_13783,N_12960);
or U14491 (N_14491,N_12066,N_12964);
nand U14492 (N_14492,N_12864,N_13086);
nor U14493 (N_14493,N_12445,N_12426);
nor U14494 (N_14494,N_12256,N_12743);
and U14495 (N_14495,N_13949,N_13453);
and U14496 (N_14496,N_13472,N_12418);
nor U14497 (N_14497,N_13887,N_13678);
nor U14498 (N_14498,N_12194,N_13820);
or U14499 (N_14499,N_13461,N_13560);
nor U14500 (N_14500,N_13910,N_12713);
nand U14501 (N_14501,N_13269,N_12024);
or U14502 (N_14502,N_12360,N_12992);
nand U14503 (N_14503,N_13032,N_12795);
xor U14504 (N_14504,N_12253,N_12742);
and U14505 (N_14505,N_12567,N_13204);
nor U14506 (N_14506,N_12227,N_13406);
nor U14507 (N_14507,N_13150,N_13692);
xor U14508 (N_14508,N_12350,N_13529);
nor U14509 (N_14509,N_12117,N_12060);
xor U14510 (N_14510,N_12643,N_12252);
nor U14511 (N_14511,N_12698,N_12670);
or U14512 (N_14512,N_13324,N_13538);
and U14513 (N_14513,N_12472,N_12103);
nor U14514 (N_14514,N_13729,N_12206);
xor U14515 (N_14515,N_12411,N_12834);
nor U14516 (N_14516,N_12777,N_13080);
nand U14517 (N_14517,N_12841,N_13211);
or U14518 (N_14518,N_12920,N_13832);
nand U14519 (N_14519,N_13328,N_12245);
or U14520 (N_14520,N_12650,N_12640);
and U14521 (N_14521,N_13266,N_12507);
nand U14522 (N_14522,N_13043,N_12150);
nor U14523 (N_14523,N_12923,N_13334);
xor U14524 (N_14524,N_13951,N_12187);
and U14525 (N_14525,N_12701,N_12233);
nor U14526 (N_14526,N_13247,N_13749);
or U14527 (N_14527,N_12011,N_12928);
and U14528 (N_14528,N_12126,N_12292);
nand U14529 (N_14529,N_13563,N_12891);
or U14530 (N_14530,N_13120,N_12474);
nor U14531 (N_14531,N_12709,N_13799);
and U14532 (N_14532,N_12785,N_12797);
nand U14533 (N_14533,N_12302,N_13823);
or U14534 (N_14534,N_13112,N_12437);
and U14535 (N_14535,N_12534,N_13394);
nand U14536 (N_14536,N_12273,N_13766);
nand U14537 (N_14537,N_13241,N_13691);
or U14538 (N_14538,N_12938,N_12790);
and U14539 (N_14539,N_12759,N_12306);
nor U14540 (N_14540,N_12521,N_13342);
nand U14541 (N_14541,N_13051,N_13265);
nor U14542 (N_14542,N_12956,N_13443);
or U14543 (N_14543,N_12685,N_13830);
nor U14544 (N_14544,N_13118,N_13196);
nor U14545 (N_14545,N_12404,N_13413);
nor U14546 (N_14546,N_12308,N_13545);
nand U14547 (N_14547,N_13372,N_12546);
and U14548 (N_14548,N_13216,N_13462);
or U14549 (N_14549,N_12182,N_12581);
and U14550 (N_14550,N_12830,N_13555);
or U14551 (N_14551,N_12686,N_12196);
and U14552 (N_14552,N_12147,N_12311);
or U14553 (N_14553,N_13037,N_12794);
and U14554 (N_14554,N_13487,N_13392);
or U14555 (N_14555,N_13235,N_13507);
nor U14556 (N_14556,N_12770,N_12550);
and U14557 (N_14557,N_12525,N_13551);
and U14558 (N_14558,N_13260,N_12088);
and U14559 (N_14559,N_13308,N_12491);
and U14560 (N_14560,N_13119,N_13223);
or U14561 (N_14561,N_13343,N_13700);
nand U14562 (N_14562,N_12539,N_12412);
and U14563 (N_14563,N_13961,N_13317);
or U14564 (N_14564,N_12489,N_13838);
nand U14565 (N_14565,N_12416,N_13559);
nand U14566 (N_14566,N_12171,N_12562);
or U14567 (N_14567,N_12595,N_13168);
or U14568 (N_14568,N_13205,N_13794);
nor U14569 (N_14569,N_13615,N_12106);
and U14570 (N_14570,N_13409,N_13971);
and U14571 (N_14571,N_13455,N_12127);
nor U14572 (N_14572,N_12294,N_13434);
nor U14573 (N_14573,N_13883,N_13055);
nor U14574 (N_14574,N_13741,N_13133);
nor U14575 (N_14575,N_12050,N_12156);
or U14576 (N_14576,N_13422,N_12933);
and U14577 (N_14577,N_12216,N_13466);
nand U14578 (N_14578,N_12590,N_12079);
or U14579 (N_14579,N_12398,N_12203);
nand U14580 (N_14580,N_12327,N_13139);
and U14581 (N_14581,N_13228,N_12339);
or U14582 (N_14582,N_12733,N_12374);
nand U14583 (N_14583,N_12955,N_13892);
and U14584 (N_14584,N_12683,N_13181);
nand U14585 (N_14585,N_13533,N_13557);
nand U14586 (N_14586,N_13464,N_12215);
nand U14587 (N_14587,N_13714,N_12135);
nand U14588 (N_14588,N_13597,N_12648);
xor U14589 (N_14589,N_13514,N_13718);
or U14590 (N_14590,N_13662,N_12572);
or U14591 (N_14591,N_13489,N_13019);
or U14592 (N_14592,N_12900,N_13646);
or U14593 (N_14593,N_12247,N_12390);
and U14594 (N_14594,N_12924,N_12869);
xor U14595 (N_14595,N_12141,N_13493);
or U14596 (N_14596,N_12129,N_12329);
or U14597 (N_14597,N_13418,N_12628);
nor U14598 (N_14598,N_13403,N_12855);
nor U14599 (N_14599,N_13039,N_12624);
and U14600 (N_14600,N_12401,N_12328);
or U14601 (N_14601,N_12090,N_13400);
nor U14602 (N_14602,N_13175,N_12035);
and U14603 (N_14603,N_12468,N_12089);
or U14604 (N_14604,N_12767,N_13727);
or U14605 (N_14605,N_13702,N_13160);
nand U14606 (N_14606,N_12626,N_13089);
nor U14607 (N_14607,N_12780,N_13939);
nand U14608 (N_14608,N_13491,N_13162);
xor U14609 (N_14609,N_13810,N_12563);
nor U14610 (N_14610,N_13925,N_12513);
nor U14611 (N_14611,N_13261,N_13280);
nand U14612 (N_14612,N_13323,N_12517);
and U14613 (N_14613,N_13854,N_12409);
nand U14614 (N_14614,N_13361,N_13556);
nor U14615 (N_14615,N_12315,N_13958);
or U14616 (N_14616,N_13349,N_12380);
nand U14617 (N_14617,N_13271,N_13607);
or U14618 (N_14618,N_13851,N_12749);
nand U14619 (N_14619,N_13420,N_12833);
or U14620 (N_14620,N_12020,N_13553);
nor U14621 (N_14621,N_13622,N_12274);
nand U14622 (N_14622,N_13358,N_13129);
or U14623 (N_14623,N_12732,N_13333);
nor U14624 (N_14624,N_12782,N_12201);
xnor U14625 (N_14625,N_13613,N_12946);
nor U14626 (N_14626,N_13233,N_12738);
or U14627 (N_14627,N_12892,N_13888);
and U14628 (N_14628,N_12668,N_12803);
nor U14629 (N_14629,N_12684,N_12712);
and U14630 (N_14630,N_13879,N_12639);
nand U14631 (N_14631,N_13987,N_13011);
nand U14632 (N_14632,N_12174,N_13398);
or U14633 (N_14633,N_13589,N_12921);
or U14634 (N_14634,N_13670,N_13352);
and U14635 (N_14635,N_13365,N_12784);
or U14636 (N_14636,N_13028,N_13008);
or U14637 (N_14637,N_13121,N_12408);
nor U14638 (N_14638,N_13852,N_13177);
nor U14639 (N_14639,N_12046,N_13865);
nand U14640 (N_14640,N_13522,N_12564);
nor U14641 (N_14641,N_13286,N_12568);
nand U14642 (N_14642,N_13436,N_12945);
nand U14643 (N_14643,N_13368,N_13639);
or U14644 (N_14644,N_12101,N_12971);
and U14645 (N_14645,N_13456,N_12044);
or U14646 (N_14646,N_12406,N_12192);
xnor U14647 (N_14647,N_13227,N_13889);
nand U14648 (N_14648,N_13083,N_13751);
nand U14649 (N_14649,N_13081,N_13759);
or U14650 (N_14650,N_13483,N_13757);
nand U14651 (N_14651,N_13885,N_13813);
nor U14652 (N_14652,N_12700,N_12321);
xor U14653 (N_14653,N_12863,N_13543);
or U14654 (N_14654,N_13554,N_13918);
and U14655 (N_14655,N_13619,N_13916);
and U14656 (N_14656,N_12081,N_12248);
and U14657 (N_14657,N_13955,N_12965);
nand U14658 (N_14658,N_13006,N_13573);
nor U14659 (N_14659,N_13357,N_13279);
and U14660 (N_14660,N_13188,N_13367);
or U14661 (N_14661,N_13102,N_13728);
xor U14662 (N_14662,N_13424,N_13752);
or U14663 (N_14663,N_13012,N_13534);
nand U14664 (N_14664,N_12175,N_12333);
and U14665 (N_14665,N_12348,N_13084);
or U14666 (N_14666,N_13636,N_13044);
xor U14667 (N_14667,N_12754,N_13459);
and U14668 (N_14668,N_13130,N_13124);
nor U14669 (N_14669,N_12338,N_13369);
or U14670 (N_14670,N_12263,N_13703);
or U14671 (N_14671,N_12297,N_12941);
and U14672 (N_14672,N_12826,N_13526);
nand U14673 (N_14673,N_12260,N_12852);
or U14674 (N_14674,N_12001,N_12415);
or U14675 (N_14675,N_13356,N_12951);
nand U14676 (N_14676,N_12688,N_12566);
and U14677 (N_14677,N_13620,N_13285);
or U14678 (N_14678,N_13414,N_12560);
and U14679 (N_14679,N_12894,N_13419);
or U14680 (N_14680,N_13506,N_12809);
nor U14681 (N_14681,N_12860,N_12258);
and U14682 (N_14682,N_13723,N_13792);
xor U14683 (N_14683,N_12573,N_13079);
xnor U14684 (N_14684,N_12587,N_13050);
nand U14685 (N_14685,N_13200,N_12039);
and U14686 (N_14686,N_12074,N_12322);
or U14687 (N_14687,N_12847,N_12565);
and U14688 (N_14688,N_13816,N_12379);
nor U14689 (N_14689,N_13167,N_13972);
or U14690 (N_14690,N_13558,N_13917);
xnor U14691 (N_14691,N_12357,N_13231);
or U14692 (N_14692,N_13648,N_13625);
xnor U14693 (N_14693,N_12953,N_13862);
and U14694 (N_14694,N_12819,N_13886);
xnor U14695 (N_14695,N_12077,N_13899);
and U14696 (N_14696,N_13606,N_13174);
or U14697 (N_14697,N_12457,N_12642);
xnor U14698 (N_14698,N_12361,N_13962);
nand U14699 (N_14699,N_12223,N_12947);
nand U14700 (N_14700,N_13963,N_13440);
and U14701 (N_14701,N_12750,N_12918);
nor U14702 (N_14702,N_12575,N_13906);
xor U14703 (N_14703,N_13219,N_13936);
nand U14704 (N_14704,N_13642,N_13621);
nand U14705 (N_14705,N_13449,N_12967);
or U14706 (N_14706,N_13726,N_12616);
and U14707 (N_14707,N_13850,N_13991);
nor U14708 (N_14708,N_13473,N_13731);
or U14709 (N_14709,N_12533,N_13500);
and U14710 (N_14710,N_12226,N_13145);
nand U14711 (N_14711,N_12211,N_13191);
nand U14712 (N_14712,N_12056,N_12319);
and U14713 (N_14713,N_12871,N_12799);
nand U14714 (N_14714,N_13915,N_12091);
and U14715 (N_14715,N_13740,N_13014);
nand U14716 (N_14716,N_12963,N_12509);
and U14717 (N_14717,N_13058,N_13417);
nor U14718 (N_14718,N_13234,N_13873);
and U14719 (N_14719,N_12985,N_13679);
nand U14720 (N_14720,N_12004,N_12368);
xor U14721 (N_14721,N_13688,N_12561);
nand U14722 (N_14722,N_13107,N_13215);
xnor U14723 (N_14723,N_13973,N_12815);
nand U14724 (N_14724,N_12221,N_12334);
and U14725 (N_14725,N_13364,N_13787);
nand U14726 (N_14726,N_13775,N_13442);
and U14727 (N_14727,N_13090,N_12105);
nand U14728 (N_14728,N_13831,N_12528);
nor U14729 (N_14729,N_13180,N_13470);
and U14730 (N_14730,N_13346,N_12007);
nand U14731 (N_14731,N_12926,N_13376);
nand U14732 (N_14732,N_12899,N_12119);
and U14733 (N_14733,N_12202,N_13716);
or U14734 (N_14734,N_13969,N_12804);
xnor U14735 (N_14735,N_12622,N_13059);
nand U14736 (N_14736,N_13366,N_13975);
nand U14737 (N_14737,N_13048,N_13934);
nand U14738 (N_14738,N_12190,N_12073);
nand U14739 (N_14739,N_12760,N_13808);
nand U14740 (N_14740,N_12059,N_13476);
or U14741 (N_14741,N_12706,N_12764);
and U14742 (N_14742,N_12776,N_12453);
or U14743 (N_14743,N_12236,N_12602);
or U14744 (N_14744,N_13194,N_12461);
nand U14745 (N_14745,N_13404,N_12362);
nand U14746 (N_14746,N_13428,N_13309);
nor U14747 (N_14747,N_12198,N_12569);
and U14748 (N_14748,N_12430,N_13721);
nand U14749 (N_14749,N_12458,N_13954);
xor U14750 (N_14750,N_13761,N_13159);
and U14751 (N_14751,N_13238,N_13651);
or U14752 (N_14752,N_13835,N_13390);
nor U14753 (N_14753,N_12974,N_12181);
xnor U14754 (N_14754,N_12138,N_12954);
and U14755 (N_14755,N_12879,N_12558);
nand U14756 (N_14756,N_13208,N_13552);
nor U14757 (N_14757,N_13941,N_13667);
nor U14758 (N_14758,N_12543,N_13698);
nor U14759 (N_14759,N_12287,N_12553);
nor U14760 (N_14760,N_12405,N_12966);
nand U14761 (N_14761,N_13999,N_12577);
nor U14762 (N_14762,N_12326,N_12911);
xnor U14763 (N_14763,N_12114,N_13132);
nor U14764 (N_14764,N_12255,N_12022);
and U14765 (N_14765,N_12469,N_12162);
nor U14766 (N_14766,N_13157,N_13480);
and U14767 (N_14767,N_13609,N_13141);
or U14768 (N_14768,N_13634,N_12071);
xor U14769 (N_14769,N_13036,N_12163);
and U14770 (N_14770,N_12862,N_12301);
or U14771 (N_14771,N_13023,N_13668);
xor U14772 (N_14772,N_12479,N_12062);
and U14773 (N_14773,N_12285,N_12080);
and U14774 (N_14774,N_12142,N_13320);
and U14775 (N_14775,N_13895,N_13445);
or U14776 (N_14776,N_13498,N_13274);
or U14777 (N_14777,N_12532,N_13682);
nor U14778 (N_14778,N_12905,N_12251);
nor U14779 (N_14779,N_13460,N_13638);
or U14780 (N_14780,N_13225,N_13447);
nor U14781 (N_14781,N_12209,N_13127);
nor U14782 (N_14782,N_13712,N_13047);
and U14783 (N_14783,N_13100,N_12337);
nor U14784 (N_14784,N_13183,N_12485);
xnor U14785 (N_14785,N_13845,N_13780);
or U14786 (N_14786,N_13675,N_12861);
and U14787 (N_14787,N_12881,N_13243);
and U14788 (N_14788,N_12186,N_12996);
nand U14789 (N_14789,N_13111,N_12346);
nand U14790 (N_14790,N_13207,N_12745);
nor U14791 (N_14791,N_13481,N_13045);
and U14792 (N_14792,N_12029,N_12288);
and U14793 (N_14793,N_13982,N_13239);
nor U14794 (N_14794,N_12831,N_12367);
and U14795 (N_14795,N_13877,N_13510);
or U14796 (N_14796,N_12139,N_13843);
or U14797 (N_14797,N_13630,N_12102);
and U14798 (N_14798,N_13665,N_12257);
nand U14799 (N_14799,N_13076,N_12269);
nor U14800 (N_14800,N_12335,N_12842);
nor U14801 (N_14801,N_12040,N_12108);
xnor U14802 (N_14802,N_13872,N_12848);
nor U14803 (N_14803,N_13592,N_13293);
and U14804 (N_14804,N_12908,N_13148);
nand U14805 (N_14805,N_13072,N_13900);
nor U14806 (N_14806,N_13389,N_13479);
nand U14807 (N_14807,N_13839,N_13311);
nand U14808 (N_14808,N_13765,N_13341);
nand U14809 (N_14809,N_13468,N_12644);
nor U14810 (N_14810,N_12403,N_12421);
nand U14811 (N_14811,N_13096,N_13020);
or U14812 (N_14812,N_13742,N_12526);
and U14813 (N_14813,N_12282,N_12032);
xor U14814 (N_14814,N_12719,N_12234);
or U14815 (N_14815,N_13199,N_13353);
nand U14816 (N_14816,N_12176,N_12728);
nand U14817 (N_14817,N_13198,N_13103);
nand U14818 (N_14818,N_13985,N_13572);
or U14819 (N_14819,N_12371,N_12343);
nor U14820 (N_14820,N_12023,N_12884);
and U14821 (N_14821,N_12446,N_13869);
nor U14822 (N_14822,N_12744,N_13565);
or U14823 (N_14823,N_13114,N_13345);
or U14824 (N_14824,N_12165,N_13024);
or U14825 (N_14825,N_12441,N_13000);
or U14826 (N_14826,N_13640,N_13907);
xnor U14827 (N_14827,N_13163,N_12376);
nand U14828 (N_14828,N_13676,N_13041);
or U14829 (N_14829,N_12191,N_13179);
nor U14830 (N_14830,N_13550,N_12490);
and U14831 (N_14831,N_12608,N_12944);
nor U14832 (N_14832,N_13763,N_12214);
xnor U14833 (N_14833,N_13193,N_13770);
and U14834 (N_14834,N_13998,N_12724);
nand U14835 (N_14835,N_12849,N_13598);
xor U14836 (N_14836,N_13513,N_12249);
or U14837 (N_14837,N_13245,N_13950);
nor U14838 (N_14838,N_13374,N_12132);
and U14839 (N_14839,N_13771,N_13291);
and U14840 (N_14840,N_12354,N_13624);
nor U14841 (N_14841,N_12038,N_13230);
and U14842 (N_14842,N_13446,N_12094);
or U14843 (N_14843,N_13065,N_12078);
xor U14844 (N_14844,N_13505,N_13743);
nand U14845 (N_14845,N_12019,N_12578);
and U14846 (N_14846,N_13075,N_13069);
nand U14847 (N_14847,N_12235,N_12242);
or U14848 (N_14848,N_13378,N_12995);
nand U14849 (N_14849,N_13828,N_12726);
xor U14850 (N_14850,N_12895,N_13337);
nand U14851 (N_14851,N_12125,N_13652);
or U14852 (N_14852,N_12484,N_12120);
xnor U14853 (N_14853,N_13791,N_13868);
xnor U14854 (N_14854,N_13884,N_12766);
xnor U14855 (N_14855,N_12820,N_13953);
nor U14856 (N_14856,N_13013,N_12948);
or U14857 (N_14857,N_12737,N_12271);
nor U14858 (N_14858,N_13612,N_13384);
xor U14859 (N_14859,N_13104,N_12220);
and U14860 (N_14860,N_12889,N_12886);
nor U14861 (N_14861,N_13457,N_13109);
or U14862 (N_14862,N_13779,N_12152);
and U14863 (N_14863,N_12332,N_13809);
nor U14864 (N_14864,N_12605,N_13030);
xnor U14865 (N_14865,N_13796,N_12659);
and U14866 (N_14866,N_12919,N_12012);
and U14867 (N_14867,N_13849,N_12487);
or U14868 (N_14868,N_13347,N_13277);
xor U14869 (N_14869,N_13284,N_12342);
xnor U14870 (N_14870,N_12772,N_12096);
or U14871 (N_14871,N_13583,N_13536);
nand U14872 (N_14872,N_13860,N_13983);
nand U14873 (N_14873,N_13940,N_12478);
and U14874 (N_14874,N_13926,N_13946);
xnor U14875 (N_14875,N_13151,N_12438);
nand U14876 (N_14876,N_12703,N_13921);
nand U14877 (N_14877,N_12399,N_13144);
and U14878 (N_14878,N_12704,N_12730);
nor U14879 (N_14879,N_12069,N_13893);
nor U14880 (N_14880,N_12674,N_13561);
nand U14881 (N_14881,N_13061,N_13738);
or U14882 (N_14882,N_12538,N_12034);
nor U14883 (N_14883,N_13818,N_13297);
or U14884 (N_14884,N_12846,N_13448);
or U14885 (N_14885,N_12455,N_12968);
nand U14886 (N_14886,N_13581,N_13430);
and U14887 (N_14887,N_13658,N_13197);
or U14888 (N_14888,N_13541,N_13784);
or U14889 (N_14889,N_13696,N_12959);
nor U14890 (N_14890,N_13056,N_12498);
and U14891 (N_14891,N_13633,N_13057);
or U14892 (N_14892,N_12857,N_13628);
or U14893 (N_14893,N_12755,N_13861);
or U14894 (N_14894,N_12916,N_12436);
nor U14895 (N_14895,N_12893,N_13465);
or U14896 (N_14896,N_12544,N_12636);
and U14897 (N_14897,N_12527,N_12903);
and U14898 (N_14898,N_12070,N_12246);
and U14899 (N_14899,N_13283,N_12798);
and U14900 (N_14900,N_13251,N_13755);
nand U14901 (N_14901,N_12691,N_13236);
nand U14902 (N_14902,N_13923,N_12729);
and U14903 (N_14903,N_12254,N_12151);
nor U14904 (N_14904,N_12758,N_13566);
and U14905 (N_14905,N_12177,N_13547);
xnor U14906 (N_14906,N_12657,N_13746);
nand U14907 (N_14907,N_13009,N_12115);
and U14908 (N_14908,N_13344,N_12395);
nor U14909 (N_14909,N_13517,N_12555);
and U14910 (N_14910,N_13515,N_12696);
nor U14911 (N_14911,N_13509,N_12483);
and U14912 (N_14912,N_12682,N_13582);
nand U14913 (N_14913,N_12502,N_12167);
nor U14914 (N_14914,N_13660,N_13143);
nand U14915 (N_14915,N_13325,N_12123);
and U14916 (N_14916,N_13595,N_12808);
xor U14917 (N_14917,N_13126,N_12612);
nor U14918 (N_14918,N_13684,N_13229);
nor U14919 (N_14919,N_13010,N_13578);
xor U14920 (N_14920,N_12085,N_12008);
and U14921 (N_14921,N_13202,N_12876);
xor U14922 (N_14922,N_13655,N_13253);
nor U14923 (N_14923,N_12312,N_13387);
and U14924 (N_14924,N_12473,N_13789);
nand U14925 (N_14925,N_12392,N_12589);
or U14926 (N_14926,N_13644,N_13206);
nor U14927 (N_14927,N_13136,N_12822);
nor U14928 (N_14928,N_12272,N_12687);
or U14929 (N_14929,N_12942,N_13909);
nor U14930 (N_14930,N_13242,N_13169);
and U14931 (N_14931,N_12283,N_13825);
and U14932 (N_14932,N_12549,N_13901);
nor U14933 (N_14933,N_12397,N_13694);
or U14934 (N_14934,N_12715,N_13546);
or U14935 (N_14935,N_13450,N_13478);
or U14936 (N_14936,N_12087,N_12769);
nor U14937 (N_14937,N_13602,N_12858);
or U14938 (N_14938,N_12396,N_13003);
nand U14939 (N_14939,N_13920,N_13876);
and U14940 (N_14940,N_12991,N_13042);
nand U14941 (N_14941,N_12897,N_13690);
and U14942 (N_14942,N_12276,N_12805);
nor U14943 (N_14943,N_13382,N_13299);
nor U14944 (N_14944,N_12711,N_12494);
nand U14945 (N_14945,N_13184,N_12977);
nand U14946 (N_14946,N_13052,N_13540);
nor U14947 (N_14947,N_12036,N_12603);
or U14948 (N_14948,N_13209,N_12907);
and U14949 (N_14949,N_12816,N_12781);
nor U14950 (N_14950,N_13590,N_13807);
nand U14951 (N_14951,N_13701,N_12161);
and U14952 (N_14952,N_12015,N_13092);
and U14953 (N_14953,N_13913,N_12917);
xnor U14954 (N_14954,N_12583,N_12925);
nor U14955 (N_14955,N_13485,N_12183);
or U14956 (N_14956,N_12364,N_12695);
and U14957 (N_14957,N_12873,N_12460);
nor U14958 (N_14958,N_13395,N_13672);
and U14959 (N_14959,N_12551,N_13040);
nand U14960 (N_14960,N_12721,N_12197);
nand U14961 (N_14961,N_13894,N_12828);
nor U14962 (N_14962,N_12718,N_12912);
and U14963 (N_14963,N_12584,N_13467);
or U14964 (N_14964,N_12224,N_13819);
xor U14965 (N_14965,N_13315,N_13988);
xor U14966 (N_14966,N_12237,N_13259);
nor U14967 (N_14967,N_13637,N_12949);
nand U14968 (N_14968,N_13282,N_13165);
nand U14969 (N_14969,N_12813,N_13411);
xnor U14970 (N_14970,N_13125,N_12637);
nor U14971 (N_14971,N_13964,N_12353);
and U14972 (N_14972,N_12481,N_13391);
and U14973 (N_14973,N_12716,N_12307);
and U14974 (N_14974,N_12910,N_12829);
and U14975 (N_14975,N_12909,N_12075);
nand U14976 (N_14976,N_13733,N_12692);
and U14977 (N_14977,N_13528,N_12281);
xnor U14978 (N_14978,N_13106,N_12279);
nand U14979 (N_14979,N_12309,N_12100);
and U14980 (N_14980,N_13593,N_13977);
nand U14981 (N_14981,N_13931,N_12449);
nand U14982 (N_14982,N_12914,N_12014);
or U14983 (N_14983,N_13758,N_12757);
or U14984 (N_14984,N_12055,N_12671);
nor U14985 (N_14985,N_13632,N_13902);
or U14986 (N_14986,N_13313,N_13093);
and U14987 (N_14987,N_13981,N_13812);
nor U14988 (N_14988,N_13407,N_12025);
or U14989 (N_14989,N_13772,N_12470);
nand U14990 (N_14990,N_12574,N_13362);
nor U14991 (N_14991,N_12638,N_12796);
nand U14992 (N_14992,N_12983,N_13192);
nor U14993 (N_14993,N_13435,N_12753);
or U14994 (N_14994,N_12694,N_13863);
and U14995 (N_14995,N_12407,N_12387);
nor U14996 (N_14996,N_13836,N_13246);
or U14997 (N_14997,N_12092,N_13154);
nand U14998 (N_14998,N_12853,N_12143);
or U14999 (N_14999,N_12239,N_12727);
or U15000 (N_15000,N_13643,N_12288);
nand U15001 (N_15001,N_12722,N_13483);
or U15002 (N_15002,N_12117,N_13370);
nand U15003 (N_15003,N_13753,N_12813);
nor U15004 (N_15004,N_13656,N_12502);
xor U15005 (N_15005,N_12770,N_12888);
nor U15006 (N_15006,N_13646,N_12324);
and U15007 (N_15007,N_12803,N_13207);
xnor U15008 (N_15008,N_13100,N_13227);
nor U15009 (N_15009,N_13914,N_12000);
nand U15010 (N_15010,N_12468,N_12875);
xnor U15011 (N_15011,N_13820,N_12673);
nor U15012 (N_15012,N_13847,N_13019);
or U15013 (N_15013,N_12496,N_13316);
nor U15014 (N_15014,N_12510,N_12643);
nor U15015 (N_15015,N_12344,N_13881);
nand U15016 (N_15016,N_13880,N_13297);
and U15017 (N_15017,N_13912,N_13293);
or U15018 (N_15018,N_13735,N_13098);
or U15019 (N_15019,N_13254,N_12293);
or U15020 (N_15020,N_13884,N_12412);
or U15021 (N_15021,N_13719,N_13422);
nor U15022 (N_15022,N_13192,N_12083);
and U15023 (N_15023,N_12311,N_13270);
and U15024 (N_15024,N_13148,N_12758);
and U15025 (N_15025,N_12176,N_12402);
nand U15026 (N_15026,N_12028,N_13218);
nor U15027 (N_15027,N_12116,N_12090);
xor U15028 (N_15028,N_12892,N_12204);
xnor U15029 (N_15029,N_12697,N_12156);
and U15030 (N_15030,N_12828,N_12623);
nand U15031 (N_15031,N_13066,N_13587);
nor U15032 (N_15032,N_12481,N_13030);
xnor U15033 (N_15033,N_13231,N_13391);
nand U15034 (N_15034,N_12348,N_13753);
xnor U15035 (N_15035,N_13398,N_13209);
nand U15036 (N_15036,N_12149,N_13799);
xnor U15037 (N_15037,N_13644,N_13800);
nor U15038 (N_15038,N_13783,N_13257);
nor U15039 (N_15039,N_13164,N_12794);
nand U15040 (N_15040,N_12991,N_12003);
xor U15041 (N_15041,N_12757,N_13855);
nor U15042 (N_15042,N_12641,N_12695);
or U15043 (N_15043,N_12970,N_12718);
nand U15044 (N_15044,N_13895,N_12049);
and U15045 (N_15045,N_13061,N_13550);
nand U15046 (N_15046,N_13182,N_12048);
and U15047 (N_15047,N_13193,N_13074);
nor U15048 (N_15048,N_12870,N_13438);
and U15049 (N_15049,N_13580,N_12850);
xnor U15050 (N_15050,N_12668,N_12817);
nand U15051 (N_15051,N_12208,N_13365);
or U15052 (N_15052,N_13235,N_12644);
xnor U15053 (N_15053,N_12345,N_13070);
or U15054 (N_15054,N_12951,N_12940);
and U15055 (N_15055,N_13847,N_12081);
nand U15056 (N_15056,N_12168,N_13321);
nor U15057 (N_15057,N_12218,N_13156);
or U15058 (N_15058,N_13398,N_12534);
nor U15059 (N_15059,N_12720,N_13816);
and U15060 (N_15060,N_12933,N_13125);
or U15061 (N_15061,N_13035,N_13693);
or U15062 (N_15062,N_12842,N_12587);
nor U15063 (N_15063,N_13997,N_12125);
nand U15064 (N_15064,N_13568,N_12900);
or U15065 (N_15065,N_12202,N_13201);
xnor U15066 (N_15066,N_12061,N_13005);
or U15067 (N_15067,N_13993,N_13940);
nand U15068 (N_15068,N_12184,N_13430);
and U15069 (N_15069,N_13637,N_12021);
xnor U15070 (N_15070,N_12397,N_12267);
nor U15071 (N_15071,N_12603,N_13264);
or U15072 (N_15072,N_12339,N_13885);
or U15073 (N_15073,N_12230,N_12760);
or U15074 (N_15074,N_13993,N_12484);
nor U15075 (N_15075,N_12184,N_12939);
or U15076 (N_15076,N_13972,N_13409);
or U15077 (N_15077,N_13240,N_12562);
nand U15078 (N_15078,N_12532,N_13926);
nor U15079 (N_15079,N_12834,N_13463);
xnor U15080 (N_15080,N_12564,N_13328);
nand U15081 (N_15081,N_13141,N_13915);
and U15082 (N_15082,N_13942,N_12221);
or U15083 (N_15083,N_12294,N_13437);
and U15084 (N_15084,N_13779,N_13328);
and U15085 (N_15085,N_12322,N_13684);
nand U15086 (N_15086,N_12265,N_12325);
and U15087 (N_15087,N_13241,N_13962);
and U15088 (N_15088,N_12259,N_13668);
or U15089 (N_15089,N_12154,N_12210);
or U15090 (N_15090,N_13429,N_13721);
xor U15091 (N_15091,N_13048,N_12428);
or U15092 (N_15092,N_13855,N_12079);
nand U15093 (N_15093,N_12201,N_13499);
and U15094 (N_15094,N_12343,N_12162);
nor U15095 (N_15095,N_13016,N_12393);
nand U15096 (N_15096,N_13385,N_12208);
or U15097 (N_15097,N_13669,N_12388);
nand U15098 (N_15098,N_12798,N_13756);
or U15099 (N_15099,N_13378,N_13775);
and U15100 (N_15100,N_12138,N_13225);
nor U15101 (N_15101,N_12383,N_13289);
xnor U15102 (N_15102,N_13260,N_12857);
nor U15103 (N_15103,N_12727,N_13814);
or U15104 (N_15104,N_12118,N_13514);
or U15105 (N_15105,N_13779,N_13652);
or U15106 (N_15106,N_12916,N_13802);
or U15107 (N_15107,N_12273,N_13423);
and U15108 (N_15108,N_13441,N_12625);
and U15109 (N_15109,N_12514,N_13427);
or U15110 (N_15110,N_13081,N_13337);
nand U15111 (N_15111,N_12048,N_13843);
nand U15112 (N_15112,N_12084,N_12790);
and U15113 (N_15113,N_13941,N_12459);
nand U15114 (N_15114,N_12528,N_12279);
or U15115 (N_15115,N_12974,N_13476);
and U15116 (N_15116,N_12314,N_12746);
nand U15117 (N_15117,N_12918,N_13909);
nand U15118 (N_15118,N_13118,N_13582);
nor U15119 (N_15119,N_12277,N_12876);
nand U15120 (N_15120,N_12314,N_13493);
or U15121 (N_15121,N_13734,N_13549);
or U15122 (N_15122,N_13263,N_13085);
or U15123 (N_15123,N_13297,N_13066);
xnor U15124 (N_15124,N_12407,N_12422);
and U15125 (N_15125,N_13648,N_12572);
xnor U15126 (N_15126,N_12308,N_13722);
and U15127 (N_15127,N_12061,N_12945);
and U15128 (N_15128,N_13871,N_12155);
nor U15129 (N_15129,N_12006,N_12823);
or U15130 (N_15130,N_13213,N_12286);
nor U15131 (N_15131,N_12984,N_13774);
and U15132 (N_15132,N_12785,N_12793);
nand U15133 (N_15133,N_13452,N_12809);
nand U15134 (N_15134,N_13197,N_12365);
nand U15135 (N_15135,N_12956,N_12512);
nor U15136 (N_15136,N_12877,N_13936);
nor U15137 (N_15137,N_12823,N_13352);
nor U15138 (N_15138,N_13526,N_13522);
and U15139 (N_15139,N_12519,N_12637);
nand U15140 (N_15140,N_13062,N_12919);
and U15141 (N_15141,N_13110,N_12638);
and U15142 (N_15142,N_12779,N_12157);
nand U15143 (N_15143,N_12302,N_12410);
or U15144 (N_15144,N_12508,N_13625);
and U15145 (N_15145,N_13128,N_12140);
xnor U15146 (N_15146,N_13241,N_12151);
xnor U15147 (N_15147,N_13984,N_12990);
and U15148 (N_15148,N_12621,N_12567);
nand U15149 (N_15149,N_13026,N_13316);
nand U15150 (N_15150,N_12130,N_13010);
or U15151 (N_15151,N_13032,N_13465);
nor U15152 (N_15152,N_12451,N_12524);
xor U15153 (N_15153,N_13367,N_12164);
xor U15154 (N_15154,N_13490,N_12677);
and U15155 (N_15155,N_13227,N_13689);
nand U15156 (N_15156,N_13613,N_13566);
xor U15157 (N_15157,N_13112,N_13246);
nand U15158 (N_15158,N_13913,N_12788);
or U15159 (N_15159,N_12493,N_12625);
or U15160 (N_15160,N_13661,N_13333);
nor U15161 (N_15161,N_13432,N_12574);
nor U15162 (N_15162,N_13026,N_13113);
nand U15163 (N_15163,N_12692,N_13510);
nor U15164 (N_15164,N_12238,N_12254);
xor U15165 (N_15165,N_13872,N_13130);
nand U15166 (N_15166,N_12346,N_12662);
and U15167 (N_15167,N_13908,N_12110);
or U15168 (N_15168,N_12735,N_12042);
and U15169 (N_15169,N_13686,N_13927);
nand U15170 (N_15170,N_13629,N_12287);
and U15171 (N_15171,N_12826,N_12895);
nor U15172 (N_15172,N_12344,N_12291);
and U15173 (N_15173,N_12118,N_12930);
nor U15174 (N_15174,N_13177,N_12959);
xor U15175 (N_15175,N_12501,N_12366);
nor U15176 (N_15176,N_13923,N_12916);
nand U15177 (N_15177,N_13334,N_12539);
nor U15178 (N_15178,N_12574,N_13291);
nand U15179 (N_15179,N_13538,N_12451);
and U15180 (N_15180,N_12021,N_13545);
or U15181 (N_15181,N_13553,N_12874);
xor U15182 (N_15182,N_13025,N_13804);
nor U15183 (N_15183,N_12579,N_13284);
and U15184 (N_15184,N_12341,N_12526);
nand U15185 (N_15185,N_13951,N_12400);
nand U15186 (N_15186,N_12859,N_12906);
nor U15187 (N_15187,N_12164,N_13946);
nand U15188 (N_15188,N_13965,N_13663);
or U15189 (N_15189,N_12513,N_13763);
and U15190 (N_15190,N_12627,N_13317);
nor U15191 (N_15191,N_12790,N_13985);
or U15192 (N_15192,N_12871,N_12465);
nand U15193 (N_15193,N_12821,N_13141);
xor U15194 (N_15194,N_12216,N_13236);
or U15195 (N_15195,N_13584,N_13855);
or U15196 (N_15196,N_13236,N_12774);
or U15197 (N_15197,N_13650,N_13670);
xnor U15198 (N_15198,N_12648,N_12300);
and U15199 (N_15199,N_13405,N_13775);
and U15200 (N_15200,N_12746,N_13844);
or U15201 (N_15201,N_12329,N_12228);
or U15202 (N_15202,N_13078,N_12805);
and U15203 (N_15203,N_12340,N_12628);
nor U15204 (N_15204,N_13967,N_13532);
and U15205 (N_15205,N_13542,N_12886);
or U15206 (N_15206,N_13753,N_13508);
or U15207 (N_15207,N_12293,N_13475);
nor U15208 (N_15208,N_13929,N_13684);
or U15209 (N_15209,N_12731,N_13891);
nor U15210 (N_15210,N_12940,N_13575);
nand U15211 (N_15211,N_12368,N_12561);
or U15212 (N_15212,N_12085,N_12132);
and U15213 (N_15213,N_12059,N_13293);
or U15214 (N_15214,N_13282,N_13767);
and U15215 (N_15215,N_13324,N_12357);
nor U15216 (N_15216,N_13888,N_12569);
nand U15217 (N_15217,N_12858,N_12979);
or U15218 (N_15218,N_12208,N_13063);
or U15219 (N_15219,N_13765,N_12790);
and U15220 (N_15220,N_13876,N_13174);
nand U15221 (N_15221,N_13441,N_13264);
or U15222 (N_15222,N_12919,N_13002);
or U15223 (N_15223,N_13294,N_12702);
or U15224 (N_15224,N_12913,N_12879);
nand U15225 (N_15225,N_13033,N_13717);
or U15226 (N_15226,N_12928,N_13577);
nor U15227 (N_15227,N_13997,N_12506);
xor U15228 (N_15228,N_12435,N_12209);
nor U15229 (N_15229,N_13000,N_13182);
and U15230 (N_15230,N_13212,N_12683);
and U15231 (N_15231,N_12631,N_13891);
or U15232 (N_15232,N_12270,N_12854);
nor U15233 (N_15233,N_13076,N_13213);
xnor U15234 (N_15234,N_12972,N_13288);
nor U15235 (N_15235,N_13235,N_12116);
nor U15236 (N_15236,N_13638,N_12157);
or U15237 (N_15237,N_12162,N_13292);
nor U15238 (N_15238,N_13027,N_12160);
and U15239 (N_15239,N_13242,N_12323);
nand U15240 (N_15240,N_12585,N_13261);
and U15241 (N_15241,N_13871,N_12279);
nor U15242 (N_15242,N_12714,N_12576);
nor U15243 (N_15243,N_12930,N_13142);
nand U15244 (N_15244,N_12813,N_12386);
and U15245 (N_15245,N_12465,N_13228);
and U15246 (N_15246,N_12707,N_12941);
or U15247 (N_15247,N_12837,N_12513);
nand U15248 (N_15248,N_12809,N_13848);
nand U15249 (N_15249,N_13085,N_12961);
or U15250 (N_15250,N_12378,N_12857);
xor U15251 (N_15251,N_13069,N_13648);
and U15252 (N_15252,N_13819,N_13440);
and U15253 (N_15253,N_13499,N_12416);
nand U15254 (N_15254,N_13665,N_13049);
nand U15255 (N_15255,N_13262,N_12888);
nor U15256 (N_15256,N_12757,N_12006);
nand U15257 (N_15257,N_12065,N_12907);
or U15258 (N_15258,N_12083,N_12891);
nand U15259 (N_15259,N_12665,N_12424);
nand U15260 (N_15260,N_12410,N_12063);
nand U15261 (N_15261,N_13813,N_12330);
xnor U15262 (N_15262,N_13921,N_13714);
nor U15263 (N_15263,N_13368,N_13166);
nor U15264 (N_15264,N_13625,N_13622);
or U15265 (N_15265,N_12623,N_13985);
and U15266 (N_15266,N_12441,N_12936);
and U15267 (N_15267,N_12971,N_12064);
and U15268 (N_15268,N_13402,N_12932);
and U15269 (N_15269,N_13774,N_13640);
or U15270 (N_15270,N_13300,N_13931);
and U15271 (N_15271,N_12031,N_12048);
nor U15272 (N_15272,N_13573,N_13804);
nor U15273 (N_15273,N_13982,N_13772);
nand U15274 (N_15274,N_12365,N_12447);
or U15275 (N_15275,N_13558,N_13364);
nand U15276 (N_15276,N_12210,N_13555);
and U15277 (N_15277,N_12993,N_12585);
nand U15278 (N_15278,N_13582,N_12996);
xnor U15279 (N_15279,N_13755,N_13744);
and U15280 (N_15280,N_13330,N_13154);
and U15281 (N_15281,N_12087,N_12675);
and U15282 (N_15282,N_13330,N_13980);
nand U15283 (N_15283,N_12675,N_13257);
nand U15284 (N_15284,N_13433,N_12177);
nor U15285 (N_15285,N_13528,N_13720);
nand U15286 (N_15286,N_12761,N_13728);
nand U15287 (N_15287,N_12734,N_13977);
nor U15288 (N_15288,N_13937,N_13192);
or U15289 (N_15289,N_12053,N_13566);
or U15290 (N_15290,N_12893,N_12383);
nor U15291 (N_15291,N_13952,N_12208);
and U15292 (N_15292,N_12793,N_13633);
nor U15293 (N_15293,N_13653,N_13835);
or U15294 (N_15294,N_13485,N_12731);
nand U15295 (N_15295,N_12007,N_13718);
and U15296 (N_15296,N_13432,N_12077);
or U15297 (N_15297,N_13977,N_12496);
and U15298 (N_15298,N_12403,N_12112);
xor U15299 (N_15299,N_13464,N_13999);
or U15300 (N_15300,N_13548,N_13008);
and U15301 (N_15301,N_12129,N_12701);
nand U15302 (N_15302,N_13139,N_13806);
or U15303 (N_15303,N_12686,N_12727);
nor U15304 (N_15304,N_13483,N_13175);
xnor U15305 (N_15305,N_12836,N_13702);
or U15306 (N_15306,N_12757,N_12145);
and U15307 (N_15307,N_12023,N_13597);
or U15308 (N_15308,N_12521,N_13376);
nor U15309 (N_15309,N_13550,N_12346);
or U15310 (N_15310,N_13652,N_13846);
and U15311 (N_15311,N_13428,N_12880);
nor U15312 (N_15312,N_12586,N_12086);
or U15313 (N_15313,N_13102,N_12140);
and U15314 (N_15314,N_13608,N_13495);
xor U15315 (N_15315,N_12402,N_12123);
nor U15316 (N_15316,N_12413,N_13221);
nand U15317 (N_15317,N_12267,N_13341);
or U15318 (N_15318,N_12942,N_12750);
nor U15319 (N_15319,N_13223,N_13728);
xor U15320 (N_15320,N_13652,N_12984);
xor U15321 (N_15321,N_12254,N_13285);
or U15322 (N_15322,N_12618,N_12702);
nand U15323 (N_15323,N_13751,N_13998);
nand U15324 (N_15324,N_12281,N_13517);
nor U15325 (N_15325,N_12489,N_13899);
or U15326 (N_15326,N_12626,N_12267);
nand U15327 (N_15327,N_13304,N_13721);
and U15328 (N_15328,N_12613,N_12146);
nor U15329 (N_15329,N_12787,N_13339);
nand U15330 (N_15330,N_13502,N_13725);
and U15331 (N_15331,N_12849,N_12963);
and U15332 (N_15332,N_13836,N_12338);
or U15333 (N_15333,N_12602,N_12502);
nor U15334 (N_15334,N_12668,N_12694);
nand U15335 (N_15335,N_13594,N_13068);
or U15336 (N_15336,N_13118,N_12906);
nand U15337 (N_15337,N_13996,N_13852);
or U15338 (N_15338,N_13210,N_13301);
nor U15339 (N_15339,N_13304,N_13014);
and U15340 (N_15340,N_12189,N_12348);
nor U15341 (N_15341,N_13067,N_12236);
nor U15342 (N_15342,N_12909,N_13876);
xnor U15343 (N_15343,N_13283,N_12822);
or U15344 (N_15344,N_13797,N_13153);
and U15345 (N_15345,N_12688,N_13298);
nor U15346 (N_15346,N_13583,N_12419);
nand U15347 (N_15347,N_13614,N_13749);
xor U15348 (N_15348,N_13964,N_13467);
or U15349 (N_15349,N_13891,N_12603);
nand U15350 (N_15350,N_13645,N_12710);
or U15351 (N_15351,N_12117,N_12701);
or U15352 (N_15352,N_13988,N_13507);
or U15353 (N_15353,N_13429,N_12278);
nand U15354 (N_15354,N_13274,N_13471);
xor U15355 (N_15355,N_12370,N_12759);
or U15356 (N_15356,N_13079,N_12116);
or U15357 (N_15357,N_13818,N_12710);
nor U15358 (N_15358,N_13499,N_13881);
and U15359 (N_15359,N_12203,N_12050);
nand U15360 (N_15360,N_13670,N_12998);
and U15361 (N_15361,N_13475,N_12504);
and U15362 (N_15362,N_12692,N_12738);
nand U15363 (N_15363,N_12687,N_13480);
xor U15364 (N_15364,N_12780,N_13773);
xnor U15365 (N_15365,N_13492,N_12080);
or U15366 (N_15366,N_13229,N_12524);
and U15367 (N_15367,N_12615,N_13997);
and U15368 (N_15368,N_12636,N_12111);
or U15369 (N_15369,N_12636,N_12409);
xor U15370 (N_15370,N_13300,N_13962);
nor U15371 (N_15371,N_13285,N_12844);
nand U15372 (N_15372,N_13597,N_12323);
and U15373 (N_15373,N_13476,N_12277);
or U15374 (N_15374,N_13790,N_12254);
or U15375 (N_15375,N_12932,N_12917);
or U15376 (N_15376,N_13442,N_13221);
and U15377 (N_15377,N_12887,N_13687);
and U15378 (N_15378,N_13634,N_13047);
nor U15379 (N_15379,N_13357,N_12455);
nand U15380 (N_15380,N_13683,N_13392);
and U15381 (N_15381,N_12912,N_12411);
xor U15382 (N_15382,N_12939,N_13293);
nor U15383 (N_15383,N_12260,N_13168);
nand U15384 (N_15384,N_12702,N_13857);
nor U15385 (N_15385,N_12471,N_13448);
or U15386 (N_15386,N_13036,N_12022);
nor U15387 (N_15387,N_13928,N_13566);
nand U15388 (N_15388,N_13240,N_13753);
nand U15389 (N_15389,N_12120,N_13260);
and U15390 (N_15390,N_12673,N_13293);
and U15391 (N_15391,N_12640,N_13325);
or U15392 (N_15392,N_12391,N_13788);
and U15393 (N_15393,N_13555,N_13453);
xor U15394 (N_15394,N_13381,N_13032);
nand U15395 (N_15395,N_13243,N_13532);
nor U15396 (N_15396,N_13708,N_13229);
and U15397 (N_15397,N_12696,N_12924);
nand U15398 (N_15398,N_12091,N_13626);
or U15399 (N_15399,N_13180,N_13615);
and U15400 (N_15400,N_12510,N_12047);
or U15401 (N_15401,N_13638,N_13477);
and U15402 (N_15402,N_12940,N_13622);
nor U15403 (N_15403,N_12008,N_12862);
nand U15404 (N_15404,N_12733,N_12890);
nand U15405 (N_15405,N_12740,N_13730);
nand U15406 (N_15406,N_13549,N_12023);
nand U15407 (N_15407,N_12594,N_12725);
nand U15408 (N_15408,N_12515,N_13117);
and U15409 (N_15409,N_12347,N_13063);
xor U15410 (N_15410,N_12403,N_12925);
or U15411 (N_15411,N_13700,N_13173);
xnor U15412 (N_15412,N_13598,N_12364);
nand U15413 (N_15413,N_13814,N_12780);
nor U15414 (N_15414,N_13663,N_13647);
and U15415 (N_15415,N_13315,N_13244);
nor U15416 (N_15416,N_13266,N_13523);
or U15417 (N_15417,N_13747,N_12825);
nand U15418 (N_15418,N_12679,N_13970);
nand U15419 (N_15419,N_12907,N_12897);
and U15420 (N_15420,N_12424,N_13451);
or U15421 (N_15421,N_13009,N_12957);
and U15422 (N_15422,N_12417,N_12066);
nor U15423 (N_15423,N_12795,N_12877);
nand U15424 (N_15424,N_12043,N_13331);
or U15425 (N_15425,N_12647,N_12257);
nand U15426 (N_15426,N_12177,N_13819);
nand U15427 (N_15427,N_12397,N_13722);
or U15428 (N_15428,N_12904,N_13955);
nor U15429 (N_15429,N_13591,N_13063);
and U15430 (N_15430,N_13648,N_13277);
nand U15431 (N_15431,N_13890,N_12848);
xnor U15432 (N_15432,N_12380,N_12059);
nor U15433 (N_15433,N_13770,N_12744);
and U15434 (N_15434,N_12897,N_12576);
or U15435 (N_15435,N_13783,N_12353);
or U15436 (N_15436,N_12080,N_12241);
nand U15437 (N_15437,N_12634,N_12437);
nor U15438 (N_15438,N_12559,N_12274);
or U15439 (N_15439,N_12073,N_12726);
xnor U15440 (N_15440,N_12442,N_12784);
nand U15441 (N_15441,N_12865,N_12574);
or U15442 (N_15442,N_12845,N_13506);
nand U15443 (N_15443,N_13366,N_13837);
nand U15444 (N_15444,N_12929,N_12421);
and U15445 (N_15445,N_13552,N_13024);
or U15446 (N_15446,N_13388,N_13321);
or U15447 (N_15447,N_13993,N_12228);
nor U15448 (N_15448,N_13770,N_12091);
and U15449 (N_15449,N_12390,N_13756);
nand U15450 (N_15450,N_13472,N_13587);
or U15451 (N_15451,N_13487,N_12571);
nor U15452 (N_15452,N_13820,N_12615);
nand U15453 (N_15453,N_12265,N_13996);
xnor U15454 (N_15454,N_12948,N_12139);
or U15455 (N_15455,N_12593,N_13178);
or U15456 (N_15456,N_13883,N_13446);
and U15457 (N_15457,N_13962,N_12573);
nor U15458 (N_15458,N_12843,N_13637);
and U15459 (N_15459,N_13216,N_12909);
and U15460 (N_15460,N_13482,N_13703);
nand U15461 (N_15461,N_13058,N_13373);
nand U15462 (N_15462,N_13350,N_13345);
and U15463 (N_15463,N_12257,N_12835);
xnor U15464 (N_15464,N_13489,N_12024);
or U15465 (N_15465,N_12908,N_13666);
nand U15466 (N_15466,N_13688,N_13012);
or U15467 (N_15467,N_12969,N_12871);
nor U15468 (N_15468,N_12573,N_13825);
nand U15469 (N_15469,N_13371,N_12242);
or U15470 (N_15470,N_12804,N_13919);
nor U15471 (N_15471,N_13980,N_12158);
and U15472 (N_15472,N_13629,N_13835);
or U15473 (N_15473,N_12587,N_13090);
or U15474 (N_15474,N_13367,N_13209);
xor U15475 (N_15475,N_13968,N_12725);
and U15476 (N_15476,N_12891,N_12458);
and U15477 (N_15477,N_12949,N_12998);
and U15478 (N_15478,N_12867,N_12775);
xor U15479 (N_15479,N_12907,N_12207);
or U15480 (N_15480,N_13628,N_13130);
and U15481 (N_15481,N_12265,N_13958);
and U15482 (N_15482,N_13433,N_13630);
xor U15483 (N_15483,N_12229,N_12800);
and U15484 (N_15484,N_12651,N_12801);
nand U15485 (N_15485,N_13519,N_12230);
or U15486 (N_15486,N_12412,N_12444);
or U15487 (N_15487,N_12508,N_12806);
nand U15488 (N_15488,N_13418,N_13537);
nor U15489 (N_15489,N_12474,N_13914);
and U15490 (N_15490,N_12336,N_12672);
or U15491 (N_15491,N_13496,N_12727);
or U15492 (N_15492,N_12544,N_13517);
nand U15493 (N_15493,N_12946,N_12035);
and U15494 (N_15494,N_13022,N_13288);
or U15495 (N_15495,N_13177,N_12957);
nand U15496 (N_15496,N_12942,N_12458);
xor U15497 (N_15497,N_12389,N_12974);
and U15498 (N_15498,N_13135,N_12556);
nand U15499 (N_15499,N_13003,N_12691);
or U15500 (N_15500,N_13051,N_12530);
and U15501 (N_15501,N_12037,N_13578);
nand U15502 (N_15502,N_13547,N_12648);
nand U15503 (N_15503,N_12395,N_12165);
xor U15504 (N_15504,N_13491,N_13766);
nor U15505 (N_15505,N_12778,N_13746);
nor U15506 (N_15506,N_12240,N_13701);
xor U15507 (N_15507,N_13645,N_13691);
nand U15508 (N_15508,N_13027,N_13489);
or U15509 (N_15509,N_12882,N_12533);
nand U15510 (N_15510,N_13521,N_13164);
nand U15511 (N_15511,N_13737,N_12215);
nor U15512 (N_15512,N_13827,N_13136);
xor U15513 (N_15513,N_13089,N_12022);
nand U15514 (N_15514,N_12231,N_13883);
nor U15515 (N_15515,N_13198,N_13840);
or U15516 (N_15516,N_13292,N_12070);
nand U15517 (N_15517,N_12700,N_13130);
xnor U15518 (N_15518,N_12945,N_12846);
nor U15519 (N_15519,N_12212,N_12773);
nor U15520 (N_15520,N_13792,N_12420);
and U15521 (N_15521,N_13594,N_12684);
or U15522 (N_15522,N_12870,N_13626);
or U15523 (N_15523,N_13172,N_13527);
and U15524 (N_15524,N_12058,N_12467);
nor U15525 (N_15525,N_12961,N_12342);
and U15526 (N_15526,N_12719,N_12586);
nor U15527 (N_15527,N_12831,N_13236);
xnor U15528 (N_15528,N_12093,N_12458);
nand U15529 (N_15529,N_13548,N_13974);
and U15530 (N_15530,N_13843,N_13515);
nor U15531 (N_15531,N_12251,N_13305);
nand U15532 (N_15532,N_12527,N_12666);
nand U15533 (N_15533,N_12155,N_12130);
nand U15534 (N_15534,N_13011,N_12998);
or U15535 (N_15535,N_13448,N_12232);
xnor U15536 (N_15536,N_12137,N_13826);
nor U15537 (N_15537,N_12109,N_12987);
or U15538 (N_15538,N_13682,N_12668);
nor U15539 (N_15539,N_12953,N_12625);
nor U15540 (N_15540,N_13816,N_12053);
xor U15541 (N_15541,N_12917,N_12722);
or U15542 (N_15542,N_13036,N_12274);
nor U15543 (N_15543,N_13526,N_13963);
nor U15544 (N_15544,N_13828,N_13691);
nand U15545 (N_15545,N_13960,N_12284);
nand U15546 (N_15546,N_13313,N_12098);
xnor U15547 (N_15547,N_12393,N_13351);
xnor U15548 (N_15548,N_12978,N_13756);
and U15549 (N_15549,N_12650,N_13508);
or U15550 (N_15550,N_13887,N_12857);
and U15551 (N_15551,N_12894,N_13930);
and U15552 (N_15552,N_13357,N_13096);
and U15553 (N_15553,N_12063,N_13045);
or U15554 (N_15554,N_12064,N_12174);
nor U15555 (N_15555,N_12451,N_12902);
nand U15556 (N_15556,N_12901,N_13661);
nand U15557 (N_15557,N_13698,N_12935);
or U15558 (N_15558,N_13645,N_13693);
nand U15559 (N_15559,N_12606,N_13137);
xnor U15560 (N_15560,N_13238,N_12484);
and U15561 (N_15561,N_12924,N_12170);
or U15562 (N_15562,N_12943,N_12312);
and U15563 (N_15563,N_12752,N_13614);
nor U15564 (N_15564,N_12906,N_12458);
and U15565 (N_15565,N_12082,N_12087);
or U15566 (N_15566,N_13093,N_12225);
xnor U15567 (N_15567,N_13353,N_12653);
and U15568 (N_15568,N_12291,N_12626);
nor U15569 (N_15569,N_12916,N_12357);
or U15570 (N_15570,N_13575,N_12858);
nor U15571 (N_15571,N_13092,N_13695);
or U15572 (N_15572,N_12545,N_13836);
and U15573 (N_15573,N_12893,N_13948);
nor U15574 (N_15574,N_12504,N_13682);
nand U15575 (N_15575,N_13515,N_12318);
or U15576 (N_15576,N_12218,N_12371);
nor U15577 (N_15577,N_12975,N_12118);
nor U15578 (N_15578,N_13990,N_12090);
and U15579 (N_15579,N_13889,N_13138);
nand U15580 (N_15580,N_12114,N_12345);
xor U15581 (N_15581,N_13841,N_12779);
and U15582 (N_15582,N_12017,N_13385);
nor U15583 (N_15583,N_12207,N_12192);
nand U15584 (N_15584,N_13513,N_13853);
nand U15585 (N_15585,N_12210,N_12636);
nor U15586 (N_15586,N_12852,N_12737);
or U15587 (N_15587,N_13640,N_13708);
or U15588 (N_15588,N_12576,N_13915);
nand U15589 (N_15589,N_12400,N_12190);
and U15590 (N_15590,N_12507,N_12299);
nand U15591 (N_15591,N_12288,N_12557);
nor U15592 (N_15592,N_12110,N_13984);
nand U15593 (N_15593,N_12534,N_13026);
or U15594 (N_15594,N_13507,N_12734);
and U15595 (N_15595,N_13023,N_12894);
and U15596 (N_15596,N_12857,N_13709);
and U15597 (N_15597,N_13618,N_13587);
nor U15598 (N_15598,N_13614,N_13940);
nor U15599 (N_15599,N_13323,N_13489);
nor U15600 (N_15600,N_13116,N_13568);
nor U15601 (N_15601,N_13920,N_13992);
and U15602 (N_15602,N_13003,N_13417);
nand U15603 (N_15603,N_13611,N_12092);
and U15604 (N_15604,N_13123,N_13993);
nor U15605 (N_15605,N_12085,N_12279);
nor U15606 (N_15606,N_12909,N_13362);
nand U15607 (N_15607,N_12945,N_13296);
or U15608 (N_15608,N_12843,N_12573);
or U15609 (N_15609,N_12239,N_13108);
nand U15610 (N_15610,N_13371,N_12531);
xor U15611 (N_15611,N_13468,N_12054);
and U15612 (N_15612,N_13218,N_13592);
and U15613 (N_15613,N_13570,N_12584);
nand U15614 (N_15614,N_12685,N_13810);
nand U15615 (N_15615,N_12636,N_12032);
and U15616 (N_15616,N_13058,N_13297);
and U15617 (N_15617,N_12731,N_12257);
nor U15618 (N_15618,N_13692,N_13094);
nor U15619 (N_15619,N_13929,N_13012);
nor U15620 (N_15620,N_13904,N_13171);
or U15621 (N_15621,N_13168,N_13092);
and U15622 (N_15622,N_12959,N_12766);
nor U15623 (N_15623,N_13402,N_12870);
and U15624 (N_15624,N_13977,N_13702);
nand U15625 (N_15625,N_13061,N_13240);
nand U15626 (N_15626,N_13538,N_12869);
or U15627 (N_15627,N_12549,N_12676);
nor U15628 (N_15628,N_13898,N_12335);
nand U15629 (N_15629,N_13235,N_12922);
xor U15630 (N_15630,N_12347,N_13613);
xnor U15631 (N_15631,N_13592,N_12650);
xor U15632 (N_15632,N_12480,N_12849);
nand U15633 (N_15633,N_13662,N_12538);
xor U15634 (N_15634,N_13797,N_12111);
and U15635 (N_15635,N_12092,N_13996);
nor U15636 (N_15636,N_12811,N_13228);
nor U15637 (N_15637,N_12458,N_13559);
xor U15638 (N_15638,N_13904,N_12754);
xnor U15639 (N_15639,N_13797,N_13530);
xnor U15640 (N_15640,N_13032,N_12511);
or U15641 (N_15641,N_13579,N_12104);
nand U15642 (N_15642,N_13676,N_12566);
nor U15643 (N_15643,N_13424,N_12046);
and U15644 (N_15644,N_13320,N_13399);
or U15645 (N_15645,N_12609,N_13109);
or U15646 (N_15646,N_12305,N_13778);
nor U15647 (N_15647,N_12289,N_12782);
nor U15648 (N_15648,N_13095,N_13825);
and U15649 (N_15649,N_13734,N_13121);
xor U15650 (N_15650,N_12572,N_12864);
xor U15651 (N_15651,N_13920,N_13420);
or U15652 (N_15652,N_12148,N_12128);
xnor U15653 (N_15653,N_13084,N_12898);
or U15654 (N_15654,N_13469,N_12020);
and U15655 (N_15655,N_13845,N_12514);
nand U15656 (N_15656,N_13077,N_12795);
nand U15657 (N_15657,N_13750,N_13903);
or U15658 (N_15658,N_13576,N_13090);
nor U15659 (N_15659,N_13901,N_13489);
nand U15660 (N_15660,N_12552,N_12727);
nor U15661 (N_15661,N_13618,N_13570);
or U15662 (N_15662,N_12540,N_12420);
xnor U15663 (N_15663,N_13780,N_13963);
nand U15664 (N_15664,N_13981,N_12521);
nand U15665 (N_15665,N_13216,N_13221);
or U15666 (N_15666,N_12959,N_13117);
and U15667 (N_15667,N_13335,N_12500);
xor U15668 (N_15668,N_12805,N_12173);
nand U15669 (N_15669,N_13519,N_13295);
xor U15670 (N_15670,N_13285,N_13125);
xnor U15671 (N_15671,N_13298,N_12854);
or U15672 (N_15672,N_12604,N_13685);
and U15673 (N_15673,N_13925,N_13743);
or U15674 (N_15674,N_12184,N_12320);
nor U15675 (N_15675,N_12239,N_13540);
nor U15676 (N_15676,N_12404,N_12276);
and U15677 (N_15677,N_12583,N_12920);
nand U15678 (N_15678,N_13351,N_13429);
xnor U15679 (N_15679,N_12499,N_13881);
nand U15680 (N_15680,N_13895,N_12398);
and U15681 (N_15681,N_13866,N_13673);
or U15682 (N_15682,N_12503,N_13667);
nor U15683 (N_15683,N_12386,N_12739);
or U15684 (N_15684,N_13179,N_13276);
or U15685 (N_15685,N_13274,N_12576);
xor U15686 (N_15686,N_12890,N_12618);
nand U15687 (N_15687,N_13317,N_12272);
nor U15688 (N_15688,N_13582,N_12767);
or U15689 (N_15689,N_13147,N_13203);
nor U15690 (N_15690,N_13717,N_12660);
nor U15691 (N_15691,N_13982,N_13829);
or U15692 (N_15692,N_13276,N_13272);
or U15693 (N_15693,N_12236,N_12806);
nor U15694 (N_15694,N_12551,N_13673);
and U15695 (N_15695,N_13520,N_12808);
nand U15696 (N_15696,N_13662,N_12121);
xor U15697 (N_15697,N_12280,N_13161);
and U15698 (N_15698,N_13597,N_12368);
and U15699 (N_15699,N_13296,N_13040);
nor U15700 (N_15700,N_12160,N_13927);
or U15701 (N_15701,N_13005,N_12736);
nor U15702 (N_15702,N_13815,N_13758);
nor U15703 (N_15703,N_12644,N_12389);
and U15704 (N_15704,N_13364,N_12269);
and U15705 (N_15705,N_13280,N_13880);
and U15706 (N_15706,N_13815,N_13873);
nor U15707 (N_15707,N_13872,N_13539);
nor U15708 (N_15708,N_13265,N_13252);
or U15709 (N_15709,N_13715,N_13956);
or U15710 (N_15710,N_13651,N_12464);
nor U15711 (N_15711,N_12653,N_13650);
nor U15712 (N_15712,N_13792,N_12194);
nor U15713 (N_15713,N_12302,N_12192);
nand U15714 (N_15714,N_13737,N_13577);
nand U15715 (N_15715,N_12487,N_12662);
nand U15716 (N_15716,N_13517,N_13537);
xor U15717 (N_15717,N_12696,N_13076);
nand U15718 (N_15718,N_13994,N_13895);
and U15719 (N_15719,N_13726,N_13566);
nor U15720 (N_15720,N_12274,N_13755);
xnor U15721 (N_15721,N_12017,N_12964);
or U15722 (N_15722,N_13149,N_13868);
nand U15723 (N_15723,N_12711,N_12714);
nor U15724 (N_15724,N_13878,N_12982);
or U15725 (N_15725,N_13455,N_13723);
nand U15726 (N_15726,N_12532,N_12667);
and U15727 (N_15727,N_12919,N_13659);
nand U15728 (N_15728,N_13542,N_13797);
and U15729 (N_15729,N_13666,N_13185);
and U15730 (N_15730,N_13515,N_13426);
and U15731 (N_15731,N_13829,N_13820);
and U15732 (N_15732,N_12819,N_12950);
nand U15733 (N_15733,N_12246,N_12007);
and U15734 (N_15734,N_12435,N_12369);
and U15735 (N_15735,N_13773,N_12027);
xor U15736 (N_15736,N_13543,N_13361);
or U15737 (N_15737,N_13683,N_12239);
nor U15738 (N_15738,N_13215,N_12180);
nor U15739 (N_15739,N_12709,N_13431);
xnor U15740 (N_15740,N_13396,N_12830);
nor U15741 (N_15741,N_12809,N_12453);
xor U15742 (N_15742,N_12154,N_13691);
or U15743 (N_15743,N_13329,N_13288);
nor U15744 (N_15744,N_13268,N_12384);
nor U15745 (N_15745,N_13061,N_12827);
or U15746 (N_15746,N_13053,N_12633);
and U15747 (N_15747,N_13508,N_12539);
nand U15748 (N_15748,N_12520,N_12909);
and U15749 (N_15749,N_13147,N_13444);
nand U15750 (N_15750,N_12103,N_12821);
and U15751 (N_15751,N_12746,N_13325);
nor U15752 (N_15752,N_12357,N_12820);
nand U15753 (N_15753,N_13246,N_13613);
nor U15754 (N_15754,N_13690,N_12591);
or U15755 (N_15755,N_13387,N_12618);
or U15756 (N_15756,N_12899,N_12707);
and U15757 (N_15757,N_13315,N_12285);
xor U15758 (N_15758,N_13526,N_13169);
or U15759 (N_15759,N_13036,N_12924);
and U15760 (N_15760,N_13776,N_12793);
or U15761 (N_15761,N_12666,N_12322);
nand U15762 (N_15762,N_13334,N_13792);
xor U15763 (N_15763,N_13634,N_13162);
nor U15764 (N_15764,N_13247,N_12582);
xor U15765 (N_15765,N_13645,N_12501);
and U15766 (N_15766,N_12034,N_12278);
nor U15767 (N_15767,N_13509,N_13508);
nand U15768 (N_15768,N_12548,N_13900);
and U15769 (N_15769,N_13635,N_13082);
xor U15770 (N_15770,N_13676,N_12991);
or U15771 (N_15771,N_12953,N_13109);
nor U15772 (N_15772,N_12390,N_13484);
or U15773 (N_15773,N_13142,N_12259);
nor U15774 (N_15774,N_13163,N_13342);
nor U15775 (N_15775,N_12339,N_13163);
or U15776 (N_15776,N_12382,N_13839);
nand U15777 (N_15777,N_13483,N_12919);
and U15778 (N_15778,N_13425,N_13831);
xor U15779 (N_15779,N_13699,N_12285);
nand U15780 (N_15780,N_13546,N_12944);
nand U15781 (N_15781,N_12289,N_13279);
xor U15782 (N_15782,N_13815,N_12715);
or U15783 (N_15783,N_12180,N_13927);
nor U15784 (N_15784,N_12999,N_13916);
and U15785 (N_15785,N_12817,N_12216);
or U15786 (N_15786,N_13288,N_12336);
nor U15787 (N_15787,N_13507,N_13421);
nor U15788 (N_15788,N_12697,N_13823);
or U15789 (N_15789,N_13736,N_13071);
and U15790 (N_15790,N_13159,N_13693);
and U15791 (N_15791,N_12404,N_12221);
xor U15792 (N_15792,N_13286,N_13202);
nand U15793 (N_15793,N_13170,N_12681);
nand U15794 (N_15794,N_13271,N_12531);
xor U15795 (N_15795,N_12372,N_13047);
nand U15796 (N_15796,N_13045,N_12678);
or U15797 (N_15797,N_12675,N_12239);
nand U15798 (N_15798,N_12932,N_12516);
nor U15799 (N_15799,N_13007,N_12183);
and U15800 (N_15800,N_12905,N_12512);
xnor U15801 (N_15801,N_12170,N_12545);
or U15802 (N_15802,N_12682,N_12324);
nor U15803 (N_15803,N_12744,N_12251);
or U15804 (N_15804,N_12684,N_13267);
nand U15805 (N_15805,N_12738,N_12373);
or U15806 (N_15806,N_13532,N_13391);
or U15807 (N_15807,N_12710,N_12590);
nor U15808 (N_15808,N_12529,N_12804);
xnor U15809 (N_15809,N_13271,N_12545);
and U15810 (N_15810,N_12688,N_12618);
nand U15811 (N_15811,N_12586,N_13968);
and U15812 (N_15812,N_13397,N_12221);
and U15813 (N_15813,N_13162,N_12618);
or U15814 (N_15814,N_12204,N_13037);
xnor U15815 (N_15815,N_12599,N_13159);
xnor U15816 (N_15816,N_13507,N_13659);
or U15817 (N_15817,N_12712,N_12554);
or U15818 (N_15818,N_12850,N_13597);
and U15819 (N_15819,N_12023,N_13106);
or U15820 (N_15820,N_13897,N_13570);
and U15821 (N_15821,N_13221,N_13799);
nor U15822 (N_15822,N_12142,N_12809);
xnor U15823 (N_15823,N_12322,N_12181);
nand U15824 (N_15824,N_13919,N_12478);
or U15825 (N_15825,N_12173,N_12263);
xnor U15826 (N_15826,N_13414,N_12577);
nand U15827 (N_15827,N_13184,N_13616);
or U15828 (N_15828,N_12264,N_12194);
or U15829 (N_15829,N_13687,N_13859);
or U15830 (N_15830,N_12765,N_13678);
nor U15831 (N_15831,N_13915,N_13803);
and U15832 (N_15832,N_13678,N_12285);
nand U15833 (N_15833,N_12440,N_13081);
nor U15834 (N_15834,N_12972,N_12364);
nand U15835 (N_15835,N_13986,N_12428);
or U15836 (N_15836,N_13926,N_13707);
nor U15837 (N_15837,N_13289,N_12646);
nand U15838 (N_15838,N_13197,N_12457);
nand U15839 (N_15839,N_13076,N_13466);
nand U15840 (N_15840,N_13630,N_12677);
xnor U15841 (N_15841,N_13191,N_12893);
or U15842 (N_15842,N_12463,N_12824);
and U15843 (N_15843,N_13062,N_12172);
nand U15844 (N_15844,N_13025,N_12252);
or U15845 (N_15845,N_12800,N_12237);
nand U15846 (N_15846,N_13483,N_13353);
or U15847 (N_15847,N_12412,N_13735);
or U15848 (N_15848,N_13550,N_12997);
or U15849 (N_15849,N_13031,N_13449);
nor U15850 (N_15850,N_12344,N_13378);
or U15851 (N_15851,N_13684,N_12883);
or U15852 (N_15852,N_12909,N_12339);
and U15853 (N_15853,N_13952,N_12821);
and U15854 (N_15854,N_12524,N_13014);
nand U15855 (N_15855,N_13969,N_12401);
nand U15856 (N_15856,N_13290,N_13523);
or U15857 (N_15857,N_12858,N_12521);
and U15858 (N_15858,N_13878,N_13112);
nand U15859 (N_15859,N_12417,N_13985);
nor U15860 (N_15860,N_12413,N_13120);
nor U15861 (N_15861,N_12679,N_13894);
xnor U15862 (N_15862,N_13768,N_13165);
or U15863 (N_15863,N_12434,N_13679);
nor U15864 (N_15864,N_13958,N_13113);
and U15865 (N_15865,N_12108,N_12861);
and U15866 (N_15866,N_12434,N_13992);
or U15867 (N_15867,N_13853,N_13998);
nand U15868 (N_15868,N_13771,N_13141);
xnor U15869 (N_15869,N_13890,N_13880);
nand U15870 (N_15870,N_13329,N_12786);
or U15871 (N_15871,N_13613,N_12943);
and U15872 (N_15872,N_12709,N_12668);
nor U15873 (N_15873,N_13274,N_12907);
nand U15874 (N_15874,N_13563,N_13110);
nor U15875 (N_15875,N_12696,N_13716);
nor U15876 (N_15876,N_13311,N_12395);
xnor U15877 (N_15877,N_12739,N_13686);
nor U15878 (N_15878,N_13879,N_12315);
nor U15879 (N_15879,N_12089,N_13735);
and U15880 (N_15880,N_13639,N_13924);
xor U15881 (N_15881,N_12749,N_13424);
or U15882 (N_15882,N_12562,N_12342);
nor U15883 (N_15883,N_13494,N_12898);
nor U15884 (N_15884,N_12149,N_12944);
and U15885 (N_15885,N_12407,N_12886);
nand U15886 (N_15886,N_13691,N_12559);
nand U15887 (N_15887,N_13929,N_13105);
and U15888 (N_15888,N_13312,N_13654);
nand U15889 (N_15889,N_12685,N_13212);
nand U15890 (N_15890,N_12138,N_13626);
nor U15891 (N_15891,N_12821,N_12693);
and U15892 (N_15892,N_12829,N_13246);
nor U15893 (N_15893,N_12514,N_13170);
nor U15894 (N_15894,N_12944,N_13596);
nor U15895 (N_15895,N_12503,N_12296);
and U15896 (N_15896,N_12434,N_12065);
or U15897 (N_15897,N_13986,N_12900);
or U15898 (N_15898,N_12917,N_13384);
nand U15899 (N_15899,N_12892,N_12191);
nor U15900 (N_15900,N_13872,N_12685);
and U15901 (N_15901,N_12879,N_12307);
or U15902 (N_15902,N_12962,N_13203);
and U15903 (N_15903,N_12681,N_13977);
nand U15904 (N_15904,N_13744,N_13283);
or U15905 (N_15905,N_12752,N_13891);
nand U15906 (N_15906,N_13417,N_13044);
nor U15907 (N_15907,N_12023,N_12477);
xor U15908 (N_15908,N_12077,N_12314);
nor U15909 (N_15909,N_13348,N_12910);
or U15910 (N_15910,N_12268,N_12893);
nand U15911 (N_15911,N_13582,N_12984);
nand U15912 (N_15912,N_12978,N_13987);
nor U15913 (N_15913,N_13368,N_12222);
or U15914 (N_15914,N_12803,N_12997);
or U15915 (N_15915,N_12931,N_12060);
or U15916 (N_15916,N_13933,N_13757);
and U15917 (N_15917,N_13178,N_12678);
or U15918 (N_15918,N_12656,N_13074);
xnor U15919 (N_15919,N_12166,N_13622);
xnor U15920 (N_15920,N_13574,N_13030);
nand U15921 (N_15921,N_12481,N_13914);
or U15922 (N_15922,N_12757,N_12900);
xor U15923 (N_15923,N_13950,N_12586);
nor U15924 (N_15924,N_12956,N_13556);
nand U15925 (N_15925,N_12346,N_12864);
nand U15926 (N_15926,N_12050,N_13299);
or U15927 (N_15927,N_13822,N_12236);
nand U15928 (N_15928,N_13572,N_12115);
nand U15929 (N_15929,N_13734,N_12634);
nor U15930 (N_15930,N_12005,N_12504);
nor U15931 (N_15931,N_12756,N_12842);
and U15932 (N_15932,N_13916,N_12496);
nor U15933 (N_15933,N_12911,N_13056);
nor U15934 (N_15934,N_13922,N_13158);
nor U15935 (N_15935,N_13761,N_13496);
xnor U15936 (N_15936,N_13768,N_12071);
nand U15937 (N_15937,N_12962,N_12208);
xnor U15938 (N_15938,N_13297,N_12983);
nor U15939 (N_15939,N_12192,N_12216);
and U15940 (N_15940,N_12947,N_13916);
and U15941 (N_15941,N_13699,N_12630);
or U15942 (N_15942,N_13553,N_12674);
and U15943 (N_15943,N_13468,N_12932);
xnor U15944 (N_15944,N_13306,N_13628);
or U15945 (N_15945,N_13263,N_12530);
and U15946 (N_15946,N_12277,N_13976);
or U15947 (N_15947,N_12467,N_13709);
nand U15948 (N_15948,N_13152,N_13094);
nor U15949 (N_15949,N_12346,N_13787);
xor U15950 (N_15950,N_12388,N_12810);
nor U15951 (N_15951,N_13941,N_12794);
or U15952 (N_15952,N_13534,N_13093);
and U15953 (N_15953,N_12157,N_13425);
nor U15954 (N_15954,N_13603,N_12972);
nand U15955 (N_15955,N_13905,N_13843);
nand U15956 (N_15956,N_12971,N_13580);
or U15957 (N_15957,N_13735,N_12870);
nand U15958 (N_15958,N_12426,N_13756);
nand U15959 (N_15959,N_12417,N_12119);
nor U15960 (N_15960,N_12357,N_13984);
or U15961 (N_15961,N_13789,N_13134);
and U15962 (N_15962,N_13513,N_13539);
nand U15963 (N_15963,N_12917,N_13097);
nand U15964 (N_15964,N_12511,N_12691);
or U15965 (N_15965,N_12816,N_13797);
and U15966 (N_15966,N_13440,N_13968);
nor U15967 (N_15967,N_13036,N_12318);
nand U15968 (N_15968,N_13481,N_13511);
xnor U15969 (N_15969,N_13308,N_13639);
and U15970 (N_15970,N_12189,N_13171);
and U15971 (N_15971,N_13590,N_13214);
nand U15972 (N_15972,N_13316,N_12210);
or U15973 (N_15973,N_12850,N_13016);
nand U15974 (N_15974,N_12546,N_12250);
or U15975 (N_15975,N_12287,N_12940);
nand U15976 (N_15976,N_12888,N_13785);
and U15977 (N_15977,N_12125,N_12932);
nand U15978 (N_15978,N_13776,N_12501);
nand U15979 (N_15979,N_13922,N_12685);
or U15980 (N_15980,N_13182,N_12160);
nor U15981 (N_15981,N_12247,N_13800);
nand U15982 (N_15982,N_13545,N_12873);
and U15983 (N_15983,N_12098,N_12072);
nor U15984 (N_15984,N_13282,N_13021);
and U15985 (N_15985,N_12574,N_12618);
and U15986 (N_15986,N_13876,N_13964);
and U15987 (N_15987,N_12239,N_12682);
nor U15988 (N_15988,N_12035,N_12002);
nand U15989 (N_15989,N_12769,N_12172);
and U15990 (N_15990,N_12887,N_12603);
and U15991 (N_15991,N_12312,N_13551);
and U15992 (N_15992,N_13448,N_12712);
and U15993 (N_15993,N_12768,N_13715);
and U15994 (N_15994,N_12276,N_13244);
nor U15995 (N_15995,N_12102,N_12519);
nand U15996 (N_15996,N_13643,N_13000);
xor U15997 (N_15997,N_12209,N_12729);
nor U15998 (N_15998,N_12406,N_12353);
and U15999 (N_15999,N_13796,N_13635);
or U16000 (N_16000,N_14528,N_15763);
or U16001 (N_16001,N_14781,N_14938);
and U16002 (N_16002,N_15647,N_14981);
nor U16003 (N_16003,N_14130,N_14026);
and U16004 (N_16004,N_14106,N_15029);
nand U16005 (N_16005,N_14114,N_14457);
nand U16006 (N_16006,N_15752,N_14933);
nand U16007 (N_16007,N_14629,N_14850);
and U16008 (N_16008,N_14198,N_15629);
or U16009 (N_16009,N_15312,N_15194);
xor U16010 (N_16010,N_15540,N_15987);
nand U16011 (N_16011,N_15329,N_15601);
nand U16012 (N_16012,N_15280,N_14823);
or U16013 (N_16013,N_15444,N_15301);
xor U16014 (N_16014,N_14094,N_14014);
or U16015 (N_16015,N_14223,N_14082);
or U16016 (N_16016,N_14243,N_14421);
nor U16017 (N_16017,N_15972,N_14076);
or U16018 (N_16018,N_15900,N_15579);
nand U16019 (N_16019,N_15798,N_14408);
xnor U16020 (N_16020,N_14202,N_15710);
nor U16021 (N_16021,N_15176,N_14530);
and U16022 (N_16022,N_14755,N_15567);
or U16023 (N_16023,N_14095,N_14443);
nor U16024 (N_16024,N_14277,N_15143);
nor U16025 (N_16025,N_15907,N_15469);
and U16026 (N_16026,N_14455,N_15576);
and U16027 (N_16027,N_15220,N_14839);
or U16028 (N_16028,N_15980,N_15273);
and U16029 (N_16029,N_14797,N_15451);
xnor U16030 (N_16030,N_15209,N_15111);
or U16031 (N_16031,N_15470,N_15170);
nand U16032 (N_16032,N_14716,N_15914);
nand U16033 (N_16033,N_15373,N_15284);
nand U16034 (N_16034,N_15453,N_14438);
or U16035 (N_16035,N_15124,N_14205);
nor U16036 (N_16036,N_14520,N_15838);
and U16037 (N_16037,N_15774,N_14749);
xor U16038 (N_16038,N_15298,N_14779);
nor U16039 (N_16039,N_14939,N_14853);
xor U16040 (N_16040,N_15251,N_14852);
and U16041 (N_16041,N_14306,N_15345);
nor U16042 (N_16042,N_15331,N_14843);
nor U16043 (N_16043,N_14739,N_15504);
nor U16044 (N_16044,N_14167,N_14038);
nor U16045 (N_16045,N_15589,N_14045);
and U16046 (N_16046,N_15719,N_14638);
or U16047 (N_16047,N_14290,N_15533);
and U16048 (N_16048,N_14023,N_15125);
nor U16049 (N_16049,N_14169,N_15510);
nand U16050 (N_16050,N_15463,N_15782);
and U16051 (N_16051,N_15435,N_14654);
nor U16052 (N_16052,N_15982,N_14664);
nand U16053 (N_16053,N_15321,N_15546);
or U16054 (N_16054,N_15711,N_15458);
nor U16055 (N_16055,N_14774,N_14371);
nand U16056 (N_16056,N_14342,N_15011);
nand U16057 (N_16057,N_15702,N_14656);
nand U16058 (N_16058,N_14985,N_14281);
or U16059 (N_16059,N_14357,N_15423);
and U16060 (N_16060,N_14419,N_15722);
or U16061 (N_16061,N_15252,N_15572);
or U16062 (N_16062,N_15202,N_14002);
and U16063 (N_16063,N_14524,N_15607);
nand U16064 (N_16064,N_15799,N_14297);
or U16065 (N_16065,N_14212,N_15267);
xnor U16066 (N_16066,N_15067,N_15317);
xnor U16067 (N_16067,N_15055,N_15214);
or U16068 (N_16068,N_15633,N_15908);
nand U16069 (N_16069,N_14775,N_15159);
and U16070 (N_16070,N_14517,N_14148);
xor U16071 (N_16071,N_15367,N_15855);
nor U16072 (N_16072,N_14879,N_14177);
or U16073 (N_16073,N_14888,N_15857);
or U16074 (N_16074,N_14617,N_14583);
or U16075 (N_16075,N_15790,N_14838);
nand U16076 (N_16076,N_14450,N_15179);
and U16077 (N_16077,N_14253,N_15973);
and U16078 (N_16078,N_15115,N_15324);
nand U16079 (N_16079,N_14526,N_15081);
nand U16080 (N_16080,N_15825,N_14559);
or U16081 (N_16081,N_14782,N_14780);
nand U16082 (N_16082,N_15609,N_14941);
or U16083 (N_16083,N_15613,N_15048);
or U16084 (N_16084,N_15729,N_14914);
and U16085 (N_16085,N_15526,N_15764);
and U16086 (N_16086,N_14927,N_14074);
and U16087 (N_16087,N_15287,N_14633);
and U16088 (N_16088,N_14066,N_15460);
nand U16089 (N_16089,N_15571,N_14579);
and U16090 (N_16090,N_14112,N_14407);
and U16091 (N_16091,N_14433,N_14098);
nand U16092 (N_16092,N_15657,N_14859);
nor U16093 (N_16093,N_15932,N_14931);
nor U16094 (N_16094,N_15052,N_14372);
nor U16095 (N_16095,N_15901,N_14562);
and U16096 (N_16096,N_15320,N_15690);
nor U16097 (N_16097,N_15920,N_15664);
xor U16098 (N_16098,N_14005,N_14195);
or U16099 (N_16099,N_15046,N_15683);
nor U16100 (N_16100,N_15065,N_14035);
nand U16101 (N_16101,N_15006,N_15465);
nor U16102 (N_16102,N_15930,N_15557);
nor U16103 (N_16103,N_15285,N_14245);
or U16104 (N_16104,N_14511,N_14204);
nand U16105 (N_16105,N_14635,N_15314);
nor U16106 (N_16106,N_14685,N_14875);
nor U16107 (N_16107,N_14668,N_14851);
nand U16108 (N_16108,N_14261,N_14976);
or U16109 (N_16109,N_14464,N_14418);
nand U16110 (N_16110,N_14601,N_14948);
and U16111 (N_16111,N_14896,N_15655);
nor U16112 (N_16112,N_14891,N_14145);
xor U16113 (N_16113,N_14570,N_14550);
nand U16114 (N_16114,N_15130,N_14993);
nand U16115 (N_16115,N_15080,N_14764);
and U16116 (N_16116,N_14961,N_14734);
or U16117 (N_16117,N_15021,N_15534);
and U16118 (N_16118,N_15337,N_14847);
or U16119 (N_16119,N_15759,N_15161);
or U16120 (N_16120,N_14122,N_14574);
and U16121 (N_16121,N_14725,N_14730);
nor U16122 (N_16122,N_14756,N_14238);
nand U16123 (N_16123,N_15456,N_14679);
and U16124 (N_16124,N_15955,N_15559);
nand U16125 (N_16125,N_14793,N_14150);
nor U16126 (N_16126,N_14310,N_15926);
and U16127 (N_16127,N_14867,N_15139);
nand U16128 (N_16128,N_15007,N_14251);
nor U16129 (N_16129,N_15902,N_15186);
and U16130 (N_16130,N_15461,N_14485);
and U16131 (N_16131,N_14828,N_15054);
or U16132 (N_16132,N_14950,N_14370);
nor U16133 (N_16133,N_14631,N_14747);
nor U16134 (N_16134,N_14615,N_14028);
xnor U16135 (N_16135,N_15598,N_14237);
nand U16136 (N_16136,N_15019,N_14271);
and U16137 (N_16137,N_14326,N_15586);
or U16138 (N_16138,N_15568,N_14362);
or U16139 (N_16139,N_14584,N_15307);
or U16140 (N_16140,N_15207,N_14701);
or U16141 (N_16141,N_14568,N_15233);
nor U16142 (N_16142,N_15163,N_15483);
or U16143 (N_16143,N_14270,N_15529);
nor U16144 (N_16144,N_14665,N_15308);
xnor U16145 (N_16145,N_15695,N_15403);
nor U16146 (N_16146,N_14576,N_15993);
or U16147 (N_16147,N_15532,N_15409);
and U16148 (N_16148,N_14022,N_15994);
or U16149 (N_16149,N_14467,N_15374);
nor U16150 (N_16150,N_14489,N_15553);
or U16151 (N_16151,N_14115,N_15262);
or U16152 (N_16152,N_15821,N_15478);
xor U16153 (N_16153,N_14795,N_15666);
nor U16154 (N_16154,N_15911,N_14469);
or U16155 (N_16155,N_14391,N_15661);
or U16156 (N_16156,N_14406,N_14534);
nand U16157 (N_16157,N_15783,N_14249);
nor U16158 (N_16158,N_14994,N_14415);
xor U16159 (N_16159,N_15728,N_14540);
nor U16160 (N_16160,N_15610,N_14432);
nand U16161 (N_16161,N_14936,N_15667);
nand U16162 (N_16162,N_14283,N_14055);
nor U16163 (N_16163,N_14211,N_14872);
nand U16164 (N_16164,N_15358,N_14302);
and U16165 (N_16165,N_14762,N_14091);
and U16166 (N_16166,N_15032,N_15175);
or U16167 (N_16167,N_14296,N_14322);
xnor U16168 (N_16168,N_15346,N_15261);
nand U16169 (N_16169,N_14116,N_15462);
and U16170 (N_16170,N_14179,N_15140);
nand U16171 (N_16171,N_14539,N_15241);
and U16172 (N_16172,N_14693,N_14063);
nand U16173 (N_16173,N_15889,N_15891);
nand U16174 (N_16174,N_15943,N_14364);
xor U16175 (N_16175,N_14324,N_14710);
nand U16176 (N_16176,N_14643,N_15810);
nor U16177 (N_16177,N_14493,N_15039);
or U16178 (N_16178,N_14378,N_14811);
nand U16179 (N_16179,N_15584,N_14806);
nand U16180 (N_16180,N_15995,N_15103);
or U16181 (N_16181,N_15068,N_15523);
nand U16182 (N_16182,N_14307,N_15548);
and U16183 (N_16183,N_15508,N_15935);
xor U16184 (N_16184,N_15873,N_15269);
nand U16185 (N_16185,N_14057,N_15757);
xor U16186 (N_16186,N_15593,N_14620);
or U16187 (N_16187,N_14299,N_14887);
and U16188 (N_16188,N_14712,N_15834);
xor U16189 (N_16189,N_14904,N_15187);
nor U16190 (N_16190,N_15615,N_14325);
or U16191 (N_16191,N_15828,N_15389);
and U16192 (N_16192,N_15845,N_14155);
nand U16193 (N_16193,N_15998,N_15477);
or U16194 (N_16194,N_14841,N_15225);
or U16195 (N_16195,N_15354,N_14247);
or U16196 (N_16196,N_15942,N_14572);
nor U16197 (N_16197,N_15182,N_15105);
or U16198 (N_16198,N_14604,N_14801);
nor U16199 (N_16199,N_14442,N_14889);
nand U16200 (N_16200,N_15419,N_15991);
nand U16201 (N_16201,N_15335,N_14153);
or U16202 (N_16202,N_14273,N_14869);
nor U16203 (N_16203,N_15650,N_14695);
nor U16204 (N_16204,N_14717,N_14567);
or U16205 (N_16205,N_15392,N_14836);
nand U16206 (N_16206,N_14451,N_15372);
nor U16207 (N_16207,N_14566,N_14514);
and U16208 (N_16208,N_15753,N_14462);
nand U16209 (N_16209,N_14110,N_14918);
nor U16210 (N_16210,N_15652,N_14741);
or U16211 (N_16211,N_14009,N_15506);
and U16212 (N_16212,N_14974,N_14949);
xor U16213 (N_16213,N_14292,N_14963);
or U16214 (N_16214,N_14006,N_15405);
nor U16215 (N_16215,N_14365,N_15224);
nor U16216 (N_16216,N_14424,N_14760);
nand U16217 (N_16217,N_15659,N_15122);
nand U16218 (N_16218,N_14487,N_14895);
nor U16219 (N_16219,N_15236,N_15137);
nand U16220 (N_16220,N_15814,N_14481);
nand U16221 (N_16221,N_14124,N_15573);
and U16222 (N_16222,N_14655,N_14414);
or U16223 (N_16223,N_14845,N_15371);
or U16224 (N_16224,N_14886,N_15760);
nor U16225 (N_16225,N_14625,N_15575);
and U16226 (N_16226,N_15671,N_15274);
or U16227 (N_16227,N_14533,N_14977);
nor U16228 (N_16228,N_14405,N_14446);
and U16229 (N_16229,N_15512,N_15867);
or U16230 (N_16230,N_15906,N_15294);
xnor U16231 (N_16231,N_14587,N_15809);
xor U16232 (N_16232,N_14348,N_14930);
nor U16233 (N_16233,N_15616,N_15746);
and U16234 (N_16234,N_15921,N_15758);
or U16235 (N_16235,N_14649,N_15196);
or U16236 (N_16236,N_14017,N_15502);
nor U16237 (N_16237,N_14700,N_15201);
nor U16238 (N_16238,N_14355,N_14968);
nor U16239 (N_16239,N_15747,N_14666);
or U16240 (N_16240,N_14784,N_15235);
nor U16241 (N_16241,N_14294,N_15905);
xor U16242 (N_16242,N_14909,N_15596);
nor U16243 (N_16243,N_14436,N_14863);
and U16244 (N_16244,N_15387,N_15248);
or U16245 (N_16245,N_15428,N_15913);
nor U16246 (N_16246,N_15933,N_15802);
and U16247 (N_16247,N_14804,N_14316);
nor U16248 (N_16248,N_14382,N_14135);
nand U16249 (N_16249,N_15471,N_15524);
nor U16250 (N_16250,N_14965,N_15624);
and U16251 (N_16251,N_14975,N_15058);
nor U16252 (N_16252,N_15434,N_15846);
nor U16253 (N_16253,N_15852,N_15736);
or U16254 (N_16254,N_15513,N_14547);
and U16255 (N_16255,N_14537,N_14794);
or U16256 (N_16256,N_15396,N_15792);
nand U16257 (N_16257,N_14934,N_15896);
and U16258 (N_16258,N_15592,N_14726);
nor U16259 (N_16259,N_15075,N_15594);
and U16260 (N_16260,N_14815,N_14293);
and U16261 (N_16261,N_15494,N_15992);
and U16262 (N_16262,N_14042,N_14551);
and U16263 (N_16263,N_14754,N_15341);
or U16264 (N_16264,N_14343,N_14377);
or U16265 (N_16265,N_14422,N_14905);
and U16266 (N_16266,N_14721,N_15964);
or U16267 (N_16267,N_15833,N_14787);
and U16268 (N_16268,N_14192,N_14921);
or U16269 (N_16269,N_14692,N_15884);
nor U16270 (N_16270,N_15378,N_14291);
and U16271 (N_16271,N_15511,N_15611);
nand U16272 (N_16272,N_14230,N_14672);
nand U16273 (N_16273,N_14733,N_15042);
nand U16274 (N_16274,N_15221,N_15129);
nand U16275 (N_16275,N_14379,N_15436);
and U16276 (N_16276,N_14241,N_15218);
and U16277 (N_16277,N_14627,N_14546);
xor U16278 (N_16278,N_14552,N_14103);
nand U16279 (N_16279,N_15489,N_15687);
nand U16280 (N_16280,N_15355,N_15574);
nor U16281 (N_16281,N_14353,N_15041);
nand U16282 (N_16282,N_15643,N_15986);
nand U16283 (N_16283,N_14070,N_14099);
or U16284 (N_16284,N_14830,N_14813);
or U16285 (N_16285,N_15984,N_14681);
and U16286 (N_16286,N_14501,N_14108);
and U16287 (N_16287,N_14286,N_15530);
nand U16288 (N_16288,N_15850,N_15204);
and U16289 (N_16289,N_14608,N_14588);
nor U16290 (N_16290,N_15569,N_15038);
and U16291 (N_16291,N_15626,N_14460);
and U16292 (N_16292,N_15599,N_15027);
nand U16293 (N_16293,N_14705,N_15953);
nand U16294 (N_16294,N_15543,N_15727);
xor U16295 (N_16295,N_15895,N_14820);
nor U16296 (N_16296,N_14262,N_14553);
or U16297 (N_16297,N_14252,N_15432);
nand U16298 (N_16298,N_14164,N_15198);
or U16299 (N_16299,N_15768,N_14288);
nor U16300 (N_16300,N_14102,N_15253);
nor U16301 (N_16301,N_14036,N_14728);
or U16302 (N_16302,N_14519,N_15679);
nand U16303 (N_16303,N_14234,N_15558);
nand U16304 (N_16304,N_14007,N_15726);
and U16305 (N_16305,N_15836,N_15564);
nor U16306 (N_16306,N_15674,N_15565);
and U16307 (N_16307,N_15842,N_14531);
nand U16308 (N_16308,N_14248,N_15527);
nor U16309 (N_16309,N_15244,N_14492);
and U16310 (N_16310,N_15051,N_15088);
or U16311 (N_16311,N_14833,N_14671);
xor U16312 (N_16312,N_15591,N_15493);
and U16313 (N_16313,N_14956,N_15577);
nor U16314 (N_16314,N_14603,N_15542);
nor U16315 (N_16315,N_14605,N_14789);
nor U16316 (N_16316,N_14769,N_15990);
or U16317 (N_16317,N_15254,N_14136);
nand U16318 (N_16318,N_14829,N_15627);
nand U16319 (N_16319,N_15823,N_14313);
nand U16320 (N_16320,N_15397,N_14004);
and U16321 (N_16321,N_15874,N_15297);
or U16322 (N_16322,N_15222,N_15794);
and U16323 (N_16323,N_14011,N_14101);
nand U16324 (N_16324,N_15965,N_14500);
or U16325 (N_16325,N_15136,N_15875);
nand U16326 (N_16326,N_14621,N_15631);
nor U16327 (N_16327,N_15438,N_15215);
or U16328 (N_16328,N_14242,N_15488);
xnor U16329 (N_16329,N_15581,N_14885);
and U16330 (N_16330,N_15277,N_15816);
or U16331 (N_16331,N_14221,N_14233);
nor U16332 (N_16332,N_14864,N_15339);
nand U16333 (N_16333,N_14352,N_15872);
nor U16334 (N_16334,N_14630,N_14439);
nor U16335 (N_16335,N_15074,N_15500);
and U16336 (N_16336,N_14020,N_14600);
or U16337 (N_16337,N_14923,N_15089);
nor U16338 (N_16338,N_15474,N_14510);
nor U16339 (N_16339,N_15820,N_15279);
and U16340 (N_16340,N_15383,N_14118);
and U16341 (N_16341,N_15151,N_14137);
xnor U16342 (N_16342,N_14381,N_15732);
or U16343 (N_16343,N_15535,N_14881);
nand U16344 (N_16344,N_15888,N_14545);
nand U16345 (N_16345,N_15446,N_14062);
or U16346 (N_16346,N_14339,N_15352);
xor U16347 (N_16347,N_15501,N_15484);
nor U16348 (N_16348,N_14081,N_14276);
nand U16349 (N_16349,N_14997,N_15743);
nand U16350 (N_16350,N_14097,N_14384);
or U16351 (N_16351,N_14704,N_14235);
or U16352 (N_16352,N_14127,N_14901);
and U16353 (N_16353,N_14799,N_15158);
nand U16354 (N_16354,N_14910,N_15417);
nand U16355 (N_16355,N_14972,N_15516);
nand U16356 (N_16356,N_15549,N_14999);
and U16357 (N_16357,N_14622,N_15881);
nor U16358 (N_16358,N_14465,N_15045);
nand U16359 (N_16359,N_15439,N_14945);
nand U16360 (N_16360,N_14295,N_15865);
and U16361 (N_16361,N_14088,N_15924);
nand U16362 (N_16362,N_15134,N_15879);
nand U16363 (N_16363,N_15721,N_15398);
and U16364 (N_16364,N_14722,N_15013);
or U16365 (N_16365,N_14808,N_14474);
nor U16366 (N_16366,N_14490,N_14340);
or U16367 (N_16367,N_14554,N_15166);
xnor U16368 (N_16368,N_14947,N_14639);
nor U16369 (N_16369,N_14428,N_14334);
nor U16370 (N_16370,N_15983,N_15288);
nand U16371 (N_16371,N_15937,N_15227);
and U16372 (N_16372,N_14516,N_14527);
nand U16373 (N_16373,N_15947,N_14134);
and U16374 (N_16374,N_15399,N_14440);
and U16375 (N_16375,N_14079,N_15360);
nand U16376 (N_16376,N_15328,N_15603);
xnor U16377 (N_16377,N_14185,N_15773);
nand U16378 (N_16378,N_15377,N_14987);
and U16379 (N_16379,N_14031,N_14816);
nand U16380 (N_16380,N_15681,N_15276);
nor U16381 (N_16381,N_14937,N_15442);
nor U16382 (N_16382,N_14731,N_15044);
or U16383 (N_16383,N_14080,N_14093);
or U16384 (N_16384,N_15651,N_14351);
nor U16385 (N_16385,N_14188,N_15580);
and U16386 (N_16386,N_15272,N_15375);
or U16387 (N_16387,N_15738,N_14647);
nor U16388 (N_16388,N_14819,N_15467);
xnor U16389 (N_16389,N_15000,N_15265);
and U16390 (N_16390,N_15796,N_14250);
xor U16391 (N_16391,N_15518,N_15079);
or U16392 (N_16392,N_15049,N_14935);
nor U16393 (N_16393,N_14040,N_14049);
xnor U16394 (N_16394,N_15514,N_14626);
nand U16395 (N_16395,N_15334,N_14577);
nand U16396 (N_16396,N_15152,N_15084);
or U16397 (N_16397,N_15441,N_15795);
nand U16398 (N_16398,N_14129,N_14345);
and U16399 (N_16399,N_14254,N_14398);
xor U16400 (N_16400,N_15754,N_14318);
and U16401 (N_16401,N_14111,N_15211);
and U16402 (N_16402,N_15713,N_14506);
or U16403 (N_16403,N_15856,N_15357);
or U16404 (N_16404,N_15365,N_15862);
and U16405 (N_16405,N_14542,N_15015);
nor U16406 (N_16406,N_14767,N_14019);
and U16407 (N_16407,N_15939,N_15155);
or U16408 (N_16408,N_15885,N_14711);
nand U16409 (N_16409,N_15952,N_14375);
nand U16410 (N_16410,N_15223,N_14441);
nor U16411 (N_16411,N_14709,N_14954);
nor U16412 (N_16412,N_14162,N_15242);
or U16413 (N_16413,N_15927,N_14911);
and U16414 (N_16414,N_14659,N_14012);
nor U16415 (N_16415,N_14266,N_14663);
nand U16416 (N_16416,N_15061,N_15876);
nor U16417 (N_16417,N_15425,N_14209);
nand U16418 (N_16418,N_14525,N_15040);
nor U16419 (N_16419,N_15778,N_14367);
and U16420 (N_16420,N_14386,N_15326);
nor U16421 (N_16421,N_15800,N_14100);
or U16422 (N_16422,N_15035,N_14876);
and U16423 (N_16423,N_15141,N_14959);
or U16424 (N_16424,N_15154,N_14676);
xnor U16425 (N_16425,N_15641,N_14561);
nor U16426 (N_16426,N_14256,N_15482);
nand U16427 (N_16427,N_14873,N_15336);
nand U16428 (N_16428,N_15391,N_14894);
xor U16429 (N_16429,N_15948,N_15466);
nor U16430 (N_16430,N_14812,N_14176);
nand U16431 (N_16431,N_15751,N_15424);
nor U16432 (N_16432,N_15296,N_14897);
nor U16433 (N_16433,N_15473,N_15184);
nand U16434 (N_16434,N_15101,N_14278);
nand U16435 (N_16435,N_14996,N_15765);
and U16436 (N_16436,N_14890,N_15827);
xnor U16437 (N_16437,N_14791,N_14646);
and U16438 (N_16438,N_15539,N_15413);
or U16439 (N_16439,N_15545,N_14580);
nor U16440 (N_16440,N_15497,N_15407);
nor U16441 (N_16441,N_14092,N_15106);
or U16442 (N_16442,N_14174,N_15491);
nand U16443 (N_16443,N_15412,N_14602);
and U16444 (N_16444,N_14182,N_14010);
xor U16445 (N_16445,N_15071,N_15400);
nand U16446 (N_16446,N_15509,N_14321);
nand U16447 (N_16447,N_15022,N_14499);
nand U16448 (N_16448,N_15431,N_15646);
or U16449 (N_16449,N_14466,N_14708);
and U16450 (N_16450,N_15234,N_14047);
nand U16451 (N_16451,N_15472,N_14715);
or U16452 (N_16452,N_14087,N_15619);
and U16453 (N_16453,N_15975,N_14724);
or U16454 (N_16454,N_14113,N_14215);
nor U16455 (N_16455,N_14750,N_14311);
or U16456 (N_16456,N_14745,N_14758);
nand U16457 (N_16457,N_14282,N_15805);
nand U16458 (N_16458,N_15685,N_14856);
xnor U16459 (N_16459,N_15043,N_14016);
and U16460 (N_16460,N_14470,N_15078);
and U16461 (N_16461,N_14482,N_14193);
and U16462 (N_16462,N_14657,N_14648);
nand U16463 (N_16463,N_15481,N_14158);
nand U16464 (N_16464,N_15343,N_15979);
nor U16465 (N_16465,N_14171,N_14684);
nand U16466 (N_16466,N_14803,N_15133);
nand U16467 (N_16467,N_14569,N_14800);
and U16468 (N_16468,N_15528,N_14571);
and U16469 (N_16469,N_15742,N_15978);
nand U16470 (N_16470,N_15109,N_14970);
xnor U16471 (N_16471,N_15904,N_15031);
and U16472 (N_16472,N_15748,N_14727);
nand U16473 (N_16473,N_14998,N_15402);
or U16474 (N_16474,N_14857,N_14163);
nand U16475 (N_16475,N_14990,N_14585);
nand U16476 (N_16476,N_14319,N_14926);
nand U16477 (N_16477,N_15718,N_14677);
nand U16478 (N_16478,N_15693,N_15969);
or U16479 (N_16479,N_15232,N_14360);
or U16480 (N_16480,N_14397,N_14642);
nor U16481 (N_16481,N_14907,N_14479);
and U16482 (N_16482,N_14928,N_14444);
or U16483 (N_16483,N_14300,N_15408);
xnor U16484 (N_16484,N_14984,N_15686);
or U16485 (N_16485,N_14374,N_15996);
nand U16486 (N_16486,N_14389,N_14688);
nand U16487 (N_16487,N_15496,N_14641);
nor U16488 (N_16488,N_14686,N_14880);
nor U16489 (N_16489,N_15390,N_15418);
xnor U16490 (N_16490,N_15429,N_14925);
and U16491 (N_16491,N_15578,N_14971);
or U16492 (N_16492,N_15437,N_15788);
or U16493 (N_16493,N_14073,N_14330);
nand U16494 (N_16494,N_14771,N_14368);
and U16495 (N_16495,N_15771,N_15113);
or U16496 (N_16496,N_14008,N_14753);
or U16497 (N_16497,N_15789,N_15180);
and U16498 (N_16498,N_15583,N_14840);
and U16499 (N_16499,N_15127,N_15289);
nand U16500 (N_16500,N_14480,N_15776);
xnor U16501 (N_16501,N_14149,N_15156);
xor U16502 (N_16502,N_15537,N_15108);
and U16503 (N_16503,N_14738,N_15490);
xnor U16504 (N_16504,N_14025,N_15637);
nor U16505 (N_16505,N_14618,N_14636);
xor U16506 (N_16506,N_15636,N_15295);
nor U16507 (N_16507,N_14394,N_15291);
or U16508 (N_16508,N_15709,N_14868);
nand U16509 (N_16509,N_14964,N_15138);
and U16510 (N_16510,N_15427,N_14592);
xnor U16511 (N_16511,N_14052,N_14349);
or U16512 (N_16512,N_15199,N_14224);
nand U16513 (N_16513,N_14298,N_14471);
or U16514 (N_16514,N_15844,N_15803);
nand U16515 (N_16515,N_15604,N_14141);
and U16516 (N_16516,N_15062,N_14117);
or U16517 (N_16517,N_15450,N_15547);
or U16518 (N_16518,N_15600,N_15395);
or U16519 (N_16519,N_14744,N_15150);
or U16520 (N_16520,N_14225,N_14431);
nand U16521 (N_16521,N_14953,N_14314);
nor U16522 (N_16522,N_14913,N_14898);
nand U16523 (N_16523,N_14995,N_15311);
nand U16524 (N_16524,N_14043,N_14982);
nand U16525 (N_16525,N_14218,N_14142);
nor U16526 (N_16526,N_15585,N_15333);
xor U16527 (N_16527,N_15791,N_14463);
and U16528 (N_16528,N_15877,N_14054);
xnor U16529 (N_16529,N_15142,N_14255);
nand U16530 (N_16530,N_14757,N_15476);
nand U16531 (N_16531,N_14199,N_15880);
xor U16532 (N_16532,N_14032,N_14495);
and U16533 (N_16533,N_15531,N_15443);
or U16534 (N_16534,N_15669,N_15912);
or U16535 (N_16535,N_15714,N_14827);
nand U16536 (N_16536,N_14240,N_14320);
nor U16537 (N_16537,N_15264,N_14069);
or U16538 (N_16538,N_14846,N_14826);
and U16539 (N_16539,N_15614,N_14736);
nor U16540 (N_16540,N_15183,N_14268);
nand U16541 (N_16541,N_15544,N_15837);
or U16542 (N_16542,N_14578,N_14143);
nor U16543 (N_16543,N_15822,N_15977);
nand U16544 (N_16544,N_15734,N_15005);
nor U16545 (N_16545,N_14652,N_14883);
nor U16546 (N_16546,N_14582,N_15960);
and U16547 (N_16547,N_14770,N_15492);
nand U16548 (N_16548,N_15486,N_14358);
nor U16549 (N_16549,N_15323,N_15612);
and U16550 (N_16550,N_14056,N_14834);
or U16551 (N_16551,N_15416,N_14257);
nand U16552 (N_16552,N_14067,N_14598);
xor U16553 (N_16553,N_15869,N_15552);
and U16554 (N_16554,N_14454,N_15099);
nor U16555 (N_16555,N_14315,N_15406);
xor U16556 (N_16556,N_14409,N_14597);
and U16557 (N_16557,N_15642,N_14698);
and U16558 (N_16558,N_15974,N_15070);
and U16559 (N_16559,N_14327,N_15682);
nor U16560 (N_16560,N_14037,N_14194);
nand U16561 (N_16561,N_15831,N_14125);
nand U16562 (N_16562,N_14874,N_15093);
and U16563 (N_16563,N_14152,N_15247);
nor U16564 (N_16564,N_15047,N_15639);
nand U16565 (N_16565,N_14402,N_14427);
or U16566 (N_16566,N_14878,N_14144);
nand U16567 (N_16567,N_15772,N_15195);
nor U16568 (N_16568,N_15230,N_15766);
and U16569 (N_16569,N_15730,N_14104);
nand U16570 (N_16570,N_15203,N_15366);
or U16571 (N_16571,N_14208,N_15426);
or U16572 (N_16572,N_15917,N_15243);
xor U16573 (N_16573,N_14624,N_14476);
nand U16574 (N_16574,N_14396,N_14557);
or U16575 (N_16575,N_14497,N_15325);
and U16576 (N_16576,N_15369,N_14448);
nand U16577 (N_16577,N_14541,N_14051);
or U16578 (N_16578,N_14549,N_15522);
and U16579 (N_16579,N_14536,N_14210);
and U16580 (N_16580,N_15167,N_14206);
and U16581 (N_16581,N_14729,N_15258);
xnor U16582 (N_16582,N_14675,N_15344);
nand U16583 (N_16583,N_15673,N_15121);
or U16584 (N_16584,N_14356,N_15193);
or U16585 (N_16585,N_15009,N_14658);
or U16586 (N_16586,N_15237,N_14763);
nor U16587 (N_16587,N_14866,N_14369);
or U16588 (N_16588,N_14591,N_14969);
xnor U16589 (N_16589,N_14560,N_14259);
nand U16590 (N_16590,N_14346,N_15306);
xnor U16591 (N_16591,N_14899,N_15025);
or U16592 (N_16592,N_15801,N_15787);
nor U16593 (N_16593,N_15563,N_14473);
and U16594 (N_16594,N_15818,N_15020);
nor U16595 (N_16595,N_14186,N_14416);
and U16596 (N_16596,N_14983,N_15382);
and U16597 (N_16597,N_14967,N_15340);
nand U16598 (N_16598,N_14445,N_14599);
nand U16599 (N_16599,N_14399,N_15767);
and U16600 (N_16600,N_15864,N_15832);
nor U16601 (N_16601,N_15468,N_14609);
nand U16602 (N_16602,N_14048,N_14287);
or U16603 (N_16603,N_14912,N_14619);
or U16604 (N_16604,N_14929,N_15703);
or U16605 (N_16605,N_14714,N_15929);
nand U16606 (N_16606,N_14376,N_15675);
nor U16607 (N_16607,N_14558,N_15870);
and U16608 (N_16608,N_14777,N_15892);
or U16609 (N_16609,N_14279,N_15961);
nor U16610 (N_16610,N_15554,N_14417);
nand U16611 (N_16611,N_15098,N_15922);
nor U16612 (N_16612,N_15966,N_15036);
nor U16613 (N_16613,N_15784,N_14944);
nor U16614 (N_16614,N_15268,N_15658);
and U16615 (N_16615,N_14229,N_15004);
or U16616 (N_16616,N_15342,N_14824);
and U16617 (N_16617,N_15410,N_14449);
and U16618 (N_16618,N_15648,N_15894);
and U16619 (N_16619,N_14090,N_15001);
nor U16620 (N_16620,N_14496,N_14046);
nand U16621 (N_16621,N_15475,N_14844);
and U16622 (N_16622,N_15541,N_15452);
nor U16623 (N_16623,N_14946,N_14940);
and U16624 (N_16624,N_15016,N_15059);
nand U16625 (N_16625,N_14157,N_14870);
xnor U16626 (N_16626,N_14264,N_15663);
or U16627 (N_16627,N_15330,N_14691);
and U16628 (N_16628,N_14821,N_14030);
and U16629 (N_16629,N_14222,N_15119);
and U16630 (N_16630,N_15689,N_15697);
nor U16631 (N_16631,N_14674,N_14640);
nand U16632 (N_16632,N_15077,N_15645);
nand U16633 (N_16633,N_15495,N_15404);
nand U16634 (N_16634,N_14978,N_14075);
or U16635 (N_16635,N_15621,N_14882);
nand U16636 (N_16636,N_15916,N_14980);
nor U16637 (N_16637,N_15804,N_14900);
nand U16638 (N_16638,N_15245,N_14044);
and U16639 (N_16639,N_14461,N_15174);
nand U16640 (N_16640,N_15775,N_14213);
nand U16641 (N_16641,N_15128,N_15480);
and U16642 (N_16642,N_15786,N_15259);
xnor U16643 (N_16643,N_14121,N_14083);
nand U16644 (N_16644,N_14350,N_14139);
or U16645 (N_16645,N_14077,N_14084);
nand U16646 (N_16646,N_15023,N_15793);
and U16647 (N_16647,N_15735,N_15076);
nand U16648 (N_16648,N_14932,N_15851);
nand U16649 (N_16649,N_15676,N_15854);
nand U16650 (N_16650,N_14543,N_14029);
or U16651 (N_16651,N_14848,N_14258);
and U16652 (N_16652,N_14329,N_15897);
and U16653 (N_16653,N_15275,N_14660);
nor U16654 (N_16654,N_15126,N_14786);
nand U16655 (N_16655,N_14126,N_14347);
and U16656 (N_16656,N_14284,N_14060);
nand U16657 (N_16657,N_15750,N_14942);
or U16658 (N_16658,N_14304,N_14565);
nand U16659 (N_16659,N_15380,N_14373);
and U16660 (N_16660,N_14702,N_14159);
nand U16661 (N_16661,N_15954,N_14263);
or U16662 (N_16662,N_14387,N_15420);
nor U16663 (N_16663,N_14860,N_14761);
or U16664 (N_16664,N_14331,N_14131);
and U16665 (N_16665,N_14231,N_14902);
or U16666 (N_16666,N_15797,N_15886);
and U16667 (N_16667,N_14274,N_15957);
and U16668 (N_16668,N_15808,N_15445);
nor U16669 (N_16669,N_14015,N_14140);
nand U16670 (N_16670,N_15063,N_15840);
nor U16671 (N_16671,N_14751,N_15769);
and U16672 (N_16672,N_15172,N_15632);
and U16673 (N_16673,N_15988,N_15363);
nor U16674 (N_16674,N_15144,N_14586);
nand U16675 (N_16675,N_14027,N_15379);
or U16676 (N_16676,N_14041,N_14706);
and U16677 (N_16677,N_14548,N_14285);
or U16678 (N_16678,N_14556,N_15347);
nor U16679 (N_16679,N_15597,N_14798);
and U16680 (N_16680,N_14743,N_15560);
xnor U16681 (N_16681,N_14456,N_15082);
and U16682 (N_16682,N_15293,N_14919);
or U16683 (N_16683,N_14523,N_15026);
and U16684 (N_16684,N_15871,N_14338);
nor U16685 (N_16685,N_15622,N_15240);
or U16686 (N_16686,N_14594,N_14564);
or U16687 (N_16687,N_14128,N_15740);
nor U16688 (N_16688,N_14768,N_14917);
and U16689 (N_16689,N_14515,N_15388);
nand U16690 (N_16690,N_14244,N_14168);
and U16691 (N_16691,N_14522,N_14458);
nor U16692 (N_16692,N_14226,N_14958);
nor U16693 (N_16693,N_14535,N_14483);
xnor U16694 (N_16694,N_15860,N_15858);
nor U16695 (N_16695,N_15485,N_15359);
nand U16696 (N_16696,N_15694,N_14333);
and U16697 (N_16697,N_15835,N_14922);
and U16698 (N_16698,N_14239,N_14190);
nand U16699 (N_16699,N_14924,N_14401);
nand U16700 (N_16700,N_15944,N_15286);
or U16701 (N_16701,N_14614,N_14344);
nor U16702 (N_16702,N_15069,N_15517);
nand U16703 (N_16703,N_15630,N_15351);
xnor U16704 (N_16704,N_15919,N_14246);
nand U16705 (N_16705,N_15556,N_14687);
or U16706 (N_16706,N_15010,N_15120);
and U16707 (N_16707,N_14109,N_15605);
or U16708 (N_16708,N_15190,N_15744);
or U16709 (N_16709,N_15309,N_14673);
or U16710 (N_16710,N_14228,N_14071);
nand U16711 (N_16711,N_14165,N_15206);
and U16712 (N_16712,N_15692,N_14988);
or U16713 (N_16713,N_15507,N_14593);
nor U16714 (N_16714,N_15018,N_14986);
and U16715 (N_16715,N_14065,N_14507);
nand U16716 (N_16716,N_14596,N_15181);
xnor U16717 (N_16717,N_14459,N_15210);
nand U16718 (N_16718,N_14871,N_14039);
xnor U16719 (N_16719,N_15191,N_14404);
nand U16720 (N_16720,N_14280,N_14512);
or U16721 (N_16721,N_14392,N_15859);
and U16722 (N_16722,N_14184,N_14699);
or U16723 (N_16723,N_14575,N_15092);
xor U16724 (N_16724,N_15164,N_15724);
and U16725 (N_16725,N_14468,N_15118);
and U16726 (N_16726,N_14064,N_14503);
nor U16727 (N_16727,N_14498,N_14175);
and U16728 (N_16728,N_14138,N_15457);
or U16729 (N_16729,N_15266,N_15316);
and U16730 (N_16730,N_14423,N_14903);
or U16731 (N_16731,N_15770,N_14380);
nor U16732 (N_16732,N_15050,N_15700);
or U16733 (N_16733,N_15918,N_14265);
nand U16734 (N_16734,N_15440,N_15160);
or U16735 (N_16735,N_14689,N_14383);
and U16736 (N_16736,N_15205,N_15094);
and U16737 (N_16737,N_15157,N_14426);
and U16738 (N_16738,N_14260,N_15411);
or U16739 (N_16739,N_15525,N_15086);
and U16740 (N_16740,N_14275,N_15684);
nand U16741 (N_16741,N_14332,N_14214);
and U16742 (N_16742,N_15848,N_14410);
and U16743 (N_16743,N_14532,N_14359);
nand U16744 (N_16744,N_15386,N_15318);
and U16745 (N_16745,N_15135,N_15903);
or U16746 (N_16746,N_15590,N_15910);
xnor U16747 (N_16747,N_14154,N_15811);
nand U16748 (N_16748,N_15656,N_15826);
and U16749 (N_16749,N_14341,N_14991);
nor U16750 (N_16750,N_14737,N_14892);
nor U16751 (N_16751,N_14862,N_14908);
nand U16752 (N_16752,N_15212,N_14484);
nor U16753 (N_16753,N_14678,N_14865);
nand U16754 (N_16754,N_14628,N_14354);
and U16755 (N_16755,N_15893,N_15950);
nor U16756 (N_16756,N_15561,N_15332);
xnor U16757 (N_16757,N_15649,N_15899);
or U16758 (N_16758,N_14682,N_15401);
and U16759 (N_16759,N_15100,N_14788);
and U16760 (N_16760,N_14107,N_15304);
and U16761 (N_16761,N_15853,N_14309);
nand U16762 (N_16762,N_15946,N_14395);
nand U16763 (N_16763,N_14632,N_14033);
or U16764 (N_16764,N_15956,N_15219);
nand U16765 (N_16765,N_15229,N_14759);
or U16766 (N_16766,N_14783,N_15385);
nor U16767 (N_16767,N_15459,N_15665);
and U16768 (N_16768,N_15699,N_15890);
and U16769 (N_16769,N_15701,N_14955);
nand U16770 (N_16770,N_14683,N_15008);
xor U16771 (N_16771,N_14217,N_14403);
nand U16772 (N_16772,N_14835,N_15017);
nor U16773 (N_16773,N_14200,N_14667);
and U16774 (N_16774,N_15238,N_14173);
xor U16775 (N_16775,N_15231,N_14573);
and U16776 (N_16776,N_15189,N_15520);
nor U16777 (N_16777,N_14400,N_15595);
nor U16778 (N_16778,N_15550,N_14078);
nor U16779 (N_16779,N_15741,N_15361);
nand U16780 (N_16780,N_14544,N_14272);
nand U16781 (N_16781,N_15064,N_15239);
xor U16782 (N_16782,N_14581,N_14412);
nor U16783 (N_16783,N_15807,N_14502);
or U16784 (N_16784,N_15839,N_15618);
and U16785 (N_16785,N_14059,N_14120);
nor U16786 (N_16786,N_14323,N_15117);
and U16787 (N_16787,N_15310,N_14068);
or U16788 (N_16788,N_14822,N_14096);
xor U16789 (N_16789,N_14809,N_15883);
nor U16790 (N_16790,N_15635,N_15691);
nor U16791 (N_16791,N_15780,N_14453);
and U16792 (N_16792,N_14623,N_14452);
nand U16793 (N_16793,N_14773,N_14644);
nand U16794 (N_16794,N_15349,N_15938);
nand U16795 (N_16795,N_15123,N_14616);
or U16796 (N_16796,N_15003,N_14203);
and U16797 (N_16797,N_14723,N_15305);
xnor U16798 (N_16798,N_15455,N_14160);
and U16799 (N_16799,N_14219,N_15415);
and U16800 (N_16800,N_15634,N_15102);
nand U16801 (N_16801,N_15246,N_14920);
nand U16802 (N_16802,N_14707,N_14740);
or U16803 (N_16803,N_15755,N_15761);
xor U16804 (N_16804,N_15327,N_14752);
or U16805 (N_16805,N_14861,N_14429);
nand U16806 (N_16806,N_14018,N_14792);
nand U16807 (N_16807,N_15348,N_15981);
nand U16808 (N_16808,N_14661,N_14818);
or U16809 (N_16809,N_15072,N_14611);
and U16810 (N_16810,N_15866,N_15302);
nor U16811 (N_16811,N_14189,N_15968);
and U16812 (N_16812,N_14960,N_15096);
xor U16813 (N_16813,N_14884,N_15781);
nand U16814 (N_16814,N_15959,N_15706);
or U16815 (N_16815,N_14952,N_15464);
or U16816 (N_16816,N_14207,N_15281);
nand U16817 (N_16817,N_14713,N_14187);
or U16818 (N_16818,N_15414,N_15934);
xnor U16819 (N_16819,N_14475,N_15898);
and U16820 (N_16820,N_14696,N_15723);
and U16821 (N_16821,N_15085,N_15271);
nand U16822 (N_16822,N_14504,N_15249);
nand U16823 (N_16823,N_14312,N_15720);
or U16824 (N_16824,N_15014,N_15654);
or U16825 (N_16825,N_14509,N_14434);
nor U16826 (N_16826,N_15999,N_15519);
nand U16827 (N_16827,N_14831,N_14606);
nand U16828 (N_16828,N_14146,N_14003);
or U16829 (N_16829,N_14430,N_15815);
or U16830 (N_16830,N_15364,N_15091);
nand U16831 (N_16831,N_15733,N_15278);
or U16832 (N_16832,N_14653,N_15132);
or U16833 (N_16833,N_14232,N_14563);
xnor U16834 (N_16834,N_15034,N_15989);
nand U16835 (N_16835,N_14772,N_14893);
nand U16836 (N_16836,N_14001,N_14719);
xnor U16837 (N_16837,N_14220,N_15087);
nand U16838 (N_16838,N_14201,N_15503);
nand U16839 (N_16839,N_14317,N_15192);
or U16840 (N_16840,N_15290,N_14979);
or U16841 (N_16841,N_15454,N_14785);
or U16842 (N_16842,N_15422,N_14303);
nor U16843 (N_16843,N_14058,N_14807);
nor U16844 (N_16844,N_15928,N_14590);
nand U16845 (N_16845,N_15963,N_15762);
and U16846 (N_16846,N_14435,N_15588);
and U16847 (N_16847,N_14610,N_15970);
nor U16848 (N_16848,N_15270,N_14170);
and U16849 (N_16849,N_15940,N_15263);
and U16850 (N_16850,N_15057,N_15012);
nor U16851 (N_16851,N_15498,N_14651);
and U16852 (N_16852,N_15256,N_15712);
nor U16853 (N_16853,N_15028,N_15644);
or U16854 (N_16854,N_15499,N_15945);
nor U16855 (N_16855,N_15678,N_15356);
or U16856 (N_16856,N_15696,N_14181);
or U16857 (N_16857,N_15620,N_14178);
and U16858 (N_16858,N_14388,N_15602);
nor U16859 (N_16859,N_15217,N_15824);
nand U16860 (N_16860,N_15073,N_15131);
and U16861 (N_16861,N_15677,N_14486);
nand U16862 (N_16862,N_15878,N_14776);
nand U16863 (N_16863,N_14805,N_15056);
or U16864 (N_16864,N_14742,N_15145);
or U16865 (N_16865,N_15255,N_14973);
nand U16866 (N_16866,N_14842,N_15739);
and U16867 (N_16867,N_15941,N_15381);
and U16868 (N_16868,N_15725,N_15208);
or U16869 (N_16869,N_15967,N_14943);
xor U16870 (N_16870,N_14494,N_15104);
nand U16871 (N_16871,N_15812,N_15228);
or U16872 (N_16872,N_15149,N_15169);
nor U16873 (N_16873,N_14832,N_15779);
and U16874 (N_16874,N_14746,N_15882);
and U16875 (N_16875,N_15707,N_15147);
nor U16876 (N_16876,N_14669,N_14849);
or U16877 (N_16877,N_15188,N_15958);
nor U16878 (N_16878,N_15704,N_14437);
or U16879 (N_16879,N_15315,N_15165);
or U16880 (N_16880,N_14962,N_15162);
nand U16881 (N_16881,N_15737,N_15756);
nand U16882 (N_16882,N_15024,N_14595);
and U16883 (N_16883,N_15053,N_15606);
and U16884 (N_16884,N_15817,N_15628);
and U16885 (N_16885,N_14197,N_15002);
and U16886 (N_16886,N_14810,N_15173);
or U16887 (N_16887,N_15260,N_15608);
nor U16888 (N_16888,N_15653,N_14589);
and U16889 (N_16889,N_15110,N_14337);
or U16890 (N_16890,N_14013,N_15562);
nand U16891 (N_16891,N_15171,N_15213);
or U16892 (N_16892,N_15863,N_14236);
nor U16893 (N_16893,N_14670,N_15430);
and U16894 (N_16894,N_15861,N_15698);
and U16895 (N_16895,N_14951,N_14086);
nand U16896 (N_16896,N_14814,N_15148);
nand U16897 (N_16897,N_14790,N_15322);
or U16898 (N_16898,N_15097,N_15303);
nor U16899 (N_16899,N_14072,N_14478);
nand U16900 (N_16900,N_14637,N_14413);
nor U16901 (N_16901,N_15587,N_15376);
nand U16902 (N_16902,N_15112,N_14697);
or U16903 (N_16903,N_15368,N_15449);
nor U16904 (N_16904,N_15688,N_15931);
nand U16905 (N_16905,N_14390,N_15841);
or U16906 (N_16906,N_15299,N_14877);
nor U16907 (N_16907,N_14366,N_14508);
nor U16908 (N_16908,N_15868,N_14105);
nor U16909 (N_16909,N_14488,N_14050);
or U16910 (N_16910,N_14966,N_15448);
and U16911 (N_16911,N_14662,N_14690);
xor U16912 (N_16912,N_14301,N_15200);
or U16913 (N_16913,N_15949,N_14085);
nor U16914 (N_16914,N_15849,N_14855);
and U16915 (N_16915,N_14650,N_14308);
or U16916 (N_16916,N_15433,N_15976);
xnor U16917 (N_16917,N_14680,N_14447);
nand U16918 (N_16918,N_14061,N_15370);
nand U16919 (N_16919,N_14858,N_14363);
nor U16920 (N_16920,N_14735,N_14491);
and U16921 (N_16921,N_14538,N_15951);
nor U16922 (N_16922,N_15623,N_14161);
xor U16923 (N_16923,N_15715,N_14132);
nand U16924 (N_16924,N_14172,N_15083);
and U16925 (N_16925,N_15717,N_15350);
xnor U16926 (N_16926,N_15090,N_15107);
nand U16927 (N_16927,N_15806,N_14607);
and U16928 (N_16928,N_14748,N_14720);
and U16929 (N_16929,N_15116,N_15909);
nor U16930 (N_16930,N_15250,N_15668);
and U16931 (N_16931,N_15936,N_14147);
and U16932 (N_16932,N_15257,N_15479);
xor U16933 (N_16933,N_14183,N_14267);
and U16934 (N_16934,N_15394,N_15037);
nand U16935 (N_16935,N_14718,N_15177);
nand U16936 (N_16936,N_14645,N_15813);
nor U16937 (N_16937,N_14053,N_15282);
or U16938 (N_16938,N_15421,N_15515);
and U16939 (N_16939,N_14335,N_15197);
or U16940 (N_16940,N_14906,N_14119);
nor U16941 (N_16941,N_14505,N_14612);
nor U16942 (N_16942,N_15670,N_15971);
and U16943 (N_16943,N_15060,N_14305);
nand U16944 (N_16944,N_15353,N_15095);
and U16945 (N_16945,N_15300,N_14196);
and U16946 (N_16946,N_15570,N_15985);
and U16947 (N_16947,N_15185,N_15915);
and U16948 (N_16948,N_14778,N_14825);
xor U16949 (N_16949,N_14000,N_14385);
nor U16950 (N_16950,N_15997,N_15226);
or U16951 (N_16951,N_14289,N_15292);
or U16952 (N_16952,N_14992,N_14151);
and U16953 (N_16953,N_14472,N_15843);
nor U16954 (N_16954,N_15830,N_15283);
and U16955 (N_16955,N_15033,N_14425);
nand U16956 (N_16956,N_15705,N_14123);
nand U16957 (N_16957,N_15566,N_15962);
nor U16958 (N_16958,N_14765,N_14328);
and U16959 (N_16959,N_15551,N_15146);
or U16960 (N_16960,N_15582,N_15785);
nor U16961 (N_16961,N_15777,N_14613);
and U16962 (N_16962,N_14854,N_15313);
or U16963 (N_16963,N_15178,N_14916);
or U16964 (N_16964,N_14915,N_14732);
nor U16965 (N_16965,N_15716,N_15521);
nor U16966 (N_16966,N_14513,N_14529);
nor U16967 (N_16967,N_15819,N_14336);
xor U16968 (N_16968,N_14156,N_15731);
and U16969 (N_16969,N_15640,N_14477);
and U16970 (N_16970,N_15393,N_15708);
and U16971 (N_16971,N_15066,N_15887);
nand U16972 (N_16972,N_14555,N_15925);
xor U16973 (N_16973,N_14021,N_15662);
and U16974 (N_16974,N_14227,N_14393);
nand U16975 (N_16975,N_14180,N_15625);
or U16976 (N_16976,N_15923,N_15114);
or U16977 (N_16977,N_15680,N_15745);
or U16978 (N_16978,N_14837,N_15660);
and U16979 (N_16979,N_15216,N_14518);
and U16980 (N_16980,N_15447,N_14133);
or U16981 (N_16981,N_15536,N_14411);
xor U16982 (N_16982,N_14802,N_14269);
and U16983 (N_16983,N_14034,N_14796);
xnor U16984 (N_16984,N_14024,N_15638);
or U16985 (N_16985,N_15505,N_14694);
nand U16986 (N_16986,N_15153,N_14361);
xnor U16987 (N_16987,N_15168,N_15617);
xnor U16988 (N_16988,N_15362,N_15555);
nand U16989 (N_16989,N_14191,N_14703);
xnor U16990 (N_16990,N_14634,N_14766);
and U16991 (N_16991,N_15030,N_15338);
nand U16992 (N_16992,N_14216,N_14521);
or U16993 (N_16993,N_15487,N_15319);
nor U16994 (N_16994,N_15847,N_14989);
nor U16995 (N_16995,N_14166,N_14089);
xnor U16996 (N_16996,N_14817,N_15672);
and U16997 (N_16997,N_14420,N_15538);
nand U16998 (N_16998,N_15384,N_15749);
nand U16999 (N_16999,N_14957,N_15829);
nand U17000 (N_17000,N_15642,N_15001);
or U17001 (N_17001,N_15953,N_15093);
nand U17002 (N_17002,N_14562,N_14613);
xnor U17003 (N_17003,N_15684,N_14866);
xor U17004 (N_17004,N_15686,N_15323);
and U17005 (N_17005,N_14647,N_14261);
and U17006 (N_17006,N_14779,N_14195);
or U17007 (N_17007,N_15040,N_15729);
and U17008 (N_17008,N_14903,N_15767);
or U17009 (N_17009,N_14407,N_14818);
nor U17010 (N_17010,N_15955,N_14818);
or U17011 (N_17011,N_14293,N_15023);
or U17012 (N_17012,N_14167,N_14237);
nor U17013 (N_17013,N_15916,N_15310);
or U17014 (N_17014,N_15026,N_15110);
nor U17015 (N_17015,N_15235,N_14657);
xnor U17016 (N_17016,N_14690,N_14821);
nor U17017 (N_17017,N_14208,N_15133);
and U17018 (N_17018,N_15029,N_15237);
nor U17019 (N_17019,N_15013,N_15461);
and U17020 (N_17020,N_14280,N_14316);
or U17021 (N_17021,N_14621,N_14355);
or U17022 (N_17022,N_14330,N_15944);
nor U17023 (N_17023,N_14392,N_14262);
and U17024 (N_17024,N_15513,N_14419);
or U17025 (N_17025,N_14235,N_15171);
or U17026 (N_17026,N_14128,N_15172);
and U17027 (N_17027,N_14676,N_14583);
or U17028 (N_17028,N_14427,N_15578);
nand U17029 (N_17029,N_14503,N_15269);
nor U17030 (N_17030,N_14203,N_15727);
or U17031 (N_17031,N_14057,N_15332);
and U17032 (N_17032,N_14273,N_15698);
nand U17033 (N_17033,N_14538,N_15226);
and U17034 (N_17034,N_15741,N_15870);
xor U17035 (N_17035,N_15801,N_15563);
or U17036 (N_17036,N_14773,N_14755);
nand U17037 (N_17037,N_14549,N_14970);
xnor U17038 (N_17038,N_15440,N_14355);
nand U17039 (N_17039,N_15404,N_14022);
nor U17040 (N_17040,N_15849,N_14992);
and U17041 (N_17041,N_14650,N_14478);
or U17042 (N_17042,N_14920,N_15400);
or U17043 (N_17043,N_14532,N_15101);
xor U17044 (N_17044,N_14072,N_15175);
nor U17045 (N_17045,N_14672,N_15605);
or U17046 (N_17046,N_15947,N_15877);
nand U17047 (N_17047,N_15813,N_15484);
nand U17048 (N_17048,N_15644,N_14976);
and U17049 (N_17049,N_15483,N_14942);
or U17050 (N_17050,N_15840,N_15980);
and U17051 (N_17051,N_14145,N_15619);
nand U17052 (N_17052,N_14333,N_14978);
nor U17053 (N_17053,N_14673,N_14111);
or U17054 (N_17054,N_15312,N_14818);
xnor U17055 (N_17055,N_14769,N_15508);
or U17056 (N_17056,N_15471,N_15265);
nor U17057 (N_17057,N_14787,N_15410);
xnor U17058 (N_17058,N_15033,N_14498);
nor U17059 (N_17059,N_14062,N_14303);
nand U17060 (N_17060,N_14147,N_14210);
nor U17061 (N_17061,N_15591,N_15154);
nor U17062 (N_17062,N_15518,N_14109);
xor U17063 (N_17063,N_15763,N_15536);
or U17064 (N_17064,N_14017,N_14678);
xor U17065 (N_17065,N_15482,N_15466);
or U17066 (N_17066,N_14277,N_14041);
nor U17067 (N_17067,N_15444,N_14139);
nand U17068 (N_17068,N_15093,N_14628);
nor U17069 (N_17069,N_15919,N_15565);
nor U17070 (N_17070,N_14481,N_15075);
and U17071 (N_17071,N_14871,N_14040);
nor U17072 (N_17072,N_14045,N_15802);
nor U17073 (N_17073,N_14300,N_14246);
or U17074 (N_17074,N_15833,N_15158);
or U17075 (N_17075,N_14240,N_15819);
or U17076 (N_17076,N_14793,N_15837);
and U17077 (N_17077,N_14733,N_14504);
nor U17078 (N_17078,N_15699,N_15371);
nor U17079 (N_17079,N_15224,N_14107);
nand U17080 (N_17080,N_14810,N_14540);
nand U17081 (N_17081,N_15291,N_15100);
and U17082 (N_17082,N_14906,N_15110);
and U17083 (N_17083,N_14658,N_15629);
or U17084 (N_17084,N_15989,N_15151);
nand U17085 (N_17085,N_15053,N_14035);
or U17086 (N_17086,N_15095,N_15629);
xor U17087 (N_17087,N_14168,N_15299);
nand U17088 (N_17088,N_14742,N_14566);
and U17089 (N_17089,N_14545,N_15205);
and U17090 (N_17090,N_15704,N_14313);
and U17091 (N_17091,N_14793,N_14674);
or U17092 (N_17092,N_15854,N_15836);
xor U17093 (N_17093,N_15048,N_15595);
nor U17094 (N_17094,N_15552,N_15338);
nand U17095 (N_17095,N_15701,N_15409);
nand U17096 (N_17096,N_15618,N_15123);
nand U17097 (N_17097,N_15523,N_14317);
nor U17098 (N_17098,N_15837,N_15182);
nor U17099 (N_17099,N_15054,N_14599);
and U17100 (N_17100,N_14644,N_15978);
or U17101 (N_17101,N_15648,N_14182);
or U17102 (N_17102,N_15397,N_15470);
or U17103 (N_17103,N_14812,N_14576);
nand U17104 (N_17104,N_14680,N_14454);
and U17105 (N_17105,N_15141,N_15212);
or U17106 (N_17106,N_14390,N_14350);
nor U17107 (N_17107,N_15701,N_15510);
nand U17108 (N_17108,N_14430,N_14823);
nor U17109 (N_17109,N_14745,N_14828);
or U17110 (N_17110,N_15464,N_15063);
nor U17111 (N_17111,N_15728,N_15601);
nor U17112 (N_17112,N_14770,N_14795);
and U17113 (N_17113,N_15431,N_15212);
and U17114 (N_17114,N_15894,N_14105);
nand U17115 (N_17115,N_14031,N_15282);
and U17116 (N_17116,N_14551,N_14360);
or U17117 (N_17117,N_14485,N_14921);
and U17118 (N_17118,N_14509,N_15623);
nand U17119 (N_17119,N_15185,N_15348);
nor U17120 (N_17120,N_15430,N_15378);
and U17121 (N_17121,N_14796,N_15845);
and U17122 (N_17122,N_14246,N_15832);
or U17123 (N_17123,N_14841,N_15703);
or U17124 (N_17124,N_14467,N_15008);
or U17125 (N_17125,N_15113,N_15041);
nor U17126 (N_17126,N_14751,N_15451);
nor U17127 (N_17127,N_14775,N_14635);
nor U17128 (N_17128,N_15010,N_14865);
and U17129 (N_17129,N_14830,N_14150);
nor U17130 (N_17130,N_15669,N_15871);
nor U17131 (N_17131,N_14375,N_15011);
nor U17132 (N_17132,N_14951,N_15350);
and U17133 (N_17133,N_15544,N_14880);
or U17134 (N_17134,N_15071,N_15074);
or U17135 (N_17135,N_15280,N_14041);
nand U17136 (N_17136,N_15830,N_15226);
nor U17137 (N_17137,N_14084,N_15232);
nand U17138 (N_17138,N_15232,N_14722);
or U17139 (N_17139,N_15243,N_14725);
and U17140 (N_17140,N_14999,N_14107);
nor U17141 (N_17141,N_15993,N_14458);
or U17142 (N_17142,N_14261,N_14663);
or U17143 (N_17143,N_14619,N_15299);
or U17144 (N_17144,N_15470,N_15945);
and U17145 (N_17145,N_14174,N_14748);
nor U17146 (N_17146,N_14872,N_14200);
nor U17147 (N_17147,N_14166,N_14552);
nand U17148 (N_17148,N_15735,N_14186);
nand U17149 (N_17149,N_14066,N_15837);
or U17150 (N_17150,N_15839,N_14197);
xor U17151 (N_17151,N_15072,N_15922);
or U17152 (N_17152,N_14335,N_14995);
and U17153 (N_17153,N_15256,N_14878);
nand U17154 (N_17154,N_15883,N_15793);
and U17155 (N_17155,N_14910,N_15331);
or U17156 (N_17156,N_14342,N_15104);
nand U17157 (N_17157,N_14586,N_14529);
or U17158 (N_17158,N_15369,N_15802);
nor U17159 (N_17159,N_15593,N_15701);
and U17160 (N_17160,N_14303,N_14560);
nor U17161 (N_17161,N_15561,N_14586);
or U17162 (N_17162,N_15910,N_15955);
nand U17163 (N_17163,N_14410,N_14031);
or U17164 (N_17164,N_14901,N_14164);
nand U17165 (N_17165,N_14792,N_15332);
nand U17166 (N_17166,N_14218,N_14854);
nand U17167 (N_17167,N_14798,N_15799);
nand U17168 (N_17168,N_14167,N_14084);
xor U17169 (N_17169,N_14293,N_15232);
and U17170 (N_17170,N_15775,N_14616);
nand U17171 (N_17171,N_15008,N_15802);
nand U17172 (N_17172,N_15915,N_15516);
nor U17173 (N_17173,N_15186,N_14680);
and U17174 (N_17174,N_15694,N_14117);
xnor U17175 (N_17175,N_14563,N_15134);
and U17176 (N_17176,N_14668,N_14446);
or U17177 (N_17177,N_14759,N_15645);
nor U17178 (N_17178,N_15184,N_14152);
and U17179 (N_17179,N_15989,N_14356);
nand U17180 (N_17180,N_14548,N_15580);
nor U17181 (N_17181,N_14468,N_14051);
and U17182 (N_17182,N_15014,N_15751);
and U17183 (N_17183,N_14966,N_14827);
nand U17184 (N_17184,N_14952,N_14366);
and U17185 (N_17185,N_14419,N_14836);
and U17186 (N_17186,N_14572,N_14581);
nor U17187 (N_17187,N_14792,N_15796);
or U17188 (N_17188,N_14068,N_14940);
nand U17189 (N_17189,N_14174,N_14129);
or U17190 (N_17190,N_14137,N_15218);
and U17191 (N_17191,N_15664,N_15314);
nand U17192 (N_17192,N_15805,N_15417);
or U17193 (N_17193,N_14695,N_15345);
and U17194 (N_17194,N_15649,N_14496);
nor U17195 (N_17195,N_15126,N_14703);
and U17196 (N_17196,N_15387,N_15434);
nand U17197 (N_17197,N_14114,N_14878);
nand U17198 (N_17198,N_15036,N_14834);
and U17199 (N_17199,N_15309,N_14895);
or U17200 (N_17200,N_14023,N_15792);
nor U17201 (N_17201,N_14815,N_15005);
or U17202 (N_17202,N_14860,N_15082);
nor U17203 (N_17203,N_15418,N_14017);
nor U17204 (N_17204,N_15923,N_14708);
xnor U17205 (N_17205,N_14904,N_14052);
nand U17206 (N_17206,N_15412,N_15081);
nand U17207 (N_17207,N_15212,N_15069);
nor U17208 (N_17208,N_15554,N_14510);
xnor U17209 (N_17209,N_15065,N_15557);
and U17210 (N_17210,N_14610,N_15589);
and U17211 (N_17211,N_14931,N_14773);
xor U17212 (N_17212,N_14552,N_15289);
nand U17213 (N_17213,N_14324,N_14002);
nor U17214 (N_17214,N_14702,N_15865);
nor U17215 (N_17215,N_14113,N_14135);
nor U17216 (N_17216,N_14343,N_15539);
nor U17217 (N_17217,N_15582,N_14379);
nand U17218 (N_17218,N_15392,N_15742);
or U17219 (N_17219,N_15338,N_15187);
xor U17220 (N_17220,N_14126,N_15688);
xnor U17221 (N_17221,N_14597,N_14251);
nand U17222 (N_17222,N_15426,N_15065);
or U17223 (N_17223,N_14863,N_14908);
nor U17224 (N_17224,N_14697,N_14252);
nand U17225 (N_17225,N_15051,N_15270);
and U17226 (N_17226,N_14392,N_14609);
xor U17227 (N_17227,N_15319,N_15743);
and U17228 (N_17228,N_14208,N_14724);
nor U17229 (N_17229,N_15467,N_15870);
and U17230 (N_17230,N_15133,N_14242);
and U17231 (N_17231,N_14701,N_14139);
nor U17232 (N_17232,N_14614,N_14781);
and U17233 (N_17233,N_15893,N_14639);
and U17234 (N_17234,N_15297,N_14671);
or U17235 (N_17235,N_15983,N_14406);
nor U17236 (N_17236,N_15284,N_15892);
and U17237 (N_17237,N_14468,N_15191);
nand U17238 (N_17238,N_15986,N_15650);
and U17239 (N_17239,N_15059,N_14145);
and U17240 (N_17240,N_15947,N_15857);
nor U17241 (N_17241,N_15570,N_14428);
xnor U17242 (N_17242,N_14541,N_14535);
nor U17243 (N_17243,N_14610,N_15806);
xnor U17244 (N_17244,N_15499,N_15339);
and U17245 (N_17245,N_14689,N_15020);
nand U17246 (N_17246,N_14169,N_14231);
and U17247 (N_17247,N_15594,N_14412);
nor U17248 (N_17248,N_14246,N_15096);
or U17249 (N_17249,N_14324,N_14941);
and U17250 (N_17250,N_15543,N_15820);
and U17251 (N_17251,N_15324,N_15110);
nor U17252 (N_17252,N_15358,N_14454);
nor U17253 (N_17253,N_15123,N_15350);
or U17254 (N_17254,N_15943,N_15128);
or U17255 (N_17255,N_14313,N_14195);
nor U17256 (N_17256,N_15604,N_14864);
or U17257 (N_17257,N_14332,N_15013);
nand U17258 (N_17258,N_14522,N_14778);
nand U17259 (N_17259,N_15046,N_14759);
nor U17260 (N_17260,N_14696,N_15244);
and U17261 (N_17261,N_14727,N_15313);
and U17262 (N_17262,N_14640,N_14605);
nand U17263 (N_17263,N_15502,N_14886);
nor U17264 (N_17264,N_15025,N_14253);
or U17265 (N_17265,N_15247,N_14930);
and U17266 (N_17266,N_15697,N_15768);
nor U17267 (N_17267,N_14039,N_15730);
nor U17268 (N_17268,N_15891,N_14042);
xor U17269 (N_17269,N_15098,N_15254);
nor U17270 (N_17270,N_14913,N_15136);
nor U17271 (N_17271,N_15054,N_14409);
xnor U17272 (N_17272,N_15398,N_14182);
and U17273 (N_17273,N_15104,N_14924);
nor U17274 (N_17274,N_14890,N_15778);
nand U17275 (N_17275,N_14142,N_14298);
nor U17276 (N_17276,N_15555,N_14231);
or U17277 (N_17277,N_14332,N_15223);
or U17278 (N_17278,N_14954,N_14172);
or U17279 (N_17279,N_14836,N_14443);
or U17280 (N_17280,N_14847,N_14930);
nand U17281 (N_17281,N_14860,N_14746);
and U17282 (N_17282,N_15408,N_14314);
or U17283 (N_17283,N_14864,N_14364);
or U17284 (N_17284,N_15523,N_14895);
or U17285 (N_17285,N_15142,N_14950);
nor U17286 (N_17286,N_14998,N_14123);
xor U17287 (N_17287,N_15651,N_14170);
nand U17288 (N_17288,N_14184,N_14394);
or U17289 (N_17289,N_15834,N_14414);
and U17290 (N_17290,N_15919,N_15968);
and U17291 (N_17291,N_15180,N_14807);
nor U17292 (N_17292,N_14507,N_14785);
nand U17293 (N_17293,N_14603,N_15985);
nor U17294 (N_17294,N_15494,N_15254);
nor U17295 (N_17295,N_14062,N_14603);
nand U17296 (N_17296,N_15716,N_14363);
or U17297 (N_17297,N_15847,N_14710);
or U17298 (N_17298,N_14831,N_14829);
or U17299 (N_17299,N_15142,N_14513);
and U17300 (N_17300,N_15300,N_14784);
nand U17301 (N_17301,N_15798,N_15747);
xnor U17302 (N_17302,N_14731,N_15298);
nand U17303 (N_17303,N_14032,N_14111);
and U17304 (N_17304,N_14435,N_15265);
nor U17305 (N_17305,N_14678,N_15454);
nand U17306 (N_17306,N_14765,N_14757);
and U17307 (N_17307,N_15700,N_15745);
nor U17308 (N_17308,N_14634,N_14426);
nor U17309 (N_17309,N_15047,N_14392);
and U17310 (N_17310,N_15164,N_14930);
or U17311 (N_17311,N_15028,N_15553);
nor U17312 (N_17312,N_14775,N_14981);
nor U17313 (N_17313,N_14390,N_14154);
nor U17314 (N_17314,N_14941,N_15803);
xor U17315 (N_17315,N_14828,N_14341);
nand U17316 (N_17316,N_15835,N_14860);
nor U17317 (N_17317,N_14906,N_14347);
or U17318 (N_17318,N_15708,N_14948);
or U17319 (N_17319,N_15523,N_15520);
nor U17320 (N_17320,N_14108,N_15932);
nor U17321 (N_17321,N_15980,N_14705);
xor U17322 (N_17322,N_14508,N_15636);
or U17323 (N_17323,N_14216,N_14352);
or U17324 (N_17324,N_15988,N_14095);
nor U17325 (N_17325,N_15680,N_15917);
nand U17326 (N_17326,N_15493,N_14216);
and U17327 (N_17327,N_15035,N_15141);
and U17328 (N_17328,N_15055,N_15870);
or U17329 (N_17329,N_14468,N_15363);
nor U17330 (N_17330,N_14964,N_14949);
nand U17331 (N_17331,N_14990,N_15412);
nor U17332 (N_17332,N_15496,N_14690);
xnor U17333 (N_17333,N_14513,N_15650);
and U17334 (N_17334,N_15205,N_15861);
or U17335 (N_17335,N_15872,N_14522);
nand U17336 (N_17336,N_14018,N_14563);
nor U17337 (N_17337,N_14631,N_14352);
and U17338 (N_17338,N_15712,N_15610);
nor U17339 (N_17339,N_14265,N_15398);
or U17340 (N_17340,N_15254,N_14811);
nor U17341 (N_17341,N_15749,N_14632);
nor U17342 (N_17342,N_14313,N_15223);
or U17343 (N_17343,N_15755,N_14063);
nand U17344 (N_17344,N_15340,N_15251);
or U17345 (N_17345,N_15027,N_15504);
or U17346 (N_17346,N_14095,N_15989);
nor U17347 (N_17347,N_14493,N_14958);
or U17348 (N_17348,N_14156,N_14044);
or U17349 (N_17349,N_14695,N_14082);
or U17350 (N_17350,N_14338,N_15531);
nor U17351 (N_17351,N_14175,N_14107);
nor U17352 (N_17352,N_15898,N_15706);
or U17353 (N_17353,N_14699,N_15294);
nor U17354 (N_17354,N_14275,N_15217);
nor U17355 (N_17355,N_14327,N_15320);
or U17356 (N_17356,N_14216,N_15571);
nand U17357 (N_17357,N_15959,N_15956);
nand U17358 (N_17358,N_14747,N_14923);
xnor U17359 (N_17359,N_14695,N_14377);
nand U17360 (N_17360,N_15721,N_15083);
nand U17361 (N_17361,N_14112,N_15604);
or U17362 (N_17362,N_15900,N_14539);
and U17363 (N_17363,N_14422,N_15099);
nor U17364 (N_17364,N_15448,N_14730);
nor U17365 (N_17365,N_15087,N_15119);
xnor U17366 (N_17366,N_15806,N_15566);
xor U17367 (N_17367,N_15224,N_14209);
nand U17368 (N_17368,N_14353,N_14244);
nor U17369 (N_17369,N_14157,N_14499);
xnor U17370 (N_17370,N_14111,N_15158);
nor U17371 (N_17371,N_14114,N_15647);
nor U17372 (N_17372,N_14860,N_14462);
nand U17373 (N_17373,N_14529,N_14077);
xor U17374 (N_17374,N_15711,N_15398);
and U17375 (N_17375,N_15120,N_14760);
nor U17376 (N_17376,N_14740,N_15263);
or U17377 (N_17377,N_14053,N_15526);
or U17378 (N_17378,N_14871,N_14977);
or U17379 (N_17379,N_15053,N_14692);
and U17380 (N_17380,N_15970,N_14880);
nand U17381 (N_17381,N_15261,N_15695);
nor U17382 (N_17382,N_15162,N_14744);
nand U17383 (N_17383,N_15409,N_14024);
nand U17384 (N_17384,N_15768,N_15535);
nand U17385 (N_17385,N_15140,N_15725);
nor U17386 (N_17386,N_14752,N_14946);
nand U17387 (N_17387,N_14252,N_15344);
nand U17388 (N_17388,N_15758,N_15598);
nand U17389 (N_17389,N_15453,N_15169);
nand U17390 (N_17390,N_15639,N_15553);
nor U17391 (N_17391,N_14599,N_15355);
nand U17392 (N_17392,N_14385,N_15326);
or U17393 (N_17393,N_15810,N_15587);
or U17394 (N_17394,N_15326,N_15243);
and U17395 (N_17395,N_14164,N_14689);
nand U17396 (N_17396,N_14314,N_14704);
or U17397 (N_17397,N_14211,N_14273);
nor U17398 (N_17398,N_15225,N_14152);
and U17399 (N_17399,N_14112,N_14843);
nor U17400 (N_17400,N_14847,N_15147);
or U17401 (N_17401,N_15429,N_14555);
nor U17402 (N_17402,N_14121,N_15418);
nand U17403 (N_17403,N_14978,N_14072);
nor U17404 (N_17404,N_14230,N_15204);
and U17405 (N_17405,N_15861,N_14935);
or U17406 (N_17406,N_15444,N_15100);
nand U17407 (N_17407,N_15361,N_15658);
xor U17408 (N_17408,N_14523,N_15978);
or U17409 (N_17409,N_15385,N_14824);
or U17410 (N_17410,N_15904,N_14319);
and U17411 (N_17411,N_14599,N_15627);
nor U17412 (N_17412,N_14394,N_14257);
or U17413 (N_17413,N_14161,N_15078);
and U17414 (N_17414,N_15476,N_15115);
nand U17415 (N_17415,N_15480,N_15812);
nor U17416 (N_17416,N_14718,N_14759);
and U17417 (N_17417,N_14055,N_14511);
nand U17418 (N_17418,N_14528,N_14670);
nand U17419 (N_17419,N_14875,N_15175);
and U17420 (N_17420,N_15264,N_15798);
nand U17421 (N_17421,N_14020,N_15966);
nor U17422 (N_17422,N_14314,N_15042);
nand U17423 (N_17423,N_15732,N_14099);
nor U17424 (N_17424,N_14789,N_14630);
nand U17425 (N_17425,N_14329,N_14821);
nand U17426 (N_17426,N_14104,N_15351);
or U17427 (N_17427,N_15651,N_15886);
or U17428 (N_17428,N_14931,N_15814);
and U17429 (N_17429,N_15331,N_14717);
nand U17430 (N_17430,N_15484,N_15841);
nor U17431 (N_17431,N_14649,N_15300);
nand U17432 (N_17432,N_15341,N_14561);
or U17433 (N_17433,N_14164,N_15813);
and U17434 (N_17434,N_14496,N_15968);
or U17435 (N_17435,N_14225,N_14667);
xor U17436 (N_17436,N_15449,N_14381);
or U17437 (N_17437,N_15422,N_14967);
nor U17438 (N_17438,N_14262,N_15255);
and U17439 (N_17439,N_14048,N_14906);
nand U17440 (N_17440,N_14355,N_14525);
and U17441 (N_17441,N_15076,N_14968);
or U17442 (N_17442,N_14200,N_15823);
and U17443 (N_17443,N_15760,N_14390);
or U17444 (N_17444,N_14898,N_15378);
nand U17445 (N_17445,N_14543,N_15069);
nand U17446 (N_17446,N_15763,N_14845);
xnor U17447 (N_17447,N_15557,N_14698);
nand U17448 (N_17448,N_14245,N_15796);
and U17449 (N_17449,N_14248,N_15712);
nor U17450 (N_17450,N_14051,N_15191);
nor U17451 (N_17451,N_15626,N_14142);
nand U17452 (N_17452,N_15253,N_14236);
and U17453 (N_17453,N_14643,N_15470);
or U17454 (N_17454,N_14346,N_15606);
or U17455 (N_17455,N_15309,N_14152);
nor U17456 (N_17456,N_15841,N_15079);
nor U17457 (N_17457,N_14505,N_15947);
nand U17458 (N_17458,N_14347,N_15450);
or U17459 (N_17459,N_15194,N_15122);
xnor U17460 (N_17460,N_15341,N_14240);
nor U17461 (N_17461,N_14004,N_15521);
nor U17462 (N_17462,N_14916,N_15668);
or U17463 (N_17463,N_15187,N_14487);
nor U17464 (N_17464,N_14421,N_15866);
nand U17465 (N_17465,N_15172,N_14199);
nand U17466 (N_17466,N_14288,N_14199);
nor U17467 (N_17467,N_14554,N_14645);
or U17468 (N_17468,N_15637,N_14643);
or U17469 (N_17469,N_15561,N_15512);
or U17470 (N_17470,N_14125,N_14674);
nor U17471 (N_17471,N_14550,N_15553);
nand U17472 (N_17472,N_14501,N_15687);
nand U17473 (N_17473,N_15664,N_14039);
nor U17474 (N_17474,N_14004,N_15727);
xor U17475 (N_17475,N_14485,N_14236);
nand U17476 (N_17476,N_15218,N_15815);
or U17477 (N_17477,N_15975,N_14124);
nor U17478 (N_17478,N_15684,N_14774);
or U17479 (N_17479,N_14882,N_15758);
and U17480 (N_17480,N_15407,N_14152);
xor U17481 (N_17481,N_15993,N_14499);
nor U17482 (N_17482,N_14280,N_15605);
or U17483 (N_17483,N_15172,N_14866);
nor U17484 (N_17484,N_14648,N_15290);
nor U17485 (N_17485,N_15645,N_14025);
nand U17486 (N_17486,N_14400,N_15859);
nand U17487 (N_17487,N_15743,N_14919);
and U17488 (N_17488,N_14309,N_14300);
and U17489 (N_17489,N_14609,N_14218);
and U17490 (N_17490,N_15711,N_15793);
nor U17491 (N_17491,N_14262,N_14067);
nor U17492 (N_17492,N_15105,N_14630);
nand U17493 (N_17493,N_15912,N_15159);
nand U17494 (N_17494,N_15035,N_15107);
nand U17495 (N_17495,N_15457,N_14429);
and U17496 (N_17496,N_15209,N_15637);
and U17497 (N_17497,N_14117,N_14814);
and U17498 (N_17498,N_15259,N_15856);
nor U17499 (N_17499,N_14835,N_15880);
and U17500 (N_17500,N_14910,N_14902);
or U17501 (N_17501,N_14263,N_15256);
and U17502 (N_17502,N_15831,N_14340);
and U17503 (N_17503,N_14840,N_14707);
or U17504 (N_17504,N_14432,N_14864);
or U17505 (N_17505,N_15500,N_14502);
nor U17506 (N_17506,N_14547,N_14823);
nor U17507 (N_17507,N_15807,N_14889);
nand U17508 (N_17508,N_15838,N_15093);
nor U17509 (N_17509,N_15506,N_15193);
nand U17510 (N_17510,N_14938,N_14303);
and U17511 (N_17511,N_15991,N_14629);
nor U17512 (N_17512,N_15823,N_14657);
nand U17513 (N_17513,N_14232,N_14098);
xnor U17514 (N_17514,N_15154,N_15466);
and U17515 (N_17515,N_14206,N_15641);
xnor U17516 (N_17516,N_14111,N_14036);
or U17517 (N_17517,N_15058,N_14214);
nand U17518 (N_17518,N_14827,N_14483);
xor U17519 (N_17519,N_14870,N_14516);
nand U17520 (N_17520,N_14350,N_14896);
nor U17521 (N_17521,N_15165,N_14258);
nand U17522 (N_17522,N_14699,N_14166);
nand U17523 (N_17523,N_14915,N_14058);
nor U17524 (N_17524,N_15137,N_15704);
or U17525 (N_17525,N_15281,N_14787);
or U17526 (N_17526,N_15214,N_15320);
and U17527 (N_17527,N_14480,N_15256);
nor U17528 (N_17528,N_15003,N_15286);
nand U17529 (N_17529,N_15990,N_15626);
or U17530 (N_17530,N_15067,N_15979);
and U17531 (N_17531,N_15126,N_14524);
nand U17532 (N_17532,N_14372,N_14788);
and U17533 (N_17533,N_15663,N_14796);
xor U17534 (N_17534,N_14982,N_14508);
xor U17535 (N_17535,N_15612,N_15366);
or U17536 (N_17536,N_14311,N_15912);
or U17537 (N_17537,N_15850,N_15104);
nor U17538 (N_17538,N_15182,N_15826);
nand U17539 (N_17539,N_14290,N_14528);
nand U17540 (N_17540,N_14357,N_15726);
and U17541 (N_17541,N_14479,N_14316);
nand U17542 (N_17542,N_14105,N_15765);
xor U17543 (N_17543,N_14697,N_15323);
nor U17544 (N_17544,N_15815,N_15271);
nand U17545 (N_17545,N_15285,N_15619);
or U17546 (N_17546,N_15025,N_15881);
nor U17547 (N_17547,N_15459,N_15829);
nand U17548 (N_17548,N_14177,N_14651);
or U17549 (N_17549,N_15154,N_14612);
nor U17550 (N_17550,N_14379,N_15753);
xnor U17551 (N_17551,N_15774,N_15123);
nand U17552 (N_17552,N_14641,N_14710);
and U17553 (N_17553,N_14845,N_14134);
or U17554 (N_17554,N_15188,N_14191);
nor U17555 (N_17555,N_15942,N_14163);
xor U17556 (N_17556,N_14887,N_14881);
or U17557 (N_17557,N_14389,N_15207);
and U17558 (N_17558,N_14058,N_15586);
nand U17559 (N_17559,N_15274,N_14378);
nand U17560 (N_17560,N_15628,N_14538);
nand U17561 (N_17561,N_15150,N_15798);
nand U17562 (N_17562,N_15927,N_15708);
nand U17563 (N_17563,N_15639,N_14291);
nand U17564 (N_17564,N_15031,N_14863);
or U17565 (N_17565,N_15448,N_15402);
and U17566 (N_17566,N_15551,N_15350);
nor U17567 (N_17567,N_15236,N_14374);
nor U17568 (N_17568,N_14315,N_15037);
xor U17569 (N_17569,N_15213,N_14123);
nand U17570 (N_17570,N_15472,N_14109);
or U17571 (N_17571,N_14491,N_15196);
xnor U17572 (N_17572,N_14015,N_14638);
and U17573 (N_17573,N_14004,N_15330);
and U17574 (N_17574,N_14651,N_14471);
nand U17575 (N_17575,N_14401,N_15074);
or U17576 (N_17576,N_15726,N_15144);
or U17577 (N_17577,N_14101,N_15778);
nand U17578 (N_17578,N_14903,N_14228);
or U17579 (N_17579,N_15343,N_15219);
nor U17580 (N_17580,N_15658,N_15382);
or U17581 (N_17581,N_15769,N_14143);
nand U17582 (N_17582,N_15107,N_14812);
nor U17583 (N_17583,N_14390,N_15446);
and U17584 (N_17584,N_15626,N_14531);
xnor U17585 (N_17585,N_14122,N_14069);
xnor U17586 (N_17586,N_14346,N_15349);
nand U17587 (N_17587,N_15606,N_15028);
nand U17588 (N_17588,N_15747,N_14216);
nor U17589 (N_17589,N_14283,N_15167);
or U17590 (N_17590,N_14103,N_15274);
or U17591 (N_17591,N_15533,N_14331);
nand U17592 (N_17592,N_14700,N_14001);
nor U17593 (N_17593,N_15728,N_15991);
xnor U17594 (N_17594,N_15081,N_14532);
or U17595 (N_17595,N_14244,N_14822);
nor U17596 (N_17596,N_15680,N_15804);
nor U17597 (N_17597,N_14773,N_14603);
nand U17598 (N_17598,N_14534,N_15422);
or U17599 (N_17599,N_14018,N_15008);
nor U17600 (N_17600,N_14601,N_15710);
nand U17601 (N_17601,N_14367,N_14484);
or U17602 (N_17602,N_14269,N_15997);
nor U17603 (N_17603,N_15860,N_14133);
and U17604 (N_17604,N_14646,N_14644);
and U17605 (N_17605,N_15737,N_14253);
nor U17606 (N_17606,N_14251,N_14374);
or U17607 (N_17607,N_15213,N_14195);
nor U17608 (N_17608,N_14501,N_14808);
or U17609 (N_17609,N_15127,N_15526);
nand U17610 (N_17610,N_14130,N_15823);
or U17611 (N_17611,N_15210,N_14688);
nor U17612 (N_17612,N_14029,N_14035);
nand U17613 (N_17613,N_15059,N_15873);
and U17614 (N_17614,N_14572,N_14967);
nor U17615 (N_17615,N_15678,N_14467);
or U17616 (N_17616,N_15354,N_15864);
nor U17617 (N_17617,N_14635,N_15847);
or U17618 (N_17618,N_14890,N_14895);
xor U17619 (N_17619,N_14246,N_15213);
nand U17620 (N_17620,N_14973,N_15446);
nand U17621 (N_17621,N_14621,N_15799);
nor U17622 (N_17622,N_14219,N_14624);
or U17623 (N_17623,N_15656,N_15788);
or U17624 (N_17624,N_15204,N_14576);
and U17625 (N_17625,N_15806,N_14528);
nand U17626 (N_17626,N_14689,N_14941);
or U17627 (N_17627,N_15160,N_14823);
nand U17628 (N_17628,N_14336,N_15572);
and U17629 (N_17629,N_15530,N_15215);
xor U17630 (N_17630,N_14775,N_14885);
nor U17631 (N_17631,N_14441,N_15832);
xnor U17632 (N_17632,N_14472,N_15695);
and U17633 (N_17633,N_14856,N_14779);
nand U17634 (N_17634,N_14725,N_14975);
nand U17635 (N_17635,N_14518,N_14804);
and U17636 (N_17636,N_15218,N_14373);
xnor U17637 (N_17637,N_15314,N_14221);
and U17638 (N_17638,N_15366,N_14017);
and U17639 (N_17639,N_15847,N_15104);
nor U17640 (N_17640,N_15308,N_15922);
xor U17641 (N_17641,N_15737,N_14830);
and U17642 (N_17642,N_14230,N_14865);
xor U17643 (N_17643,N_14450,N_15568);
and U17644 (N_17644,N_15696,N_15780);
nor U17645 (N_17645,N_14084,N_15896);
xor U17646 (N_17646,N_14192,N_14418);
xor U17647 (N_17647,N_15644,N_15018);
nand U17648 (N_17648,N_14931,N_14049);
and U17649 (N_17649,N_14680,N_14732);
or U17650 (N_17650,N_15141,N_15061);
and U17651 (N_17651,N_15419,N_15776);
nor U17652 (N_17652,N_15081,N_14729);
nor U17653 (N_17653,N_14602,N_15435);
xor U17654 (N_17654,N_14584,N_14113);
and U17655 (N_17655,N_14796,N_14367);
or U17656 (N_17656,N_14959,N_14480);
and U17657 (N_17657,N_15639,N_15986);
and U17658 (N_17658,N_14363,N_15113);
or U17659 (N_17659,N_15043,N_14596);
nand U17660 (N_17660,N_15965,N_15188);
and U17661 (N_17661,N_15763,N_14909);
nor U17662 (N_17662,N_14658,N_15576);
nand U17663 (N_17663,N_14884,N_15754);
or U17664 (N_17664,N_15327,N_15338);
nor U17665 (N_17665,N_14806,N_14473);
nor U17666 (N_17666,N_14706,N_14553);
and U17667 (N_17667,N_15085,N_14407);
nand U17668 (N_17668,N_14798,N_14553);
nor U17669 (N_17669,N_14030,N_15731);
xor U17670 (N_17670,N_15106,N_15474);
and U17671 (N_17671,N_15889,N_15162);
xor U17672 (N_17672,N_15660,N_14920);
nor U17673 (N_17673,N_15206,N_14188);
nand U17674 (N_17674,N_15273,N_15955);
or U17675 (N_17675,N_14785,N_15307);
nor U17676 (N_17676,N_14143,N_15953);
nor U17677 (N_17677,N_14725,N_15770);
xnor U17678 (N_17678,N_14667,N_14223);
and U17679 (N_17679,N_14762,N_15894);
xor U17680 (N_17680,N_15882,N_14171);
nand U17681 (N_17681,N_14819,N_14861);
or U17682 (N_17682,N_14103,N_14523);
and U17683 (N_17683,N_14566,N_15752);
nand U17684 (N_17684,N_15116,N_14923);
and U17685 (N_17685,N_14068,N_14794);
or U17686 (N_17686,N_15463,N_14153);
nand U17687 (N_17687,N_15795,N_14456);
or U17688 (N_17688,N_15134,N_15516);
nand U17689 (N_17689,N_15942,N_15755);
nand U17690 (N_17690,N_15806,N_14296);
xor U17691 (N_17691,N_14289,N_14790);
nand U17692 (N_17692,N_14654,N_14366);
or U17693 (N_17693,N_15645,N_14190);
nor U17694 (N_17694,N_15360,N_15886);
nand U17695 (N_17695,N_14198,N_15506);
nor U17696 (N_17696,N_14764,N_14596);
xor U17697 (N_17697,N_14002,N_14295);
nand U17698 (N_17698,N_15995,N_14595);
nand U17699 (N_17699,N_15526,N_15267);
and U17700 (N_17700,N_15875,N_14821);
nor U17701 (N_17701,N_14113,N_14538);
nor U17702 (N_17702,N_15516,N_14992);
and U17703 (N_17703,N_15223,N_14000);
nor U17704 (N_17704,N_15718,N_15420);
xnor U17705 (N_17705,N_15708,N_15470);
or U17706 (N_17706,N_15041,N_14608);
or U17707 (N_17707,N_15240,N_15758);
or U17708 (N_17708,N_15889,N_14112);
and U17709 (N_17709,N_15754,N_14327);
nand U17710 (N_17710,N_15992,N_15522);
nor U17711 (N_17711,N_14246,N_14701);
nor U17712 (N_17712,N_14879,N_14363);
or U17713 (N_17713,N_14565,N_15111);
nor U17714 (N_17714,N_15289,N_15585);
nor U17715 (N_17715,N_14414,N_15520);
nor U17716 (N_17716,N_14780,N_14223);
nand U17717 (N_17717,N_14657,N_14273);
nand U17718 (N_17718,N_14357,N_15808);
nor U17719 (N_17719,N_15268,N_14572);
nor U17720 (N_17720,N_15545,N_14175);
xnor U17721 (N_17721,N_15077,N_15917);
or U17722 (N_17722,N_14006,N_14644);
nor U17723 (N_17723,N_14851,N_15880);
nand U17724 (N_17724,N_15333,N_15897);
or U17725 (N_17725,N_15427,N_15327);
nor U17726 (N_17726,N_15916,N_14718);
and U17727 (N_17727,N_15295,N_14756);
xnor U17728 (N_17728,N_14552,N_15440);
nor U17729 (N_17729,N_15223,N_14757);
and U17730 (N_17730,N_14138,N_15660);
nand U17731 (N_17731,N_15419,N_15660);
nand U17732 (N_17732,N_15426,N_14958);
nor U17733 (N_17733,N_15423,N_14164);
nand U17734 (N_17734,N_14376,N_15264);
nand U17735 (N_17735,N_15024,N_15314);
nand U17736 (N_17736,N_14603,N_14622);
nor U17737 (N_17737,N_15158,N_14775);
nor U17738 (N_17738,N_14050,N_14468);
nand U17739 (N_17739,N_14209,N_15548);
nand U17740 (N_17740,N_14320,N_14180);
or U17741 (N_17741,N_14472,N_14622);
xor U17742 (N_17742,N_15489,N_14092);
and U17743 (N_17743,N_14245,N_14175);
and U17744 (N_17744,N_15916,N_14586);
xor U17745 (N_17745,N_14000,N_14011);
nand U17746 (N_17746,N_14895,N_14154);
nor U17747 (N_17747,N_15534,N_15529);
xor U17748 (N_17748,N_14077,N_15966);
nand U17749 (N_17749,N_15406,N_15817);
nor U17750 (N_17750,N_15924,N_15310);
or U17751 (N_17751,N_15737,N_14251);
nand U17752 (N_17752,N_14754,N_15107);
nor U17753 (N_17753,N_14160,N_15093);
nand U17754 (N_17754,N_15289,N_15197);
nor U17755 (N_17755,N_14413,N_14978);
and U17756 (N_17756,N_14401,N_14233);
nand U17757 (N_17757,N_14311,N_14898);
and U17758 (N_17758,N_15645,N_14883);
xnor U17759 (N_17759,N_15931,N_15995);
or U17760 (N_17760,N_14431,N_15398);
nor U17761 (N_17761,N_15778,N_14237);
nand U17762 (N_17762,N_15168,N_14685);
and U17763 (N_17763,N_15221,N_14536);
nor U17764 (N_17764,N_15119,N_14159);
nand U17765 (N_17765,N_14156,N_15522);
and U17766 (N_17766,N_14076,N_14471);
nor U17767 (N_17767,N_14262,N_15931);
or U17768 (N_17768,N_14522,N_15908);
nand U17769 (N_17769,N_15619,N_14160);
nor U17770 (N_17770,N_15817,N_14063);
xor U17771 (N_17771,N_15203,N_15853);
nor U17772 (N_17772,N_14222,N_15665);
and U17773 (N_17773,N_14492,N_15171);
or U17774 (N_17774,N_15038,N_14162);
or U17775 (N_17775,N_14707,N_15166);
or U17776 (N_17776,N_15816,N_14911);
nand U17777 (N_17777,N_14480,N_15673);
nand U17778 (N_17778,N_15945,N_15589);
xnor U17779 (N_17779,N_15164,N_14416);
and U17780 (N_17780,N_15913,N_14172);
nor U17781 (N_17781,N_15728,N_14089);
xnor U17782 (N_17782,N_14584,N_15670);
xnor U17783 (N_17783,N_14470,N_15750);
nor U17784 (N_17784,N_15073,N_14635);
or U17785 (N_17785,N_15615,N_14518);
and U17786 (N_17786,N_14132,N_15994);
and U17787 (N_17787,N_14870,N_15863);
xnor U17788 (N_17788,N_15723,N_14315);
or U17789 (N_17789,N_14109,N_15833);
nor U17790 (N_17790,N_15600,N_14781);
nor U17791 (N_17791,N_14201,N_15140);
or U17792 (N_17792,N_15197,N_14389);
nand U17793 (N_17793,N_15053,N_15671);
nor U17794 (N_17794,N_14720,N_15623);
or U17795 (N_17795,N_15560,N_14117);
nor U17796 (N_17796,N_15824,N_14265);
or U17797 (N_17797,N_14027,N_14196);
or U17798 (N_17798,N_14916,N_15331);
and U17799 (N_17799,N_15247,N_15950);
xnor U17800 (N_17800,N_15992,N_14007);
nand U17801 (N_17801,N_14242,N_14286);
xor U17802 (N_17802,N_14130,N_15469);
or U17803 (N_17803,N_14858,N_15164);
nor U17804 (N_17804,N_15921,N_14484);
and U17805 (N_17805,N_15250,N_14730);
and U17806 (N_17806,N_14262,N_14589);
or U17807 (N_17807,N_14864,N_15516);
or U17808 (N_17808,N_14384,N_15465);
nor U17809 (N_17809,N_14281,N_15684);
nand U17810 (N_17810,N_15812,N_14720);
nor U17811 (N_17811,N_14556,N_15924);
nor U17812 (N_17812,N_15098,N_15678);
and U17813 (N_17813,N_15966,N_14537);
and U17814 (N_17814,N_15584,N_14606);
nor U17815 (N_17815,N_14295,N_15690);
or U17816 (N_17816,N_15567,N_15022);
xor U17817 (N_17817,N_15827,N_15243);
nand U17818 (N_17818,N_14725,N_15785);
nand U17819 (N_17819,N_14841,N_15538);
xor U17820 (N_17820,N_15221,N_14588);
xnor U17821 (N_17821,N_15509,N_14007);
and U17822 (N_17822,N_14148,N_15599);
and U17823 (N_17823,N_15695,N_15033);
nor U17824 (N_17824,N_14356,N_14107);
nor U17825 (N_17825,N_15500,N_15018);
nand U17826 (N_17826,N_14068,N_14994);
or U17827 (N_17827,N_14934,N_14438);
nor U17828 (N_17828,N_15348,N_15552);
or U17829 (N_17829,N_14328,N_15343);
xor U17830 (N_17830,N_15114,N_15674);
nand U17831 (N_17831,N_15787,N_15462);
or U17832 (N_17832,N_15782,N_15023);
nand U17833 (N_17833,N_15380,N_15303);
nand U17834 (N_17834,N_15294,N_14849);
or U17835 (N_17835,N_14876,N_14873);
nand U17836 (N_17836,N_14279,N_14975);
or U17837 (N_17837,N_14892,N_15673);
nand U17838 (N_17838,N_15624,N_15791);
nor U17839 (N_17839,N_14957,N_14625);
or U17840 (N_17840,N_14589,N_15546);
or U17841 (N_17841,N_14610,N_14839);
nand U17842 (N_17842,N_14954,N_14573);
and U17843 (N_17843,N_15861,N_14315);
and U17844 (N_17844,N_14800,N_15211);
nand U17845 (N_17845,N_14854,N_15979);
and U17846 (N_17846,N_14887,N_14496);
or U17847 (N_17847,N_14387,N_14340);
or U17848 (N_17848,N_15085,N_14486);
nor U17849 (N_17849,N_15653,N_15374);
or U17850 (N_17850,N_14790,N_14412);
nand U17851 (N_17851,N_14600,N_14675);
or U17852 (N_17852,N_14259,N_15628);
and U17853 (N_17853,N_14468,N_15747);
nor U17854 (N_17854,N_15055,N_14626);
and U17855 (N_17855,N_15948,N_14538);
nor U17856 (N_17856,N_15473,N_15164);
and U17857 (N_17857,N_14026,N_14307);
nand U17858 (N_17858,N_14154,N_15669);
or U17859 (N_17859,N_15409,N_15069);
and U17860 (N_17860,N_14248,N_15831);
and U17861 (N_17861,N_14718,N_15910);
nor U17862 (N_17862,N_15166,N_15944);
nor U17863 (N_17863,N_15733,N_15421);
xnor U17864 (N_17864,N_14104,N_14125);
and U17865 (N_17865,N_14013,N_14436);
nand U17866 (N_17866,N_14536,N_15134);
nor U17867 (N_17867,N_14788,N_14561);
or U17868 (N_17868,N_15291,N_15117);
and U17869 (N_17869,N_15159,N_14336);
and U17870 (N_17870,N_15714,N_14779);
or U17871 (N_17871,N_15225,N_15323);
or U17872 (N_17872,N_14480,N_15541);
xnor U17873 (N_17873,N_15677,N_15179);
and U17874 (N_17874,N_14599,N_14278);
and U17875 (N_17875,N_14118,N_14191);
nand U17876 (N_17876,N_15363,N_15832);
nor U17877 (N_17877,N_15182,N_14929);
nand U17878 (N_17878,N_15137,N_15759);
nor U17879 (N_17879,N_14457,N_15512);
and U17880 (N_17880,N_15307,N_14166);
and U17881 (N_17881,N_15873,N_14163);
nand U17882 (N_17882,N_14637,N_15506);
nor U17883 (N_17883,N_15829,N_14356);
and U17884 (N_17884,N_14340,N_15079);
and U17885 (N_17885,N_14983,N_15161);
nand U17886 (N_17886,N_15058,N_15844);
or U17887 (N_17887,N_14318,N_14837);
nor U17888 (N_17888,N_15879,N_15386);
xnor U17889 (N_17889,N_14431,N_14849);
or U17890 (N_17890,N_15973,N_14748);
or U17891 (N_17891,N_15239,N_15887);
nand U17892 (N_17892,N_15906,N_15378);
nand U17893 (N_17893,N_14761,N_14057);
or U17894 (N_17894,N_14477,N_14978);
and U17895 (N_17895,N_14357,N_14549);
xnor U17896 (N_17896,N_14646,N_14336);
or U17897 (N_17897,N_15030,N_14070);
nand U17898 (N_17898,N_15307,N_15711);
and U17899 (N_17899,N_15771,N_14095);
and U17900 (N_17900,N_14583,N_14983);
and U17901 (N_17901,N_15210,N_15007);
nor U17902 (N_17902,N_14281,N_14729);
nor U17903 (N_17903,N_14040,N_15539);
nand U17904 (N_17904,N_15421,N_14619);
nand U17905 (N_17905,N_15287,N_14967);
or U17906 (N_17906,N_15603,N_15619);
and U17907 (N_17907,N_15059,N_15286);
nor U17908 (N_17908,N_15696,N_15800);
or U17909 (N_17909,N_14539,N_15090);
xnor U17910 (N_17910,N_15390,N_15589);
and U17911 (N_17911,N_15260,N_15210);
xor U17912 (N_17912,N_15562,N_14639);
nor U17913 (N_17913,N_14198,N_14120);
nand U17914 (N_17914,N_14033,N_15695);
or U17915 (N_17915,N_15538,N_15923);
or U17916 (N_17916,N_14054,N_14675);
nor U17917 (N_17917,N_14394,N_15778);
xor U17918 (N_17918,N_14376,N_14855);
or U17919 (N_17919,N_14908,N_14361);
nand U17920 (N_17920,N_15990,N_14199);
nor U17921 (N_17921,N_15623,N_14156);
or U17922 (N_17922,N_15110,N_15039);
nand U17923 (N_17923,N_14415,N_15169);
and U17924 (N_17924,N_14734,N_14579);
nand U17925 (N_17925,N_14641,N_15683);
and U17926 (N_17926,N_14774,N_15288);
nor U17927 (N_17927,N_14879,N_14137);
nor U17928 (N_17928,N_15262,N_14889);
nor U17929 (N_17929,N_14168,N_15900);
or U17930 (N_17930,N_15253,N_14338);
or U17931 (N_17931,N_14926,N_15933);
nor U17932 (N_17932,N_14506,N_15937);
xor U17933 (N_17933,N_15430,N_15960);
nor U17934 (N_17934,N_15902,N_15492);
nor U17935 (N_17935,N_15720,N_15469);
or U17936 (N_17936,N_14781,N_15565);
or U17937 (N_17937,N_14358,N_14670);
and U17938 (N_17938,N_14303,N_14821);
or U17939 (N_17939,N_15886,N_14333);
xnor U17940 (N_17940,N_14113,N_14035);
nor U17941 (N_17941,N_14883,N_15302);
nor U17942 (N_17942,N_15727,N_15204);
and U17943 (N_17943,N_14180,N_15712);
nand U17944 (N_17944,N_15092,N_14707);
nand U17945 (N_17945,N_14232,N_15297);
nor U17946 (N_17946,N_14122,N_14471);
or U17947 (N_17947,N_15720,N_14624);
nand U17948 (N_17948,N_14451,N_15458);
nand U17949 (N_17949,N_15400,N_15815);
nand U17950 (N_17950,N_14994,N_14147);
nor U17951 (N_17951,N_15999,N_15661);
or U17952 (N_17952,N_15642,N_15612);
nand U17953 (N_17953,N_14052,N_15232);
or U17954 (N_17954,N_14698,N_14013);
nand U17955 (N_17955,N_15414,N_14333);
nand U17956 (N_17956,N_14241,N_14263);
nor U17957 (N_17957,N_15429,N_15153);
and U17958 (N_17958,N_15397,N_15779);
and U17959 (N_17959,N_14011,N_14453);
nand U17960 (N_17960,N_14081,N_15340);
or U17961 (N_17961,N_15436,N_14659);
or U17962 (N_17962,N_15757,N_14197);
nand U17963 (N_17963,N_14974,N_15397);
and U17964 (N_17964,N_14422,N_14589);
nor U17965 (N_17965,N_15040,N_14184);
xnor U17966 (N_17966,N_14158,N_15261);
or U17967 (N_17967,N_15770,N_15366);
nand U17968 (N_17968,N_14946,N_15065);
and U17969 (N_17969,N_14164,N_14642);
and U17970 (N_17970,N_15480,N_14511);
or U17971 (N_17971,N_15924,N_14714);
nand U17972 (N_17972,N_14879,N_14823);
and U17973 (N_17973,N_14215,N_14385);
or U17974 (N_17974,N_15141,N_15566);
and U17975 (N_17975,N_14866,N_15016);
nand U17976 (N_17976,N_15108,N_14952);
nor U17977 (N_17977,N_15249,N_14118);
and U17978 (N_17978,N_14044,N_15242);
and U17979 (N_17979,N_14643,N_14685);
nand U17980 (N_17980,N_15805,N_15983);
nor U17981 (N_17981,N_14350,N_14468);
and U17982 (N_17982,N_14952,N_14666);
or U17983 (N_17983,N_14456,N_14746);
xor U17984 (N_17984,N_14401,N_15492);
and U17985 (N_17985,N_14939,N_15166);
and U17986 (N_17986,N_14442,N_15043);
xor U17987 (N_17987,N_14358,N_14371);
nor U17988 (N_17988,N_14993,N_14300);
nand U17989 (N_17989,N_14668,N_14431);
nand U17990 (N_17990,N_14910,N_15321);
or U17991 (N_17991,N_14537,N_15370);
nor U17992 (N_17992,N_14739,N_15253);
or U17993 (N_17993,N_15567,N_14420);
or U17994 (N_17994,N_14239,N_14376);
xor U17995 (N_17995,N_14725,N_14362);
nand U17996 (N_17996,N_15557,N_14056);
and U17997 (N_17997,N_15129,N_14113);
nor U17998 (N_17998,N_15072,N_15445);
xor U17999 (N_17999,N_14653,N_14579);
nand U18000 (N_18000,N_16395,N_17389);
nor U18001 (N_18001,N_17843,N_17499);
or U18002 (N_18002,N_17083,N_16702);
and U18003 (N_18003,N_16649,N_16766);
and U18004 (N_18004,N_17889,N_16075);
nand U18005 (N_18005,N_16475,N_17610);
nand U18006 (N_18006,N_17922,N_16682);
and U18007 (N_18007,N_17804,N_17576);
nor U18008 (N_18008,N_17482,N_17050);
nor U18009 (N_18009,N_17598,N_16963);
and U18010 (N_18010,N_17793,N_16518);
nor U18011 (N_18011,N_16814,N_17017);
xnor U18012 (N_18012,N_16374,N_17696);
nor U18013 (N_18013,N_16293,N_17081);
xnor U18014 (N_18014,N_17084,N_17591);
and U18015 (N_18015,N_16866,N_16451);
xnor U18016 (N_18016,N_17559,N_17519);
xnor U18017 (N_18017,N_17725,N_16332);
nand U18018 (N_18018,N_16225,N_17495);
nand U18019 (N_18019,N_16193,N_16940);
or U18020 (N_18020,N_17269,N_16662);
or U18021 (N_18021,N_17551,N_16288);
nand U18022 (N_18022,N_16961,N_16260);
or U18023 (N_18023,N_17208,N_17644);
nor U18024 (N_18024,N_17563,N_17865);
xor U18025 (N_18025,N_16049,N_16465);
and U18026 (N_18026,N_17789,N_17851);
nor U18027 (N_18027,N_17254,N_17618);
or U18028 (N_18028,N_16815,N_17409);
nor U18029 (N_18029,N_16037,N_17419);
xor U18030 (N_18030,N_16411,N_17461);
and U18031 (N_18031,N_17221,N_17981);
and U18032 (N_18032,N_16852,N_17999);
and U18033 (N_18033,N_16915,N_16425);
nand U18034 (N_18034,N_16651,N_17196);
and U18035 (N_18035,N_17022,N_17051);
xnor U18036 (N_18036,N_16665,N_17752);
and U18037 (N_18037,N_17677,N_17354);
nand U18038 (N_18038,N_16675,N_16842);
nor U18039 (N_18039,N_16116,N_16474);
nor U18040 (N_18040,N_16093,N_17270);
nor U18041 (N_18041,N_16464,N_16657);
nand U18042 (N_18042,N_17806,N_16946);
and U18043 (N_18043,N_17187,N_17853);
nand U18044 (N_18044,N_16357,N_16132);
and U18045 (N_18045,N_16984,N_16389);
and U18046 (N_18046,N_17894,N_16631);
nor U18047 (N_18047,N_16032,N_16066);
nor U18048 (N_18048,N_17932,N_16558);
nor U18049 (N_18049,N_17881,N_17708);
nand U18050 (N_18050,N_16292,N_17417);
or U18051 (N_18051,N_17567,N_16811);
nor U18052 (N_18052,N_17204,N_16568);
nor U18053 (N_18053,N_16047,N_16711);
xnor U18054 (N_18054,N_17227,N_16868);
xor U18055 (N_18055,N_17327,N_16186);
and U18056 (N_18056,N_16385,N_17823);
and U18057 (N_18057,N_16752,N_17260);
nand U18058 (N_18058,N_17935,N_17684);
nor U18059 (N_18059,N_17537,N_17010);
or U18060 (N_18060,N_16031,N_16264);
and U18061 (N_18061,N_17021,N_16044);
nand U18062 (N_18062,N_17357,N_17788);
xor U18063 (N_18063,N_17780,N_16504);
and U18064 (N_18064,N_17513,N_17163);
nor U18065 (N_18065,N_16400,N_16883);
nand U18066 (N_18066,N_16211,N_17186);
and U18067 (N_18067,N_17517,N_16621);
nand U18068 (N_18068,N_16479,N_17747);
and U18069 (N_18069,N_17678,N_16561);
nor U18070 (N_18070,N_17383,N_17681);
nor U18071 (N_18071,N_17338,N_16535);
xor U18072 (N_18072,N_17261,N_17278);
nor U18073 (N_18073,N_17697,N_17300);
nand U18074 (N_18074,N_17984,N_17997);
xor U18075 (N_18075,N_16166,N_16542);
xor U18076 (N_18076,N_16096,N_17957);
nor U18077 (N_18077,N_17818,N_16845);
or U18078 (N_18078,N_17710,N_17469);
nand U18079 (N_18079,N_16019,N_16900);
or U18080 (N_18080,N_16202,N_17873);
and U18081 (N_18081,N_16333,N_17103);
nand U18082 (N_18082,N_16959,N_16945);
and U18083 (N_18083,N_17245,N_17168);
nand U18084 (N_18084,N_16549,N_17514);
xor U18085 (N_18085,N_16496,N_16063);
or U18086 (N_18086,N_17579,N_16003);
nor U18087 (N_18087,N_17509,N_17866);
nor U18088 (N_18088,N_17146,N_17352);
nand U18089 (N_18089,N_17962,N_16403);
and U18090 (N_18090,N_16458,N_16001);
xnor U18091 (N_18091,N_17369,N_17939);
nor U18092 (N_18092,N_17448,N_17869);
nor U18093 (N_18093,N_17458,N_17914);
and U18094 (N_18094,N_17407,N_16301);
and U18095 (N_18095,N_17573,N_16689);
nand U18096 (N_18096,N_17402,N_17488);
nor U18097 (N_18097,N_16080,N_17016);
nor U18098 (N_18098,N_16365,N_17284);
and U18099 (N_18099,N_16499,N_16509);
nand U18100 (N_18100,N_16402,N_17189);
and U18101 (N_18101,N_16950,N_16567);
and U18102 (N_18102,N_17496,N_16862);
or U18103 (N_18103,N_17463,N_17941);
or U18104 (N_18104,N_16776,N_17413);
or U18105 (N_18105,N_16557,N_16299);
nand U18106 (N_18106,N_16199,N_16935);
nor U18107 (N_18107,N_17828,N_17005);
nand U18108 (N_18108,N_17795,N_16459);
nand U18109 (N_18109,N_16204,N_17213);
nor U18110 (N_18110,N_17777,N_17632);
nor U18111 (N_18111,N_16909,N_16009);
or U18112 (N_18112,N_16516,N_17476);
nor U18113 (N_18113,N_17716,N_17497);
or U18114 (N_18114,N_17673,N_17113);
nand U18115 (N_18115,N_17165,N_17190);
and U18116 (N_18116,N_17515,N_17283);
or U18117 (N_18117,N_16074,N_16762);
nor U18118 (N_18118,N_16248,N_17958);
or U18119 (N_18119,N_17114,N_16358);
or U18120 (N_18120,N_16577,N_16198);
nand U18121 (N_18121,N_16515,N_16599);
nand U18122 (N_18122,N_17698,N_16180);
and U18123 (N_18123,N_17919,N_17439);
and U18124 (N_18124,N_17875,N_16169);
xor U18125 (N_18125,N_17808,N_16369);
and U18126 (N_18126,N_16798,N_17794);
nand U18127 (N_18127,N_16636,N_16175);
and U18128 (N_18128,N_17290,N_16467);
nand U18129 (N_18129,N_17832,N_16927);
and U18130 (N_18130,N_17368,N_17129);
nand U18131 (N_18131,N_16489,N_16065);
nor U18132 (N_18132,N_17315,N_16786);
or U18133 (N_18133,N_16258,N_17220);
and U18134 (N_18134,N_16121,N_16789);
nand U18135 (N_18135,N_16000,N_17304);
nor U18136 (N_18136,N_17266,N_16746);
nor U18137 (N_18137,N_16763,N_16566);
and U18138 (N_18138,N_16912,N_17403);
nand U18139 (N_18139,N_16684,N_16036);
nor U18140 (N_18140,N_17735,N_17655);
xnor U18141 (N_18141,N_16462,N_16871);
nand U18142 (N_18142,N_16254,N_16415);
nand U18143 (N_18143,N_16807,N_16017);
or U18144 (N_18144,N_17161,N_16751);
nand U18145 (N_18145,N_17344,N_17271);
or U18146 (N_18146,N_17728,N_16781);
nand U18147 (N_18147,N_17322,N_17756);
or U18148 (N_18148,N_17111,N_17264);
nand U18149 (N_18149,N_16461,N_17019);
and U18150 (N_18150,N_17240,N_17790);
nor U18151 (N_18151,N_16068,N_17700);
and U18152 (N_18152,N_16004,N_17621);
and U18153 (N_18153,N_16229,N_17947);
or U18154 (N_18154,N_16448,N_16905);
nand U18155 (N_18155,N_16717,N_16362);
nand U18156 (N_18156,N_17105,N_16768);
nor U18157 (N_18157,N_17243,N_17842);
or U18158 (N_18158,N_17432,N_16368);
nand U18159 (N_18159,N_16942,N_17726);
nor U18160 (N_18160,N_16218,N_17769);
nand U18161 (N_18161,N_16092,N_17709);
nor U18162 (N_18162,N_16081,N_16339);
and U18163 (N_18163,N_16405,N_17142);
or U18164 (N_18164,N_16994,N_17032);
or U18165 (N_18165,N_16147,N_16988);
nor U18166 (N_18166,N_17241,N_16351);
nand U18167 (N_18167,N_16686,N_17042);
nor U18168 (N_18168,N_16491,N_17000);
and U18169 (N_18169,N_17502,N_16409);
nor U18170 (N_18170,N_17041,N_17233);
or U18171 (N_18171,N_17702,N_16290);
or U18172 (N_18172,N_16094,N_16315);
or U18173 (N_18173,N_17393,N_17454);
nor U18174 (N_18174,N_16976,N_16646);
or U18175 (N_18175,N_16250,N_16124);
nor U18176 (N_18176,N_17028,N_17167);
or U18177 (N_18177,N_16157,N_17924);
or U18178 (N_18178,N_16624,N_16226);
and U18179 (N_18179,N_16817,N_16178);
and U18180 (N_18180,N_17137,N_16050);
or U18181 (N_18181,N_17738,N_16452);
nand U18182 (N_18182,N_16142,N_17316);
nor U18183 (N_18183,N_16213,N_17277);
and U18184 (N_18184,N_17377,N_17792);
nand U18185 (N_18185,N_16914,N_17372);
or U18186 (N_18186,N_16140,N_17412);
nand U18187 (N_18187,N_16281,N_17065);
and U18188 (N_18188,N_16043,N_17001);
and U18189 (N_18189,N_17172,N_16920);
nor U18190 (N_18190,N_17874,N_17649);
nor U18191 (N_18191,N_17141,N_17852);
or U18192 (N_18192,N_16583,N_17427);
and U18193 (N_18193,N_16934,N_17486);
nor U18194 (N_18194,N_17311,N_17151);
nor U18195 (N_18195,N_16222,N_16628);
nand U18196 (N_18196,N_17973,N_16341);
xnor U18197 (N_18197,N_16471,N_17477);
nand U18198 (N_18198,N_16972,N_16062);
or U18199 (N_18199,N_17934,N_17855);
or U18200 (N_18200,N_17029,N_16256);
or U18201 (N_18201,N_17665,N_17094);
or U18202 (N_18202,N_16363,N_16980);
and U18203 (N_18203,N_17931,N_17586);
and U18204 (N_18204,N_16591,N_17671);
or U18205 (N_18205,N_16579,N_17720);
xnor U18206 (N_18206,N_17596,N_16174);
nand U18207 (N_18207,N_16408,N_16782);
nor U18208 (N_18208,N_17078,N_17195);
nand U18209 (N_18209,N_16478,N_16687);
and U18210 (N_18210,N_17787,N_16632);
nand U18211 (N_18211,N_17468,N_16604);
and U18212 (N_18212,N_17009,N_17149);
nor U18213 (N_18213,N_17930,N_16623);
or U18214 (N_18214,N_17159,N_17560);
or U18215 (N_18215,N_16601,N_16273);
or U18216 (N_18216,N_16843,N_16476);
or U18217 (N_18217,N_16445,N_16681);
or U18218 (N_18218,N_17179,N_16446);
and U18219 (N_18219,N_16838,N_16308);
or U18220 (N_18220,N_17288,N_16261);
or U18221 (N_18221,N_17653,N_17031);
nand U18222 (N_18222,N_17859,N_17951);
and U18223 (N_18223,N_16525,N_16795);
or U18224 (N_18224,N_16565,N_17332);
and U18225 (N_18225,N_17492,N_16192);
nand U18226 (N_18226,N_17569,N_16569);
nand U18227 (N_18227,N_16406,N_16699);
and U18228 (N_18228,N_16421,N_17723);
nand U18229 (N_18229,N_17211,N_17191);
xnor U18230 (N_18230,N_16418,N_16680);
nor U18231 (N_18231,N_16955,N_17478);
nand U18232 (N_18232,N_17830,N_17512);
and U18233 (N_18233,N_16997,N_16110);
xor U18234 (N_18234,N_17764,N_17088);
or U18235 (N_18235,N_16442,N_16943);
or U18236 (N_18236,N_16748,N_17637);
nand U18237 (N_18237,N_16791,N_16519);
nor U18238 (N_18238,N_16171,N_16241);
nor U18239 (N_18239,N_17394,N_17494);
and U18240 (N_18240,N_16833,N_16770);
nor U18241 (N_18241,N_16939,N_17916);
xor U18242 (N_18242,N_17157,N_17376);
or U18243 (N_18243,N_16867,N_17026);
and U18244 (N_18244,N_17046,N_16750);
or U18245 (N_18245,N_17169,N_17504);
and U18246 (N_18246,N_17385,N_17136);
or U18247 (N_18247,N_17093,N_17438);
nand U18248 (N_18248,N_16006,N_17824);
and U18249 (N_18249,N_16122,N_16373);
nand U18250 (N_18250,N_16644,N_16777);
nand U18251 (N_18251,N_17132,N_16126);
and U18252 (N_18252,N_17647,N_17742);
and U18253 (N_18253,N_16506,N_16787);
or U18254 (N_18254,N_16576,N_16424);
nand U18255 (N_18255,N_17308,N_16309);
nand U18256 (N_18256,N_16806,N_17500);
xor U18257 (N_18257,N_16376,N_17143);
or U18258 (N_18258,N_16528,N_17614);
or U18259 (N_18259,N_17858,N_17802);
or U18260 (N_18260,N_16613,N_16554);
or U18261 (N_18261,N_17058,N_16804);
or U18262 (N_18262,N_17971,N_16257);
and U18263 (N_18263,N_16145,N_16371);
nor U18264 (N_18264,N_17908,N_17783);
or U18265 (N_18265,N_17236,N_16419);
and U18266 (N_18266,N_16349,N_17127);
or U18267 (N_18267,N_16191,N_16234);
nand U18268 (N_18268,N_17231,N_17007);
nor U18269 (N_18269,N_17328,N_17302);
and U18270 (N_18270,N_17133,N_17526);
or U18271 (N_18271,N_17856,N_17306);
and U18272 (N_18272,N_17654,N_17685);
and U18273 (N_18273,N_17218,N_17964);
and U18274 (N_18274,N_16978,N_16018);
and U18275 (N_18275,N_17917,N_17037);
nand U18276 (N_18276,N_16130,N_17774);
and U18277 (N_18277,N_17651,N_17730);
and U18278 (N_18278,N_16352,N_17287);
and U18279 (N_18279,N_17834,N_17837);
nand U18280 (N_18280,N_16923,N_16873);
or U18281 (N_18281,N_16117,N_17566);
and U18282 (N_18282,N_16099,N_17667);
nor U18283 (N_18283,N_17929,N_17734);
nand U18284 (N_18284,N_16429,N_16189);
or U18285 (N_18285,N_17238,N_16056);
nor U18286 (N_18286,N_17472,N_17880);
xnor U18287 (N_18287,N_16823,N_16648);
xnor U18288 (N_18288,N_17295,N_16654);
nor U18289 (N_18289,N_16297,N_16188);
xor U18290 (N_18290,N_17555,N_16020);
and U18291 (N_18291,N_16219,N_17979);
nor U18292 (N_18292,N_16025,N_17839);
nand U18293 (N_18293,N_17571,N_16713);
xnor U18294 (N_18294,N_17663,N_17550);
or U18295 (N_18295,N_16906,N_17814);
or U18296 (N_18296,N_16187,N_16853);
nand U18297 (N_18297,N_16598,N_17303);
nand U18298 (N_18298,N_17467,N_17912);
nor U18299 (N_18299,N_17099,N_17066);
and U18300 (N_18300,N_16220,N_17617);
nand U18301 (N_18301,N_17572,N_17252);
nand U18302 (N_18302,N_17362,N_16876);
and U18303 (N_18303,N_17313,N_16740);
nor U18304 (N_18304,N_16589,N_17622);
xor U18305 (N_18305,N_17247,N_16443);
or U18306 (N_18306,N_17225,N_17582);
and U18307 (N_18307,N_17992,N_16718);
xnor U18308 (N_18308,N_17520,N_16008);
nor U18309 (N_18309,N_16359,N_17707);
nor U18310 (N_18310,N_17092,N_16435);
nand U18311 (N_18311,N_16179,N_17404);
xnor U18312 (N_18312,N_16221,N_16055);
nor U18313 (N_18313,N_17845,N_16857);
nand U18314 (N_18314,N_17670,N_17396);
or U18315 (N_18315,N_16139,N_16394);
nor U18316 (N_18316,N_17718,N_17692);
and U18317 (N_18317,N_16771,N_16283);
and U18318 (N_18318,N_17453,N_17753);
or U18319 (N_18319,N_16505,N_16327);
xor U18320 (N_18320,N_16154,N_16494);
nand U18321 (N_18321,N_16597,N_17237);
xnor U18322 (N_18322,N_17075,N_16076);
and U18323 (N_18323,N_16274,N_17498);
nand U18324 (N_18324,N_17330,N_17988);
nand U18325 (N_18325,N_16730,N_16266);
or U18326 (N_18326,N_16820,N_16911);
or U18327 (N_18327,N_17864,N_17184);
or U18328 (N_18328,N_17722,N_16846);
and U18329 (N_18329,N_16670,N_17397);
nor U18330 (N_18330,N_16760,N_16412);
or U18331 (N_18331,N_17620,N_17547);
nor U18332 (N_18332,N_16397,N_16432);
nor U18333 (N_18333,N_17907,N_16749);
xnor U18334 (N_18334,N_16655,N_16739);
or U18335 (N_18335,N_17549,N_17181);
nand U18336 (N_18336,N_16916,N_16625);
and U18337 (N_18337,N_16836,N_17324);
nor U18338 (N_18338,N_16511,N_17222);
or U18339 (N_18339,N_16812,N_16534);
or U18340 (N_18340,N_17194,N_16305);
and U18341 (N_18341,N_16706,N_16658);
and U18342 (N_18342,N_17175,N_16156);
and U18343 (N_18343,N_16469,N_16490);
and U18344 (N_18344,N_17536,N_16433);
and U18345 (N_18345,N_16919,N_16536);
nand U18346 (N_18346,N_16615,N_17969);
nor U18347 (N_18347,N_17705,N_16249);
nand U18348 (N_18348,N_16855,N_16279);
nand U18349 (N_18349,N_17188,N_17786);
nor U18350 (N_18350,N_17612,N_16200);
and U18351 (N_18351,N_16078,N_17493);
and U18352 (N_18352,N_16247,N_16493);
or U18353 (N_18353,N_17033,N_16324);
nand U18354 (N_18354,N_16380,N_17391);
xor U18355 (N_18355,N_17895,N_16829);
nor U18356 (N_18356,N_17750,N_16141);
and U18357 (N_18357,N_16162,N_17664);
and U18358 (N_18358,N_16246,N_17018);
or U18359 (N_18359,N_16639,N_17317);
nand U18360 (N_18360,N_16059,N_17460);
nand U18361 (N_18361,N_17535,N_17381);
nand U18362 (N_18362,N_16058,N_16010);
nand U18363 (N_18363,N_17721,N_16100);
and U18364 (N_18364,N_17430,N_17963);
nor U18365 (N_18365,N_17740,N_16118);
and U18366 (N_18366,N_17603,N_16585);
nand U18367 (N_18367,N_17212,N_17599);
and U18368 (N_18368,N_16693,N_16340);
or U18369 (N_18369,N_17158,N_17867);
or U18370 (N_18370,N_16860,N_17539);
and U18371 (N_18371,N_16431,N_17055);
nand U18372 (N_18372,N_16390,N_16386);
nand U18373 (N_18373,N_17980,N_16965);
and U18374 (N_18374,N_16932,N_16630);
nor U18375 (N_18375,N_17455,N_16127);
nand U18376 (N_18376,N_16553,N_16284);
nor U18377 (N_18377,N_17418,N_16237);
nor U18378 (N_18378,N_16137,N_17027);
and U18379 (N_18379,N_17624,N_16456);
and U18380 (N_18380,N_17887,N_17982);
xnor U18381 (N_18381,N_17145,N_17443);
nand U18382 (N_18382,N_17544,N_16951);
nand U18383 (N_18383,N_17100,N_16353);
nor U18384 (N_18384,N_17784,N_17457);
and U18385 (N_18385,N_17049,N_17246);
and U18386 (N_18386,N_17810,N_16588);
nand U18387 (N_18387,N_17329,N_16120);
nand U18388 (N_18388,N_17531,N_16272);
and U18389 (N_18389,N_17226,N_16769);
nand U18390 (N_18390,N_17672,N_17897);
xnor U18391 (N_18391,N_16270,N_16331);
and U18392 (N_18392,N_17841,N_16837);
nand U18393 (N_18393,N_17868,N_17680);
nor U18394 (N_18394,N_17761,N_16600);
and U18395 (N_18395,N_16593,N_16023);
and U18396 (N_18396,N_17643,N_16404);
nor U18397 (N_18397,N_17619,N_16007);
and U18398 (N_18398,N_17844,N_17886);
nor U18399 (N_18399,N_17004,N_17959);
nand U18400 (N_18400,N_16354,N_17054);
and U18401 (N_18401,N_17592,N_16129);
nand U18402 (N_18402,N_17117,N_17870);
and U18403 (N_18403,N_17452,N_16841);
nand U18404 (N_18404,N_16714,N_17905);
nand U18405 (N_18405,N_17089,N_16381);
nand U18406 (N_18406,N_17057,N_17206);
or U18407 (N_18407,N_16011,N_17416);
nand U18408 (N_18408,N_16463,N_17578);
xor U18409 (N_18409,N_17255,N_16572);
nand U18410 (N_18410,N_16969,N_17609);
nor U18411 (N_18411,N_16885,N_17339);
and U18412 (N_18412,N_16231,N_17331);
nand U18413 (N_18413,N_16796,N_17428);
and U18414 (N_18414,N_17147,N_16538);
nor U18415 (N_18415,N_16529,N_17077);
nand U18416 (N_18416,N_17694,N_16227);
nor U18417 (N_18417,N_17527,N_16849);
nor U18418 (N_18418,N_16500,N_17589);
or U18419 (N_18419,N_17938,N_16620);
xor U18420 (N_18420,N_17119,N_16485);
nand U18421 (N_18421,N_17139,N_16695);
nand U18422 (N_18422,N_17584,N_17178);
or U18423 (N_18423,N_16015,N_16286);
nand U18424 (N_18424,N_16437,N_17203);
and U18425 (N_18425,N_16197,N_16098);
nor U18426 (N_18426,N_16450,N_17470);
nand U18427 (N_18427,N_17965,N_16556);
and U18428 (N_18428,N_17465,N_17661);
nor U18429 (N_18429,N_17879,N_17820);
nand U18430 (N_18430,N_16958,N_17076);
or U18431 (N_18431,N_17479,N_17898);
nor U18432 (N_18432,N_17892,N_17604);
and U18433 (N_18433,N_16552,N_16524);
nand U18434 (N_18434,N_17501,N_16115);
nor U18435 (N_18435,N_17193,N_17371);
nand U18436 (N_18436,N_16338,N_16575);
nand U18437 (N_18437,N_17768,N_17030);
and U18438 (N_18438,N_17634,N_16701);
or U18439 (N_18439,N_17767,N_16560);
and U18440 (N_18440,N_17164,N_16652);
and U18441 (N_18441,N_16077,N_16797);
nor U18442 (N_18442,N_16304,N_17909);
xor U18443 (N_18443,N_16586,N_16278);
or U18444 (N_18444,N_16671,N_16828);
or U18445 (N_18445,N_17543,N_17002);
or U18446 (N_18446,N_17781,N_17390);
and U18447 (N_18447,N_17286,N_16236);
nand U18448 (N_18448,N_17760,N_17778);
nand U18449 (N_18449,N_17253,N_16563);
or U18450 (N_18450,N_16087,N_17309);
or U18451 (N_18451,N_17860,N_17575);
and U18452 (N_18452,N_16269,N_17862);
nand U18453 (N_18453,N_16998,N_17926);
and U18454 (N_18454,N_17131,N_17952);
xor U18455 (N_18455,N_16238,N_17360);
and U18456 (N_18456,N_16112,N_17518);
nor U18457 (N_18457,N_17216,N_16195);
nand U18458 (N_18458,N_17878,N_17524);
or U18459 (N_18459,N_16230,N_17809);
nand U18460 (N_18460,N_16048,N_16877);
or U18461 (N_18461,N_16460,N_16893);
xnor U18462 (N_18462,N_16417,N_16131);
or U18463 (N_18463,N_17408,N_16207);
and U18464 (N_18464,N_17706,N_16033);
and U18465 (N_18465,N_16161,N_17154);
xor U18466 (N_18466,N_16133,N_16948);
nor U18467 (N_18467,N_17395,N_17405);
or U18468 (N_18468,N_16578,N_16881);
nor U18469 (N_18469,N_16741,N_16974);
xor U18470 (N_18470,N_16026,N_17949);
nor U18471 (N_18471,N_16878,N_17420);
and U18472 (N_18472,N_17485,N_17574);
or U18473 (N_18473,N_16674,N_16869);
nand U18474 (N_18474,N_17995,N_17993);
nor U18475 (N_18475,N_16143,N_16989);
and U18476 (N_18476,N_17207,N_17557);
nand U18477 (N_18477,N_17558,N_17148);
or U18478 (N_18478,N_16737,N_17732);
or U18479 (N_18479,N_16642,N_16985);
nor U18480 (N_18480,N_16892,N_16864);
nor U18481 (N_18481,N_16172,N_17384);
nor U18482 (N_18482,N_17588,N_17060);
nand U18483 (N_18483,N_16082,N_17024);
nor U18484 (N_18484,N_16407,N_17298);
or U18485 (N_18485,N_17293,N_17364);
nand U18486 (N_18486,N_16992,N_16910);
nand U18487 (N_18487,N_16975,N_17090);
nor U18488 (N_18488,N_17484,N_16393);
nor U18489 (N_18489,N_17101,N_17325);
nor U18490 (N_18490,N_16612,N_16167);
and U18491 (N_18491,N_16858,N_17961);
nor U18492 (N_18492,N_17365,N_16986);
nand U18493 (N_18493,N_17974,N_17883);
and U18494 (N_18494,N_17890,N_16183);
nand U18495 (N_18495,N_16678,N_17776);
nand U18496 (N_18496,N_16716,N_16067);
nand U18497 (N_18497,N_16822,N_16870);
and U18498 (N_18498,N_16801,N_17955);
and U18499 (N_18499,N_17899,N_17507);
xnor U18500 (N_18500,N_16382,N_16208);
xnor U18501 (N_18501,N_16850,N_16816);
and U18502 (N_18502,N_17200,N_17773);
or U18503 (N_18503,N_17442,N_17739);
or U18504 (N_18504,N_17490,N_16103);
and U18505 (N_18505,N_17410,N_17013);
nand U18506 (N_18506,N_17102,N_16917);
and U18507 (N_18507,N_16773,N_17511);
nor U18508 (N_18508,N_16164,N_17259);
and U18509 (N_18509,N_16396,N_17805);
and U18510 (N_18510,N_17215,N_17280);
nor U18511 (N_18511,N_16420,N_17944);
nand U18512 (N_18512,N_17345,N_17893);
or U18513 (N_18513,N_16303,N_17782);
xnor U18514 (N_18514,N_17421,N_16908);
nor U18515 (N_18515,N_17450,N_16155);
or U18516 (N_18516,N_17977,N_17625);
or U18517 (N_18517,N_16398,N_17333);
or U18518 (N_18518,N_16736,N_17817);
and U18519 (N_18519,N_16571,N_16983);
and U18520 (N_18520,N_16125,N_16255);
xnor U18521 (N_18521,N_16165,N_17491);
nor U18522 (N_18522,N_17967,N_17605);
or U18523 (N_18523,N_16617,N_16051);
and U18524 (N_18524,N_16498,N_16979);
and U18525 (N_18525,N_16083,N_17921);
nand U18526 (N_18526,N_16999,N_17160);
or U18527 (N_18527,N_16401,N_17462);
and U18528 (N_18528,N_16772,N_17848);
and U18529 (N_18529,N_16243,N_16774);
and U18530 (N_18530,N_17424,N_17234);
and U18531 (N_18531,N_17434,N_17440);
or U18532 (N_18532,N_16527,N_17927);
or U18533 (N_18533,N_17626,N_17257);
or U18534 (N_18534,N_16423,N_16618);
nor U18535 (N_18535,N_16921,N_17801);
nand U18536 (N_18536,N_17445,N_17202);
nand U18537 (N_18537,N_16323,N_16326);
nand U18538 (N_18538,N_17177,N_16874);
or U18539 (N_18539,N_17972,N_17745);
nor U18540 (N_18540,N_16523,N_17530);
and U18541 (N_18541,N_17068,N_16594);
or U18542 (N_18542,N_16793,N_16851);
nand U18543 (N_18543,N_17265,N_16719);
xor U18544 (N_18544,N_17289,N_16562);
and U18545 (N_18545,N_17640,N_17067);
nand U18546 (N_18546,N_16217,N_16756);
or U18547 (N_18547,N_17456,N_17256);
nor U18548 (N_18548,N_16410,N_16805);
nand U18549 (N_18549,N_17044,N_17945);
xnor U18550 (N_18550,N_16872,N_17449);
or U18551 (N_18551,N_16439,N_16555);
xor U18552 (N_18552,N_17648,N_17249);
nand U18553 (N_18553,N_16271,N_16991);
xnor U18554 (N_18554,N_17884,N_16449);
nand U18555 (N_18555,N_16930,N_16627);
and U18556 (N_18556,N_17754,N_16660);
or U18557 (N_18557,N_16024,N_17447);
nand U18558 (N_18558,N_17350,N_16030);
and U18559 (N_18559,N_17933,N_16809);
nor U18560 (N_18560,N_17174,N_16416);
nand U18561 (N_18561,N_17091,N_16735);
and U18562 (N_18562,N_16106,N_17292);
xnor U18563 (N_18563,N_17095,N_16703);
or U18564 (N_18564,N_17370,N_16477);
or U18565 (N_18565,N_17398,N_17281);
nor U18566 (N_18566,N_17791,N_16302);
nand U18567 (N_18567,N_17082,N_16573);
nand U18568 (N_18568,N_17960,N_16244);
or U18569 (N_18569,N_16602,N_17087);
nor U18570 (N_18570,N_17748,N_16319);
nor U18571 (N_18571,N_16788,N_16582);
nand U18572 (N_18572,N_16497,N_16513);
xor U18573 (N_18573,N_17915,N_17314);
nor U18574 (N_18574,N_16289,N_16884);
or U18575 (N_18575,N_16214,N_17657);
nand U18576 (N_18576,N_17594,N_17629);
nor U18577 (N_18577,N_17765,N_16223);
and U18578 (N_18578,N_16673,N_16531);
or U18579 (N_18579,N_16073,N_16337);
nor U18580 (N_18580,N_17244,N_17863);
and U18581 (N_18581,N_16123,N_17639);
nand U18582 (N_18582,N_16831,N_17719);
or U18583 (N_18583,N_17552,N_17533);
nand U18584 (N_18584,N_17435,N_17601);
and U18585 (N_18585,N_17180,N_17473);
and U18586 (N_18586,N_16184,N_17699);
or U18587 (N_18587,N_16216,N_16700);
nor U18588 (N_18588,N_16635,N_17990);
and U18589 (N_18589,N_16013,N_17274);
nor U18590 (N_18590,N_16607,N_17606);
nor U18591 (N_18591,N_17996,N_16827);
and U18592 (N_18592,N_16267,N_16813);
xor U18593 (N_18593,N_17666,N_17297);
and U18594 (N_18594,N_16375,N_16848);
or U18595 (N_18595,N_16611,N_16265);
and U18596 (N_18596,N_16709,N_16818);
nor U18597 (N_18597,N_17210,N_16775);
xnor U18598 (N_18598,N_16522,N_16095);
and U18599 (N_18599,N_17779,N_16794);
nand U18600 (N_18600,N_17849,N_17251);
and U18601 (N_18601,N_17353,N_16743);
or U18602 (N_18602,N_16928,N_16894);
nand U18603 (N_18603,N_17691,N_17436);
and U18604 (N_18604,N_17737,N_16532);
nand U18605 (N_18605,N_16960,N_16160);
nor U18606 (N_18606,N_16224,N_16715);
nand U18607 (N_18607,N_17656,N_16486);
nand U18608 (N_18608,N_17831,N_17998);
and U18609 (N_18609,N_16440,N_17235);
nand U18610 (N_18610,N_16366,N_17942);
nor U18611 (N_18611,N_17762,N_16206);
or U18612 (N_18612,N_16344,N_16987);
and U18613 (N_18613,N_17217,N_16859);
nand U18614 (N_18614,N_16483,N_17846);
nand U18615 (N_18615,N_16296,N_16539);
nor U18616 (N_18616,N_17185,N_16757);
and U18617 (N_18617,N_17627,N_17920);
nand U18618 (N_18618,N_17382,N_16725);
nor U18619 (N_18619,N_17925,N_17712);
nand U18620 (N_18620,N_16968,N_16668);
nand U18621 (N_18621,N_16543,N_17039);
nand U18622 (N_18622,N_17122,N_17937);
or U18623 (N_18623,N_16564,N_17975);
nor U18624 (N_18624,N_16645,N_16704);
nor U18625 (N_18625,N_16661,N_16252);
or U18626 (N_18626,N_16379,N_17106);
nand U18627 (N_18627,N_17607,N_17061);
nand U18628 (N_18628,N_16287,N_16669);
nor U18629 (N_18629,N_16079,N_16196);
nor U18630 (N_18630,N_16038,N_17910);
nand U18631 (N_18631,N_17401,N_16101);
or U18632 (N_18632,N_17323,N_17541);
nand U18633 (N_18633,N_17043,N_16856);
nor U18634 (N_18634,N_17636,N_17351);
nand U18635 (N_18635,N_17803,N_17561);
nor U18636 (N_18636,N_16294,N_17770);
or U18637 (N_18637,N_17826,N_17534);
nand U18638 (N_18638,N_17638,N_16792);
and U18639 (N_18639,N_17688,N_16102);
and U18640 (N_18640,N_16508,N_17714);
nor U18641 (N_18641,N_16731,N_17441);
nor U18642 (N_18642,N_17562,N_17936);
nand U18643 (N_18643,N_16936,N_16107);
nor U18644 (N_18644,N_16259,N_16526);
and U18645 (N_18645,N_16482,N_17506);
nor U18646 (N_18646,N_17197,N_16320);
or U18647 (N_18647,N_17523,N_16104);
and U18648 (N_18648,N_16039,N_17276);
and U18649 (N_18649,N_16898,N_16314);
nand U18650 (N_18650,N_17829,N_16559);
nand U18651 (N_18651,N_16753,N_16399);
nor U18652 (N_18652,N_17568,N_16041);
nor U18653 (N_18653,N_16712,N_17827);
and U18654 (N_18654,N_16392,N_17976);
and U18655 (N_18655,N_17669,N_17069);
nand U18656 (N_18656,N_17471,N_16785);
nand U18657 (N_18657,N_17785,N_17144);
nor U18658 (N_18658,N_17047,N_16938);
and U18659 (N_18659,N_16929,N_16918);
and U18660 (N_18660,N_17367,N_17816);
or U18661 (N_18661,N_16427,N_17464);
nand U18662 (N_18662,N_16925,N_17318);
or U18663 (N_18663,N_17736,N_16580);
or U18664 (N_18664,N_17411,N_16388);
nor U18665 (N_18665,N_16370,N_17036);
nor U18666 (N_18666,N_17230,N_17319);
and U18667 (N_18667,N_16436,N_17918);
and U18668 (N_18668,N_17630,N_16481);
and U18669 (N_18669,N_17150,N_17020);
and U18670 (N_18670,N_16880,N_16734);
or U18671 (N_18671,N_17219,N_16723);
or U18672 (N_18672,N_16210,N_17433);
and U18673 (N_18673,N_16054,N_16666);
nand U18674 (N_18674,N_17668,N_16176);
nor U18675 (N_18675,N_16492,N_17733);
xnor U18676 (N_18676,N_17349,N_16097);
xor U18677 (N_18677,N_17299,N_17483);
xor U18678 (N_18678,N_17112,N_16981);
and U18679 (N_18679,N_17891,N_16313);
nor U18680 (N_18680,N_16587,N_16378);
nand U18681 (N_18681,N_16907,N_17214);
nand U18682 (N_18682,N_16487,N_16891);
nor U18683 (N_18683,N_17115,N_17425);
and U18684 (N_18684,N_16707,N_16596);
xnor U18685 (N_18685,N_16937,N_16825);
or U18686 (N_18686,N_16606,N_16614);
and U18687 (N_18687,N_16071,N_17911);
xor U18688 (N_18688,N_17755,N_16276);
or U18689 (N_18689,N_16205,N_17358);
or U18690 (N_18690,N_16336,N_16956);
nor U18691 (N_18691,N_16643,N_16158);
or U18692 (N_18692,N_17156,N_17275);
nand U18693 (N_18693,N_17746,N_16342);
or U18694 (N_18694,N_17540,N_16190);
or U18695 (N_18695,N_17052,N_16765);
nand U18696 (N_18696,N_17532,N_16933);
xnor U18697 (N_18697,N_16840,N_17038);
nor U18698 (N_18698,N_17134,N_16311);
and U18699 (N_18699,N_17064,N_16824);
xor U18700 (N_18700,N_16034,N_17854);
nand U18701 (N_18701,N_16890,N_16904);
nand U18702 (N_18702,N_17948,N_16454);
and U18703 (N_18703,N_16113,N_16810);
and U18704 (N_18704,N_16064,N_17813);
or U18705 (N_18705,N_16619,N_17356);
nand U18706 (N_18706,N_17741,N_16902);
or U18707 (N_18707,N_17577,N_16239);
nor U18708 (N_18708,N_17679,N_16819);
or U18709 (N_18709,N_16924,N_16088);
and U18710 (N_18710,N_16316,N_16967);
nor U18711 (N_18711,N_16347,N_17650);
or U18712 (N_18712,N_16533,N_17380);
nor U18713 (N_18713,N_16727,N_17763);
nor U18714 (N_18714,N_17480,N_17056);
nor U18715 (N_18715,N_16537,N_16228);
or U18716 (N_18716,N_16052,N_16422);
xor U18717 (N_18717,N_17285,N_17913);
nor U18718 (N_18718,N_17340,N_16153);
and U18719 (N_18719,N_17267,N_16135);
nand U18720 (N_18720,N_17528,N_17565);
xnor U18721 (N_18721,N_17602,N_17729);
nor U18722 (N_18722,N_16745,N_17183);
or U18723 (N_18723,N_17045,N_17994);
and U18724 (N_18724,N_17758,N_16488);
and U18725 (N_18725,N_17759,N_17521);
nand U18726 (N_18726,N_17953,N_17727);
nor U18727 (N_18727,N_17173,N_16605);
or U18728 (N_18728,N_16330,N_17675);
and U18729 (N_18729,N_17250,N_16212);
or U18730 (N_18730,N_17882,N_16306);
xnor U18731 (N_18731,N_17262,N_17232);
and U18732 (N_18732,N_16982,N_17110);
or U18733 (N_18733,N_17120,N_16691);
and U18734 (N_18734,N_16185,N_16949);
and U18735 (N_18735,N_17954,N_17107);
xor U18736 (N_18736,N_16803,N_17968);
nand U18737 (N_18737,N_16042,N_17775);
or U18738 (N_18738,N_17062,N_17807);
xor U18739 (N_18739,N_16761,N_17310);
and U18740 (N_18740,N_17335,N_16590);
nor U18741 (N_18741,N_17652,N_17564);
or U18742 (N_18742,N_17034,N_16973);
or U18743 (N_18743,N_16780,N_16046);
or U18744 (N_18744,N_17711,N_17943);
nand U18745 (N_18745,N_17548,N_16990);
and U18746 (N_18746,N_16138,N_17140);
nor U18747 (N_18747,N_16414,N_16667);
nand U18748 (N_18748,N_17554,N_16830);
or U18749 (N_18749,N_17124,N_17850);
nor U18750 (N_18750,N_17108,N_17481);
and U18751 (N_18751,N_16447,N_16194);
xnor U18752 (N_18752,N_16470,N_16321);
or U18753 (N_18753,N_17073,N_17155);
and U18754 (N_18754,N_16895,N_16372);
and U18755 (N_18755,N_17683,N_17258);
and U18756 (N_18756,N_16387,N_17374);
nand U18757 (N_18757,N_16086,N_17006);
nor U18758 (N_18758,N_17902,N_17361);
or U18759 (N_18759,N_16148,N_16609);
nand U18760 (N_18760,N_16799,N_16650);
and U18761 (N_18761,N_16692,N_17014);
and U18762 (N_18762,N_16134,N_16501);
nand U18763 (N_18763,N_17983,N_17166);
or U18764 (N_18764,N_16683,N_16209);
nand U18765 (N_18765,N_16455,N_17703);
xor U18766 (N_18766,N_17812,N_17799);
or U18767 (N_18767,N_17611,N_17487);
and U18768 (N_18768,N_17701,N_16663);
or U18769 (N_18769,N_17388,N_17201);
and U18770 (N_18770,N_16710,N_17966);
nor U18771 (N_18771,N_16641,N_16325);
and U18772 (N_18772,N_17048,N_16726);
nor U18773 (N_18773,N_17595,N_17751);
nor U18774 (N_18774,N_16177,N_16720);
nand U18775 (N_18775,N_16783,N_16441);
and U18776 (N_18776,N_16732,N_17633);
and U18777 (N_18777,N_16897,N_17348);
nor U18778 (N_18778,N_17928,N_17597);
xor U18779 (N_18779,N_16510,N_16659);
nor U18780 (N_18780,N_17545,N_17320);
or U18781 (N_18781,N_16755,N_16865);
or U18782 (N_18782,N_17825,N_16150);
or U18783 (N_18783,N_16729,N_17205);
or U18784 (N_18784,N_17008,N_16152);
or U18785 (N_18785,N_17126,N_16343);
nor U18786 (N_18786,N_16215,N_17035);
and U18787 (N_18787,N_17321,N_16854);
or U18788 (N_18788,N_16335,N_17646);
nand U18789 (N_18789,N_16672,N_17431);
nor U18790 (N_18790,N_17242,N_16355);
nand U18791 (N_18791,N_16861,N_16014);
or U18792 (N_18792,N_17847,N_16964);
and U18793 (N_18793,N_17542,N_17466);
and U18794 (N_18794,N_17176,N_16061);
nor U18795 (N_18795,N_16626,N_16426);
or U18796 (N_18796,N_17985,N_16291);
nor U18797 (N_18797,N_17422,N_17940);
nor U18798 (N_18798,N_17097,N_17040);
and U18799 (N_18799,N_16438,N_17687);
nor U18800 (N_18800,N_16944,N_17693);
nor U18801 (N_18801,N_16502,N_17400);
nor U18802 (N_18802,N_16457,N_16495);
nand U18803 (N_18803,N_16367,N_17423);
and U18804 (N_18804,N_16334,N_17263);
or U18805 (N_18805,N_17861,N_16090);
xor U18806 (N_18806,N_16738,N_17121);
and U18807 (N_18807,N_17363,N_16653);
and U18808 (N_18808,N_17341,N_16733);
xor U18809 (N_18809,N_17334,N_17098);
or U18810 (N_18810,N_16754,N_16995);
and U18811 (N_18811,N_17888,N_16784);
xnor U18812 (N_18812,N_16002,N_17766);
nor U18813 (N_18813,N_16012,N_16808);
xnor U18814 (N_18814,N_17885,N_17387);
and U18815 (N_18815,N_16610,N_17489);
or U18816 (N_18816,N_16941,N_17104);
nor U18817 (N_18817,N_17326,N_17583);
or U18818 (N_18818,N_17689,N_16391);
and U18819 (N_18819,N_17135,N_16581);
nor U18820 (N_18820,N_17138,N_17109);
and U18821 (N_18821,N_16574,N_16993);
or U18822 (N_18822,N_17628,N_17015);
nor U18823 (N_18823,N_16584,N_16947);
or U18824 (N_18824,N_16957,N_16970);
xor U18825 (N_18825,N_17901,N_17118);
and U18826 (N_18826,N_16790,N_16111);
nor U18827 (N_18827,N_17616,N_17970);
or U18828 (N_18828,N_17871,N_16119);
and U18829 (N_18829,N_16453,N_16821);
or U18830 (N_18830,N_16280,N_16603);
or U18831 (N_18831,N_16182,N_17744);
xnor U18832 (N_18832,N_16903,N_17273);
and U18833 (N_18833,N_17771,N_16677);
or U18834 (N_18834,N_17170,N_17923);
or U18835 (N_18835,N_17359,N_16232);
nand U18836 (N_18836,N_16688,N_17198);
or U18837 (N_18837,N_16899,N_17130);
nand U18838 (N_18838,N_17294,N_17414);
or U18839 (N_18839,N_16310,N_16022);
or U18840 (N_18840,N_16879,N_16697);
or U18841 (N_18841,N_16383,N_17717);
nand U18842 (N_18842,N_17635,N_16728);
nor U18843 (N_18843,N_17570,N_17503);
nand U18844 (N_18844,N_16962,N_16690);
nand U18845 (N_18845,N_17116,N_17342);
and U18846 (N_18846,N_16705,N_16484);
nor U18847 (N_18847,N_17312,N_16656);
nand U18848 (N_18848,N_17248,N_16834);
and U18849 (N_18849,N_16759,N_17590);
nor U18850 (N_18850,N_16282,N_17366);
and U18851 (N_18851,N_17896,N_16312);
nand U18852 (N_18852,N_16570,N_17877);
nor U18853 (N_18853,N_17608,N_17631);
or U18854 (N_18854,N_17529,N_16886);
or U18855 (N_18855,N_17192,N_17343);
nor U18856 (N_18856,N_17704,N_16245);
and U18857 (N_18857,N_17713,N_16971);
nor U18858 (N_18858,N_17695,N_17991);
and U18859 (N_18859,N_17593,N_17798);
or U18860 (N_18860,N_16826,N_16128);
xor U18861 (N_18861,N_17429,N_16679);
and U18862 (N_18862,N_17373,N_17836);
nor U18863 (N_18863,N_17437,N_16413);
xnor U18864 (N_18864,N_17346,N_16545);
or U18865 (N_18865,N_16168,N_16295);
nand U18866 (N_18866,N_16507,N_16027);
xor U18867 (N_18867,N_16240,N_16345);
xor U18868 (N_18868,N_16616,N_16546);
or U18869 (N_18869,N_17642,N_16045);
nor U18870 (N_18870,N_17386,N_16040);
xor U18871 (N_18871,N_17228,N_17645);
and U18872 (N_18872,N_17096,N_16285);
or U18873 (N_18873,N_17378,N_16889);
and U18874 (N_18874,N_17162,N_17600);
nor U18875 (N_18875,N_16035,N_16913);
nand U18876 (N_18876,N_17223,N_17392);
nor U18877 (N_18877,N_16664,N_16053);
nor U18878 (N_18878,N_17615,N_17796);
nor U18879 (N_18879,N_16638,N_16863);
nor U18880 (N_18880,N_16444,N_17835);
or U18881 (N_18881,N_17682,N_16235);
nand U18882 (N_18882,N_16263,N_17229);
and U18883 (N_18883,N_17072,N_16778);
and U18884 (N_18884,N_17797,N_16996);
nand U18885 (N_18885,N_17659,N_17171);
or U18886 (N_18886,N_17510,N_17749);
xnor U18887 (N_18887,N_17282,N_16360);
or U18888 (N_18888,N_16521,N_17538);
nor U18889 (N_18889,N_17399,N_17989);
and U18890 (N_18890,N_17153,N_17903);
xnor U18891 (N_18891,N_17811,N_17279);
nor U18892 (N_18892,N_16698,N_16722);
xnor U18893 (N_18893,N_16203,N_17516);
nand U18894 (N_18894,N_16468,N_16802);
xnor U18895 (N_18895,N_16430,N_16472);
nor U18896 (N_18896,N_16028,N_17585);
or U18897 (N_18897,N_17070,N_17641);
xor U18898 (N_18898,N_17125,N_16262);
nor U18899 (N_18899,N_16694,N_17426);
and U18900 (N_18900,N_17347,N_17724);
nand U18901 (N_18901,N_16779,N_16647);
and U18902 (N_18902,N_16514,N_17686);
or U18903 (N_18903,N_17838,N_16544);
and U18904 (N_18904,N_16084,N_16541);
and U18905 (N_18905,N_16146,N_16633);
nand U18906 (N_18906,N_17580,N_16512);
or U18907 (N_18907,N_17086,N_17209);
nand U18908 (N_18908,N_17546,N_17581);
nor U18909 (N_18909,N_16637,N_16428);
and U18910 (N_18910,N_16070,N_16307);
nand U18911 (N_18911,N_16181,N_17815);
nor U18912 (N_18912,N_16520,N_17003);
nand U18913 (N_18913,N_16300,N_17085);
nor U18914 (N_18914,N_17199,N_17587);
or U18915 (N_18915,N_17307,N_17553);
xnor U18916 (N_18916,N_16473,N_17152);
or U18917 (N_18917,N_16242,N_17946);
or U18918 (N_18918,N_17662,N_17950);
or U18919 (N_18919,N_17012,N_17355);
or U18920 (N_18920,N_16747,N_17444);
nand U18921 (N_18921,N_17079,N_17336);
or U18922 (N_18922,N_16547,N_16548);
nand U18923 (N_18923,N_16896,N_16057);
nand U18924 (N_18924,N_16348,N_16888);
nor U18925 (N_18925,N_17819,N_17900);
nand U18926 (N_18926,N_16275,N_16835);
or U18927 (N_18927,N_17556,N_17080);
and U18928 (N_18928,N_17291,N_17857);
nor U18929 (N_18929,N_17011,N_17525);
xor U18930 (N_18930,N_16592,N_16163);
nand U18931 (N_18931,N_16021,N_16144);
nor U18932 (N_18932,N_17840,N_17063);
or U18933 (N_18933,N_17071,N_17978);
nand U18934 (N_18934,N_16016,N_16800);
or U18935 (N_18935,N_17379,N_16072);
nand U18936 (N_18936,N_16364,N_16109);
nand U18937 (N_18937,N_17025,N_17772);
nand U18938 (N_18938,N_17182,N_16356);
or U18939 (N_18939,N_17956,N_16350);
nor U18940 (N_18940,N_16480,N_16268);
nand U18941 (N_18941,N_16384,N_16839);
nor U18942 (N_18942,N_16151,N_17800);
or U18943 (N_18943,N_16091,N_17872);
xnor U18944 (N_18944,N_16954,N_17059);
nand U18945 (N_18945,N_17053,N_17474);
and U18946 (N_18946,N_17272,N_16721);
nor U18947 (N_18947,N_16742,N_16764);
nand U18948 (N_18948,N_16233,N_17690);
nand U18949 (N_18949,N_17239,N_17821);
and U18950 (N_18950,N_16434,N_16540);
or U18951 (N_18951,N_16640,N_17904);
xnor U18952 (N_18952,N_17305,N_17715);
nor U18953 (N_18953,N_16882,N_16317);
nor U18954 (N_18954,N_16329,N_16361);
nand U18955 (N_18955,N_17757,N_17822);
nor U18956 (N_18956,N_16685,N_16875);
nand U18957 (N_18957,N_16977,N_16346);
nand U18958 (N_18958,N_17128,N_17674);
nand U18959 (N_18959,N_16724,N_17676);
or U18960 (N_18960,N_17505,N_16622);
or U18961 (N_18961,N_17023,N_16551);
or U18962 (N_18962,N_16887,N_16744);
nor U18963 (N_18963,N_17268,N_16377);
and U18964 (N_18964,N_16298,N_16105);
nor U18965 (N_18965,N_16966,N_17224);
nand U18966 (N_18966,N_16149,N_16696);
nor U18967 (N_18967,N_16277,N_16173);
or U18968 (N_18968,N_17522,N_16608);
and U18969 (N_18969,N_16676,N_17833);
and U18970 (N_18970,N_16253,N_16595);
nand U18971 (N_18971,N_16318,N_17296);
nor U18972 (N_18972,N_17508,N_16159);
nor U18973 (N_18973,N_17123,N_16517);
nand U18974 (N_18974,N_17459,N_16060);
nand U18975 (N_18975,N_16926,N_16089);
nor U18976 (N_18976,N_16029,N_17475);
and U18977 (N_18977,N_16844,N_17987);
or U18978 (N_18978,N_16530,N_17337);
and U18979 (N_18979,N_16201,N_16136);
or U18980 (N_18980,N_17731,N_16952);
or U18981 (N_18981,N_16953,N_17623);
nor U18982 (N_18982,N_17074,N_16629);
nor U18983 (N_18983,N_16901,N_17986);
or U18984 (N_18984,N_16847,N_16931);
nand U18985 (N_18985,N_16069,N_16328);
nor U18986 (N_18986,N_17613,N_16758);
nand U18987 (N_18987,N_16503,N_17658);
nand U18988 (N_18988,N_16634,N_16085);
nand U18989 (N_18989,N_16550,N_17906);
or U18990 (N_18990,N_16108,N_16170);
nand U18991 (N_18991,N_17301,N_17375);
nor U18992 (N_18992,N_16466,N_17876);
nand U18993 (N_18993,N_17415,N_16251);
and U18994 (N_18994,N_16767,N_16708);
and U18995 (N_18995,N_17446,N_17660);
nor U18996 (N_18996,N_17743,N_16832);
and U18997 (N_18997,N_17451,N_16322);
nand U18998 (N_18998,N_16114,N_17406);
or U18999 (N_18999,N_16005,N_16922);
nor U19000 (N_19000,N_16997,N_16719);
nand U19001 (N_19001,N_16623,N_16227);
nand U19002 (N_19002,N_16117,N_17841);
nand U19003 (N_19003,N_17937,N_16820);
and U19004 (N_19004,N_17631,N_17027);
nand U19005 (N_19005,N_16260,N_16241);
or U19006 (N_19006,N_17804,N_17933);
or U19007 (N_19007,N_17406,N_17933);
and U19008 (N_19008,N_17944,N_17469);
or U19009 (N_19009,N_17589,N_17459);
nor U19010 (N_19010,N_17734,N_16403);
and U19011 (N_19011,N_17834,N_17452);
nor U19012 (N_19012,N_16770,N_16159);
and U19013 (N_19013,N_16608,N_17781);
nor U19014 (N_19014,N_16476,N_16660);
or U19015 (N_19015,N_16543,N_17959);
or U19016 (N_19016,N_16581,N_17348);
nor U19017 (N_19017,N_17922,N_16099);
or U19018 (N_19018,N_17853,N_17189);
and U19019 (N_19019,N_17512,N_17395);
xor U19020 (N_19020,N_17900,N_16883);
or U19021 (N_19021,N_16668,N_16056);
nand U19022 (N_19022,N_17717,N_16631);
and U19023 (N_19023,N_16661,N_16134);
nand U19024 (N_19024,N_17322,N_17209);
or U19025 (N_19025,N_16152,N_17529);
or U19026 (N_19026,N_16856,N_17682);
and U19027 (N_19027,N_16315,N_17925);
nand U19028 (N_19028,N_17777,N_17504);
nand U19029 (N_19029,N_17781,N_17755);
or U19030 (N_19030,N_16525,N_16737);
or U19031 (N_19031,N_17812,N_17703);
nor U19032 (N_19032,N_16275,N_16223);
nand U19033 (N_19033,N_17291,N_17495);
nor U19034 (N_19034,N_16410,N_16861);
nand U19035 (N_19035,N_17648,N_17604);
nor U19036 (N_19036,N_17896,N_16426);
and U19037 (N_19037,N_17298,N_16361);
nand U19038 (N_19038,N_16614,N_16919);
xor U19039 (N_19039,N_16743,N_17777);
or U19040 (N_19040,N_16586,N_16118);
and U19041 (N_19041,N_17593,N_16900);
nand U19042 (N_19042,N_16424,N_17259);
and U19043 (N_19043,N_16718,N_16661);
xor U19044 (N_19044,N_17658,N_17822);
nor U19045 (N_19045,N_16771,N_16712);
and U19046 (N_19046,N_16373,N_16846);
or U19047 (N_19047,N_16696,N_16670);
nand U19048 (N_19048,N_16921,N_17143);
and U19049 (N_19049,N_17584,N_16786);
or U19050 (N_19050,N_16091,N_17665);
nor U19051 (N_19051,N_16646,N_16546);
nor U19052 (N_19052,N_16202,N_17101);
nor U19053 (N_19053,N_17800,N_16612);
and U19054 (N_19054,N_17750,N_16904);
nor U19055 (N_19055,N_17694,N_17992);
or U19056 (N_19056,N_17283,N_17427);
nand U19057 (N_19057,N_16440,N_16712);
and U19058 (N_19058,N_16692,N_17836);
xor U19059 (N_19059,N_16740,N_17199);
nor U19060 (N_19060,N_17543,N_17452);
nor U19061 (N_19061,N_16213,N_16503);
nand U19062 (N_19062,N_17942,N_16629);
xnor U19063 (N_19063,N_17747,N_16787);
or U19064 (N_19064,N_16015,N_16832);
nand U19065 (N_19065,N_16405,N_16015);
or U19066 (N_19066,N_17923,N_16977);
or U19067 (N_19067,N_17682,N_16861);
nand U19068 (N_19068,N_17433,N_16179);
and U19069 (N_19069,N_17624,N_17467);
nor U19070 (N_19070,N_17811,N_16689);
nor U19071 (N_19071,N_17398,N_17667);
or U19072 (N_19072,N_17351,N_17943);
or U19073 (N_19073,N_17216,N_16556);
nand U19074 (N_19074,N_16823,N_16909);
nor U19075 (N_19075,N_16210,N_16734);
nand U19076 (N_19076,N_16851,N_16205);
or U19077 (N_19077,N_17226,N_16404);
nor U19078 (N_19078,N_17821,N_17405);
or U19079 (N_19079,N_16576,N_16137);
or U19080 (N_19080,N_17133,N_17622);
xor U19081 (N_19081,N_16687,N_17726);
or U19082 (N_19082,N_16368,N_16952);
and U19083 (N_19083,N_17316,N_16108);
nor U19084 (N_19084,N_17688,N_17476);
nand U19085 (N_19085,N_17214,N_16731);
and U19086 (N_19086,N_16192,N_16679);
and U19087 (N_19087,N_17769,N_16826);
or U19088 (N_19088,N_17935,N_17916);
nand U19089 (N_19089,N_16718,N_16512);
nor U19090 (N_19090,N_16663,N_17197);
nand U19091 (N_19091,N_17655,N_17932);
nor U19092 (N_19092,N_17027,N_16916);
or U19093 (N_19093,N_17605,N_16498);
nand U19094 (N_19094,N_16088,N_16413);
xnor U19095 (N_19095,N_17105,N_17016);
nand U19096 (N_19096,N_17822,N_17430);
nand U19097 (N_19097,N_17681,N_16718);
and U19098 (N_19098,N_17525,N_16751);
and U19099 (N_19099,N_17039,N_17066);
nor U19100 (N_19100,N_17690,N_16584);
or U19101 (N_19101,N_17229,N_17977);
nand U19102 (N_19102,N_16972,N_16250);
or U19103 (N_19103,N_16892,N_16531);
nand U19104 (N_19104,N_17575,N_16434);
and U19105 (N_19105,N_16343,N_16266);
nor U19106 (N_19106,N_17627,N_17543);
and U19107 (N_19107,N_16308,N_16760);
xor U19108 (N_19108,N_16532,N_17551);
and U19109 (N_19109,N_16264,N_17186);
nand U19110 (N_19110,N_16808,N_16748);
and U19111 (N_19111,N_16461,N_16526);
nand U19112 (N_19112,N_16168,N_16845);
nand U19113 (N_19113,N_16591,N_16223);
and U19114 (N_19114,N_17471,N_16041);
nand U19115 (N_19115,N_16603,N_17108);
or U19116 (N_19116,N_16723,N_16264);
xor U19117 (N_19117,N_16911,N_16747);
and U19118 (N_19118,N_17015,N_17384);
xnor U19119 (N_19119,N_17835,N_17385);
and U19120 (N_19120,N_17795,N_17652);
xor U19121 (N_19121,N_17676,N_17043);
xor U19122 (N_19122,N_16041,N_17015);
nor U19123 (N_19123,N_16857,N_17492);
or U19124 (N_19124,N_16067,N_16259);
or U19125 (N_19125,N_16440,N_17916);
or U19126 (N_19126,N_16680,N_16007);
and U19127 (N_19127,N_16451,N_16678);
or U19128 (N_19128,N_17359,N_17762);
nand U19129 (N_19129,N_17325,N_17750);
nor U19130 (N_19130,N_16193,N_16282);
nand U19131 (N_19131,N_17448,N_16332);
xnor U19132 (N_19132,N_16239,N_16277);
xnor U19133 (N_19133,N_16286,N_17846);
and U19134 (N_19134,N_16239,N_16203);
and U19135 (N_19135,N_17588,N_16858);
nor U19136 (N_19136,N_17709,N_16118);
or U19137 (N_19137,N_16446,N_17527);
and U19138 (N_19138,N_17239,N_17262);
and U19139 (N_19139,N_17497,N_17241);
nor U19140 (N_19140,N_16289,N_16949);
nor U19141 (N_19141,N_17888,N_17570);
nor U19142 (N_19142,N_17874,N_16305);
nor U19143 (N_19143,N_16864,N_16370);
and U19144 (N_19144,N_17799,N_17294);
or U19145 (N_19145,N_17261,N_17606);
or U19146 (N_19146,N_16071,N_16839);
nand U19147 (N_19147,N_16176,N_17153);
nand U19148 (N_19148,N_17027,N_17378);
or U19149 (N_19149,N_17606,N_16925);
or U19150 (N_19150,N_16916,N_17407);
or U19151 (N_19151,N_17589,N_16921);
nand U19152 (N_19152,N_16504,N_16328);
and U19153 (N_19153,N_16904,N_17113);
and U19154 (N_19154,N_17457,N_16479);
nor U19155 (N_19155,N_17896,N_16713);
or U19156 (N_19156,N_17890,N_17102);
xor U19157 (N_19157,N_17846,N_17784);
nor U19158 (N_19158,N_16294,N_17945);
and U19159 (N_19159,N_16670,N_17928);
nand U19160 (N_19160,N_16029,N_17650);
nand U19161 (N_19161,N_17829,N_17418);
and U19162 (N_19162,N_17686,N_17383);
or U19163 (N_19163,N_16269,N_17736);
and U19164 (N_19164,N_17552,N_17325);
or U19165 (N_19165,N_16241,N_16932);
nand U19166 (N_19166,N_16397,N_16333);
nor U19167 (N_19167,N_16858,N_16313);
nand U19168 (N_19168,N_16904,N_17518);
or U19169 (N_19169,N_17717,N_17800);
and U19170 (N_19170,N_16318,N_17388);
nor U19171 (N_19171,N_16125,N_16568);
nand U19172 (N_19172,N_16659,N_16626);
nor U19173 (N_19173,N_16326,N_16101);
nor U19174 (N_19174,N_17315,N_17810);
and U19175 (N_19175,N_17808,N_17701);
and U19176 (N_19176,N_16417,N_16270);
nor U19177 (N_19177,N_16712,N_17638);
nand U19178 (N_19178,N_17173,N_16881);
nor U19179 (N_19179,N_17182,N_16407);
and U19180 (N_19180,N_17018,N_16728);
or U19181 (N_19181,N_17062,N_17185);
or U19182 (N_19182,N_16067,N_16012);
nor U19183 (N_19183,N_17637,N_16168);
xnor U19184 (N_19184,N_17961,N_17936);
and U19185 (N_19185,N_16211,N_17102);
nand U19186 (N_19186,N_17750,N_17393);
or U19187 (N_19187,N_17255,N_16381);
nand U19188 (N_19188,N_17395,N_16894);
nand U19189 (N_19189,N_16937,N_16275);
or U19190 (N_19190,N_16504,N_16426);
or U19191 (N_19191,N_17993,N_16201);
nand U19192 (N_19192,N_16446,N_16890);
nor U19193 (N_19193,N_17649,N_17445);
and U19194 (N_19194,N_17428,N_16850);
or U19195 (N_19195,N_16658,N_17671);
or U19196 (N_19196,N_17858,N_17443);
or U19197 (N_19197,N_17554,N_16517);
and U19198 (N_19198,N_16110,N_17399);
nor U19199 (N_19199,N_16420,N_17377);
or U19200 (N_19200,N_17991,N_16023);
nand U19201 (N_19201,N_17310,N_17283);
nor U19202 (N_19202,N_16275,N_16444);
and U19203 (N_19203,N_16471,N_16868);
or U19204 (N_19204,N_16673,N_17690);
nor U19205 (N_19205,N_16817,N_16226);
nand U19206 (N_19206,N_17467,N_16291);
or U19207 (N_19207,N_17921,N_16791);
nor U19208 (N_19208,N_17194,N_16551);
and U19209 (N_19209,N_17348,N_17967);
nand U19210 (N_19210,N_17077,N_17604);
nand U19211 (N_19211,N_17280,N_16170);
or U19212 (N_19212,N_16297,N_16090);
nor U19213 (N_19213,N_17993,N_17508);
nor U19214 (N_19214,N_16094,N_16554);
or U19215 (N_19215,N_16010,N_16694);
or U19216 (N_19216,N_16260,N_16617);
or U19217 (N_19217,N_16247,N_17362);
nand U19218 (N_19218,N_17975,N_16082);
and U19219 (N_19219,N_17701,N_17405);
nand U19220 (N_19220,N_17626,N_17308);
nor U19221 (N_19221,N_16344,N_16932);
and U19222 (N_19222,N_17477,N_17620);
nor U19223 (N_19223,N_17817,N_17814);
and U19224 (N_19224,N_16506,N_17046);
or U19225 (N_19225,N_16149,N_17754);
or U19226 (N_19226,N_17923,N_17912);
nand U19227 (N_19227,N_16499,N_16602);
xor U19228 (N_19228,N_16218,N_17463);
and U19229 (N_19229,N_16078,N_16907);
or U19230 (N_19230,N_16484,N_17449);
and U19231 (N_19231,N_17092,N_16786);
and U19232 (N_19232,N_17725,N_17147);
or U19233 (N_19233,N_17557,N_17568);
or U19234 (N_19234,N_17083,N_16285);
or U19235 (N_19235,N_17483,N_17025);
or U19236 (N_19236,N_17158,N_17023);
or U19237 (N_19237,N_17627,N_17368);
or U19238 (N_19238,N_16461,N_16854);
or U19239 (N_19239,N_16253,N_17940);
or U19240 (N_19240,N_16303,N_17266);
nor U19241 (N_19241,N_16648,N_16748);
nor U19242 (N_19242,N_17365,N_17939);
nand U19243 (N_19243,N_17613,N_16870);
or U19244 (N_19244,N_16225,N_17365);
and U19245 (N_19245,N_16057,N_17635);
nand U19246 (N_19246,N_17345,N_17844);
and U19247 (N_19247,N_17941,N_16848);
nor U19248 (N_19248,N_16861,N_16129);
xnor U19249 (N_19249,N_16373,N_16838);
or U19250 (N_19250,N_16544,N_16818);
or U19251 (N_19251,N_16755,N_17494);
or U19252 (N_19252,N_16696,N_17411);
nand U19253 (N_19253,N_17109,N_16374);
nand U19254 (N_19254,N_17341,N_16645);
nor U19255 (N_19255,N_17502,N_17442);
or U19256 (N_19256,N_16759,N_16502);
and U19257 (N_19257,N_17534,N_17867);
nand U19258 (N_19258,N_17937,N_16561);
xnor U19259 (N_19259,N_17191,N_17962);
or U19260 (N_19260,N_17226,N_17797);
nand U19261 (N_19261,N_17366,N_17007);
or U19262 (N_19262,N_16260,N_17341);
and U19263 (N_19263,N_17896,N_17954);
or U19264 (N_19264,N_17689,N_17807);
nor U19265 (N_19265,N_17757,N_17333);
xnor U19266 (N_19266,N_16281,N_17056);
nand U19267 (N_19267,N_16757,N_17098);
nor U19268 (N_19268,N_17976,N_17892);
and U19269 (N_19269,N_17481,N_16478);
nor U19270 (N_19270,N_16007,N_17592);
nor U19271 (N_19271,N_17554,N_17876);
and U19272 (N_19272,N_17432,N_17897);
nand U19273 (N_19273,N_16749,N_16086);
nand U19274 (N_19274,N_16013,N_16737);
xor U19275 (N_19275,N_17842,N_16960);
and U19276 (N_19276,N_16256,N_17323);
nor U19277 (N_19277,N_16136,N_16865);
xnor U19278 (N_19278,N_16007,N_17528);
and U19279 (N_19279,N_16481,N_16055);
nand U19280 (N_19280,N_16932,N_17652);
nand U19281 (N_19281,N_17106,N_16847);
nand U19282 (N_19282,N_16858,N_17627);
or U19283 (N_19283,N_16715,N_16285);
xnor U19284 (N_19284,N_16720,N_17055);
and U19285 (N_19285,N_16185,N_16758);
and U19286 (N_19286,N_16398,N_16359);
xnor U19287 (N_19287,N_17718,N_17154);
or U19288 (N_19288,N_17016,N_17100);
or U19289 (N_19289,N_16256,N_16219);
nand U19290 (N_19290,N_17385,N_16147);
and U19291 (N_19291,N_17429,N_16325);
and U19292 (N_19292,N_16817,N_17593);
nor U19293 (N_19293,N_17345,N_17427);
nand U19294 (N_19294,N_16195,N_17673);
or U19295 (N_19295,N_16619,N_16666);
nand U19296 (N_19296,N_16666,N_17224);
and U19297 (N_19297,N_17593,N_16323);
xor U19298 (N_19298,N_16978,N_17866);
and U19299 (N_19299,N_17898,N_17333);
nand U19300 (N_19300,N_16108,N_17431);
and U19301 (N_19301,N_17896,N_17689);
and U19302 (N_19302,N_17196,N_17910);
xnor U19303 (N_19303,N_17552,N_17420);
or U19304 (N_19304,N_17207,N_17647);
nor U19305 (N_19305,N_17199,N_16533);
or U19306 (N_19306,N_16230,N_16401);
nor U19307 (N_19307,N_17661,N_16243);
and U19308 (N_19308,N_17184,N_17031);
and U19309 (N_19309,N_17959,N_16308);
nor U19310 (N_19310,N_16208,N_17120);
and U19311 (N_19311,N_17526,N_16503);
nand U19312 (N_19312,N_17444,N_17076);
nand U19313 (N_19313,N_17175,N_16072);
nand U19314 (N_19314,N_17205,N_17504);
nor U19315 (N_19315,N_16470,N_16890);
and U19316 (N_19316,N_16214,N_16882);
nor U19317 (N_19317,N_16285,N_17994);
and U19318 (N_19318,N_16309,N_16938);
nor U19319 (N_19319,N_16347,N_16340);
xor U19320 (N_19320,N_16146,N_17665);
or U19321 (N_19321,N_17830,N_16675);
and U19322 (N_19322,N_17920,N_16265);
xnor U19323 (N_19323,N_16509,N_16326);
nand U19324 (N_19324,N_17449,N_17588);
nand U19325 (N_19325,N_17004,N_16832);
nand U19326 (N_19326,N_16105,N_17484);
and U19327 (N_19327,N_17378,N_17872);
or U19328 (N_19328,N_17866,N_16728);
nor U19329 (N_19329,N_17844,N_17609);
nand U19330 (N_19330,N_17676,N_17037);
nand U19331 (N_19331,N_16567,N_16406);
and U19332 (N_19332,N_16849,N_16250);
nand U19333 (N_19333,N_16773,N_16441);
and U19334 (N_19334,N_16379,N_16815);
or U19335 (N_19335,N_17651,N_17777);
nor U19336 (N_19336,N_17697,N_17322);
and U19337 (N_19337,N_17469,N_16214);
or U19338 (N_19338,N_17310,N_17225);
nand U19339 (N_19339,N_16367,N_16311);
nor U19340 (N_19340,N_17862,N_16776);
nor U19341 (N_19341,N_17763,N_16848);
nor U19342 (N_19342,N_16939,N_16167);
nand U19343 (N_19343,N_17622,N_17056);
or U19344 (N_19344,N_16066,N_16632);
and U19345 (N_19345,N_16555,N_16945);
or U19346 (N_19346,N_16695,N_16528);
xor U19347 (N_19347,N_16309,N_16805);
nor U19348 (N_19348,N_17368,N_17593);
nand U19349 (N_19349,N_16162,N_17751);
and U19350 (N_19350,N_17563,N_17160);
xnor U19351 (N_19351,N_16083,N_17372);
and U19352 (N_19352,N_17820,N_16998);
nand U19353 (N_19353,N_17542,N_17511);
or U19354 (N_19354,N_17667,N_17195);
nand U19355 (N_19355,N_17372,N_16569);
nand U19356 (N_19356,N_17842,N_17493);
nor U19357 (N_19357,N_16346,N_17159);
nand U19358 (N_19358,N_16764,N_17707);
and U19359 (N_19359,N_17567,N_17304);
or U19360 (N_19360,N_17615,N_17633);
nand U19361 (N_19361,N_17200,N_16105);
nor U19362 (N_19362,N_17476,N_16889);
and U19363 (N_19363,N_17094,N_16607);
nand U19364 (N_19364,N_17418,N_17604);
and U19365 (N_19365,N_16833,N_17171);
or U19366 (N_19366,N_17870,N_17978);
nor U19367 (N_19367,N_16711,N_17500);
nand U19368 (N_19368,N_17187,N_17432);
or U19369 (N_19369,N_16850,N_16078);
nor U19370 (N_19370,N_16658,N_17001);
xnor U19371 (N_19371,N_17715,N_16262);
xor U19372 (N_19372,N_17273,N_17712);
nor U19373 (N_19373,N_16845,N_16609);
xor U19374 (N_19374,N_17739,N_17783);
xnor U19375 (N_19375,N_17751,N_16490);
nor U19376 (N_19376,N_17649,N_16070);
or U19377 (N_19377,N_17480,N_17209);
nand U19378 (N_19378,N_17748,N_16978);
nand U19379 (N_19379,N_17264,N_17424);
nand U19380 (N_19380,N_17623,N_17840);
and U19381 (N_19381,N_17575,N_16335);
nor U19382 (N_19382,N_17547,N_16906);
nand U19383 (N_19383,N_17876,N_17428);
nor U19384 (N_19384,N_16035,N_16663);
nor U19385 (N_19385,N_17606,N_16486);
nand U19386 (N_19386,N_16999,N_17172);
and U19387 (N_19387,N_17221,N_17803);
nor U19388 (N_19388,N_16239,N_16415);
nor U19389 (N_19389,N_17538,N_17956);
nor U19390 (N_19390,N_17550,N_17958);
xor U19391 (N_19391,N_17565,N_17247);
and U19392 (N_19392,N_17670,N_17632);
and U19393 (N_19393,N_16838,N_16790);
nor U19394 (N_19394,N_16650,N_16762);
nor U19395 (N_19395,N_16013,N_17268);
or U19396 (N_19396,N_17761,N_16662);
nand U19397 (N_19397,N_17383,N_17243);
nand U19398 (N_19398,N_17185,N_17217);
xnor U19399 (N_19399,N_17117,N_16633);
xor U19400 (N_19400,N_17444,N_17560);
nand U19401 (N_19401,N_17808,N_16424);
nand U19402 (N_19402,N_17194,N_17133);
nand U19403 (N_19403,N_17622,N_17127);
nand U19404 (N_19404,N_16123,N_17717);
nor U19405 (N_19405,N_16147,N_17044);
or U19406 (N_19406,N_17746,N_16005);
or U19407 (N_19407,N_16103,N_17901);
or U19408 (N_19408,N_17730,N_16814);
or U19409 (N_19409,N_17080,N_16768);
nor U19410 (N_19410,N_17913,N_16882);
nor U19411 (N_19411,N_17980,N_17986);
nor U19412 (N_19412,N_17813,N_17911);
and U19413 (N_19413,N_17387,N_17347);
or U19414 (N_19414,N_17751,N_16494);
and U19415 (N_19415,N_17878,N_16727);
or U19416 (N_19416,N_16313,N_16885);
and U19417 (N_19417,N_16655,N_17493);
nor U19418 (N_19418,N_17374,N_17795);
xnor U19419 (N_19419,N_17378,N_16492);
nand U19420 (N_19420,N_16953,N_16525);
nand U19421 (N_19421,N_16538,N_17808);
and U19422 (N_19422,N_16047,N_16927);
nor U19423 (N_19423,N_17080,N_17549);
and U19424 (N_19424,N_17936,N_17600);
nor U19425 (N_19425,N_16641,N_17780);
nand U19426 (N_19426,N_17161,N_16631);
and U19427 (N_19427,N_16848,N_16960);
or U19428 (N_19428,N_16167,N_16044);
and U19429 (N_19429,N_16103,N_16094);
nor U19430 (N_19430,N_17441,N_17638);
nand U19431 (N_19431,N_17330,N_16359);
and U19432 (N_19432,N_17934,N_17432);
or U19433 (N_19433,N_17442,N_17760);
nand U19434 (N_19434,N_17412,N_17913);
xnor U19435 (N_19435,N_16747,N_16282);
nand U19436 (N_19436,N_16727,N_17521);
and U19437 (N_19437,N_16958,N_17387);
and U19438 (N_19438,N_17432,N_16451);
or U19439 (N_19439,N_17463,N_17820);
xor U19440 (N_19440,N_16588,N_16496);
nand U19441 (N_19441,N_17720,N_17499);
or U19442 (N_19442,N_16347,N_16588);
nand U19443 (N_19443,N_17436,N_16157);
or U19444 (N_19444,N_16057,N_16294);
and U19445 (N_19445,N_17352,N_16288);
and U19446 (N_19446,N_17522,N_16927);
nand U19447 (N_19447,N_17957,N_17908);
nand U19448 (N_19448,N_16554,N_17401);
xnor U19449 (N_19449,N_17242,N_17103);
xor U19450 (N_19450,N_16217,N_17926);
xnor U19451 (N_19451,N_16178,N_16336);
nand U19452 (N_19452,N_17581,N_16688);
nor U19453 (N_19453,N_17351,N_17242);
or U19454 (N_19454,N_16967,N_16267);
and U19455 (N_19455,N_17132,N_16790);
or U19456 (N_19456,N_16238,N_16054);
nor U19457 (N_19457,N_17306,N_17648);
nor U19458 (N_19458,N_16692,N_17476);
and U19459 (N_19459,N_16763,N_16923);
xor U19460 (N_19460,N_16247,N_17018);
nor U19461 (N_19461,N_16051,N_17343);
nor U19462 (N_19462,N_17705,N_17914);
and U19463 (N_19463,N_17778,N_17728);
and U19464 (N_19464,N_17330,N_17759);
nand U19465 (N_19465,N_17887,N_17111);
and U19466 (N_19466,N_17654,N_16405);
or U19467 (N_19467,N_17992,N_16067);
nand U19468 (N_19468,N_16654,N_16935);
or U19469 (N_19469,N_16894,N_16061);
nand U19470 (N_19470,N_17366,N_17107);
nand U19471 (N_19471,N_16361,N_17939);
or U19472 (N_19472,N_17068,N_16660);
nor U19473 (N_19473,N_17197,N_16145);
nand U19474 (N_19474,N_16359,N_17733);
or U19475 (N_19475,N_17122,N_16956);
and U19476 (N_19476,N_16360,N_16970);
or U19477 (N_19477,N_17389,N_16313);
or U19478 (N_19478,N_16197,N_17538);
nor U19479 (N_19479,N_17578,N_16283);
nand U19480 (N_19480,N_17337,N_16986);
nor U19481 (N_19481,N_17548,N_17727);
nand U19482 (N_19482,N_17464,N_17206);
or U19483 (N_19483,N_17132,N_17104);
nor U19484 (N_19484,N_16320,N_17764);
and U19485 (N_19485,N_17297,N_16021);
and U19486 (N_19486,N_16156,N_17615);
nor U19487 (N_19487,N_16426,N_17197);
or U19488 (N_19488,N_17255,N_17516);
or U19489 (N_19489,N_16187,N_16185);
and U19490 (N_19490,N_17532,N_17947);
xor U19491 (N_19491,N_17917,N_17762);
and U19492 (N_19492,N_16947,N_17786);
nand U19493 (N_19493,N_17675,N_17923);
nor U19494 (N_19494,N_17789,N_16761);
nor U19495 (N_19495,N_17343,N_16009);
nand U19496 (N_19496,N_16025,N_16287);
and U19497 (N_19497,N_17981,N_17984);
nor U19498 (N_19498,N_16596,N_16053);
nor U19499 (N_19499,N_17265,N_17886);
or U19500 (N_19500,N_16941,N_16525);
xnor U19501 (N_19501,N_16501,N_16342);
nand U19502 (N_19502,N_17261,N_17827);
nand U19503 (N_19503,N_16867,N_16144);
xnor U19504 (N_19504,N_17577,N_16445);
nand U19505 (N_19505,N_17553,N_16907);
nand U19506 (N_19506,N_17616,N_17697);
nor U19507 (N_19507,N_17629,N_16982);
xor U19508 (N_19508,N_16116,N_17005);
or U19509 (N_19509,N_17127,N_17270);
xor U19510 (N_19510,N_16614,N_16330);
or U19511 (N_19511,N_17751,N_16404);
nand U19512 (N_19512,N_16248,N_17178);
or U19513 (N_19513,N_16576,N_16439);
nand U19514 (N_19514,N_17929,N_16540);
and U19515 (N_19515,N_17852,N_16717);
nor U19516 (N_19516,N_16735,N_17622);
or U19517 (N_19517,N_17357,N_17866);
or U19518 (N_19518,N_17596,N_17348);
nor U19519 (N_19519,N_16529,N_16804);
nor U19520 (N_19520,N_16138,N_16276);
nand U19521 (N_19521,N_17664,N_16453);
nor U19522 (N_19522,N_17490,N_16538);
nand U19523 (N_19523,N_16994,N_17353);
nand U19524 (N_19524,N_17416,N_17114);
nand U19525 (N_19525,N_17283,N_16951);
nor U19526 (N_19526,N_17884,N_17356);
nor U19527 (N_19527,N_16576,N_17092);
nor U19528 (N_19528,N_16568,N_16388);
and U19529 (N_19529,N_16920,N_17706);
nor U19530 (N_19530,N_16618,N_17513);
nand U19531 (N_19531,N_17116,N_17784);
xor U19532 (N_19532,N_16668,N_17394);
and U19533 (N_19533,N_17965,N_16689);
or U19534 (N_19534,N_17643,N_17057);
or U19535 (N_19535,N_16278,N_17661);
and U19536 (N_19536,N_16787,N_16381);
nand U19537 (N_19537,N_16636,N_17734);
nor U19538 (N_19538,N_17178,N_16102);
nor U19539 (N_19539,N_17307,N_16523);
nand U19540 (N_19540,N_16471,N_16897);
or U19541 (N_19541,N_16132,N_17279);
xnor U19542 (N_19542,N_16615,N_17200);
and U19543 (N_19543,N_17725,N_16757);
and U19544 (N_19544,N_16303,N_17259);
or U19545 (N_19545,N_17125,N_17465);
nand U19546 (N_19546,N_17186,N_16416);
or U19547 (N_19547,N_17892,N_16559);
or U19548 (N_19548,N_17872,N_17975);
nor U19549 (N_19549,N_17126,N_16458);
nor U19550 (N_19550,N_17443,N_17291);
or U19551 (N_19551,N_16882,N_16348);
and U19552 (N_19552,N_17134,N_16486);
and U19553 (N_19553,N_17706,N_16097);
and U19554 (N_19554,N_17558,N_17081);
nand U19555 (N_19555,N_16457,N_16571);
nand U19556 (N_19556,N_17441,N_17505);
nor U19557 (N_19557,N_16640,N_16143);
and U19558 (N_19558,N_16485,N_17677);
nor U19559 (N_19559,N_17826,N_17181);
nand U19560 (N_19560,N_17018,N_17056);
and U19561 (N_19561,N_17409,N_16322);
nor U19562 (N_19562,N_17913,N_16629);
and U19563 (N_19563,N_16087,N_17986);
and U19564 (N_19564,N_17714,N_16086);
and U19565 (N_19565,N_17653,N_17291);
nor U19566 (N_19566,N_17424,N_17184);
or U19567 (N_19567,N_17105,N_17470);
nor U19568 (N_19568,N_17048,N_17676);
nand U19569 (N_19569,N_17992,N_16908);
xor U19570 (N_19570,N_17953,N_16649);
nand U19571 (N_19571,N_16480,N_16305);
nand U19572 (N_19572,N_16458,N_17766);
nor U19573 (N_19573,N_17836,N_17903);
or U19574 (N_19574,N_17723,N_17730);
nand U19575 (N_19575,N_16126,N_17483);
nand U19576 (N_19576,N_16817,N_17565);
nand U19577 (N_19577,N_16556,N_17029);
or U19578 (N_19578,N_17844,N_17073);
nand U19579 (N_19579,N_17089,N_17932);
and U19580 (N_19580,N_17259,N_16410);
or U19581 (N_19581,N_17679,N_17866);
and U19582 (N_19582,N_17997,N_17236);
or U19583 (N_19583,N_17627,N_16525);
and U19584 (N_19584,N_17615,N_16622);
nand U19585 (N_19585,N_16491,N_16532);
nand U19586 (N_19586,N_17494,N_16146);
or U19587 (N_19587,N_16903,N_17199);
xnor U19588 (N_19588,N_17758,N_17985);
or U19589 (N_19589,N_17171,N_17894);
nor U19590 (N_19590,N_17968,N_17030);
or U19591 (N_19591,N_17425,N_17327);
nand U19592 (N_19592,N_16141,N_17482);
or U19593 (N_19593,N_17935,N_16039);
nor U19594 (N_19594,N_16240,N_17741);
or U19595 (N_19595,N_17295,N_16403);
nand U19596 (N_19596,N_17620,N_17092);
nor U19597 (N_19597,N_17127,N_16121);
and U19598 (N_19598,N_16684,N_17438);
nor U19599 (N_19599,N_17169,N_17806);
nor U19600 (N_19600,N_16741,N_16865);
nor U19601 (N_19601,N_17386,N_17864);
nor U19602 (N_19602,N_17576,N_17546);
or U19603 (N_19603,N_16430,N_17062);
nor U19604 (N_19604,N_16113,N_16867);
or U19605 (N_19605,N_16487,N_17714);
nand U19606 (N_19606,N_16353,N_17852);
nand U19607 (N_19607,N_16797,N_16495);
nand U19608 (N_19608,N_16053,N_17882);
nor U19609 (N_19609,N_16382,N_16855);
xor U19610 (N_19610,N_16280,N_17882);
and U19611 (N_19611,N_16844,N_16112);
and U19612 (N_19612,N_16557,N_17900);
nand U19613 (N_19613,N_17606,N_17785);
nand U19614 (N_19614,N_17486,N_17595);
and U19615 (N_19615,N_17006,N_16860);
or U19616 (N_19616,N_17363,N_16987);
and U19617 (N_19617,N_16052,N_17444);
nor U19618 (N_19618,N_16847,N_16295);
and U19619 (N_19619,N_16204,N_17458);
and U19620 (N_19620,N_16573,N_16261);
and U19621 (N_19621,N_17380,N_17213);
or U19622 (N_19622,N_17628,N_16372);
or U19623 (N_19623,N_16222,N_16325);
and U19624 (N_19624,N_17293,N_17061);
and U19625 (N_19625,N_16909,N_16065);
nor U19626 (N_19626,N_16908,N_16630);
nor U19627 (N_19627,N_17095,N_16854);
nand U19628 (N_19628,N_17140,N_17200);
nor U19629 (N_19629,N_17587,N_17298);
nand U19630 (N_19630,N_17517,N_17647);
and U19631 (N_19631,N_17865,N_16855);
xor U19632 (N_19632,N_17172,N_17064);
or U19633 (N_19633,N_17553,N_17008);
nor U19634 (N_19634,N_16146,N_17767);
nand U19635 (N_19635,N_17506,N_17203);
and U19636 (N_19636,N_16233,N_17045);
nor U19637 (N_19637,N_16896,N_17595);
and U19638 (N_19638,N_17307,N_17859);
and U19639 (N_19639,N_17088,N_17984);
nand U19640 (N_19640,N_16373,N_16001);
nor U19641 (N_19641,N_17478,N_17552);
xor U19642 (N_19642,N_17584,N_17756);
and U19643 (N_19643,N_16823,N_17665);
xor U19644 (N_19644,N_17150,N_16536);
and U19645 (N_19645,N_17359,N_16204);
and U19646 (N_19646,N_17064,N_17028);
or U19647 (N_19647,N_17446,N_17891);
or U19648 (N_19648,N_16241,N_16610);
nand U19649 (N_19649,N_16812,N_17702);
or U19650 (N_19650,N_17641,N_16197);
or U19651 (N_19651,N_16623,N_16521);
and U19652 (N_19652,N_16096,N_17462);
or U19653 (N_19653,N_16517,N_17599);
or U19654 (N_19654,N_16711,N_16931);
and U19655 (N_19655,N_17468,N_17430);
nand U19656 (N_19656,N_16324,N_16677);
or U19657 (N_19657,N_16244,N_17177);
and U19658 (N_19658,N_16389,N_17857);
nor U19659 (N_19659,N_17055,N_17694);
or U19660 (N_19660,N_16497,N_17063);
nand U19661 (N_19661,N_17841,N_16540);
xor U19662 (N_19662,N_16871,N_17337);
or U19663 (N_19663,N_17122,N_16155);
and U19664 (N_19664,N_17435,N_16001);
xor U19665 (N_19665,N_16553,N_17621);
nor U19666 (N_19666,N_16333,N_17903);
nand U19667 (N_19667,N_17838,N_16656);
or U19668 (N_19668,N_16896,N_16895);
or U19669 (N_19669,N_17499,N_17139);
nand U19670 (N_19670,N_16801,N_16460);
and U19671 (N_19671,N_16026,N_17751);
or U19672 (N_19672,N_17001,N_16171);
or U19673 (N_19673,N_17480,N_17768);
or U19674 (N_19674,N_17183,N_17828);
nand U19675 (N_19675,N_16485,N_16183);
nand U19676 (N_19676,N_16279,N_16829);
or U19677 (N_19677,N_17676,N_17084);
xnor U19678 (N_19678,N_17705,N_16352);
nand U19679 (N_19679,N_17607,N_17511);
nand U19680 (N_19680,N_16940,N_16076);
or U19681 (N_19681,N_16736,N_16364);
and U19682 (N_19682,N_17239,N_17034);
nor U19683 (N_19683,N_16161,N_16892);
or U19684 (N_19684,N_16857,N_17259);
nor U19685 (N_19685,N_17572,N_17287);
or U19686 (N_19686,N_16096,N_17381);
nand U19687 (N_19687,N_16672,N_16504);
nand U19688 (N_19688,N_16923,N_16517);
or U19689 (N_19689,N_16202,N_16910);
nand U19690 (N_19690,N_16685,N_17935);
nand U19691 (N_19691,N_16761,N_17003);
and U19692 (N_19692,N_17018,N_17655);
nand U19693 (N_19693,N_16917,N_17926);
and U19694 (N_19694,N_16476,N_17269);
and U19695 (N_19695,N_17581,N_17399);
nand U19696 (N_19696,N_16110,N_17352);
nand U19697 (N_19697,N_17683,N_16273);
nand U19698 (N_19698,N_17786,N_17222);
nand U19699 (N_19699,N_16542,N_16996);
or U19700 (N_19700,N_17737,N_16922);
nand U19701 (N_19701,N_17756,N_17076);
xnor U19702 (N_19702,N_16671,N_16020);
and U19703 (N_19703,N_16891,N_17144);
nand U19704 (N_19704,N_17361,N_16814);
nand U19705 (N_19705,N_17705,N_16421);
nor U19706 (N_19706,N_17600,N_16368);
nand U19707 (N_19707,N_16940,N_17127);
xnor U19708 (N_19708,N_16975,N_17535);
nand U19709 (N_19709,N_17019,N_16766);
and U19710 (N_19710,N_16681,N_16606);
or U19711 (N_19711,N_16653,N_16437);
nand U19712 (N_19712,N_16667,N_16901);
or U19713 (N_19713,N_16904,N_16810);
and U19714 (N_19714,N_17549,N_17353);
nor U19715 (N_19715,N_17581,N_17609);
or U19716 (N_19716,N_17929,N_17631);
nor U19717 (N_19717,N_16757,N_16238);
and U19718 (N_19718,N_17187,N_16143);
and U19719 (N_19719,N_17327,N_17123);
nor U19720 (N_19720,N_16855,N_16357);
xnor U19721 (N_19721,N_16639,N_17021);
and U19722 (N_19722,N_16680,N_16992);
nand U19723 (N_19723,N_16473,N_16788);
nor U19724 (N_19724,N_17092,N_17273);
nand U19725 (N_19725,N_17320,N_17472);
and U19726 (N_19726,N_17840,N_16679);
or U19727 (N_19727,N_17141,N_16188);
and U19728 (N_19728,N_16725,N_17010);
nor U19729 (N_19729,N_16500,N_17475);
nor U19730 (N_19730,N_17553,N_17778);
and U19731 (N_19731,N_17690,N_17051);
or U19732 (N_19732,N_17081,N_16570);
and U19733 (N_19733,N_16738,N_16921);
nand U19734 (N_19734,N_17644,N_16294);
or U19735 (N_19735,N_17554,N_17526);
and U19736 (N_19736,N_17912,N_17067);
nor U19737 (N_19737,N_17525,N_17565);
and U19738 (N_19738,N_17700,N_16535);
nand U19739 (N_19739,N_16513,N_17112);
nand U19740 (N_19740,N_16524,N_17389);
or U19741 (N_19741,N_16171,N_16129);
nand U19742 (N_19742,N_17103,N_16356);
or U19743 (N_19743,N_17180,N_17719);
nand U19744 (N_19744,N_16948,N_17871);
and U19745 (N_19745,N_16392,N_16699);
nand U19746 (N_19746,N_17655,N_17275);
nor U19747 (N_19747,N_16161,N_17316);
nor U19748 (N_19748,N_16827,N_16126);
or U19749 (N_19749,N_17414,N_16035);
or U19750 (N_19750,N_17187,N_17400);
nor U19751 (N_19751,N_16063,N_17217);
and U19752 (N_19752,N_17296,N_16740);
or U19753 (N_19753,N_16819,N_17919);
xor U19754 (N_19754,N_16512,N_16332);
or U19755 (N_19755,N_16658,N_16932);
or U19756 (N_19756,N_16641,N_17389);
and U19757 (N_19757,N_17022,N_16705);
or U19758 (N_19758,N_17112,N_17916);
and U19759 (N_19759,N_17845,N_16151);
and U19760 (N_19760,N_16411,N_16629);
nand U19761 (N_19761,N_17290,N_16968);
nand U19762 (N_19762,N_17097,N_17194);
and U19763 (N_19763,N_16335,N_17170);
nor U19764 (N_19764,N_17798,N_16694);
nand U19765 (N_19765,N_16172,N_17173);
nor U19766 (N_19766,N_16676,N_17096);
and U19767 (N_19767,N_17372,N_17666);
or U19768 (N_19768,N_16643,N_16036);
or U19769 (N_19769,N_16450,N_17431);
and U19770 (N_19770,N_16781,N_17530);
and U19771 (N_19771,N_17568,N_17313);
and U19772 (N_19772,N_17256,N_16522);
and U19773 (N_19773,N_16127,N_17498);
nor U19774 (N_19774,N_16587,N_16522);
nand U19775 (N_19775,N_16826,N_17275);
nor U19776 (N_19776,N_16113,N_17492);
nor U19777 (N_19777,N_17249,N_16346);
and U19778 (N_19778,N_16313,N_16327);
and U19779 (N_19779,N_16263,N_16881);
nor U19780 (N_19780,N_16466,N_17145);
and U19781 (N_19781,N_16895,N_17405);
nor U19782 (N_19782,N_16436,N_17584);
nand U19783 (N_19783,N_16377,N_17909);
nor U19784 (N_19784,N_17863,N_17633);
or U19785 (N_19785,N_17675,N_16485);
or U19786 (N_19786,N_17811,N_16663);
and U19787 (N_19787,N_17516,N_16690);
or U19788 (N_19788,N_17240,N_16364);
nor U19789 (N_19789,N_17114,N_16643);
and U19790 (N_19790,N_17305,N_16958);
nand U19791 (N_19791,N_16167,N_17267);
or U19792 (N_19792,N_16920,N_17336);
nor U19793 (N_19793,N_16533,N_17486);
or U19794 (N_19794,N_17354,N_16283);
nand U19795 (N_19795,N_17302,N_16423);
xnor U19796 (N_19796,N_17543,N_16587);
or U19797 (N_19797,N_16706,N_16690);
or U19798 (N_19798,N_16722,N_17675);
nand U19799 (N_19799,N_17978,N_16707);
nand U19800 (N_19800,N_16687,N_16731);
nor U19801 (N_19801,N_16675,N_17506);
nand U19802 (N_19802,N_17052,N_16479);
nand U19803 (N_19803,N_16373,N_16491);
and U19804 (N_19804,N_16470,N_17626);
or U19805 (N_19805,N_17479,N_16689);
and U19806 (N_19806,N_17698,N_17887);
xor U19807 (N_19807,N_17601,N_16803);
and U19808 (N_19808,N_16255,N_17842);
nor U19809 (N_19809,N_16143,N_16882);
xor U19810 (N_19810,N_17914,N_16057);
nand U19811 (N_19811,N_16259,N_17793);
and U19812 (N_19812,N_17506,N_16173);
or U19813 (N_19813,N_17201,N_17007);
and U19814 (N_19814,N_17902,N_17529);
xnor U19815 (N_19815,N_17646,N_17570);
and U19816 (N_19816,N_17568,N_16617);
or U19817 (N_19817,N_16137,N_17564);
or U19818 (N_19818,N_17770,N_16419);
and U19819 (N_19819,N_16706,N_17570);
or U19820 (N_19820,N_16917,N_17332);
and U19821 (N_19821,N_17459,N_17089);
or U19822 (N_19822,N_17262,N_17055);
and U19823 (N_19823,N_17694,N_17643);
nor U19824 (N_19824,N_17870,N_17320);
nand U19825 (N_19825,N_16119,N_17012);
nor U19826 (N_19826,N_16173,N_16538);
nor U19827 (N_19827,N_16306,N_16777);
nor U19828 (N_19828,N_17272,N_16432);
nor U19829 (N_19829,N_16045,N_17723);
and U19830 (N_19830,N_16579,N_17873);
or U19831 (N_19831,N_16801,N_17831);
nand U19832 (N_19832,N_17645,N_17300);
and U19833 (N_19833,N_16641,N_16284);
nand U19834 (N_19834,N_17193,N_17599);
nand U19835 (N_19835,N_16497,N_16584);
or U19836 (N_19836,N_17277,N_17989);
xnor U19837 (N_19837,N_17992,N_17200);
or U19838 (N_19838,N_17214,N_17191);
nor U19839 (N_19839,N_16145,N_16048);
nor U19840 (N_19840,N_17693,N_16581);
and U19841 (N_19841,N_16575,N_17719);
xnor U19842 (N_19842,N_16627,N_17997);
or U19843 (N_19843,N_17370,N_17027);
nand U19844 (N_19844,N_17489,N_17486);
and U19845 (N_19845,N_16761,N_16714);
and U19846 (N_19846,N_17058,N_16744);
or U19847 (N_19847,N_16876,N_16056);
and U19848 (N_19848,N_16415,N_16425);
xor U19849 (N_19849,N_16060,N_17035);
nand U19850 (N_19850,N_16639,N_16906);
or U19851 (N_19851,N_16882,N_17049);
or U19852 (N_19852,N_16939,N_17207);
nand U19853 (N_19853,N_17916,N_16491);
or U19854 (N_19854,N_16078,N_17131);
or U19855 (N_19855,N_17084,N_16830);
xnor U19856 (N_19856,N_17995,N_17702);
nor U19857 (N_19857,N_16067,N_17269);
and U19858 (N_19858,N_16186,N_17229);
nand U19859 (N_19859,N_17603,N_17848);
or U19860 (N_19860,N_16936,N_17504);
nor U19861 (N_19861,N_16319,N_16040);
nand U19862 (N_19862,N_16600,N_16123);
nor U19863 (N_19863,N_16376,N_16820);
and U19864 (N_19864,N_17877,N_16465);
or U19865 (N_19865,N_17017,N_16896);
and U19866 (N_19866,N_17795,N_16818);
or U19867 (N_19867,N_16632,N_17893);
nor U19868 (N_19868,N_17508,N_17772);
and U19869 (N_19869,N_17914,N_16354);
and U19870 (N_19870,N_16226,N_17404);
nand U19871 (N_19871,N_17779,N_17043);
nor U19872 (N_19872,N_17438,N_17987);
and U19873 (N_19873,N_17771,N_16163);
and U19874 (N_19874,N_17583,N_17528);
or U19875 (N_19875,N_17676,N_16482);
and U19876 (N_19876,N_17484,N_16925);
and U19877 (N_19877,N_17909,N_16140);
and U19878 (N_19878,N_16850,N_17087);
nor U19879 (N_19879,N_16212,N_16556);
and U19880 (N_19880,N_17852,N_17694);
or U19881 (N_19881,N_17565,N_16594);
or U19882 (N_19882,N_17555,N_17663);
and U19883 (N_19883,N_17578,N_17396);
nand U19884 (N_19884,N_17048,N_16168);
or U19885 (N_19885,N_17322,N_16568);
and U19886 (N_19886,N_17942,N_16382);
nand U19887 (N_19887,N_17984,N_17790);
nand U19888 (N_19888,N_17770,N_16541);
nand U19889 (N_19889,N_17563,N_16500);
or U19890 (N_19890,N_16154,N_17762);
or U19891 (N_19891,N_16709,N_17307);
nor U19892 (N_19892,N_17405,N_16938);
and U19893 (N_19893,N_17478,N_17668);
nor U19894 (N_19894,N_16665,N_17300);
and U19895 (N_19895,N_17321,N_17983);
nand U19896 (N_19896,N_16491,N_17158);
nor U19897 (N_19897,N_16181,N_16121);
and U19898 (N_19898,N_16985,N_16828);
xor U19899 (N_19899,N_17391,N_17303);
xnor U19900 (N_19900,N_16506,N_17310);
nand U19901 (N_19901,N_17939,N_16725);
or U19902 (N_19902,N_17959,N_17706);
xnor U19903 (N_19903,N_16319,N_16920);
and U19904 (N_19904,N_17564,N_16838);
nor U19905 (N_19905,N_17993,N_17747);
xor U19906 (N_19906,N_17676,N_16045);
nand U19907 (N_19907,N_17128,N_17634);
nand U19908 (N_19908,N_17759,N_16724);
nand U19909 (N_19909,N_16049,N_16122);
and U19910 (N_19910,N_17954,N_16598);
nand U19911 (N_19911,N_17312,N_17005);
or U19912 (N_19912,N_17240,N_17295);
nor U19913 (N_19913,N_16944,N_16522);
nand U19914 (N_19914,N_17611,N_17686);
or U19915 (N_19915,N_16939,N_16350);
nand U19916 (N_19916,N_17618,N_16681);
and U19917 (N_19917,N_17828,N_17921);
and U19918 (N_19918,N_17606,N_17414);
nor U19919 (N_19919,N_16821,N_16129);
or U19920 (N_19920,N_16738,N_16060);
and U19921 (N_19921,N_17978,N_16153);
nand U19922 (N_19922,N_17529,N_17041);
nand U19923 (N_19923,N_17436,N_17224);
or U19924 (N_19924,N_17730,N_16521);
nor U19925 (N_19925,N_16374,N_17590);
and U19926 (N_19926,N_17297,N_16243);
nand U19927 (N_19927,N_16978,N_16855);
or U19928 (N_19928,N_16857,N_16224);
or U19929 (N_19929,N_16938,N_16839);
nand U19930 (N_19930,N_16868,N_16406);
or U19931 (N_19931,N_17928,N_16851);
or U19932 (N_19932,N_16696,N_16533);
nand U19933 (N_19933,N_17551,N_17273);
xor U19934 (N_19934,N_16045,N_16160);
or U19935 (N_19935,N_16037,N_16196);
nand U19936 (N_19936,N_16111,N_17385);
or U19937 (N_19937,N_17216,N_17827);
nand U19938 (N_19938,N_17503,N_16656);
nand U19939 (N_19939,N_17080,N_17990);
nor U19940 (N_19940,N_17183,N_17877);
or U19941 (N_19941,N_16857,N_16712);
xor U19942 (N_19942,N_16100,N_16207);
and U19943 (N_19943,N_16980,N_16883);
or U19944 (N_19944,N_17501,N_17867);
or U19945 (N_19945,N_17334,N_17145);
xnor U19946 (N_19946,N_16555,N_16012);
and U19947 (N_19947,N_17187,N_17196);
or U19948 (N_19948,N_16982,N_16416);
or U19949 (N_19949,N_16959,N_17530);
nor U19950 (N_19950,N_16645,N_16501);
nor U19951 (N_19951,N_16687,N_17716);
nor U19952 (N_19952,N_16611,N_17515);
or U19953 (N_19953,N_17347,N_16743);
nand U19954 (N_19954,N_16047,N_17385);
nand U19955 (N_19955,N_17496,N_16023);
or U19956 (N_19956,N_17065,N_17745);
nor U19957 (N_19957,N_17520,N_17633);
xnor U19958 (N_19958,N_16550,N_17753);
and U19959 (N_19959,N_16676,N_16941);
nor U19960 (N_19960,N_16171,N_17154);
or U19961 (N_19961,N_17753,N_17850);
nor U19962 (N_19962,N_16666,N_16639);
nor U19963 (N_19963,N_16118,N_17817);
nor U19964 (N_19964,N_17911,N_16273);
and U19965 (N_19965,N_17809,N_17859);
nand U19966 (N_19966,N_16533,N_16990);
or U19967 (N_19967,N_16477,N_17094);
nand U19968 (N_19968,N_17552,N_16744);
or U19969 (N_19969,N_17196,N_16691);
and U19970 (N_19970,N_17239,N_16430);
and U19971 (N_19971,N_17552,N_17116);
xnor U19972 (N_19972,N_17647,N_17960);
nor U19973 (N_19973,N_16878,N_17408);
and U19974 (N_19974,N_17689,N_17674);
or U19975 (N_19975,N_16069,N_16537);
nor U19976 (N_19976,N_16710,N_16080);
nand U19977 (N_19977,N_16126,N_17855);
and U19978 (N_19978,N_16529,N_16126);
nor U19979 (N_19979,N_16088,N_17018);
and U19980 (N_19980,N_16507,N_17053);
xor U19981 (N_19981,N_17461,N_16590);
xnor U19982 (N_19982,N_16011,N_16037);
nand U19983 (N_19983,N_16276,N_17309);
and U19984 (N_19984,N_16001,N_16394);
and U19985 (N_19985,N_17905,N_17061);
nor U19986 (N_19986,N_16739,N_16825);
and U19987 (N_19987,N_16386,N_16845);
nor U19988 (N_19988,N_17083,N_17703);
or U19989 (N_19989,N_17035,N_17040);
or U19990 (N_19990,N_16847,N_16967);
and U19991 (N_19991,N_16355,N_16615);
and U19992 (N_19992,N_16824,N_16251);
xnor U19993 (N_19993,N_17619,N_16746);
nand U19994 (N_19994,N_17440,N_16948);
or U19995 (N_19995,N_17160,N_17317);
or U19996 (N_19996,N_17504,N_17772);
nand U19997 (N_19997,N_17133,N_17726);
nand U19998 (N_19998,N_16705,N_17504);
nor U19999 (N_19999,N_17514,N_16202);
nand UO_0 (O_0,N_19020,N_18847);
nand UO_1 (O_1,N_18075,N_18803);
nand UO_2 (O_2,N_19223,N_19454);
nand UO_3 (O_3,N_19392,N_19547);
nand UO_4 (O_4,N_18351,N_18280);
nand UO_5 (O_5,N_19600,N_19049);
or UO_6 (O_6,N_19998,N_18427);
and UO_7 (O_7,N_18994,N_19302);
xor UO_8 (O_8,N_18254,N_18218);
nand UO_9 (O_9,N_19524,N_19615);
or UO_10 (O_10,N_19191,N_19339);
xnor UO_11 (O_11,N_18687,N_18603);
nor UO_12 (O_12,N_18002,N_18948);
and UO_13 (O_13,N_19437,N_18873);
and UO_14 (O_14,N_18996,N_18032);
and UO_15 (O_15,N_19019,N_19139);
nand UO_16 (O_16,N_19477,N_19542);
or UO_17 (O_17,N_19529,N_18760);
xnor UO_18 (O_18,N_19708,N_19935);
nand UO_19 (O_19,N_18058,N_18858);
xnor UO_20 (O_20,N_19250,N_18321);
nor UO_21 (O_21,N_19222,N_18885);
or UO_22 (O_22,N_19590,N_19865);
nor UO_23 (O_23,N_19902,N_19276);
or UO_24 (O_24,N_18093,N_19537);
and UO_25 (O_25,N_19093,N_19960);
nand UO_26 (O_26,N_18721,N_18616);
or UO_27 (O_27,N_18673,N_18816);
or UO_28 (O_28,N_19714,N_19499);
or UO_29 (O_29,N_19081,N_18463);
nand UO_30 (O_30,N_19480,N_19869);
or UO_31 (O_31,N_18776,N_18805);
nor UO_32 (O_32,N_18980,N_19560);
or UO_33 (O_33,N_18957,N_19980);
or UO_34 (O_34,N_18596,N_19812);
nor UO_35 (O_35,N_19182,N_19380);
and UO_36 (O_36,N_19439,N_18214);
or UO_37 (O_37,N_18380,N_18407);
nor UO_38 (O_38,N_19554,N_19654);
nor UO_39 (O_39,N_18363,N_19601);
nand UO_40 (O_40,N_18652,N_19069);
and UO_41 (O_41,N_19283,N_19984);
xnor UO_42 (O_42,N_18553,N_18126);
or UO_43 (O_43,N_18952,N_18307);
nor UO_44 (O_44,N_18099,N_19146);
nor UO_45 (O_45,N_18298,N_18774);
or UO_46 (O_46,N_19962,N_18510);
nor UO_47 (O_47,N_18864,N_19447);
nand UO_48 (O_48,N_19387,N_19238);
nand UO_49 (O_49,N_19764,N_19956);
nor UO_50 (O_50,N_19577,N_19977);
nor UO_51 (O_51,N_18743,N_18089);
and UO_52 (O_52,N_19732,N_18279);
and UO_53 (O_53,N_18076,N_19565);
nor UO_54 (O_54,N_18570,N_18162);
nor UO_55 (O_55,N_18394,N_18573);
nor UO_56 (O_56,N_18506,N_18680);
xor UO_57 (O_57,N_18170,N_18421);
and UO_58 (O_58,N_18825,N_18323);
nand UO_59 (O_59,N_19162,N_19314);
or UO_60 (O_60,N_19305,N_18887);
nor UO_61 (O_61,N_19434,N_19262);
nand UO_62 (O_62,N_18345,N_18904);
and UO_63 (O_63,N_19776,N_19011);
nor UO_64 (O_64,N_19737,N_18625);
or UO_65 (O_65,N_19493,N_19589);
or UO_66 (O_66,N_18258,N_19607);
nor UO_67 (O_67,N_18710,N_18236);
nand UO_68 (O_68,N_18921,N_18349);
nand UO_69 (O_69,N_19625,N_19694);
nand UO_70 (O_70,N_18387,N_18752);
nor UO_71 (O_71,N_19844,N_19966);
and UO_72 (O_72,N_19418,N_19648);
nand UO_73 (O_73,N_19325,N_19707);
and UO_74 (O_74,N_18003,N_19284);
nor UO_75 (O_75,N_19574,N_19065);
and UO_76 (O_76,N_19946,N_18425);
and UO_77 (O_77,N_18802,N_19239);
and UO_78 (O_78,N_19598,N_19744);
or UO_79 (O_79,N_19703,N_18841);
nor UO_80 (O_80,N_19018,N_18189);
nor UO_81 (O_81,N_19680,N_18529);
nand UO_82 (O_82,N_19346,N_18571);
nand UO_83 (O_83,N_19295,N_19123);
nand UO_84 (O_84,N_19003,N_18852);
nor UO_85 (O_85,N_19345,N_19716);
nor UO_86 (O_86,N_18967,N_18005);
nor UO_87 (O_87,N_19285,N_18508);
nor UO_88 (O_88,N_18038,N_18205);
or UO_89 (O_89,N_19997,N_19055);
nor UO_90 (O_90,N_18057,N_18013);
and UO_91 (O_91,N_19288,N_18543);
xor UO_92 (O_92,N_19396,N_19568);
nand UO_93 (O_93,N_19344,N_19487);
nand UO_94 (O_94,N_19630,N_18992);
nand UO_95 (O_95,N_18183,N_19575);
or UO_96 (O_96,N_19414,N_18991);
nor UO_97 (O_97,N_18779,N_18455);
nand UO_98 (O_98,N_19545,N_19553);
nand UO_99 (O_99,N_19635,N_19178);
nand UO_100 (O_100,N_18201,N_18191);
or UO_101 (O_101,N_19320,N_19546);
nand UO_102 (O_102,N_18954,N_19569);
xor UO_103 (O_103,N_19368,N_18821);
nor UO_104 (O_104,N_18981,N_19866);
nand UO_105 (O_105,N_18305,N_19702);
nand UO_106 (O_106,N_19689,N_18520);
and UO_107 (O_107,N_18583,N_19944);
xor UO_108 (O_108,N_19072,N_18563);
nand UO_109 (O_109,N_18857,N_19857);
xor UO_110 (O_110,N_18662,N_18737);
nor UO_111 (O_111,N_18728,N_18541);
or UO_112 (O_112,N_19053,N_18912);
and UO_113 (O_113,N_19823,N_18540);
or UO_114 (O_114,N_18224,N_19221);
nand UO_115 (O_115,N_18809,N_19544);
xnor UO_116 (O_116,N_18602,N_19909);
or UO_117 (O_117,N_19111,N_19619);
nand UO_118 (O_118,N_19083,N_18188);
or UO_119 (O_119,N_19484,N_19196);
or UO_120 (O_120,N_19006,N_19700);
nand UO_121 (O_121,N_19512,N_18064);
nand UO_122 (O_122,N_18830,N_18088);
nand UO_123 (O_123,N_19201,N_18762);
nor UO_124 (O_124,N_18273,N_19733);
nand UO_125 (O_125,N_18785,N_18295);
nor UO_126 (O_126,N_18960,N_19697);
nor UO_127 (O_127,N_18461,N_19452);
or UO_128 (O_128,N_19879,N_18084);
and UO_129 (O_129,N_18528,N_18987);
and UO_130 (O_130,N_19193,N_19331);
nand UO_131 (O_131,N_18733,N_19076);
nor UO_132 (O_132,N_18654,N_19532);
nand UO_133 (O_133,N_18990,N_19496);
or UO_134 (O_134,N_19179,N_19036);
nor UO_135 (O_135,N_19955,N_19354);
nand UO_136 (O_136,N_19969,N_18513);
or UO_137 (O_137,N_18839,N_18660);
and UO_138 (O_138,N_19292,N_18070);
nor UO_139 (O_139,N_19631,N_19849);
and UO_140 (O_140,N_19151,N_18907);
nand UO_141 (O_141,N_18634,N_19062);
xnor UO_142 (O_142,N_18937,N_18232);
nor UO_143 (O_143,N_19185,N_19819);
xnor UO_144 (O_144,N_18641,N_19032);
and UO_145 (O_145,N_19172,N_19033);
nor UO_146 (O_146,N_19726,N_18934);
nand UO_147 (O_147,N_18327,N_18524);
and UO_148 (O_148,N_19402,N_18496);
nor UO_149 (O_149,N_19850,N_18955);
and UO_150 (O_150,N_19720,N_18418);
and UO_151 (O_151,N_18889,N_18432);
and UO_152 (O_152,N_19886,N_19951);
nor UO_153 (O_153,N_19335,N_18787);
nand UO_154 (O_154,N_18333,N_18238);
nor UO_155 (O_155,N_19027,N_18286);
or UO_156 (O_156,N_18487,N_18239);
nand UO_157 (O_157,N_19161,N_19699);
and UO_158 (O_158,N_19840,N_19381);
nand UO_159 (O_159,N_19725,N_18715);
nor UO_160 (O_160,N_18691,N_18398);
or UO_161 (O_161,N_18467,N_18357);
or UO_162 (O_162,N_19564,N_19638);
nor UO_163 (O_163,N_19056,N_19551);
or UO_164 (O_164,N_18049,N_18711);
and UO_165 (O_165,N_18185,N_18574);
xnor UO_166 (O_166,N_19455,N_19306);
and UO_167 (O_167,N_18208,N_19300);
or UO_168 (O_168,N_18671,N_18036);
nor UO_169 (O_169,N_19674,N_19129);
and UO_170 (O_170,N_19023,N_18113);
nand UO_171 (O_171,N_19063,N_18290);
nand UO_172 (O_172,N_18585,N_18688);
xor UO_173 (O_173,N_18584,N_19411);
or UO_174 (O_174,N_18819,N_19957);
or UO_175 (O_175,N_19555,N_19527);
nand UO_176 (O_176,N_18669,N_19175);
or UO_177 (O_177,N_18562,N_19762);
nand UO_178 (O_178,N_19017,N_18147);
and UO_179 (O_179,N_19563,N_19649);
nand UO_180 (O_180,N_19611,N_18861);
nor UO_181 (O_181,N_19525,N_19486);
nor UO_182 (O_182,N_19746,N_19459);
nand UO_183 (O_183,N_19138,N_18423);
nor UO_184 (O_184,N_18160,N_19265);
nor UO_185 (O_185,N_19074,N_19627);
nand UO_186 (O_186,N_19667,N_19342);
or UO_187 (O_187,N_19816,N_19312);
and UO_188 (O_188,N_18791,N_18667);
and UO_189 (O_189,N_18197,N_18429);
or UO_190 (O_190,N_18374,N_18350);
and UO_191 (O_191,N_18386,N_19438);
nor UO_192 (O_192,N_19800,N_18910);
or UO_193 (O_193,N_18471,N_18092);
or UO_194 (O_194,N_18466,N_19152);
nand UO_195 (O_195,N_19307,N_19632);
nand UO_196 (O_196,N_19400,N_19675);
or UO_197 (O_197,N_18723,N_18181);
or UO_198 (O_198,N_18107,N_19571);
and UO_199 (O_199,N_18668,N_19166);
nor UO_200 (O_200,N_18203,N_19165);
nand UO_201 (O_201,N_18226,N_19263);
nand UO_202 (O_202,N_18535,N_18901);
or UO_203 (O_203,N_19573,N_18604);
or UO_204 (O_204,N_18659,N_19333);
or UO_205 (O_205,N_19478,N_19144);
nand UO_206 (O_206,N_18707,N_18447);
and UO_207 (O_207,N_19430,N_19237);
xnor UO_208 (O_208,N_18134,N_18291);
and UO_209 (O_209,N_19163,N_19405);
or UO_210 (O_210,N_19431,N_18137);
or UO_211 (O_211,N_19110,N_19082);
nand UO_212 (O_212,N_19220,N_18382);
nand UO_213 (O_213,N_19651,N_18316);
nand UO_214 (O_214,N_18590,N_19369);
nor UO_215 (O_215,N_19770,N_19806);
nand UO_216 (O_216,N_18031,N_18938);
xor UO_217 (O_217,N_19358,N_18923);
and UO_218 (O_218,N_18903,N_18995);
nand UO_219 (O_219,N_18109,N_19176);
nor UO_220 (O_220,N_19050,N_19281);
nor UO_221 (O_221,N_18138,N_19080);
or UO_222 (O_222,N_19991,N_19105);
and UO_223 (O_223,N_19410,N_19329);
nand UO_224 (O_224,N_19365,N_18909);
and UO_225 (O_225,N_19352,N_18303);
and UO_226 (O_226,N_19647,N_18699);
and UO_227 (O_227,N_19794,N_19462);
and UO_228 (O_228,N_18761,N_19024);
and UO_229 (O_229,N_19561,N_19153);
nor UO_230 (O_230,N_19739,N_19071);
and UO_231 (O_231,N_18169,N_19713);
nand UO_232 (O_232,N_19646,N_18985);
nor UO_233 (O_233,N_18220,N_19385);
xnor UO_234 (O_234,N_18542,N_19669);
nor UO_235 (O_235,N_19738,N_19880);
nor UO_236 (O_236,N_19422,N_18928);
nor UO_237 (O_237,N_19652,N_18836);
or UO_238 (O_238,N_19164,N_19058);
nand UO_239 (O_239,N_19976,N_19143);
nand UO_240 (O_240,N_18838,N_18977);
or UO_241 (O_241,N_19184,N_19192);
nor UO_242 (O_242,N_18308,N_19324);
and UO_243 (O_243,N_19847,N_18769);
nor UO_244 (O_244,N_18870,N_18338);
xnor UO_245 (O_245,N_19842,N_18856);
xnor UO_246 (O_246,N_18012,N_18034);
nor UO_247 (O_247,N_19347,N_18117);
and UO_248 (O_248,N_19258,N_18620);
nor UO_249 (O_249,N_19735,N_18505);
and UO_250 (O_250,N_19476,N_19734);
or UO_251 (O_251,N_18961,N_18749);
nand UO_252 (O_252,N_18610,N_19836);
and UO_253 (O_253,N_18566,N_18317);
nor UO_254 (O_254,N_19245,N_19883);
and UO_255 (O_255,N_19042,N_19685);
and UO_256 (O_256,N_19509,N_19046);
and UO_257 (O_257,N_19831,N_18843);
nand UO_258 (O_258,N_19323,N_19086);
or UO_259 (O_259,N_18131,N_18325);
xnor UO_260 (O_260,N_18180,N_19435);
nand UO_261 (O_261,N_19884,N_19982);
and UO_262 (O_262,N_18629,N_18678);
or UO_263 (O_263,N_19142,N_19294);
or UO_264 (O_264,N_19127,N_19595);
nand UO_265 (O_265,N_18558,N_19119);
and UO_266 (O_266,N_19197,N_19412);
and UO_267 (O_267,N_19691,N_18982);
and UO_268 (O_268,N_19906,N_19522);
nor UO_269 (O_269,N_19456,N_18219);
or UO_270 (O_270,N_18037,N_19180);
or UO_271 (O_271,N_18278,N_19892);
and UO_272 (O_272,N_19559,N_19597);
nor UO_273 (O_273,N_19827,N_18900);
nor UO_274 (O_274,N_19140,N_18240);
or UO_275 (O_275,N_18826,N_19107);
nor UO_276 (O_276,N_18265,N_19838);
and UO_277 (O_277,N_18009,N_18628);
nor UO_278 (O_278,N_19116,N_18048);
xnor UO_279 (O_279,N_18378,N_19661);
or UO_280 (O_280,N_18670,N_18007);
nor UO_281 (O_281,N_18184,N_19855);
nor UO_282 (O_282,N_19938,N_19766);
nor UO_283 (O_283,N_19684,N_18128);
and UO_284 (O_284,N_18833,N_19817);
or UO_285 (O_285,N_18582,N_18456);
nor UO_286 (O_286,N_19871,N_18972);
and UO_287 (O_287,N_19124,N_18588);
and UO_288 (O_288,N_18143,N_19623);
or UO_289 (O_289,N_18404,N_18293);
nand UO_290 (O_290,N_19633,N_19386);
nor UO_291 (O_291,N_19315,N_19132);
or UO_292 (O_292,N_18198,N_18739);
or UO_293 (O_293,N_19482,N_18063);
nand UO_294 (O_294,N_18672,N_18241);
nand UO_295 (O_295,N_18517,N_18727);
nand UO_296 (O_296,N_18800,N_19515);
nor UO_297 (O_297,N_18299,N_18477);
or UO_298 (O_298,N_19752,N_18886);
nand UO_299 (O_299,N_19867,N_18086);
or UO_300 (O_300,N_19772,N_18082);
nand UO_301 (O_301,N_19915,N_18397);
and UO_302 (O_302,N_18133,N_18726);
nor UO_303 (O_303,N_19360,N_19778);
and UO_304 (O_304,N_18194,N_18095);
and UO_305 (O_305,N_18060,N_18442);
xnor UO_306 (O_306,N_19876,N_18212);
xor UO_307 (O_307,N_18643,N_19121);
nor UO_308 (O_308,N_18569,N_18975);
xor UO_309 (O_309,N_18424,N_19461);
nor UO_310 (O_310,N_19117,N_19277);
nor UO_311 (O_311,N_19815,N_18416);
or UO_312 (O_312,N_19157,N_18789);
nor UO_313 (O_313,N_18024,N_19541);
nand UO_314 (O_314,N_19722,N_18098);
and UO_315 (O_315,N_19174,N_19814);
or UO_316 (O_316,N_19786,N_18817);
or UO_317 (O_317,N_19267,N_18073);
xnor UO_318 (O_318,N_19041,N_19147);
nand UO_319 (O_319,N_19468,N_18626);
and UO_320 (O_320,N_18896,N_18872);
and UO_321 (O_321,N_18237,N_18035);
nor UO_322 (O_322,N_18251,N_18783);
xor UO_323 (O_323,N_18915,N_18917);
and UO_324 (O_324,N_18488,N_18067);
nand UO_325 (O_325,N_19044,N_19787);
nor UO_326 (O_326,N_19286,N_18646);
and UO_327 (O_327,N_19096,N_18020);
or UO_328 (O_328,N_18877,N_18282);
or UO_329 (O_329,N_18043,N_18534);
and UO_330 (O_330,N_19665,N_19407);
nand UO_331 (O_331,N_19103,N_19204);
and UO_332 (O_332,N_18056,N_18264);
or UO_333 (O_333,N_18685,N_19624);
nand UO_334 (O_334,N_19639,N_18775);
or UO_335 (O_335,N_18249,N_18202);
nand UO_336 (O_336,N_19520,N_19941);
nor UO_337 (O_337,N_18276,N_18110);
nand UO_338 (O_338,N_19862,N_19760);
nor UO_339 (O_339,N_18755,N_19497);
and UO_340 (O_340,N_18638,N_19896);
nand UO_341 (O_341,N_18362,N_18225);
nand UO_342 (O_342,N_19255,N_19662);
nand UO_343 (O_343,N_18601,N_19846);
and UO_344 (O_344,N_19710,N_18572);
nand UO_345 (O_345,N_19719,N_18684);
or UO_346 (O_346,N_19741,N_18428);
and UO_347 (O_347,N_18178,N_19834);
xor UO_348 (O_348,N_18983,N_19471);
or UO_349 (O_349,N_19985,N_19005);
and UO_350 (O_350,N_19021,N_18068);
nor UO_351 (O_351,N_18512,N_18297);
or UO_352 (O_352,N_18469,N_19421);
and UO_353 (O_353,N_18055,N_19605);
nand UO_354 (O_354,N_19230,N_18581);
nand UO_355 (O_355,N_18700,N_19860);
or UO_356 (O_356,N_18217,N_18122);
nor UO_357 (O_357,N_18256,N_18052);
nand UO_358 (O_358,N_18621,N_18431);
or UO_359 (O_359,N_19371,N_19463);
or UO_360 (O_360,N_18340,N_19536);
or UO_361 (O_361,N_19897,N_18246);
or UO_362 (O_362,N_19535,N_18970);
nand UO_363 (O_363,N_18757,N_18161);
or UO_364 (O_364,N_18159,N_19933);
nor UO_365 (O_365,N_19367,N_19796);
nor UO_366 (O_366,N_19767,N_19895);
nor UO_367 (O_367,N_18452,N_19304);
and UO_368 (O_368,N_19492,N_19094);
and UO_369 (O_369,N_18156,N_18951);
nand UO_370 (O_370,N_18719,N_18409);
and UO_371 (O_371,N_19436,N_19531);
nand UO_372 (O_372,N_19655,N_18272);
nor UO_373 (O_373,N_19290,N_18689);
and UO_374 (O_374,N_19761,N_19303);
nand UO_375 (O_375,N_18854,N_18550);
nor UO_376 (O_376,N_19994,N_18196);
and UO_377 (O_377,N_18281,N_19183);
or UO_378 (O_378,N_19214,N_18044);
or UO_379 (O_379,N_19064,N_19246);
and UO_380 (O_380,N_19075,N_18072);
or UO_381 (O_381,N_18283,N_19350);
and UO_382 (O_382,N_19943,N_19671);
nor UO_383 (O_383,N_18085,N_18893);
or UO_384 (O_384,N_18567,N_19359);
nor UO_385 (O_385,N_19318,N_18666);
or UO_386 (O_386,N_19891,N_19446);
xor UO_387 (O_387,N_18489,N_18449);
nand UO_388 (O_388,N_19711,N_19030);
xnor UO_389 (O_389,N_18891,N_19503);
and UO_390 (O_390,N_19473,N_18511);
or UO_391 (O_391,N_19460,N_19099);
and UO_392 (O_392,N_19904,N_19500);
nor UO_393 (O_393,N_18173,N_18438);
nand UO_394 (O_394,N_18211,N_18735);
nand UO_395 (O_395,N_18328,N_19274);
and UO_396 (O_396,N_18973,N_18771);
nor UO_397 (O_397,N_18950,N_19451);
nand UO_398 (O_398,N_18412,N_18648);
nor UO_399 (O_399,N_18580,N_19807);
and UO_400 (O_400,N_18577,N_19557);
and UO_401 (O_401,N_19275,N_18978);
and UO_402 (O_402,N_18446,N_19448);
and UO_403 (O_403,N_18840,N_19298);
nor UO_404 (O_404,N_18827,N_18647);
nand UO_405 (O_405,N_19773,N_19629);
nor UO_406 (O_406,N_19781,N_18319);
nand UO_407 (O_407,N_18556,N_18618);
nand UO_408 (O_408,N_18294,N_18895);
nor UO_409 (O_409,N_18054,N_19810);
and UO_410 (O_410,N_18564,N_18121);
and UO_411 (O_411,N_19465,N_19495);
nor UO_412 (O_412,N_19321,N_18657);
nor UO_413 (O_413,N_18549,N_19219);
nand UO_414 (O_414,N_18968,N_19194);
and UO_415 (O_415,N_18863,N_19929);
and UO_416 (O_416,N_18632,N_19472);
nand UO_417 (O_417,N_19588,N_19491);
and UO_418 (O_418,N_18371,N_19785);
or UO_419 (O_419,N_18359,N_18692);
nand UO_420 (O_420,N_19606,N_19795);
or UO_421 (O_421,N_19899,N_19361);
nand UO_422 (O_422,N_19516,N_18364);
or UO_423 (O_423,N_18186,N_19640);
nand UO_424 (O_424,N_19753,N_18724);
nor UO_425 (O_425,N_19244,N_18018);
or UO_426 (O_426,N_19291,N_18554);
nor UO_427 (O_427,N_18575,N_19370);
or UO_428 (O_428,N_18120,N_19728);
or UO_429 (O_429,N_19765,N_18804);
nor UO_430 (O_430,N_18890,N_18144);
or UO_431 (O_431,N_19160,N_19521);
nor UO_432 (O_432,N_19264,N_19308);
and UO_433 (O_433,N_19363,N_19645);
nor UO_434 (O_434,N_18729,N_19596);
and UO_435 (O_435,N_18764,N_19978);
nand UO_436 (O_436,N_19609,N_18207);
nand UO_437 (O_437,N_19224,N_18751);
and UO_438 (O_438,N_19488,N_19485);
or UO_439 (O_439,N_19068,N_19348);
nand UO_440 (O_440,N_18233,N_18589);
or UO_441 (O_441,N_18686,N_19873);
nand UO_442 (O_442,N_19188,N_18940);
nor UO_443 (O_443,N_18897,N_19232);
nand UO_444 (O_444,N_19552,N_19918);
and UO_445 (O_445,N_19528,N_19864);
nand UO_446 (O_446,N_18472,N_19610);
nand UO_447 (O_447,N_19198,N_18025);
nor UO_448 (O_448,N_18112,N_19481);
and UO_449 (O_449,N_18050,N_19048);
or UO_450 (O_450,N_18087,N_19266);
or UO_451 (O_451,N_19777,N_19097);
or UO_452 (O_452,N_18959,N_19756);
or UO_453 (O_453,N_18880,N_19106);
nor UO_454 (O_454,N_19424,N_19372);
xor UO_455 (O_455,N_19170,N_18894);
and UO_456 (O_456,N_18223,N_19974);
and UO_457 (O_457,N_19877,N_18440);
nor UO_458 (O_458,N_19133,N_18344);
and UO_459 (O_459,N_19824,N_19903);
nor UO_460 (O_460,N_18027,N_18415);
and UO_461 (O_461,N_18142,N_18250);
xnor UO_462 (O_462,N_18115,N_18413);
and UO_463 (O_463,N_18742,N_19517);
nor UO_464 (O_464,N_18849,N_19205);
or UO_465 (O_465,N_18174,N_18645);
or UO_466 (O_466,N_19016,N_18405);
or UO_467 (O_467,N_18552,N_19750);
xnor UO_468 (O_468,N_19604,N_19874);
xnor UO_469 (O_469,N_18963,N_18812);
and UO_470 (O_470,N_18091,N_18094);
or UO_471 (O_471,N_18314,N_19592);
or UO_472 (O_472,N_19514,N_19658);
nand UO_473 (O_473,N_18253,N_18578);
or UO_474 (O_474,N_19681,N_19821);
or UO_475 (O_475,N_19845,N_19937);
xor UO_476 (O_476,N_18192,N_19177);
nor UO_477 (O_477,N_19243,N_19186);
or UO_478 (O_478,N_18962,N_19872);
xnor UO_479 (O_479,N_18718,N_18105);
nor UO_480 (O_480,N_19950,N_19374);
or UO_481 (O_481,N_19798,N_19695);
nand UO_482 (O_482,N_18594,N_18296);
nand UO_483 (O_483,N_19548,N_19317);
nand UO_484 (O_484,N_18557,N_19135);
nand UO_485 (O_485,N_18102,N_18015);
and UO_486 (O_486,N_19791,N_19120);
nor UO_487 (O_487,N_18451,N_18936);
xor UO_488 (O_488,N_19031,N_19051);
nand UO_489 (O_489,N_19745,N_18988);
and UO_490 (O_490,N_19268,N_18532);
nor UO_491 (O_491,N_19401,N_18911);
and UO_492 (O_492,N_19029,N_18125);
or UO_493 (O_493,N_19566,N_19926);
nand UO_494 (O_494,N_19444,N_19373);
and UO_495 (O_495,N_19077,N_18503);
or UO_496 (O_496,N_18309,N_19718);
and UO_497 (O_497,N_18304,N_19090);
nor UO_498 (O_498,N_19433,N_18644);
or UO_499 (O_499,N_18245,N_18622);
or UO_500 (O_500,N_18639,N_18650);
xnor UO_501 (O_501,N_18445,N_18615);
nand UO_502 (O_502,N_18200,N_19682);
nand UO_503 (O_503,N_19888,N_18794);
and UO_504 (O_504,N_18677,N_19853);
and UO_505 (O_505,N_18747,N_19579);
or UO_506 (O_506,N_18997,N_18734);
nand UO_507 (O_507,N_18481,N_18521);
and UO_508 (O_508,N_18053,N_18175);
and UO_509 (O_509,N_19901,N_18001);
nand UO_510 (O_510,N_18507,N_18493);
and UO_511 (O_511,N_18411,N_18260);
nor UO_512 (O_512,N_19211,N_18986);
nor UO_513 (O_513,N_19397,N_18209);
and UO_514 (O_514,N_19832,N_18712);
and UO_515 (O_515,N_18172,N_18022);
nor UO_516 (O_516,N_18215,N_18478);
and UO_517 (O_517,N_19208,N_19441);
and UO_518 (O_518,N_18016,N_19530);
and UO_519 (O_519,N_19717,N_19672);
and UO_520 (O_520,N_18470,N_18966);
nor UO_521 (O_521,N_19406,N_19567);
nor UO_522 (O_522,N_19934,N_18320);
or UO_523 (O_523,N_19173,N_19322);
xnor UO_524 (O_524,N_18656,N_19015);
or UO_525 (O_525,N_18096,N_18796);
and UO_526 (O_526,N_18019,N_18527);
nand UO_527 (O_527,N_19570,N_18842);
nand UO_528 (O_528,N_19914,N_18679);
nor UO_529 (O_529,N_19670,N_19206);
nor UO_530 (O_530,N_19078,N_18168);
nor UO_531 (O_531,N_19878,N_18484);
and UO_532 (O_532,N_19882,N_18738);
nor UO_533 (O_533,N_18066,N_19313);
or UO_534 (O_534,N_19278,N_18815);
nand UO_535 (O_535,N_19763,N_19271);
or UO_536 (O_536,N_19768,N_19964);
and UO_537 (O_537,N_19679,N_18165);
nand UO_538 (O_538,N_18081,N_18753);
and UO_539 (O_539,N_18004,N_18116);
or UO_540 (O_540,N_18605,N_18614);
xnor UO_541 (O_541,N_18697,N_18866);
nor UO_542 (O_542,N_19581,N_18922);
nor UO_543 (O_543,N_18559,N_19007);
or UO_544 (O_544,N_18586,N_19983);
or UO_545 (O_545,N_19328,N_19802);
nand UO_546 (O_546,N_18100,N_18443);
and UO_547 (O_547,N_18430,N_19820);
nand UO_548 (O_548,N_18797,N_18354);
xnor UO_549 (O_549,N_18494,N_19549);
and UO_550 (O_550,N_19822,N_19656);
and UO_551 (O_551,N_18514,N_19332);
or UO_552 (O_552,N_18612,N_19908);
nand UO_553 (O_553,N_19376,N_18933);
nor UO_554 (O_554,N_18017,N_18141);
nor UO_555 (O_555,N_18074,N_19483);
or UO_556 (O_556,N_19084,N_19508);
nor UO_557 (O_557,N_18693,N_18925);
nor UO_558 (O_558,N_19921,N_18683);
nor UO_559 (O_559,N_19043,N_19550);
nand UO_560 (O_560,N_19754,N_19602);
xnor UO_561 (O_561,N_18777,N_19693);
nand UO_562 (O_562,N_19924,N_19309);
xor UO_563 (O_563,N_19740,N_18792);
or UO_564 (O_564,N_19310,N_18059);
and UO_565 (O_565,N_19856,N_19037);
or UO_566 (O_566,N_19971,N_18336);
nor UO_567 (O_567,N_18597,N_19894);
and UO_568 (O_568,N_19972,N_18998);
nor UO_569 (O_569,N_19990,N_19505);
and UO_570 (O_570,N_18342,N_18132);
nand UO_571 (O_571,N_19098,N_19657);
and UO_572 (O_572,N_18682,N_19137);
xnor UO_573 (O_573,N_18367,N_18560);
nand UO_574 (O_574,N_18177,N_18130);
and UO_575 (O_575,N_18846,N_18935);
nor UO_576 (O_576,N_18732,N_18221);
nor UO_577 (O_577,N_19830,N_18878);
nand UO_578 (O_578,N_18906,N_18698);
nand UO_579 (O_579,N_18617,N_19498);
or UO_580 (O_580,N_18731,N_19299);
and UO_581 (O_581,N_18450,N_19704);
and UO_582 (O_582,N_18811,N_19774);
or UO_583 (O_583,N_18011,N_19925);
xor UO_584 (O_584,N_18624,N_18229);
nor UO_585 (O_585,N_19518,N_18231);
xor UO_586 (O_586,N_19900,N_18741);
nor UO_587 (O_587,N_18497,N_18145);
and UO_588 (O_588,N_19622,N_19939);
or UO_589 (O_589,N_18274,N_18918);
xnor UO_590 (O_590,N_19666,N_19408);
xor UO_591 (O_591,N_19790,N_18500);
or UO_592 (O_592,N_19203,N_18365);
or UO_593 (O_593,N_19248,N_18862);
nor UO_594 (O_594,N_18377,N_18591);
xor UO_595 (O_595,N_18665,N_19002);
xor UO_596 (O_596,N_18271,N_19663);
nand UO_597 (O_597,N_19644,N_18930);
nor UO_598 (O_598,N_19311,N_18926);
or UO_599 (O_599,N_18482,N_18913);
nor UO_600 (O_600,N_18784,N_19501);
nor UO_601 (O_601,N_18778,N_18103);
and UO_602 (O_602,N_19730,N_19026);
and UO_603 (O_603,N_19391,N_18754);
and UO_604 (O_604,N_18010,N_18400);
nor UO_605 (O_605,N_18381,N_19910);
nor UO_606 (O_606,N_19875,N_19721);
or UO_607 (O_607,N_18441,N_18725);
or UO_608 (O_608,N_18101,N_18539);
and UO_609 (O_609,N_18545,N_19930);
and UO_610 (O_610,N_18929,N_19784);
or UO_611 (O_611,N_18530,N_19678);
xor UO_612 (O_612,N_19420,N_18460);
and UO_613 (O_613,N_19355,N_19511);
or UO_614 (O_614,N_18905,N_18324);
nand UO_615 (O_615,N_18595,N_19035);
xor UO_616 (O_616,N_19234,N_19089);
nand UO_617 (O_617,N_18292,N_18318);
nor UO_618 (O_618,N_19687,N_18352);
xor UO_619 (O_619,N_19757,N_18045);
or UO_620 (O_620,N_19257,N_19189);
or UO_621 (O_621,N_19936,N_18801);
nor UO_622 (O_622,N_19583,N_18782);
nand UO_623 (O_623,N_18795,N_18547);
and UO_624 (O_624,N_19712,N_19092);
nand UO_625 (O_625,N_18396,N_19229);
or UO_626 (O_626,N_18593,N_19423);
or UO_627 (O_627,N_19398,N_19209);
xnor UO_628 (O_628,N_19008,N_18780);
and UO_629 (O_629,N_18509,N_18277);
and UO_630 (O_630,N_18640,N_19202);
or UO_631 (O_631,N_19351,N_18395);
and UO_632 (O_632,N_18690,N_19393);
and UO_633 (O_633,N_19449,N_19818);
nand UO_634 (O_634,N_19828,N_19247);
nor UO_635 (O_635,N_19156,N_19743);
nand UO_636 (O_636,N_19409,N_18867);
or UO_637 (O_637,N_18969,N_19539);
nor UO_638 (O_638,N_18631,N_19953);
xnor UO_639 (O_639,N_18078,N_18568);
and UO_640 (O_640,N_18720,N_19612);
nand UO_641 (O_641,N_19280,N_18065);
xor UO_642 (O_642,N_19057,N_18114);
nor UO_643 (O_643,N_19394,N_18457);
or UO_644 (O_644,N_18609,N_18661);
xnor UO_645 (O_645,N_18772,N_18023);
or UO_646 (O_646,N_18244,N_18956);
nand UO_647 (O_647,N_19009,N_18681);
or UO_648 (O_648,N_18814,N_18703);
and UO_649 (O_649,N_18561,N_18871);
and UO_650 (O_650,N_18964,N_19911);
or UO_651 (O_651,N_18653,N_19996);
nor UO_652 (O_652,N_18021,N_18807);
nor UO_653 (O_653,N_19253,N_18519);
and UO_654 (O_654,N_19580,N_19989);
or UO_655 (O_655,N_18322,N_18633);
nand UO_656 (O_656,N_18538,N_18879);
nand UO_657 (O_657,N_18993,N_19467);
and UO_658 (O_658,N_18392,N_19004);
and UO_659 (O_659,N_18370,N_19797);
nand UO_660 (O_660,N_18946,N_18227);
nand UO_661 (O_661,N_19949,N_19854);
xor UO_662 (O_662,N_19287,N_18171);
nor UO_663 (O_663,N_18195,N_18630);
nor UO_664 (O_664,N_18026,N_18736);
or UO_665 (O_665,N_18259,N_18786);
xnor UO_666 (O_666,N_19013,N_18153);
nand UO_667 (O_667,N_19510,N_19154);
or UO_668 (O_668,N_18375,N_18953);
nor UO_669 (O_669,N_18882,N_18941);
xnor UO_670 (O_670,N_19523,N_19954);
nor UO_671 (O_671,N_18306,N_18600);
nor UO_672 (O_672,N_18860,N_19688);
and UO_673 (O_673,N_19330,N_19145);
nor UO_674 (O_674,N_18914,N_18835);
nand UO_675 (O_675,N_19543,N_19337);
and UO_676 (O_676,N_18555,N_18368);
nor UO_677 (O_677,N_19001,N_19217);
and UO_678 (O_678,N_19723,N_18745);
or UO_679 (O_679,N_19364,N_19149);
or UO_680 (O_680,N_18190,N_18537);
nand UO_681 (O_681,N_19403,N_19826);
and UO_682 (O_682,N_19813,N_19395);
xnor UO_683 (O_683,N_18263,N_18080);
or UO_684 (O_684,N_18127,N_18820);
nand UO_685 (O_685,N_18740,N_18565);
nor UO_686 (O_686,N_18475,N_19968);
and UO_687 (O_687,N_19578,N_19356);
or UO_688 (O_688,N_18823,N_18498);
or UO_689 (O_689,N_19070,N_19585);
xor UO_690 (O_690,N_18649,N_18331);
and UO_691 (O_691,N_18204,N_19269);
nor UO_692 (O_692,N_18927,N_19226);
and UO_693 (O_693,N_19316,N_18942);
or UO_694 (O_694,N_19582,N_19620);
and UO_695 (O_695,N_18366,N_18199);
xor UO_696 (O_696,N_19963,N_19958);
or UO_697 (O_697,N_18042,N_19101);
nand UO_698 (O_698,N_18014,N_19464);
xor UO_699 (O_699,N_18465,N_19594);
and UO_700 (O_700,N_18334,N_19526);
and UO_701 (O_701,N_19724,N_19066);
or UO_702 (O_702,N_19804,N_19673);
nor UO_703 (O_703,N_18383,N_18047);
nand UO_704 (O_704,N_19045,N_19126);
nand UO_705 (O_705,N_18855,N_19025);
nor UO_706 (O_706,N_19759,N_18490);
nor UO_707 (O_707,N_19959,N_19425);
nor UO_708 (O_708,N_18810,N_18974);
nand UO_709 (O_709,N_19362,N_19375);
or UO_710 (O_710,N_18419,N_18140);
and UO_711 (O_711,N_19747,N_19889);
xor UO_712 (O_712,N_18658,N_18071);
or UO_713 (O_713,N_19837,N_19556);
nand UO_714 (O_714,N_18944,N_19378);
nor UO_715 (O_715,N_18546,N_19334);
or UO_716 (O_716,N_19047,N_18330);
nand UO_717 (O_717,N_19584,N_18129);
or UO_718 (O_718,N_18262,N_18806);
and UO_719 (O_719,N_18908,N_18790);
nor UO_720 (O_720,N_19235,N_19349);
nand UO_721 (O_721,N_19353,N_18694);
and UO_722 (O_722,N_18788,N_19506);
nor UO_723 (O_723,N_19540,N_18730);
or UO_724 (O_724,N_19965,N_19141);
or UO_725 (O_725,N_18329,N_18389);
nor UO_726 (O_726,N_18206,N_18326);
nor UO_727 (O_727,N_19642,N_19432);
nand UO_728 (O_728,N_19241,N_18417);
or UO_729 (O_729,N_19256,N_18391);
or UO_730 (O_730,N_18706,N_18123);
nor UO_731 (O_731,N_18599,N_18949);
or UO_732 (O_732,N_18388,N_19249);
and UO_733 (O_733,N_19384,N_18041);
or UO_734 (O_734,N_18437,N_19664);
or UO_735 (O_735,N_18230,N_18636);
xnor UO_736 (O_736,N_19751,N_19028);
and UO_737 (O_737,N_19775,N_18606);
nand UO_738 (O_738,N_18119,N_19470);
or UO_739 (O_739,N_19558,N_18798);
nand UO_740 (O_740,N_19272,N_18040);
nor UO_741 (O_741,N_18931,N_18676);
or UO_742 (O_742,N_19236,N_19533);
and UO_743 (O_743,N_19952,N_18883);
nand UO_744 (O_744,N_19199,N_19102);
and UO_745 (O_745,N_18248,N_19885);
or UO_746 (O_746,N_18151,N_19833);
nand UO_747 (O_747,N_18269,N_18300);
nand UO_748 (O_748,N_18756,N_19788);
nor UO_749 (O_749,N_19341,N_19706);
and UO_750 (O_750,N_19169,N_18385);
xnor UO_751 (O_751,N_19792,N_19890);
and UO_752 (O_752,N_18958,N_18108);
nand UO_753 (O_753,N_19279,N_19254);
nand UO_754 (O_754,N_18341,N_19112);
xor UO_755 (O_755,N_19181,N_18360);
or UO_756 (O_756,N_19593,N_19843);
nand UO_757 (O_757,N_19416,N_19128);
and UO_758 (O_758,N_19586,N_19799);
nand UO_759 (O_759,N_18499,N_18714);
nand UO_760 (O_760,N_18399,N_18285);
or UO_761 (O_761,N_18148,N_18448);
nor UO_762 (O_762,N_19931,N_19771);
nand UO_763 (O_763,N_18284,N_19686);
and UO_764 (O_764,N_19067,N_18104);
nand UO_765 (O_765,N_19614,N_19427);
nand UO_766 (O_766,N_18216,N_19801);
xnor UO_767 (O_767,N_18077,N_18301);
nand UO_768 (O_768,N_18458,N_19319);
xnor UO_769 (O_769,N_19366,N_18410);
nor UO_770 (O_770,N_19868,N_19227);
nand UO_771 (O_771,N_18709,N_18393);
nor UO_772 (O_772,N_19948,N_19379);
nand UO_773 (O_773,N_19088,N_18485);
or UO_774 (O_774,N_18157,N_19104);
or UO_775 (O_775,N_19336,N_19453);
or UO_776 (O_776,N_18150,N_19458);
nand UO_777 (O_777,N_18083,N_18744);
nand UO_778 (O_778,N_18551,N_18899);
xnor UO_779 (O_779,N_19940,N_19251);
or UO_780 (O_780,N_18155,N_18369);
or UO_781 (O_781,N_18302,N_18868);
or UO_782 (O_782,N_18337,N_19426);
and UO_783 (O_783,N_19599,N_19109);
nor UO_784 (O_784,N_19893,N_18675);
nand UO_785 (O_785,N_18831,N_18486);
and UO_786 (O_786,N_19637,N_19905);
nand UO_787 (O_787,N_19114,N_18943);
or UO_788 (O_788,N_18353,N_19789);
and UO_789 (O_789,N_19327,N_18459);
nand UO_790 (O_790,N_18533,N_18773);
nor UO_791 (O_791,N_19338,N_18358);
and UO_792 (O_792,N_18702,N_19301);
or UO_793 (O_793,N_18464,N_19085);
nor UO_794 (O_794,N_18837,N_18420);
nand UO_795 (O_795,N_18976,N_19442);
and UO_796 (O_796,N_19475,N_18152);
nor UO_797 (O_797,N_18916,N_18384);
nor UO_798 (O_798,N_19608,N_18971);
nor UO_799 (O_799,N_19059,N_18613);
or UO_800 (O_800,N_19626,N_18767);
xor UO_801 (O_801,N_19851,N_18888);
nand UO_802 (O_802,N_18261,N_19115);
nand UO_803 (O_803,N_18111,N_19079);
nand UO_804 (O_804,N_19296,N_19167);
nand UO_805 (O_805,N_18210,N_19100);
and UO_806 (O_806,N_18275,N_18118);
nand UO_807 (O_807,N_19932,N_19736);
xnor UO_808 (O_808,N_18476,N_18869);
xnor UO_809 (O_809,N_19404,N_18828);
or UO_810 (O_810,N_19225,N_19148);
and UO_811 (O_811,N_18166,N_18608);
and UO_812 (O_812,N_19383,N_18310);
xor UO_813 (O_813,N_19443,N_19210);
nand UO_814 (O_814,N_18453,N_19973);
nor UO_815 (O_815,N_19758,N_19616);
and UO_816 (O_816,N_18158,N_18587);
and UO_817 (O_817,N_18346,N_18818);
nand UO_818 (O_818,N_18287,N_18623);
or UO_819 (O_819,N_18920,N_18492);
or UO_820 (O_820,N_18793,N_18881);
or UO_821 (O_821,N_19995,N_19676);
nor UO_822 (O_822,N_19829,N_18234);
xnor UO_823 (O_823,N_19417,N_19215);
or UO_824 (O_824,N_19591,N_18139);
and UO_825 (O_825,N_18813,N_18829);
and UO_826 (O_826,N_18674,N_18548);
or UO_827 (O_827,N_19587,N_18579);
nor UO_828 (O_828,N_19159,N_18167);
nand UO_829 (O_829,N_18376,N_18355);
nor UO_830 (O_830,N_19389,N_18750);
and UO_831 (O_831,N_19216,N_18268);
nand UO_832 (O_832,N_19927,N_19683);
nor UO_833 (O_833,N_19942,N_18892);
nand UO_834 (O_834,N_18462,N_19171);
or UO_835 (O_835,N_19979,N_18695);
nand UO_836 (O_836,N_19504,N_19000);
nand UO_837 (O_837,N_18984,N_18255);
nor UO_838 (O_838,N_18339,N_18526);
and UO_839 (O_839,N_19780,N_19916);
or UO_840 (O_840,N_19061,N_19457);
xnor UO_841 (O_841,N_18945,N_19060);
or UO_842 (O_842,N_19668,N_19228);
nor UO_843 (O_843,N_18763,N_18876);
nor UO_844 (O_844,N_18875,N_19388);
and UO_845 (O_845,N_18222,N_18433);
nor UO_846 (O_846,N_18267,N_19783);
nand UO_847 (O_847,N_19643,N_19701);
nand UO_848 (O_848,N_19155,N_19382);
nand UO_849 (O_849,N_19988,N_18491);
and UO_850 (O_850,N_19987,N_19038);
and UO_851 (O_851,N_19692,N_18874);
nand UO_852 (O_852,N_18401,N_18704);
nand UO_853 (O_853,N_18522,N_19200);
xnor UO_854 (O_854,N_18046,N_19947);
nor UO_855 (O_855,N_19479,N_18822);
nand UO_856 (O_856,N_19913,N_19168);
and UO_857 (O_857,N_18266,N_18924);
and UO_858 (O_858,N_18474,N_19242);
xor UO_859 (O_859,N_18372,N_18663);
and UO_860 (O_860,N_18051,N_19399);
nor UO_861 (O_861,N_18598,N_18502);
nor UO_862 (O_862,N_19259,N_18781);
nor UO_863 (O_863,N_18859,N_18379);
or UO_864 (O_864,N_19628,N_19130);
xor UO_865 (O_865,N_19967,N_18193);
nand UO_866 (O_866,N_18947,N_19113);
or UO_867 (O_867,N_19961,N_19870);
or UO_868 (O_868,N_18028,N_18939);
and UO_869 (O_869,N_19195,N_19289);
nor UO_870 (O_870,N_18746,N_18637);
nand UO_871 (O_871,N_18213,N_19779);
nand UO_872 (O_872,N_18651,N_19917);
xnor UO_873 (O_873,N_18770,N_19252);
xor UO_874 (O_874,N_19534,N_18844);
and UO_875 (O_875,N_19390,N_18135);
nor UO_876 (O_876,N_19970,N_19705);
and UO_877 (O_877,N_18516,N_18435);
or UO_878 (O_878,N_19513,N_18525);
nand UO_879 (O_879,N_19131,N_19919);
and UO_880 (O_880,N_18252,N_18079);
or UO_881 (O_881,N_19034,N_18228);
nor UO_882 (O_882,N_19118,N_18402);
and UO_883 (O_883,N_19429,N_19782);
nor UO_884 (O_884,N_19010,N_18708);
and UO_885 (O_885,N_18270,N_19125);
or UO_886 (O_886,N_19731,N_18247);
or UO_887 (O_887,N_19613,N_19861);
nand UO_888 (O_888,N_18696,N_18187);
and UO_889 (O_889,N_18008,N_19920);
nand UO_890 (O_890,N_18106,N_19928);
nand UO_891 (O_891,N_18768,N_18501);
xor UO_892 (O_892,N_18426,N_18717);
nor UO_893 (O_893,N_18722,N_19187);
nand UO_894 (O_894,N_18154,N_18480);
nor UO_895 (O_895,N_19282,N_18163);
and UO_896 (O_896,N_18403,N_18436);
xor UO_897 (O_897,N_18164,N_18902);
nand UO_898 (O_898,N_18523,N_18030);
xor UO_899 (O_899,N_19095,N_19091);
or UO_900 (O_900,N_19835,N_18315);
nand UO_901 (O_901,N_19419,N_19907);
nand UO_902 (O_902,N_19450,N_19012);
nor UO_903 (O_903,N_19709,N_19636);
nand UO_904 (O_904,N_19562,N_18664);
nor UO_905 (O_905,N_18289,N_18850);
nor UO_906 (O_906,N_18919,N_18758);
or UO_907 (O_907,N_18716,N_19218);
nand UO_908 (O_908,N_18348,N_18851);
and UO_909 (O_909,N_18765,N_18701);
nand UO_910 (O_910,N_19489,N_18149);
or UO_911 (O_911,N_19809,N_18029);
nor UO_912 (O_912,N_19852,N_18627);
or UO_913 (O_913,N_19634,N_19999);
nand UO_914 (O_914,N_18468,N_19769);
nor UO_915 (O_915,N_18182,N_19022);
xor UO_916 (O_916,N_19507,N_19727);
nor UO_917 (O_917,N_18335,N_18518);
and UO_918 (O_918,N_18069,N_19863);
and UO_919 (O_919,N_19755,N_19898);
nand UO_920 (O_920,N_18408,N_19040);
nand UO_921 (O_921,N_19190,N_18361);
nor UO_922 (O_922,N_18483,N_18039);
nand UO_923 (O_923,N_19122,N_18766);
nand UO_924 (O_924,N_19136,N_19922);
nor UO_925 (O_925,N_19158,N_19603);
and UO_926 (O_926,N_18061,N_18832);
and UO_927 (O_927,N_19494,N_19808);
nor UO_928 (O_928,N_18759,N_19653);
nor UO_929 (O_929,N_18000,N_18611);
nor UO_930 (O_930,N_18748,N_19014);
or UO_931 (O_931,N_19340,N_19326);
or UO_932 (O_932,N_19297,N_19073);
or UO_933 (O_933,N_19054,N_18422);
and UO_934 (O_934,N_19975,N_19825);
or UO_935 (O_935,N_18536,N_19466);
nor UO_936 (O_936,N_18531,N_19690);
or UO_937 (O_937,N_19696,N_18454);
or UO_938 (O_938,N_18853,N_19273);
xnor UO_939 (O_939,N_19992,N_18288);
or UO_940 (O_940,N_18713,N_18635);
and UO_941 (O_941,N_18235,N_19859);
xnor UO_942 (O_942,N_19881,N_18176);
nor UO_943 (O_943,N_19659,N_18932);
nand UO_944 (O_944,N_19469,N_19923);
or UO_945 (O_945,N_19261,N_18979);
nor UO_946 (O_946,N_19377,N_18799);
or UO_947 (O_947,N_18097,N_19742);
or UO_948 (O_948,N_18347,N_19490);
nand UO_949 (O_949,N_18312,N_19811);
nor UO_950 (O_950,N_19729,N_19428);
and UO_951 (O_951,N_18356,N_19698);
nand UO_952 (O_952,N_18242,N_18824);
nand UO_953 (O_953,N_18898,N_18808);
or UO_954 (O_954,N_19839,N_18406);
and UO_955 (O_955,N_19260,N_19357);
and UO_956 (O_956,N_19660,N_19981);
or UO_957 (O_957,N_18414,N_19986);
or UO_958 (O_958,N_18642,N_18999);
nor UO_959 (O_959,N_18257,N_19502);
or UO_960 (O_960,N_19841,N_18439);
or UO_961 (O_961,N_18033,N_19233);
and UO_962 (O_962,N_19415,N_18544);
nor UO_963 (O_963,N_19945,N_19749);
xor UO_964 (O_964,N_19641,N_18343);
or UO_965 (O_965,N_19231,N_18434);
nand UO_966 (O_966,N_19440,N_18473);
or UO_967 (O_967,N_18373,N_19474);
and UO_968 (O_968,N_18655,N_18834);
nand UO_969 (O_969,N_18515,N_19650);
nor UO_970 (O_970,N_19270,N_19212);
or UO_971 (O_971,N_19621,N_18062);
xnor UO_972 (O_972,N_19618,N_18146);
or UO_973 (O_973,N_18006,N_18136);
nand UO_974 (O_974,N_18311,N_18607);
and UO_975 (O_975,N_18884,N_19343);
or UO_976 (O_976,N_18848,N_19858);
nand UO_977 (O_977,N_18495,N_18179);
nor UO_978 (O_978,N_19617,N_18845);
nand UO_979 (O_979,N_19538,N_19576);
and UO_980 (O_980,N_19108,N_19887);
nand UO_981 (O_981,N_19207,N_18313);
nor UO_982 (O_982,N_19087,N_19715);
nand UO_983 (O_983,N_18989,N_18444);
xnor UO_984 (O_984,N_19445,N_18865);
and UO_985 (O_985,N_18504,N_19039);
nand UO_986 (O_986,N_18705,N_19134);
nor UO_987 (O_987,N_18479,N_19413);
and UO_988 (O_988,N_19912,N_18332);
and UO_989 (O_989,N_19748,N_19240);
nor UO_990 (O_990,N_18124,N_19677);
nand UO_991 (O_991,N_19805,N_19803);
or UO_992 (O_992,N_18390,N_18965);
nor UO_993 (O_993,N_19052,N_19213);
or UO_994 (O_994,N_19848,N_19519);
and UO_995 (O_995,N_19793,N_19993);
and UO_996 (O_996,N_18619,N_19572);
or UO_997 (O_997,N_18592,N_18576);
and UO_998 (O_998,N_18090,N_18243);
and UO_999 (O_999,N_19293,N_19150);
nand UO_1000 (O_1000,N_18317,N_18851);
nor UO_1001 (O_1001,N_18100,N_18755);
nand UO_1002 (O_1002,N_18126,N_19122);
xnor UO_1003 (O_1003,N_19437,N_19139);
and UO_1004 (O_1004,N_19780,N_18538);
nor UO_1005 (O_1005,N_19362,N_19603);
nand UO_1006 (O_1006,N_19714,N_18458);
nor UO_1007 (O_1007,N_18034,N_18294);
xnor UO_1008 (O_1008,N_18483,N_19848);
nor UO_1009 (O_1009,N_19476,N_18235);
nor UO_1010 (O_1010,N_18485,N_19664);
nand UO_1011 (O_1011,N_19392,N_18529);
nor UO_1012 (O_1012,N_18887,N_18809);
nor UO_1013 (O_1013,N_18383,N_18268);
nor UO_1014 (O_1014,N_18150,N_18172);
or UO_1015 (O_1015,N_18512,N_19559);
xor UO_1016 (O_1016,N_18375,N_18881);
nor UO_1017 (O_1017,N_18295,N_19816);
and UO_1018 (O_1018,N_18547,N_19787);
nor UO_1019 (O_1019,N_18712,N_18363);
nor UO_1020 (O_1020,N_19134,N_18698);
nand UO_1021 (O_1021,N_19318,N_18433);
and UO_1022 (O_1022,N_19267,N_18797);
or UO_1023 (O_1023,N_18616,N_18998);
nand UO_1024 (O_1024,N_18634,N_19166);
xor UO_1025 (O_1025,N_19057,N_18854);
xor UO_1026 (O_1026,N_18000,N_19544);
and UO_1027 (O_1027,N_18643,N_18054);
and UO_1028 (O_1028,N_19024,N_19080);
nor UO_1029 (O_1029,N_18596,N_18351);
or UO_1030 (O_1030,N_19178,N_19988);
and UO_1031 (O_1031,N_19608,N_18640);
nor UO_1032 (O_1032,N_18486,N_18146);
nand UO_1033 (O_1033,N_18550,N_18279);
and UO_1034 (O_1034,N_18306,N_19852);
nand UO_1035 (O_1035,N_19731,N_18345);
nand UO_1036 (O_1036,N_18110,N_19570);
xor UO_1037 (O_1037,N_19417,N_19429);
and UO_1038 (O_1038,N_19188,N_18076);
nand UO_1039 (O_1039,N_18317,N_19359);
or UO_1040 (O_1040,N_18887,N_18320);
xnor UO_1041 (O_1041,N_18698,N_18028);
and UO_1042 (O_1042,N_18732,N_19204);
nand UO_1043 (O_1043,N_19605,N_19114);
or UO_1044 (O_1044,N_19980,N_18706);
and UO_1045 (O_1045,N_18627,N_18750);
and UO_1046 (O_1046,N_18941,N_19778);
or UO_1047 (O_1047,N_18069,N_19284);
and UO_1048 (O_1048,N_18389,N_19821);
or UO_1049 (O_1049,N_18798,N_18899);
xnor UO_1050 (O_1050,N_19645,N_18055);
xor UO_1051 (O_1051,N_18901,N_19988);
xor UO_1052 (O_1052,N_18895,N_19354);
nand UO_1053 (O_1053,N_19245,N_18667);
xor UO_1054 (O_1054,N_18106,N_19001);
or UO_1055 (O_1055,N_19893,N_19934);
and UO_1056 (O_1056,N_18689,N_19477);
nand UO_1057 (O_1057,N_18897,N_19162);
or UO_1058 (O_1058,N_19357,N_19765);
nand UO_1059 (O_1059,N_19466,N_18902);
nor UO_1060 (O_1060,N_18828,N_18036);
nor UO_1061 (O_1061,N_19956,N_19512);
nor UO_1062 (O_1062,N_19090,N_19666);
and UO_1063 (O_1063,N_19966,N_18726);
xnor UO_1064 (O_1064,N_19548,N_19402);
xnor UO_1065 (O_1065,N_19013,N_19140);
or UO_1066 (O_1066,N_18312,N_18029);
nand UO_1067 (O_1067,N_19852,N_18554);
and UO_1068 (O_1068,N_19455,N_18535);
nor UO_1069 (O_1069,N_18953,N_18554);
nor UO_1070 (O_1070,N_19588,N_18292);
nor UO_1071 (O_1071,N_19093,N_19196);
nor UO_1072 (O_1072,N_19316,N_19081);
or UO_1073 (O_1073,N_18158,N_19507);
nor UO_1074 (O_1074,N_19745,N_18467);
and UO_1075 (O_1075,N_19465,N_19481);
nor UO_1076 (O_1076,N_18364,N_18445);
or UO_1077 (O_1077,N_18883,N_18662);
nand UO_1078 (O_1078,N_18989,N_19469);
xnor UO_1079 (O_1079,N_18196,N_18915);
or UO_1080 (O_1080,N_18673,N_19919);
and UO_1081 (O_1081,N_18186,N_18169);
or UO_1082 (O_1082,N_18087,N_18216);
nor UO_1083 (O_1083,N_19914,N_19733);
and UO_1084 (O_1084,N_19496,N_19154);
and UO_1085 (O_1085,N_19120,N_18320);
nand UO_1086 (O_1086,N_18321,N_19696);
nand UO_1087 (O_1087,N_19259,N_18427);
nand UO_1088 (O_1088,N_19257,N_19960);
nor UO_1089 (O_1089,N_19690,N_18211);
or UO_1090 (O_1090,N_18249,N_19942);
nand UO_1091 (O_1091,N_19747,N_18651);
or UO_1092 (O_1092,N_18364,N_19287);
nor UO_1093 (O_1093,N_19340,N_19683);
and UO_1094 (O_1094,N_19672,N_19869);
nand UO_1095 (O_1095,N_18591,N_19823);
or UO_1096 (O_1096,N_19750,N_19043);
or UO_1097 (O_1097,N_18542,N_19153);
and UO_1098 (O_1098,N_18792,N_19397);
nor UO_1099 (O_1099,N_19991,N_19891);
xnor UO_1100 (O_1100,N_18355,N_19352);
nor UO_1101 (O_1101,N_19770,N_19511);
and UO_1102 (O_1102,N_18855,N_18461);
and UO_1103 (O_1103,N_19797,N_18596);
or UO_1104 (O_1104,N_18144,N_19002);
nor UO_1105 (O_1105,N_18900,N_19592);
or UO_1106 (O_1106,N_19861,N_19205);
or UO_1107 (O_1107,N_18965,N_19432);
nand UO_1108 (O_1108,N_18852,N_18902);
nor UO_1109 (O_1109,N_19508,N_19435);
or UO_1110 (O_1110,N_19174,N_19261);
nand UO_1111 (O_1111,N_19340,N_19976);
and UO_1112 (O_1112,N_19021,N_19024);
nor UO_1113 (O_1113,N_19075,N_18514);
and UO_1114 (O_1114,N_18919,N_18360);
and UO_1115 (O_1115,N_19533,N_19230);
nor UO_1116 (O_1116,N_18522,N_19480);
or UO_1117 (O_1117,N_18982,N_18034);
xnor UO_1118 (O_1118,N_18576,N_18738);
xor UO_1119 (O_1119,N_19809,N_19116);
nand UO_1120 (O_1120,N_19253,N_19057);
and UO_1121 (O_1121,N_19270,N_19674);
nand UO_1122 (O_1122,N_18889,N_18480);
nand UO_1123 (O_1123,N_18823,N_18857);
or UO_1124 (O_1124,N_18396,N_19668);
and UO_1125 (O_1125,N_18855,N_18417);
nor UO_1126 (O_1126,N_18666,N_18992);
and UO_1127 (O_1127,N_19863,N_19963);
and UO_1128 (O_1128,N_19521,N_18571);
nand UO_1129 (O_1129,N_18382,N_18554);
nor UO_1130 (O_1130,N_18353,N_19021);
nand UO_1131 (O_1131,N_19235,N_18418);
nor UO_1132 (O_1132,N_19171,N_18617);
xor UO_1133 (O_1133,N_18215,N_19083);
nand UO_1134 (O_1134,N_18882,N_19510);
or UO_1135 (O_1135,N_18785,N_18052);
or UO_1136 (O_1136,N_18163,N_18202);
and UO_1137 (O_1137,N_19554,N_19521);
nand UO_1138 (O_1138,N_19967,N_19425);
nor UO_1139 (O_1139,N_18134,N_18905);
nor UO_1140 (O_1140,N_19965,N_18916);
nand UO_1141 (O_1141,N_18107,N_19476);
nor UO_1142 (O_1142,N_19777,N_18935);
and UO_1143 (O_1143,N_19118,N_18863);
and UO_1144 (O_1144,N_18086,N_19787);
and UO_1145 (O_1145,N_19078,N_19119);
and UO_1146 (O_1146,N_19036,N_18880);
nand UO_1147 (O_1147,N_18719,N_18697);
nor UO_1148 (O_1148,N_18506,N_19188);
and UO_1149 (O_1149,N_18978,N_19333);
and UO_1150 (O_1150,N_19450,N_19380);
and UO_1151 (O_1151,N_19348,N_19302);
or UO_1152 (O_1152,N_19486,N_19520);
and UO_1153 (O_1153,N_19684,N_18056);
or UO_1154 (O_1154,N_18949,N_19792);
nand UO_1155 (O_1155,N_18678,N_19648);
or UO_1156 (O_1156,N_18891,N_19544);
nor UO_1157 (O_1157,N_19631,N_19749);
and UO_1158 (O_1158,N_19200,N_18591);
nor UO_1159 (O_1159,N_19837,N_18003);
nand UO_1160 (O_1160,N_19201,N_19722);
nand UO_1161 (O_1161,N_19987,N_18087);
and UO_1162 (O_1162,N_18457,N_18923);
or UO_1163 (O_1163,N_18813,N_19911);
nor UO_1164 (O_1164,N_19542,N_18275);
nor UO_1165 (O_1165,N_19929,N_19713);
nor UO_1166 (O_1166,N_18797,N_18976);
nor UO_1167 (O_1167,N_18038,N_18925);
or UO_1168 (O_1168,N_19681,N_19149);
nand UO_1169 (O_1169,N_19667,N_19905);
or UO_1170 (O_1170,N_18477,N_19311);
or UO_1171 (O_1171,N_19922,N_18862);
nor UO_1172 (O_1172,N_18054,N_18335);
nor UO_1173 (O_1173,N_18429,N_19248);
nand UO_1174 (O_1174,N_19607,N_18538);
nor UO_1175 (O_1175,N_18661,N_18628);
or UO_1176 (O_1176,N_19954,N_18561);
nand UO_1177 (O_1177,N_19407,N_19106);
and UO_1178 (O_1178,N_18497,N_19420);
and UO_1179 (O_1179,N_19246,N_19834);
nand UO_1180 (O_1180,N_19980,N_18301);
and UO_1181 (O_1181,N_19332,N_19781);
xnor UO_1182 (O_1182,N_18736,N_18507);
and UO_1183 (O_1183,N_19877,N_18542);
xnor UO_1184 (O_1184,N_18068,N_18722);
and UO_1185 (O_1185,N_18914,N_19509);
nand UO_1186 (O_1186,N_18116,N_19772);
and UO_1187 (O_1187,N_19813,N_18264);
or UO_1188 (O_1188,N_18368,N_19972);
or UO_1189 (O_1189,N_19973,N_19675);
xnor UO_1190 (O_1190,N_19529,N_19353);
nand UO_1191 (O_1191,N_18819,N_18305);
nor UO_1192 (O_1192,N_18552,N_19460);
xnor UO_1193 (O_1193,N_18528,N_19540);
nand UO_1194 (O_1194,N_19991,N_19710);
or UO_1195 (O_1195,N_18401,N_19242);
or UO_1196 (O_1196,N_19165,N_18963);
xnor UO_1197 (O_1197,N_19991,N_18239);
nor UO_1198 (O_1198,N_19194,N_19048);
nor UO_1199 (O_1199,N_18360,N_19262);
nand UO_1200 (O_1200,N_19917,N_18253);
or UO_1201 (O_1201,N_18924,N_19112);
or UO_1202 (O_1202,N_18520,N_18696);
or UO_1203 (O_1203,N_18588,N_18029);
or UO_1204 (O_1204,N_19514,N_18241);
nor UO_1205 (O_1205,N_19494,N_19447);
nor UO_1206 (O_1206,N_18000,N_19570);
nor UO_1207 (O_1207,N_18616,N_18520);
xor UO_1208 (O_1208,N_18565,N_18588);
nand UO_1209 (O_1209,N_19788,N_18723);
or UO_1210 (O_1210,N_18382,N_18078);
or UO_1211 (O_1211,N_18946,N_19539);
or UO_1212 (O_1212,N_19000,N_18794);
nor UO_1213 (O_1213,N_19589,N_18137);
and UO_1214 (O_1214,N_18422,N_19418);
and UO_1215 (O_1215,N_19346,N_19656);
nor UO_1216 (O_1216,N_19534,N_18066);
xor UO_1217 (O_1217,N_19676,N_18484);
or UO_1218 (O_1218,N_19952,N_19031);
xnor UO_1219 (O_1219,N_18055,N_18447);
nor UO_1220 (O_1220,N_18684,N_18584);
or UO_1221 (O_1221,N_19164,N_19124);
nand UO_1222 (O_1222,N_18771,N_18144);
and UO_1223 (O_1223,N_19643,N_19597);
nand UO_1224 (O_1224,N_19414,N_18763);
xor UO_1225 (O_1225,N_19066,N_18497);
or UO_1226 (O_1226,N_18975,N_18439);
nand UO_1227 (O_1227,N_19427,N_19336);
nor UO_1228 (O_1228,N_19507,N_18735);
and UO_1229 (O_1229,N_18010,N_18570);
xor UO_1230 (O_1230,N_19632,N_18283);
nand UO_1231 (O_1231,N_19604,N_19557);
or UO_1232 (O_1232,N_19028,N_18951);
and UO_1233 (O_1233,N_18686,N_19815);
nand UO_1234 (O_1234,N_19890,N_18909);
nor UO_1235 (O_1235,N_18754,N_19453);
or UO_1236 (O_1236,N_19781,N_19612);
nand UO_1237 (O_1237,N_19253,N_18083);
nor UO_1238 (O_1238,N_19267,N_19889);
or UO_1239 (O_1239,N_18184,N_19779);
nand UO_1240 (O_1240,N_18669,N_18804);
nand UO_1241 (O_1241,N_19935,N_19840);
nand UO_1242 (O_1242,N_19372,N_18102);
and UO_1243 (O_1243,N_19805,N_19928);
nor UO_1244 (O_1244,N_19190,N_19628);
or UO_1245 (O_1245,N_19072,N_19360);
or UO_1246 (O_1246,N_18697,N_18612);
and UO_1247 (O_1247,N_18260,N_19380);
nor UO_1248 (O_1248,N_18657,N_18046);
nor UO_1249 (O_1249,N_19526,N_18717);
nor UO_1250 (O_1250,N_19965,N_19501);
or UO_1251 (O_1251,N_18980,N_18743);
nor UO_1252 (O_1252,N_18885,N_18044);
nand UO_1253 (O_1253,N_19299,N_18779);
and UO_1254 (O_1254,N_19482,N_18753);
and UO_1255 (O_1255,N_18745,N_18010);
and UO_1256 (O_1256,N_19069,N_19182);
and UO_1257 (O_1257,N_18641,N_19878);
nor UO_1258 (O_1258,N_18696,N_18289);
nand UO_1259 (O_1259,N_19117,N_19639);
nor UO_1260 (O_1260,N_18147,N_19285);
and UO_1261 (O_1261,N_18299,N_19771);
nand UO_1262 (O_1262,N_18022,N_19321);
xor UO_1263 (O_1263,N_18789,N_19499);
nand UO_1264 (O_1264,N_19672,N_19266);
nor UO_1265 (O_1265,N_18902,N_19703);
and UO_1266 (O_1266,N_19297,N_18272);
nand UO_1267 (O_1267,N_19924,N_19436);
or UO_1268 (O_1268,N_18090,N_18916);
nand UO_1269 (O_1269,N_19638,N_19333);
and UO_1270 (O_1270,N_18819,N_19056);
nand UO_1271 (O_1271,N_18712,N_19374);
and UO_1272 (O_1272,N_18216,N_18426);
or UO_1273 (O_1273,N_18982,N_18118);
nand UO_1274 (O_1274,N_19519,N_18193);
or UO_1275 (O_1275,N_19710,N_18412);
nor UO_1276 (O_1276,N_18666,N_19814);
nand UO_1277 (O_1277,N_19033,N_18482);
or UO_1278 (O_1278,N_18965,N_18105);
and UO_1279 (O_1279,N_18101,N_19259);
or UO_1280 (O_1280,N_18956,N_18147);
or UO_1281 (O_1281,N_19895,N_18369);
and UO_1282 (O_1282,N_18909,N_18920);
or UO_1283 (O_1283,N_18963,N_19093);
or UO_1284 (O_1284,N_19469,N_19558);
nand UO_1285 (O_1285,N_18513,N_18128);
and UO_1286 (O_1286,N_18530,N_19696);
nand UO_1287 (O_1287,N_18912,N_19615);
nand UO_1288 (O_1288,N_18254,N_18623);
or UO_1289 (O_1289,N_19390,N_18113);
and UO_1290 (O_1290,N_18487,N_18629);
and UO_1291 (O_1291,N_18114,N_19804);
and UO_1292 (O_1292,N_18138,N_19838);
or UO_1293 (O_1293,N_18043,N_19484);
xnor UO_1294 (O_1294,N_18702,N_19284);
and UO_1295 (O_1295,N_19090,N_18803);
nand UO_1296 (O_1296,N_19460,N_18574);
and UO_1297 (O_1297,N_18304,N_18367);
and UO_1298 (O_1298,N_18886,N_18335);
or UO_1299 (O_1299,N_18617,N_18867);
nor UO_1300 (O_1300,N_18146,N_19152);
and UO_1301 (O_1301,N_19791,N_19185);
or UO_1302 (O_1302,N_18531,N_19971);
xnor UO_1303 (O_1303,N_19464,N_19655);
and UO_1304 (O_1304,N_19728,N_19608);
xnor UO_1305 (O_1305,N_19564,N_18099);
nor UO_1306 (O_1306,N_19791,N_19222);
nor UO_1307 (O_1307,N_19394,N_18516);
and UO_1308 (O_1308,N_18865,N_18730);
and UO_1309 (O_1309,N_19040,N_19502);
nand UO_1310 (O_1310,N_19564,N_18013);
nor UO_1311 (O_1311,N_18998,N_19893);
or UO_1312 (O_1312,N_18029,N_18777);
nor UO_1313 (O_1313,N_18412,N_18120);
xor UO_1314 (O_1314,N_18482,N_19491);
nand UO_1315 (O_1315,N_18486,N_19247);
or UO_1316 (O_1316,N_19875,N_19418);
nand UO_1317 (O_1317,N_18680,N_19224);
nand UO_1318 (O_1318,N_19883,N_18546);
nand UO_1319 (O_1319,N_18801,N_19492);
and UO_1320 (O_1320,N_18506,N_18998);
and UO_1321 (O_1321,N_18890,N_19348);
and UO_1322 (O_1322,N_18613,N_19264);
nor UO_1323 (O_1323,N_18486,N_18479);
nor UO_1324 (O_1324,N_18937,N_18072);
nand UO_1325 (O_1325,N_19241,N_19776);
nand UO_1326 (O_1326,N_19445,N_18797);
and UO_1327 (O_1327,N_18939,N_18410);
nand UO_1328 (O_1328,N_18612,N_19755);
or UO_1329 (O_1329,N_19706,N_18460);
nor UO_1330 (O_1330,N_18650,N_19299);
nand UO_1331 (O_1331,N_18372,N_18751);
nor UO_1332 (O_1332,N_19323,N_19761);
nand UO_1333 (O_1333,N_19144,N_19966);
nor UO_1334 (O_1334,N_18939,N_18864);
nand UO_1335 (O_1335,N_19490,N_18027);
nand UO_1336 (O_1336,N_19775,N_18377);
nor UO_1337 (O_1337,N_19848,N_19818);
and UO_1338 (O_1338,N_19736,N_18299);
or UO_1339 (O_1339,N_18679,N_18900);
nand UO_1340 (O_1340,N_18376,N_18343);
and UO_1341 (O_1341,N_18126,N_19716);
or UO_1342 (O_1342,N_18051,N_19515);
nand UO_1343 (O_1343,N_19990,N_19725);
nor UO_1344 (O_1344,N_19237,N_19624);
nor UO_1345 (O_1345,N_19955,N_18017);
nor UO_1346 (O_1346,N_18255,N_18343);
nor UO_1347 (O_1347,N_18448,N_19675);
and UO_1348 (O_1348,N_19583,N_18576);
or UO_1349 (O_1349,N_19381,N_19435);
nor UO_1350 (O_1350,N_18464,N_19754);
or UO_1351 (O_1351,N_19383,N_19551);
nand UO_1352 (O_1352,N_19400,N_18804);
nand UO_1353 (O_1353,N_18319,N_19900);
nor UO_1354 (O_1354,N_18257,N_19627);
nor UO_1355 (O_1355,N_18045,N_18003);
and UO_1356 (O_1356,N_19940,N_19322);
nand UO_1357 (O_1357,N_18910,N_18555);
and UO_1358 (O_1358,N_18369,N_19066);
nor UO_1359 (O_1359,N_18507,N_19547);
xor UO_1360 (O_1360,N_18146,N_19690);
nand UO_1361 (O_1361,N_19653,N_18154);
or UO_1362 (O_1362,N_19929,N_19256);
nor UO_1363 (O_1363,N_18906,N_19639);
xnor UO_1364 (O_1364,N_18038,N_19882);
nand UO_1365 (O_1365,N_18056,N_19836);
and UO_1366 (O_1366,N_18464,N_19488);
nand UO_1367 (O_1367,N_18562,N_19385);
or UO_1368 (O_1368,N_18797,N_19719);
and UO_1369 (O_1369,N_18297,N_18715);
nand UO_1370 (O_1370,N_19051,N_18111);
and UO_1371 (O_1371,N_18454,N_18270);
xor UO_1372 (O_1372,N_18112,N_18756);
nor UO_1373 (O_1373,N_18777,N_18974);
nand UO_1374 (O_1374,N_18864,N_19020);
and UO_1375 (O_1375,N_18325,N_19650);
nand UO_1376 (O_1376,N_19785,N_18134);
and UO_1377 (O_1377,N_18646,N_19926);
or UO_1378 (O_1378,N_18520,N_19269);
nor UO_1379 (O_1379,N_19336,N_18019);
nand UO_1380 (O_1380,N_19612,N_18317);
or UO_1381 (O_1381,N_19590,N_18861);
nand UO_1382 (O_1382,N_19176,N_18162);
nor UO_1383 (O_1383,N_18575,N_18305);
xnor UO_1384 (O_1384,N_18379,N_18798);
or UO_1385 (O_1385,N_19986,N_18701);
xnor UO_1386 (O_1386,N_19527,N_18414);
nor UO_1387 (O_1387,N_19840,N_19288);
nor UO_1388 (O_1388,N_18550,N_19608);
and UO_1389 (O_1389,N_18685,N_19460);
or UO_1390 (O_1390,N_18668,N_19271);
nor UO_1391 (O_1391,N_19292,N_18149);
nand UO_1392 (O_1392,N_18774,N_18312);
or UO_1393 (O_1393,N_19329,N_19887);
xnor UO_1394 (O_1394,N_18806,N_19874);
nand UO_1395 (O_1395,N_18197,N_19810);
nor UO_1396 (O_1396,N_18192,N_19362);
nor UO_1397 (O_1397,N_19916,N_18789);
and UO_1398 (O_1398,N_19884,N_19977);
xor UO_1399 (O_1399,N_19592,N_18075);
and UO_1400 (O_1400,N_19437,N_19171);
or UO_1401 (O_1401,N_19794,N_18639);
nand UO_1402 (O_1402,N_18699,N_19120);
nand UO_1403 (O_1403,N_18468,N_19916);
nand UO_1404 (O_1404,N_19442,N_18847);
or UO_1405 (O_1405,N_18524,N_19142);
or UO_1406 (O_1406,N_18797,N_18438);
or UO_1407 (O_1407,N_18105,N_19609);
nor UO_1408 (O_1408,N_18168,N_19208);
xnor UO_1409 (O_1409,N_18285,N_18535);
or UO_1410 (O_1410,N_18563,N_18056);
or UO_1411 (O_1411,N_18223,N_18745);
nand UO_1412 (O_1412,N_18456,N_18499);
and UO_1413 (O_1413,N_19305,N_19416);
or UO_1414 (O_1414,N_18079,N_19895);
nand UO_1415 (O_1415,N_18531,N_19315);
nor UO_1416 (O_1416,N_18479,N_18715);
or UO_1417 (O_1417,N_19250,N_18265);
nor UO_1418 (O_1418,N_19375,N_19943);
nand UO_1419 (O_1419,N_19258,N_19747);
nor UO_1420 (O_1420,N_19649,N_19480);
nor UO_1421 (O_1421,N_18054,N_18577);
or UO_1422 (O_1422,N_18822,N_18417);
nor UO_1423 (O_1423,N_19790,N_18728);
and UO_1424 (O_1424,N_18032,N_18160);
nor UO_1425 (O_1425,N_19980,N_18601);
nand UO_1426 (O_1426,N_18424,N_19776);
xnor UO_1427 (O_1427,N_19190,N_18944);
nor UO_1428 (O_1428,N_19251,N_18889);
nor UO_1429 (O_1429,N_19820,N_19483);
nand UO_1430 (O_1430,N_19207,N_19950);
or UO_1431 (O_1431,N_18314,N_19750);
nor UO_1432 (O_1432,N_18968,N_19747);
xnor UO_1433 (O_1433,N_19075,N_19237);
nand UO_1434 (O_1434,N_19801,N_19808);
and UO_1435 (O_1435,N_18654,N_18759);
or UO_1436 (O_1436,N_18998,N_18801);
nand UO_1437 (O_1437,N_19563,N_18783);
nor UO_1438 (O_1438,N_18379,N_18591);
nand UO_1439 (O_1439,N_18352,N_18442);
or UO_1440 (O_1440,N_19953,N_18089);
and UO_1441 (O_1441,N_19804,N_18048);
nand UO_1442 (O_1442,N_18348,N_18724);
nand UO_1443 (O_1443,N_19017,N_19529);
or UO_1444 (O_1444,N_18263,N_19114);
nand UO_1445 (O_1445,N_18246,N_18872);
nand UO_1446 (O_1446,N_18491,N_18419);
and UO_1447 (O_1447,N_19118,N_19326);
xor UO_1448 (O_1448,N_19822,N_19642);
nor UO_1449 (O_1449,N_19281,N_19577);
and UO_1450 (O_1450,N_19660,N_18227);
nor UO_1451 (O_1451,N_18403,N_18961);
xor UO_1452 (O_1452,N_19439,N_18849);
nand UO_1453 (O_1453,N_18717,N_18898);
or UO_1454 (O_1454,N_18131,N_18644);
nand UO_1455 (O_1455,N_18972,N_19914);
nand UO_1456 (O_1456,N_18609,N_19038);
nor UO_1457 (O_1457,N_18688,N_19767);
and UO_1458 (O_1458,N_19532,N_19694);
or UO_1459 (O_1459,N_18105,N_18762);
or UO_1460 (O_1460,N_18343,N_18742);
nor UO_1461 (O_1461,N_19843,N_18771);
nor UO_1462 (O_1462,N_19342,N_18326);
xnor UO_1463 (O_1463,N_18481,N_18929);
or UO_1464 (O_1464,N_18072,N_19446);
and UO_1465 (O_1465,N_18906,N_19633);
nor UO_1466 (O_1466,N_19959,N_18794);
nor UO_1467 (O_1467,N_18749,N_18199);
nand UO_1468 (O_1468,N_18086,N_19948);
and UO_1469 (O_1469,N_18498,N_18345);
xor UO_1470 (O_1470,N_18976,N_19836);
and UO_1471 (O_1471,N_18688,N_18234);
nand UO_1472 (O_1472,N_19521,N_18953);
xor UO_1473 (O_1473,N_19440,N_18300);
nor UO_1474 (O_1474,N_19174,N_18798);
nor UO_1475 (O_1475,N_19115,N_18993);
nand UO_1476 (O_1476,N_19976,N_19382);
nor UO_1477 (O_1477,N_19764,N_19624);
nand UO_1478 (O_1478,N_18145,N_18796);
or UO_1479 (O_1479,N_18704,N_18203);
nand UO_1480 (O_1480,N_19458,N_19957);
or UO_1481 (O_1481,N_18557,N_18213);
nand UO_1482 (O_1482,N_19047,N_19844);
and UO_1483 (O_1483,N_18421,N_19556);
nand UO_1484 (O_1484,N_18019,N_18090);
or UO_1485 (O_1485,N_18371,N_19421);
and UO_1486 (O_1486,N_19640,N_18866);
nand UO_1487 (O_1487,N_18910,N_19380);
and UO_1488 (O_1488,N_18643,N_18549);
and UO_1489 (O_1489,N_19210,N_18801);
nor UO_1490 (O_1490,N_18712,N_19213);
or UO_1491 (O_1491,N_18411,N_19159);
nor UO_1492 (O_1492,N_18563,N_19619);
or UO_1493 (O_1493,N_19918,N_19310);
nand UO_1494 (O_1494,N_18399,N_19746);
and UO_1495 (O_1495,N_19994,N_19829);
xor UO_1496 (O_1496,N_19634,N_18256);
nor UO_1497 (O_1497,N_19406,N_18868);
or UO_1498 (O_1498,N_18049,N_19424);
xor UO_1499 (O_1499,N_19549,N_19265);
xor UO_1500 (O_1500,N_18496,N_18792);
and UO_1501 (O_1501,N_19289,N_19039);
xor UO_1502 (O_1502,N_19033,N_19073);
nand UO_1503 (O_1503,N_18042,N_18298);
and UO_1504 (O_1504,N_18915,N_19769);
nor UO_1505 (O_1505,N_18031,N_19501);
xnor UO_1506 (O_1506,N_19325,N_19417);
nor UO_1507 (O_1507,N_18288,N_19048);
and UO_1508 (O_1508,N_18435,N_19814);
or UO_1509 (O_1509,N_18055,N_18898);
nand UO_1510 (O_1510,N_19457,N_19691);
xnor UO_1511 (O_1511,N_19553,N_18628);
or UO_1512 (O_1512,N_19969,N_18262);
nand UO_1513 (O_1513,N_19440,N_19624);
nand UO_1514 (O_1514,N_19109,N_18674);
or UO_1515 (O_1515,N_19298,N_19110);
nor UO_1516 (O_1516,N_19061,N_19281);
and UO_1517 (O_1517,N_19448,N_18381);
xnor UO_1518 (O_1518,N_19904,N_19166);
and UO_1519 (O_1519,N_18622,N_19418);
and UO_1520 (O_1520,N_19271,N_18682);
or UO_1521 (O_1521,N_18506,N_19980);
nor UO_1522 (O_1522,N_19592,N_19172);
or UO_1523 (O_1523,N_19935,N_19412);
xor UO_1524 (O_1524,N_19641,N_18814);
nor UO_1525 (O_1525,N_19657,N_18628);
xnor UO_1526 (O_1526,N_18186,N_19127);
and UO_1527 (O_1527,N_18742,N_19760);
nor UO_1528 (O_1528,N_19866,N_18798);
xor UO_1529 (O_1529,N_18441,N_18731);
and UO_1530 (O_1530,N_18393,N_18371);
nor UO_1531 (O_1531,N_18583,N_18411);
nand UO_1532 (O_1532,N_18399,N_18668);
and UO_1533 (O_1533,N_18030,N_18603);
or UO_1534 (O_1534,N_19713,N_18462);
nor UO_1535 (O_1535,N_19005,N_18878);
or UO_1536 (O_1536,N_18500,N_19081);
nor UO_1537 (O_1537,N_19606,N_18372);
and UO_1538 (O_1538,N_19637,N_19827);
xor UO_1539 (O_1539,N_19760,N_19508);
nand UO_1540 (O_1540,N_18448,N_19550);
or UO_1541 (O_1541,N_18444,N_18967);
and UO_1542 (O_1542,N_19408,N_18032);
or UO_1543 (O_1543,N_19840,N_19953);
nand UO_1544 (O_1544,N_18992,N_19501);
and UO_1545 (O_1545,N_19800,N_19484);
nor UO_1546 (O_1546,N_18939,N_18982);
nand UO_1547 (O_1547,N_19196,N_19300);
xnor UO_1548 (O_1548,N_19658,N_18606);
or UO_1549 (O_1549,N_18205,N_18418);
and UO_1550 (O_1550,N_18662,N_18983);
nand UO_1551 (O_1551,N_18958,N_19156);
nand UO_1552 (O_1552,N_19953,N_18635);
nor UO_1553 (O_1553,N_18435,N_18170);
nand UO_1554 (O_1554,N_18529,N_18015);
nor UO_1555 (O_1555,N_18431,N_18490);
nor UO_1556 (O_1556,N_19888,N_18223);
and UO_1557 (O_1557,N_18714,N_19370);
nand UO_1558 (O_1558,N_18975,N_18315);
nor UO_1559 (O_1559,N_18515,N_19375);
or UO_1560 (O_1560,N_19706,N_18507);
or UO_1561 (O_1561,N_19822,N_19183);
nand UO_1562 (O_1562,N_19551,N_18166);
and UO_1563 (O_1563,N_19398,N_19777);
xnor UO_1564 (O_1564,N_18737,N_18854);
or UO_1565 (O_1565,N_19289,N_19132);
or UO_1566 (O_1566,N_18945,N_18006);
nor UO_1567 (O_1567,N_18554,N_19963);
and UO_1568 (O_1568,N_18661,N_19883);
nor UO_1569 (O_1569,N_19768,N_18111);
and UO_1570 (O_1570,N_18984,N_18347);
and UO_1571 (O_1571,N_19411,N_18454);
or UO_1572 (O_1572,N_19213,N_18196);
nand UO_1573 (O_1573,N_18660,N_18069);
nor UO_1574 (O_1574,N_19337,N_18124);
nand UO_1575 (O_1575,N_18669,N_18303);
nor UO_1576 (O_1576,N_18877,N_18967);
or UO_1577 (O_1577,N_19035,N_19496);
nand UO_1578 (O_1578,N_18692,N_19471);
nor UO_1579 (O_1579,N_18711,N_19785);
and UO_1580 (O_1580,N_19273,N_18833);
or UO_1581 (O_1581,N_18532,N_18155);
nor UO_1582 (O_1582,N_18396,N_18886);
nand UO_1583 (O_1583,N_18961,N_18762);
nand UO_1584 (O_1584,N_19148,N_19224);
or UO_1585 (O_1585,N_18266,N_18446);
and UO_1586 (O_1586,N_18957,N_18126);
and UO_1587 (O_1587,N_18437,N_19699);
and UO_1588 (O_1588,N_19073,N_18415);
nand UO_1589 (O_1589,N_19698,N_18301);
and UO_1590 (O_1590,N_19728,N_18560);
nor UO_1591 (O_1591,N_19355,N_19930);
or UO_1592 (O_1592,N_18278,N_18907);
nor UO_1593 (O_1593,N_19019,N_19084);
or UO_1594 (O_1594,N_18251,N_18416);
and UO_1595 (O_1595,N_18904,N_19965);
or UO_1596 (O_1596,N_19524,N_18394);
and UO_1597 (O_1597,N_19654,N_18193);
nor UO_1598 (O_1598,N_18362,N_18361);
nand UO_1599 (O_1599,N_19909,N_18338);
or UO_1600 (O_1600,N_18993,N_18833);
and UO_1601 (O_1601,N_18166,N_18219);
xnor UO_1602 (O_1602,N_19312,N_18026);
nor UO_1603 (O_1603,N_18519,N_19639);
xnor UO_1604 (O_1604,N_18549,N_19412);
and UO_1605 (O_1605,N_19149,N_19320);
nor UO_1606 (O_1606,N_18704,N_18543);
xor UO_1607 (O_1607,N_18013,N_19077);
or UO_1608 (O_1608,N_19263,N_18031);
nand UO_1609 (O_1609,N_19579,N_18984);
and UO_1610 (O_1610,N_19659,N_18613);
and UO_1611 (O_1611,N_18374,N_18513);
nand UO_1612 (O_1612,N_19025,N_18635);
nor UO_1613 (O_1613,N_19065,N_18982);
xnor UO_1614 (O_1614,N_18239,N_18135);
and UO_1615 (O_1615,N_18792,N_19900);
nand UO_1616 (O_1616,N_19038,N_18197);
nor UO_1617 (O_1617,N_18577,N_18579);
xor UO_1618 (O_1618,N_18008,N_19907);
nand UO_1619 (O_1619,N_18122,N_19055);
xnor UO_1620 (O_1620,N_19086,N_19420);
or UO_1621 (O_1621,N_18636,N_18522);
nor UO_1622 (O_1622,N_18483,N_19235);
xnor UO_1623 (O_1623,N_19328,N_18841);
nor UO_1624 (O_1624,N_18507,N_19112);
and UO_1625 (O_1625,N_19810,N_19402);
nor UO_1626 (O_1626,N_18844,N_18010);
xor UO_1627 (O_1627,N_18727,N_19563);
nor UO_1628 (O_1628,N_19827,N_18419);
or UO_1629 (O_1629,N_18934,N_19635);
or UO_1630 (O_1630,N_18746,N_18806);
nor UO_1631 (O_1631,N_18870,N_18392);
nand UO_1632 (O_1632,N_19757,N_19267);
or UO_1633 (O_1633,N_18419,N_18170);
nor UO_1634 (O_1634,N_19511,N_18392);
or UO_1635 (O_1635,N_18915,N_18505);
nand UO_1636 (O_1636,N_19102,N_18241);
and UO_1637 (O_1637,N_18274,N_18211);
and UO_1638 (O_1638,N_19443,N_18121);
nor UO_1639 (O_1639,N_18362,N_19984);
and UO_1640 (O_1640,N_19081,N_19158);
nand UO_1641 (O_1641,N_19229,N_19515);
xor UO_1642 (O_1642,N_19616,N_18102);
or UO_1643 (O_1643,N_19819,N_19416);
and UO_1644 (O_1644,N_18221,N_19200);
xor UO_1645 (O_1645,N_18116,N_18884);
or UO_1646 (O_1646,N_19879,N_18699);
nor UO_1647 (O_1647,N_18559,N_18666);
nor UO_1648 (O_1648,N_18589,N_19255);
or UO_1649 (O_1649,N_18881,N_18450);
and UO_1650 (O_1650,N_19952,N_19263);
nand UO_1651 (O_1651,N_19345,N_19481);
nand UO_1652 (O_1652,N_18925,N_18972);
or UO_1653 (O_1653,N_18808,N_19933);
and UO_1654 (O_1654,N_19554,N_18041);
or UO_1655 (O_1655,N_18201,N_18606);
nor UO_1656 (O_1656,N_19755,N_18608);
or UO_1657 (O_1657,N_19553,N_18632);
or UO_1658 (O_1658,N_18629,N_19095);
or UO_1659 (O_1659,N_18865,N_18986);
nor UO_1660 (O_1660,N_18977,N_18150);
nor UO_1661 (O_1661,N_18637,N_18902);
or UO_1662 (O_1662,N_18783,N_19199);
nor UO_1663 (O_1663,N_19348,N_18198);
nor UO_1664 (O_1664,N_18578,N_19132);
or UO_1665 (O_1665,N_19517,N_18914);
or UO_1666 (O_1666,N_18413,N_18148);
or UO_1667 (O_1667,N_19653,N_19879);
nor UO_1668 (O_1668,N_19508,N_19670);
or UO_1669 (O_1669,N_18193,N_18344);
or UO_1670 (O_1670,N_18173,N_19665);
nor UO_1671 (O_1671,N_19540,N_19037);
nor UO_1672 (O_1672,N_19447,N_19608);
nand UO_1673 (O_1673,N_19233,N_19752);
xor UO_1674 (O_1674,N_19389,N_19373);
nand UO_1675 (O_1675,N_18142,N_18936);
or UO_1676 (O_1676,N_19747,N_19294);
and UO_1677 (O_1677,N_18554,N_18951);
or UO_1678 (O_1678,N_19009,N_19209);
or UO_1679 (O_1679,N_18430,N_19160);
and UO_1680 (O_1680,N_19326,N_19777);
and UO_1681 (O_1681,N_19896,N_18859);
nand UO_1682 (O_1682,N_19405,N_18983);
and UO_1683 (O_1683,N_18786,N_19982);
and UO_1684 (O_1684,N_18327,N_18108);
and UO_1685 (O_1685,N_18007,N_18454);
nor UO_1686 (O_1686,N_19728,N_19793);
and UO_1687 (O_1687,N_19804,N_18225);
nand UO_1688 (O_1688,N_19475,N_18155);
nand UO_1689 (O_1689,N_19554,N_19949);
and UO_1690 (O_1690,N_19399,N_19711);
nor UO_1691 (O_1691,N_18919,N_19314);
nor UO_1692 (O_1692,N_18534,N_19333);
and UO_1693 (O_1693,N_19345,N_19252);
nand UO_1694 (O_1694,N_18556,N_18208);
or UO_1695 (O_1695,N_19829,N_19954);
nor UO_1696 (O_1696,N_19212,N_19252);
xor UO_1697 (O_1697,N_18234,N_19761);
or UO_1698 (O_1698,N_19774,N_18689);
nor UO_1699 (O_1699,N_18510,N_19148);
or UO_1700 (O_1700,N_18792,N_19419);
and UO_1701 (O_1701,N_19395,N_19754);
nand UO_1702 (O_1702,N_18170,N_19431);
nor UO_1703 (O_1703,N_19529,N_18082);
and UO_1704 (O_1704,N_19350,N_18894);
nand UO_1705 (O_1705,N_18003,N_18176);
and UO_1706 (O_1706,N_18957,N_18835);
and UO_1707 (O_1707,N_18878,N_19843);
nand UO_1708 (O_1708,N_19037,N_18639);
nor UO_1709 (O_1709,N_18235,N_18584);
nand UO_1710 (O_1710,N_19133,N_18561);
xor UO_1711 (O_1711,N_18482,N_18289);
xor UO_1712 (O_1712,N_18716,N_19823);
nor UO_1713 (O_1713,N_19971,N_18683);
nand UO_1714 (O_1714,N_18960,N_18402);
or UO_1715 (O_1715,N_19701,N_18788);
nand UO_1716 (O_1716,N_19248,N_18141);
nor UO_1717 (O_1717,N_18300,N_18048);
xor UO_1718 (O_1718,N_18486,N_19646);
and UO_1719 (O_1719,N_18593,N_18992);
nor UO_1720 (O_1720,N_18405,N_19476);
and UO_1721 (O_1721,N_18776,N_18606);
xnor UO_1722 (O_1722,N_18292,N_18306);
and UO_1723 (O_1723,N_19277,N_18087);
and UO_1724 (O_1724,N_18524,N_18450);
nand UO_1725 (O_1725,N_19565,N_19148);
or UO_1726 (O_1726,N_19445,N_18533);
and UO_1727 (O_1727,N_19561,N_19471);
nor UO_1728 (O_1728,N_19281,N_18174);
or UO_1729 (O_1729,N_19754,N_18165);
nor UO_1730 (O_1730,N_19106,N_18224);
nor UO_1731 (O_1731,N_18178,N_19388);
and UO_1732 (O_1732,N_18519,N_19569);
and UO_1733 (O_1733,N_18360,N_18438);
xnor UO_1734 (O_1734,N_18088,N_19943);
and UO_1735 (O_1735,N_19031,N_18993);
xnor UO_1736 (O_1736,N_19599,N_19352);
nand UO_1737 (O_1737,N_18394,N_19446);
or UO_1738 (O_1738,N_19925,N_18379);
nand UO_1739 (O_1739,N_19934,N_19130);
nand UO_1740 (O_1740,N_18274,N_18325);
nand UO_1741 (O_1741,N_19505,N_19525);
nor UO_1742 (O_1742,N_19456,N_18474);
or UO_1743 (O_1743,N_18687,N_18776);
nor UO_1744 (O_1744,N_18181,N_19541);
or UO_1745 (O_1745,N_19965,N_18541);
nor UO_1746 (O_1746,N_18657,N_19332);
nand UO_1747 (O_1747,N_18737,N_18455);
or UO_1748 (O_1748,N_18574,N_19275);
nor UO_1749 (O_1749,N_18707,N_19737);
nor UO_1750 (O_1750,N_19556,N_19874);
and UO_1751 (O_1751,N_19509,N_18725);
nand UO_1752 (O_1752,N_18909,N_19051);
nor UO_1753 (O_1753,N_19428,N_18060);
and UO_1754 (O_1754,N_19489,N_19905);
or UO_1755 (O_1755,N_18124,N_19640);
nor UO_1756 (O_1756,N_19620,N_18405);
and UO_1757 (O_1757,N_19911,N_18624);
and UO_1758 (O_1758,N_19476,N_19593);
nand UO_1759 (O_1759,N_18468,N_19125);
and UO_1760 (O_1760,N_18199,N_19469);
nor UO_1761 (O_1761,N_19066,N_18470);
nand UO_1762 (O_1762,N_18646,N_18179);
xnor UO_1763 (O_1763,N_19391,N_19557);
nor UO_1764 (O_1764,N_18316,N_18359);
nor UO_1765 (O_1765,N_19932,N_19067);
nor UO_1766 (O_1766,N_19013,N_18831);
nor UO_1767 (O_1767,N_18184,N_18559);
nor UO_1768 (O_1768,N_19826,N_19423);
nand UO_1769 (O_1769,N_19796,N_19455);
and UO_1770 (O_1770,N_18216,N_18554);
and UO_1771 (O_1771,N_19700,N_19562);
nand UO_1772 (O_1772,N_19672,N_19871);
or UO_1773 (O_1773,N_19117,N_19608);
xor UO_1774 (O_1774,N_18314,N_19631);
and UO_1775 (O_1775,N_18336,N_18005);
xor UO_1776 (O_1776,N_18489,N_18264);
or UO_1777 (O_1777,N_19373,N_19709);
nor UO_1778 (O_1778,N_18707,N_18997);
nand UO_1779 (O_1779,N_19118,N_18626);
nand UO_1780 (O_1780,N_19374,N_18529);
and UO_1781 (O_1781,N_18561,N_18933);
and UO_1782 (O_1782,N_18578,N_18083);
nand UO_1783 (O_1783,N_18865,N_19362);
or UO_1784 (O_1784,N_19457,N_19115);
nor UO_1785 (O_1785,N_18359,N_19915);
or UO_1786 (O_1786,N_18176,N_18707);
nor UO_1787 (O_1787,N_19485,N_19932);
nor UO_1788 (O_1788,N_19226,N_18821);
and UO_1789 (O_1789,N_18130,N_18666);
nor UO_1790 (O_1790,N_18593,N_19274);
nor UO_1791 (O_1791,N_18060,N_19110);
and UO_1792 (O_1792,N_18240,N_18543);
xor UO_1793 (O_1793,N_19310,N_19745);
nor UO_1794 (O_1794,N_19190,N_19756);
nor UO_1795 (O_1795,N_18050,N_18098);
or UO_1796 (O_1796,N_19109,N_19861);
or UO_1797 (O_1797,N_18845,N_19880);
and UO_1798 (O_1798,N_19477,N_19253);
xnor UO_1799 (O_1799,N_18818,N_19956);
and UO_1800 (O_1800,N_18070,N_18492);
and UO_1801 (O_1801,N_18516,N_19002);
and UO_1802 (O_1802,N_18240,N_18669);
and UO_1803 (O_1803,N_19302,N_19793);
nor UO_1804 (O_1804,N_18315,N_18734);
nor UO_1805 (O_1805,N_18504,N_18714);
or UO_1806 (O_1806,N_19916,N_18933);
xor UO_1807 (O_1807,N_18608,N_18736);
and UO_1808 (O_1808,N_18310,N_18245);
xnor UO_1809 (O_1809,N_19222,N_18623);
nor UO_1810 (O_1810,N_18434,N_18664);
or UO_1811 (O_1811,N_18398,N_19200);
or UO_1812 (O_1812,N_18324,N_19901);
nand UO_1813 (O_1813,N_19663,N_19172);
and UO_1814 (O_1814,N_19694,N_19702);
and UO_1815 (O_1815,N_19565,N_18815);
or UO_1816 (O_1816,N_18880,N_18479);
nand UO_1817 (O_1817,N_18950,N_19798);
nand UO_1818 (O_1818,N_19851,N_19943);
nand UO_1819 (O_1819,N_18797,N_18310);
nand UO_1820 (O_1820,N_19733,N_18322);
nand UO_1821 (O_1821,N_19201,N_19857);
and UO_1822 (O_1822,N_18102,N_18985);
or UO_1823 (O_1823,N_18718,N_18206);
and UO_1824 (O_1824,N_19710,N_19177);
and UO_1825 (O_1825,N_19798,N_19589);
and UO_1826 (O_1826,N_19842,N_19991);
and UO_1827 (O_1827,N_18936,N_19157);
and UO_1828 (O_1828,N_18487,N_18929);
and UO_1829 (O_1829,N_19612,N_19155);
xor UO_1830 (O_1830,N_19048,N_19594);
nand UO_1831 (O_1831,N_18037,N_19983);
or UO_1832 (O_1832,N_18831,N_19677);
nor UO_1833 (O_1833,N_18766,N_18770);
and UO_1834 (O_1834,N_19962,N_18708);
nand UO_1835 (O_1835,N_18030,N_18491);
nor UO_1836 (O_1836,N_18653,N_18232);
nand UO_1837 (O_1837,N_18573,N_19502);
nand UO_1838 (O_1838,N_19336,N_19016);
xnor UO_1839 (O_1839,N_19177,N_19670);
nand UO_1840 (O_1840,N_18158,N_19237);
nand UO_1841 (O_1841,N_18191,N_18373);
nor UO_1842 (O_1842,N_18528,N_19199);
and UO_1843 (O_1843,N_18845,N_19587);
nor UO_1844 (O_1844,N_19621,N_19108);
and UO_1845 (O_1845,N_19508,N_19302);
or UO_1846 (O_1846,N_19983,N_18488);
xnor UO_1847 (O_1847,N_18574,N_19130);
or UO_1848 (O_1848,N_19477,N_18287);
nor UO_1849 (O_1849,N_19042,N_18442);
xnor UO_1850 (O_1850,N_19677,N_19096);
and UO_1851 (O_1851,N_19204,N_18229);
nand UO_1852 (O_1852,N_19354,N_18346);
or UO_1853 (O_1853,N_18923,N_19029);
nor UO_1854 (O_1854,N_19253,N_19125);
nand UO_1855 (O_1855,N_18206,N_19649);
nor UO_1856 (O_1856,N_19951,N_19671);
nor UO_1857 (O_1857,N_19571,N_19357);
nand UO_1858 (O_1858,N_19987,N_19989);
nor UO_1859 (O_1859,N_18387,N_19684);
and UO_1860 (O_1860,N_18190,N_18846);
or UO_1861 (O_1861,N_19328,N_19708);
or UO_1862 (O_1862,N_18862,N_18231);
nor UO_1863 (O_1863,N_18541,N_18935);
nand UO_1864 (O_1864,N_19692,N_18482);
and UO_1865 (O_1865,N_19231,N_18931);
xor UO_1866 (O_1866,N_19718,N_18065);
xnor UO_1867 (O_1867,N_19333,N_18364);
nand UO_1868 (O_1868,N_18624,N_18092);
or UO_1869 (O_1869,N_19855,N_18494);
or UO_1870 (O_1870,N_19688,N_19103);
and UO_1871 (O_1871,N_19568,N_18936);
xnor UO_1872 (O_1872,N_18194,N_18458);
and UO_1873 (O_1873,N_18460,N_18498);
or UO_1874 (O_1874,N_19807,N_18459);
nand UO_1875 (O_1875,N_18674,N_19780);
nand UO_1876 (O_1876,N_19406,N_19895);
and UO_1877 (O_1877,N_19004,N_19605);
nor UO_1878 (O_1878,N_19896,N_19715);
nor UO_1879 (O_1879,N_18986,N_18111);
nor UO_1880 (O_1880,N_19892,N_18655);
nand UO_1881 (O_1881,N_19094,N_18040);
or UO_1882 (O_1882,N_18183,N_18085);
or UO_1883 (O_1883,N_18063,N_18986);
and UO_1884 (O_1884,N_18037,N_18712);
nand UO_1885 (O_1885,N_18995,N_18762);
or UO_1886 (O_1886,N_18410,N_19629);
or UO_1887 (O_1887,N_18490,N_19450);
or UO_1888 (O_1888,N_19674,N_19260);
and UO_1889 (O_1889,N_18968,N_18683);
or UO_1890 (O_1890,N_19329,N_18333);
and UO_1891 (O_1891,N_19009,N_18347);
nand UO_1892 (O_1892,N_18999,N_19566);
nand UO_1893 (O_1893,N_18327,N_18855);
nor UO_1894 (O_1894,N_19950,N_18052);
nand UO_1895 (O_1895,N_19673,N_18002);
and UO_1896 (O_1896,N_18948,N_18190);
or UO_1897 (O_1897,N_19562,N_19524);
or UO_1898 (O_1898,N_19151,N_18176);
nand UO_1899 (O_1899,N_18746,N_18958);
nand UO_1900 (O_1900,N_19081,N_18026);
nand UO_1901 (O_1901,N_19492,N_19691);
and UO_1902 (O_1902,N_19714,N_18309);
or UO_1903 (O_1903,N_18180,N_18226);
nand UO_1904 (O_1904,N_19669,N_19047);
or UO_1905 (O_1905,N_19337,N_19744);
nor UO_1906 (O_1906,N_18666,N_19512);
or UO_1907 (O_1907,N_19787,N_19071);
nor UO_1908 (O_1908,N_18392,N_18798);
nand UO_1909 (O_1909,N_19919,N_18407);
and UO_1910 (O_1910,N_19857,N_19037);
or UO_1911 (O_1911,N_18738,N_19872);
or UO_1912 (O_1912,N_18332,N_19963);
nand UO_1913 (O_1913,N_19789,N_18895);
nand UO_1914 (O_1914,N_18322,N_18731);
nor UO_1915 (O_1915,N_18029,N_19084);
and UO_1916 (O_1916,N_19874,N_19361);
nor UO_1917 (O_1917,N_18894,N_18861);
nor UO_1918 (O_1918,N_19201,N_19471);
nand UO_1919 (O_1919,N_19930,N_19052);
or UO_1920 (O_1920,N_18451,N_18760);
nand UO_1921 (O_1921,N_18228,N_19791);
nand UO_1922 (O_1922,N_18315,N_19505);
nor UO_1923 (O_1923,N_18112,N_19047);
nand UO_1924 (O_1924,N_19935,N_19566);
and UO_1925 (O_1925,N_18842,N_19249);
and UO_1926 (O_1926,N_18523,N_18740);
nand UO_1927 (O_1927,N_19807,N_19847);
or UO_1928 (O_1928,N_18114,N_18215);
and UO_1929 (O_1929,N_18352,N_18560);
and UO_1930 (O_1930,N_19681,N_19613);
and UO_1931 (O_1931,N_19654,N_18034);
and UO_1932 (O_1932,N_18249,N_19821);
nand UO_1933 (O_1933,N_18866,N_18793);
or UO_1934 (O_1934,N_18365,N_18502);
or UO_1935 (O_1935,N_18258,N_18257);
nand UO_1936 (O_1936,N_18293,N_18638);
nor UO_1937 (O_1937,N_19817,N_18500);
nand UO_1938 (O_1938,N_19511,N_19454);
and UO_1939 (O_1939,N_19188,N_18212);
nor UO_1940 (O_1940,N_18188,N_18278);
or UO_1941 (O_1941,N_18831,N_18790);
nor UO_1942 (O_1942,N_19024,N_19515);
xor UO_1943 (O_1943,N_19549,N_18190);
xor UO_1944 (O_1944,N_19701,N_19712);
or UO_1945 (O_1945,N_18789,N_18471);
nand UO_1946 (O_1946,N_19542,N_19249);
nor UO_1947 (O_1947,N_19636,N_19737);
and UO_1948 (O_1948,N_18343,N_19339);
nand UO_1949 (O_1949,N_19353,N_18328);
nor UO_1950 (O_1950,N_18012,N_19244);
xnor UO_1951 (O_1951,N_18192,N_18191);
and UO_1952 (O_1952,N_18412,N_18804);
nand UO_1953 (O_1953,N_19865,N_19547);
xor UO_1954 (O_1954,N_18347,N_19569);
nor UO_1955 (O_1955,N_19393,N_18903);
xor UO_1956 (O_1956,N_18576,N_19441);
and UO_1957 (O_1957,N_18808,N_19185);
and UO_1958 (O_1958,N_18028,N_19146);
nor UO_1959 (O_1959,N_18857,N_18202);
or UO_1960 (O_1960,N_18746,N_18599);
nand UO_1961 (O_1961,N_18012,N_19193);
nor UO_1962 (O_1962,N_18939,N_18717);
or UO_1963 (O_1963,N_19937,N_18216);
and UO_1964 (O_1964,N_18002,N_19081);
nor UO_1965 (O_1965,N_19067,N_18972);
or UO_1966 (O_1966,N_18359,N_19464);
nand UO_1967 (O_1967,N_19503,N_19790);
and UO_1968 (O_1968,N_19122,N_19500);
or UO_1969 (O_1969,N_19429,N_18107);
xnor UO_1970 (O_1970,N_19150,N_19535);
or UO_1971 (O_1971,N_19401,N_19258);
or UO_1972 (O_1972,N_18841,N_19591);
nor UO_1973 (O_1973,N_19321,N_19950);
nor UO_1974 (O_1974,N_19167,N_18417);
nand UO_1975 (O_1975,N_19932,N_19511);
nor UO_1976 (O_1976,N_18537,N_19303);
and UO_1977 (O_1977,N_19615,N_18478);
nor UO_1978 (O_1978,N_18962,N_19090);
or UO_1979 (O_1979,N_18871,N_18689);
nand UO_1980 (O_1980,N_19401,N_18542);
nor UO_1981 (O_1981,N_18313,N_18550);
nor UO_1982 (O_1982,N_18314,N_19092);
nand UO_1983 (O_1983,N_19090,N_19230);
or UO_1984 (O_1984,N_18086,N_18289);
and UO_1985 (O_1985,N_19361,N_18540);
nand UO_1986 (O_1986,N_18347,N_18214);
nand UO_1987 (O_1987,N_19605,N_19593);
xnor UO_1988 (O_1988,N_19910,N_18832);
or UO_1989 (O_1989,N_19878,N_18765);
nand UO_1990 (O_1990,N_19911,N_18662);
or UO_1991 (O_1991,N_19589,N_19727);
and UO_1992 (O_1992,N_18462,N_19794);
nand UO_1993 (O_1993,N_18219,N_18857);
nand UO_1994 (O_1994,N_19196,N_19139);
or UO_1995 (O_1995,N_18270,N_18630);
or UO_1996 (O_1996,N_18871,N_19963);
or UO_1997 (O_1997,N_18277,N_18488);
nand UO_1998 (O_1998,N_18928,N_18378);
nand UO_1999 (O_1999,N_19549,N_19622);
and UO_2000 (O_2000,N_18919,N_18983);
nor UO_2001 (O_2001,N_19600,N_18831);
and UO_2002 (O_2002,N_19497,N_18658);
nand UO_2003 (O_2003,N_19909,N_18114);
nor UO_2004 (O_2004,N_19134,N_19679);
nand UO_2005 (O_2005,N_18479,N_19320);
and UO_2006 (O_2006,N_19096,N_19455);
nor UO_2007 (O_2007,N_18487,N_19495);
nor UO_2008 (O_2008,N_19025,N_18910);
nor UO_2009 (O_2009,N_18907,N_19578);
xnor UO_2010 (O_2010,N_18790,N_19360);
or UO_2011 (O_2011,N_18212,N_18875);
nor UO_2012 (O_2012,N_19846,N_18015);
or UO_2013 (O_2013,N_18014,N_18713);
nor UO_2014 (O_2014,N_19819,N_18112);
nor UO_2015 (O_2015,N_18069,N_19779);
or UO_2016 (O_2016,N_19747,N_18473);
and UO_2017 (O_2017,N_18615,N_19798);
and UO_2018 (O_2018,N_18809,N_18633);
nor UO_2019 (O_2019,N_19125,N_19224);
nor UO_2020 (O_2020,N_18511,N_18219);
and UO_2021 (O_2021,N_18080,N_18777);
nand UO_2022 (O_2022,N_19527,N_19216);
nor UO_2023 (O_2023,N_18687,N_18401);
nand UO_2024 (O_2024,N_18276,N_19789);
nor UO_2025 (O_2025,N_19008,N_19855);
and UO_2026 (O_2026,N_18852,N_19379);
and UO_2027 (O_2027,N_19292,N_19882);
or UO_2028 (O_2028,N_19206,N_18393);
nand UO_2029 (O_2029,N_19004,N_19887);
nand UO_2030 (O_2030,N_18168,N_19623);
nand UO_2031 (O_2031,N_18041,N_19614);
or UO_2032 (O_2032,N_19378,N_18490);
or UO_2033 (O_2033,N_18966,N_18752);
nor UO_2034 (O_2034,N_18155,N_18272);
and UO_2035 (O_2035,N_18318,N_18194);
xnor UO_2036 (O_2036,N_18999,N_19558);
and UO_2037 (O_2037,N_19206,N_19340);
or UO_2038 (O_2038,N_18978,N_18499);
nor UO_2039 (O_2039,N_18925,N_18551);
nand UO_2040 (O_2040,N_18795,N_18817);
xor UO_2041 (O_2041,N_19569,N_18661);
and UO_2042 (O_2042,N_18454,N_18823);
or UO_2043 (O_2043,N_19407,N_19037);
or UO_2044 (O_2044,N_19530,N_19852);
nand UO_2045 (O_2045,N_19598,N_18551);
nor UO_2046 (O_2046,N_18244,N_19823);
nor UO_2047 (O_2047,N_19026,N_19655);
nand UO_2048 (O_2048,N_18885,N_19596);
and UO_2049 (O_2049,N_19109,N_19445);
or UO_2050 (O_2050,N_19744,N_19099);
or UO_2051 (O_2051,N_18741,N_19347);
nand UO_2052 (O_2052,N_19174,N_18364);
nor UO_2053 (O_2053,N_19943,N_18331);
nor UO_2054 (O_2054,N_18168,N_18821);
or UO_2055 (O_2055,N_19562,N_18706);
and UO_2056 (O_2056,N_19484,N_19793);
and UO_2057 (O_2057,N_19435,N_18378);
nand UO_2058 (O_2058,N_19789,N_19949);
nand UO_2059 (O_2059,N_18889,N_19152);
nor UO_2060 (O_2060,N_19501,N_18725);
and UO_2061 (O_2061,N_18635,N_18627);
nor UO_2062 (O_2062,N_18041,N_19209);
xnor UO_2063 (O_2063,N_19363,N_18463);
nand UO_2064 (O_2064,N_19930,N_19410);
nand UO_2065 (O_2065,N_18787,N_19226);
and UO_2066 (O_2066,N_18618,N_19737);
or UO_2067 (O_2067,N_19909,N_18989);
nor UO_2068 (O_2068,N_19091,N_18711);
or UO_2069 (O_2069,N_18419,N_18692);
nor UO_2070 (O_2070,N_18494,N_18841);
nand UO_2071 (O_2071,N_19370,N_18457);
nor UO_2072 (O_2072,N_19354,N_18904);
nor UO_2073 (O_2073,N_19945,N_18911);
xor UO_2074 (O_2074,N_18404,N_18079);
or UO_2075 (O_2075,N_18140,N_19186);
and UO_2076 (O_2076,N_19062,N_19073);
or UO_2077 (O_2077,N_18191,N_18620);
and UO_2078 (O_2078,N_19456,N_18139);
or UO_2079 (O_2079,N_19743,N_19217);
nor UO_2080 (O_2080,N_18868,N_19157);
nor UO_2081 (O_2081,N_18968,N_19145);
or UO_2082 (O_2082,N_19366,N_19251);
or UO_2083 (O_2083,N_18212,N_19382);
nor UO_2084 (O_2084,N_19712,N_18018);
nand UO_2085 (O_2085,N_19186,N_19230);
and UO_2086 (O_2086,N_18054,N_19508);
nor UO_2087 (O_2087,N_19075,N_18188);
nand UO_2088 (O_2088,N_19063,N_19547);
nor UO_2089 (O_2089,N_19426,N_18493);
nor UO_2090 (O_2090,N_19045,N_18931);
nor UO_2091 (O_2091,N_19766,N_19106);
nor UO_2092 (O_2092,N_19095,N_19210);
and UO_2093 (O_2093,N_19252,N_19669);
and UO_2094 (O_2094,N_19630,N_19963);
and UO_2095 (O_2095,N_19073,N_18865);
nand UO_2096 (O_2096,N_18861,N_18588);
and UO_2097 (O_2097,N_18476,N_18197);
nor UO_2098 (O_2098,N_18333,N_19416);
nor UO_2099 (O_2099,N_18589,N_18117);
or UO_2100 (O_2100,N_18566,N_19560);
nor UO_2101 (O_2101,N_18153,N_19578);
and UO_2102 (O_2102,N_18730,N_18275);
and UO_2103 (O_2103,N_19666,N_18747);
nor UO_2104 (O_2104,N_18173,N_19859);
nor UO_2105 (O_2105,N_19441,N_18000);
or UO_2106 (O_2106,N_19403,N_18820);
or UO_2107 (O_2107,N_19016,N_18136);
nand UO_2108 (O_2108,N_18545,N_18108);
and UO_2109 (O_2109,N_18258,N_18848);
nand UO_2110 (O_2110,N_18162,N_19191);
and UO_2111 (O_2111,N_18213,N_18577);
and UO_2112 (O_2112,N_18742,N_18192);
nand UO_2113 (O_2113,N_19949,N_19682);
nor UO_2114 (O_2114,N_18242,N_19451);
nand UO_2115 (O_2115,N_19563,N_19159);
nor UO_2116 (O_2116,N_19755,N_18974);
and UO_2117 (O_2117,N_19277,N_19694);
or UO_2118 (O_2118,N_18351,N_18788);
nor UO_2119 (O_2119,N_18490,N_19312);
nand UO_2120 (O_2120,N_19123,N_18378);
and UO_2121 (O_2121,N_19173,N_19123);
nand UO_2122 (O_2122,N_18084,N_18911);
xor UO_2123 (O_2123,N_19660,N_19026);
or UO_2124 (O_2124,N_18332,N_19768);
xnor UO_2125 (O_2125,N_18769,N_19226);
nand UO_2126 (O_2126,N_19277,N_18765);
nor UO_2127 (O_2127,N_18779,N_19292);
nand UO_2128 (O_2128,N_18734,N_18739);
nand UO_2129 (O_2129,N_19797,N_19164);
nor UO_2130 (O_2130,N_18388,N_19083);
xnor UO_2131 (O_2131,N_18026,N_18091);
nand UO_2132 (O_2132,N_18733,N_19894);
nor UO_2133 (O_2133,N_19991,N_19456);
and UO_2134 (O_2134,N_19043,N_19608);
and UO_2135 (O_2135,N_18076,N_18861);
nand UO_2136 (O_2136,N_18433,N_18350);
and UO_2137 (O_2137,N_18777,N_18308);
xnor UO_2138 (O_2138,N_18849,N_19239);
and UO_2139 (O_2139,N_18725,N_19200);
nand UO_2140 (O_2140,N_18893,N_19611);
and UO_2141 (O_2141,N_18959,N_19444);
or UO_2142 (O_2142,N_18998,N_19156);
or UO_2143 (O_2143,N_18848,N_19448);
nor UO_2144 (O_2144,N_18830,N_19206);
nand UO_2145 (O_2145,N_19909,N_19317);
nand UO_2146 (O_2146,N_19782,N_18714);
and UO_2147 (O_2147,N_18603,N_18483);
nand UO_2148 (O_2148,N_18969,N_18242);
nand UO_2149 (O_2149,N_18828,N_18181);
or UO_2150 (O_2150,N_19705,N_18645);
xnor UO_2151 (O_2151,N_18544,N_19329);
xor UO_2152 (O_2152,N_18938,N_18770);
and UO_2153 (O_2153,N_19061,N_19165);
and UO_2154 (O_2154,N_19962,N_18983);
or UO_2155 (O_2155,N_19949,N_19121);
or UO_2156 (O_2156,N_18748,N_18848);
or UO_2157 (O_2157,N_18194,N_19234);
nand UO_2158 (O_2158,N_18105,N_19858);
or UO_2159 (O_2159,N_18318,N_18357);
nand UO_2160 (O_2160,N_19390,N_18162);
nand UO_2161 (O_2161,N_19508,N_18769);
and UO_2162 (O_2162,N_19403,N_18480);
nand UO_2163 (O_2163,N_19778,N_19636);
nand UO_2164 (O_2164,N_18934,N_19638);
nand UO_2165 (O_2165,N_19725,N_19037);
or UO_2166 (O_2166,N_19426,N_18182);
xor UO_2167 (O_2167,N_18934,N_19615);
and UO_2168 (O_2168,N_19669,N_19437);
nor UO_2169 (O_2169,N_19302,N_18916);
and UO_2170 (O_2170,N_18273,N_19339);
and UO_2171 (O_2171,N_19170,N_19119);
nand UO_2172 (O_2172,N_18019,N_19046);
nor UO_2173 (O_2173,N_19673,N_19602);
nor UO_2174 (O_2174,N_18179,N_18122);
nand UO_2175 (O_2175,N_19329,N_18786);
or UO_2176 (O_2176,N_19724,N_18205);
nor UO_2177 (O_2177,N_18424,N_19804);
nand UO_2178 (O_2178,N_19188,N_18692);
nand UO_2179 (O_2179,N_18164,N_18136);
and UO_2180 (O_2180,N_19186,N_18663);
or UO_2181 (O_2181,N_19444,N_18763);
nand UO_2182 (O_2182,N_19053,N_19732);
xor UO_2183 (O_2183,N_18861,N_18321);
nand UO_2184 (O_2184,N_18703,N_18179);
or UO_2185 (O_2185,N_18292,N_19515);
or UO_2186 (O_2186,N_18623,N_18610);
nand UO_2187 (O_2187,N_19018,N_19289);
nor UO_2188 (O_2188,N_19123,N_19448);
nand UO_2189 (O_2189,N_19705,N_18793);
xnor UO_2190 (O_2190,N_18791,N_18704);
and UO_2191 (O_2191,N_18562,N_18768);
nor UO_2192 (O_2192,N_18183,N_19510);
nor UO_2193 (O_2193,N_19714,N_18994);
and UO_2194 (O_2194,N_19373,N_18198);
or UO_2195 (O_2195,N_18103,N_18607);
xnor UO_2196 (O_2196,N_19257,N_19976);
nor UO_2197 (O_2197,N_18615,N_19117);
nor UO_2198 (O_2198,N_19789,N_19937);
nor UO_2199 (O_2199,N_18817,N_19392);
or UO_2200 (O_2200,N_18488,N_18502);
or UO_2201 (O_2201,N_19337,N_19406);
nand UO_2202 (O_2202,N_19698,N_18863);
nand UO_2203 (O_2203,N_18760,N_18532);
or UO_2204 (O_2204,N_19925,N_18989);
xor UO_2205 (O_2205,N_18993,N_19018);
or UO_2206 (O_2206,N_19340,N_19085);
xnor UO_2207 (O_2207,N_18358,N_18039);
and UO_2208 (O_2208,N_19733,N_18711);
and UO_2209 (O_2209,N_19062,N_18733);
nand UO_2210 (O_2210,N_19180,N_18328);
nor UO_2211 (O_2211,N_19298,N_19871);
nor UO_2212 (O_2212,N_18914,N_18071);
nand UO_2213 (O_2213,N_18918,N_18376);
nand UO_2214 (O_2214,N_18479,N_19355);
or UO_2215 (O_2215,N_19076,N_18670);
nor UO_2216 (O_2216,N_19797,N_19214);
and UO_2217 (O_2217,N_18061,N_19557);
and UO_2218 (O_2218,N_18173,N_18601);
and UO_2219 (O_2219,N_19200,N_19821);
nor UO_2220 (O_2220,N_19090,N_19528);
or UO_2221 (O_2221,N_19568,N_18143);
or UO_2222 (O_2222,N_18680,N_18333);
or UO_2223 (O_2223,N_19493,N_19412);
nand UO_2224 (O_2224,N_19331,N_18214);
or UO_2225 (O_2225,N_19932,N_18489);
nor UO_2226 (O_2226,N_18557,N_18256);
and UO_2227 (O_2227,N_19045,N_19371);
xor UO_2228 (O_2228,N_18519,N_19319);
nor UO_2229 (O_2229,N_18408,N_19006);
xor UO_2230 (O_2230,N_19569,N_18399);
xnor UO_2231 (O_2231,N_19145,N_19569);
or UO_2232 (O_2232,N_19140,N_18453);
xor UO_2233 (O_2233,N_19397,N_18127);
nor UO_2234 (O_2234,N_18772,N_18560);
nand UO_2235 (O_2235,N_18677,N_19157);
and UO_2236 (O_2236,N_18258,N_19480);
or UO_2237 (O_2237,N_18343,N_19765);
xnor UO_2238 (O_2238,N_19745,N_18129);
nand UO_2239 (O_2239,N_19895,N_18856);
nand UO_2240 (O_2240,N_19013,N_19628);
xor UO_2241 (O_2241,N_18463,N_19161);
and UO_2242 (O_2242,N_19659,N_18309);
nand UO_2243 (O_2243,N_19004,N_18926);
or UO_2244 (O_2244,N_18873,N_18158);
and UO_2245 (O_2245,N_19972,N_19761);
and UO_2246 (O_2246,N_19708,N_18066);
nor UO_2247 (O_2247,N_18047,N_18699);
nor UO_2248 (O_2248,N_18997,N_19338);
nand UO_2249 (O_2249,N_18273,N_18912);
nor UO_2250 (O_2250,N_19237,N_19163);
or UO_2251 (O_2251,N_19063,N_19820);
nand UO_2252 (O_2252,N_18706,N_19716);
or UO_2253 (O_2253,N_18370,N_19127);
nand UO_2254 (O_2254,N_19609,N_19762);
or UO_2255 (O_2255,N_18013,N_19966);
or UO_2256 (O_2256,N_19288,N_18025);
nand UO_2257 (O_2257,N_19713,N_19990);
nand UO_2258 (O_2258,N_19331,N_18322);
nor UO_2259 (O_2259,N_19138,N_18973);
nor UO_2260 (O_2260,N_19241,N_18066);
or UO_2261 (O_2261,N_19413,N_19071);
or UO_2262 (O_2262,N_18970,N_19616);
and UO_2263 (O_2263,N_19044,N_18644);
or UO_2264 (O_2264,N_18523,N_19887);
or UO_2265 (O_2265,N_18606,N_19365);
and UO_2266 (O_2266,N_18507,N_19532);
and UO_2267 (O_2267,N_19820,N_19221);
nand UO_2268 (O_2268,N_19113,N_19339);
nand UO_2269 (O_2269,N_19952,N_18440);
nand UO_2270 (O_2270,N_18879,N_18571);
or UO_2271 (O_2271,N_18349,N_19752);
xnor UO_2272 (O_2272,N_18346,N_19677);
nand UO_2273 (O_2273,N_19824,N_19722);
nor UO_2274 (O_2274,N_19119,N_19307);
nor UO_2275 (O_2275,N_19575,N_18011);
or UO_2276 (O_2276,N_18552,N_19598);
nand UO_2277 (O_2277,N_18069,N_18098);
and UO_2278 (O_2278,N_19256,N_18032);
and UO_2279 (O_2279,N_18888,N_19227);
nand UO_2280 (O_2280,N_19666,N_19639);
nor UO_2281 (O_2281,N_19151,N_18636);
and UO_2282 (O_2282,N_19415,N_19480);
nand UO_2283 (O_2283,N_18826,N_19534);
or UO_2284 (O_2284,N_19686,N_19361);
and UO_2285 (O_2285,N_19357,N_18659);
and UO_2286 (O_2286,N_19060,N_19066);
nor UO_2287 (O_2287,N_19160,N_19934);
or UO_2288 (O_2288,N_19894,N_18083);
or UO_2289 (O_2289,N_18417,N_19351);
nand UO_2290 (O_2290,N_19381,N_18558);
nand UO_2291 (O_2291,N_19419,N_19869);
or UO_2292 (O_2292,N_19393,N_19757);
or UO_2293 (O_2293,N_19509,N_18583);
or UO_2294 (O_2294,N_19773,N_18776);
and UO_2295 (O_2295,N_18066,N_18980);
nor UO_2296 (O_2296,N_19593,N_18917);
and UO_2297 (O_2297,N_19136,N_18012);
xor UO_2298 (O_2298,N_19490,N_19691);
xor UO_2299 (O_2299,N_18641,N_19654);
xor UO_2300 (O_2300,N_18876,N_19214);
nand UO_2301 (O_2301,N_19828,N_18610);
or UO_2302 (O_2302,N_18957,N_18052);
nor UO_2303 (O_2303,N_18412,N_18280);
nand UO_2304 (O_2304,N_19645,N_18351);
and UO_2305 (O_2305,N_18419,N_19984);
xor UO_2306 (O_2306,N_19435,N_19334);
or UO_2307 (O_2307,N_18333,N_18898);
and UO_2308 (O_2308,N_19491,N_19908);
and UO_2309 (O_2309,N_19775,N_18769);
nor UO_2310 (O_2310,N_18908,N_19540);
nor UO_2311 (O_2311,N_18888,N_18413);
and UO_2312 (O_2312,N_18070,N_19985);
nand UO_2313 (O_2313,N_18289,N_19044);
xnor UO_2314 (O_2314,N_19775,N_19864);
or UO_2315 (O_2315,N_18125,N_18212);
or UO_2316 (O_2316,N_19954,N_18144);
or UO_2317 (O_2317,N_18481,N_18757);
nand UO_2318 (O_2318,N_19139,N_19931);
nor UO_2319 (O_2319,N_18412,N_18127);
nand UO_2320 (O_2320,N_19327,N_19824);
xnor UO_2321 (O_2321,N_19051,N_18670);
and UO_2322 (O_2322,N_18969,N_19690);
and UO_2323 (O_2323,N_18016,N_18451);
xor UO_2324 (O_2324,N_18146,N_18516);
or UO_2325 (O_2325,N_18597,N_18428);
and UO_2326 (O_2326,N_18843,N_18083);
and UO_2327 (O_2327,N_19763,N_18619);
or UO_2328 (O_2328,N_18572,N_19714);
nand UO_2329 (O_2329,N_18716,N_19632);
nand UO_2330 (O_2330,N_19701,N_19674);
or UO_2331 (O_2331,N_19529,N_19549);
xnor UO_2332 (O_2332,N_18240,N_18437);
or UO_2333 (O_2333,N_19160,N_18055);
or UO_2334 (O_2334,N_19684,N_19939);
and UO_2335 (O_2335,N_19918,N_19015);
nor UO_2336 (O_2336,N_19872,N_18574);
and UO_2337 (O_2337,N_19559,N_18765);
and UO_2338 (O_2338,N_18468,N_18032);
nand UO_2339 (O_2339,N_19106,N_19994);
or UO_2340 (O_2340,N_18200,N_18226);
nor UO_2341 (O_2341,N_19192,N_18367);
or UO_2342 (O_2342,N_18413,N_18570);
xor UO_2343 (O_2343,N_18369,N_18373);
and UO_2344 (O_2344,N_19886,N_18287);
or UO_2345 (O_2345,N_19591,N_19128);
or UO_2346 (O_2346,N_18184,N_18832);
nand UO_2347 (O_2347,N_18837,N_19177);
nand UO_2348 (O_2348,N_18791,N_19293);
nand UO_2349 (O_2349,N_18955,N_18169);
and UO_2350 (O_2350,N_18864,N_18450);
and UO_2351 (O_2351,N_19307,N_18758);
xnor UO_2352 (O_2352,N_19455,N_18004);
or UO_2353 (O_2353,N_19448,N_19738);
nand UO_2354 (O_2354,N_18658,N_19200);
nor UO_2355 (O_2355,N_18864,N_19825);
or UO_2356 (O_2356,N_18182,N_19338);
nor UO_2357 (O_2357,N_18996,N_18313);
nand UO_2358 (O_2358,N_19960,N_19779);
nor UO_2359 (O_2359,N_18927,N_19371);
or UO_2360 (O_2360,N_18942,N_18715);
xor UO_2361 (O_2361,N_19808,N_18606);
or UO_2362 (O_2362,N_19447,N_19841);
nor UO_2363 (O_2363,N_18009,N_18725);
nand UO_2364 (O_2364,N_18192,N_18165);
and UO_2365 (O_2365,N_18645,N_19815);
nor UO_2366 (O_2366,N_19602,N_18040);
or UO_2367 (O_2367,N_19590,N_19847);
and UO_2368 (O_2368,N_19274,N_18889);
nand UO_2369 (O_2369,N_19820,N_19666);
nor UO_2370 (O_2370,N_18570,N_19484);
or UO_2371 (O_2371,N_19751,N_18014);
nor UO_2372 (O_2372,N_18332,N_18007);
nand UO_2373 (O_2373,N_19442,N_18317);
nand UO_2374 (O_2374,N_19899,N_18576);
nor UO_2375 (O_2375,N_18822,N_19270);
or UO_2376 (O_2376,N_19567,N_18143);
or UO_2377 (O_2377,N_19680,N_18025);
nand UO_2378 (O_2378,N_19526,N_19036);
and UO_2379 (O_2379,N_18482,N_19751);
and UO_2380 (O_2380,N_19535,N_19635);
or UO_2381 (O_2381,N_19537,N_19723);
and UO_2382 (O_2382,N_18556,N_18837);
nor UO_2383 (O_2383,N_19482,N_19880);
or UO_2384 (O_2384,N_19989,N_19008);
nor UO_2385 (O_2385,N_19691,N_19890);
nand UO_2386 (O_2386,N_18093,N_18059);
and UO_2387 (O_2387,N_19511,N_18590);
xnor UO_2388 (O_2388,N_18833,N_19491);
nor UO_2389 (O_2389,N_18437,N_18424);
xnor UO_2390 (O_2390,N_18086,N_18303);
nand UO_2391 (O_2391,N_19468,N_18459);
nor UO_2392 (O_2392,N_18306,N_18346);
and UO_2393 (O_2393,N_19137,N_18755);
xnor UO_2394 (O_2394,N_18750,N_18936);
and UO_2395 (O_2395,N_19118,N_19124);
nand UO_2396 (O_2396,N_18066,N_18448);
nand UO_2397 (O_2397,N_18023,N_19651);
nand UO_2398 (O_2398,N_19524,N_19546);
and UO_2399 (O_2399,N_19954,N_19289);
xnor UO_2400 (O_2400,N_19354,N_18767);
nor UO_2401 (O_2401,N_19796,N_18794);
xor UO_2402 (O_2402,N_18156,N_18165);
and UO_2403 (O_2403,N_18118,N_19294);
nand UO_2404 (O_2404,N_19516,N_19995);
and UO_2405 (O_2405,N_19111,N_19502);
or UO_2406 (O_2406,N_18412,N_19461);
nor UO_2407 (O_2407,N_19416,N_18321);
and UO_2408 (O_2408,N_19627,N_18974);
nand UO_2409 (O_2409,N_19013,N_19531);
nand UO_2410 (O_2410,N_19670,N_19183);
or UO_2411 (O_2411,N_19996,N_18836);
nor UO_2412 (O_2412,N_18777,N_19665);
or UO_2413 (O_2413,N_18776,N_19884);
or UO_2414 (O_2414,N_19188,N_18548);
or UO_2415 (O_2415,N_18200,N_19632);
and UO_2416 (O_2416,N_18773,N_18452);
and UO_2417 (O_2417,N_19664,N_18379);
nand UO_2418 (O_2418,N_19143,N_19647);
and UO_2419 (O_2419,N_19385,N_19957);
and UO_2420 (O_2420,N_18789,N_18402);
and UO_2421 (O_2421,N_19749,N_19032);
or UO_2422 (O_2422,N_18140,N_18678);
nor UO_2423 (O_2423,N_18977,N_18760);
nor UO_2424 (O_2424,N_19204,N_18191);
or UO_2425 (O_2425,N_18968,N_19818);
nand UO_2426 (O_2426,N_18414,N_18301);
nor UO_2427 (O_2427,N_18122,N_19865);
nand UO_2428 (O_2428,N_18692,N_19561);
or UO_2429 (O_2429,N_18253,N_18520);
or UO_2430 (O_2430,N_19171,N_18973);
nor UO_2431 (O_2431,N_19691,N_18104);
and UO_2432 (O_2432,N_19338,N_18019);
and UO_2433 (O_2433,N_19953,N_19034);
nor UO_2434 (O_2434,N_19633,N_19016);
or UO_2435 (O_2435,N_18086,N_19586);
nand UO_2436 (O_2436,N_18190,N_19984);
and UO_2437 (O_2437,N_19901,N_19073);
nor UO_2438 (O_2438,N_19175,N_18821);
nor UO_2439 (O_2439,N_19607,N_19219);
and UO_2440 (O_2440,N_19590,N_18991);
xor UO_2441 (O_2441,N_18424,N_19801);
nor UO_2442 (O_2442,N_19921,N_19659);
and UO_2443 (O_2443,N_19761,N_18488);
or UO_2444 (O_2444,N_18330,N_19850);
nand UO_2445 (O_2445,N_18858,N_18705);
and UO_2446 (O_2446,N_18932,N_19881);
nand UO_2447 (O_2447,N_19991,N_18222);
or UO_2448 (O_2448,N_18275,N_19809);
and UO_2449 (O_2449,N_19990,N_18187);
or UO_2450 (O_2450,N_18598,N_18023);
nand UO_2451 (O_2451,N_19022,N_18677);
nor UO_2452 (O_2452,N_18346,N_18547);
and UO_2453 (O_2453,N_19856,N_19368);
nand UO_2454 (O_2454,N_18991,N_19473);
and UO_2455 (O_2455,N_19888,N_18213);
nand UO_2456 (O_2456,N_19780,N_18977);
and UO_2457 (O_2457,N_18494,N_19588);
nor UO_2458 (O_2458,N_19414,N_19808);
nor UO_2459 (O_2459,N_19415,N_18573);
or UO_2460 (O_2460,N_19399,N_18144);
nor UO_2461 (O_2461,N_18055,N_19643);
nor UO_2462 (O_2462,N_19463,N_19760);
nor UO_2463 (O_2463,N_19782,N_19887);
nor UO_2464 (O_2464,N_18284,N_18236);
or UO_2465 (O_2465,N_18108,N_18117);
nor UO_2466 (O_2466,N_19284,N_18261);
or UO_2467 (O_2467,N_18441,N_18975);
and UO_2468 (O_2468,N_19981,N_18064);
nor UO_2469 (O_2469,N_18491,N_19128);
nor UO_2470 (O_2470,N_19499,N_18220);
nand UO_2471 (O_2471,N_19997,N_19117);
or UO_2472 (O_2472,N_19424,N_19091);
nor UO_2473 (O_2473,N_19431,N_19428);
xor UO_2474 (O_2474,N_19778,N_18825);
nor UO_2475 (O_2475,N_19640,N_19922);
xor UO_2476 (O_2476,N_19906,N_19699);
and UO_2477 (O_2477,N_18784,N_18441);
nor UO_2478 (O_2478,N_19247,N_18854);
or UO_2479 (O_2479,N_19965,N_18278);
and UO_2480 (O_2480,N_19490,N_19004);
nand UO_2481 (O_2481,N_19061,N_19045);
nand UO_2482 (O_2482,N_18003,N_19930);
xor UO_2483 (O_2483,N_19496,N_18322);
nor UO_2484 (O_2484,N_19922,N_18717);
nor UO_2485 (O_2485,N_18846,N_19582);
nor UO_2486 (O_2486,N_19524,N_19367);
nor UO_2487 (O_2487,N_18716,N_19687);
nand UO_2488 (O_2488,N_18620,N_18129);
nand UO_2489 (O_2489,N_18386,N_18771);
or UO_2490 (O_2490,N_18044,N_19891);
nor UO_2491 (O_2491,N_19791,N_19165);
xnor UO_2492 (O_2492,N_18820,N_18427);
or UO_2493 (O_2493,N_18283,N_19084);
and UO_2494 (O_2494,N_18460,N_19850);
or UO_2495 (O_2495,N_18431,N_18842);
nand UO_2496 (O_2496,N_18300,N_19705);
or UO_2497 (O_2497,N_19488,N_18116);
or UO_2498 (O_2498,N_18051,N_18981);
nand UO_2499 (O_2499,N_18663,N_18364);
endmodule