module basic_500_3000_500_50_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_484,In_492);
nand U1 (N_1,In_25,In_289);
and U2 (N_2,In_78,In_325);
nand U3 (N_3,In_20,In_442);
nand U4 (N_4,In_114,In_276);
and U5 (N_5,In_39,In_118);
nor U6 (N_6,In_439,In_188);
nor U7 (N_7,In_416,In_191);
or U8 (N_8,In_221,In_213);
nor U9 (N_9,In_125,In_391);
or U10 (N_10,In_23,In_8);
and U11 (N_11,In_367,In_7);
or U12 (N_12,In_79,In_243);
and U13 (N_13,In_219,In_486);
nand U14 (N_14,In_313,In_324);
nor U15 (N_15,In_207,In_88);
nor U16 (N_16,In_393,In_175);
and U17 (N_17,In_444,In_346);
or U18 (N_18,In_69,In_285);
nand U19 (N_19,In_269,In_495);
nand U20 (N_20,In_326,In_310);
and U21 (N_21,In_38,In_198);
nand U22 (N_22,In_372,In_132);
nand U23 (N_23,In_124,In_447);
nor U24 (N_24,In_499,In_111);
or U25 (N_25,In_57,In_344);
or U26 (N_26,In_151,In_275);
and U27 (N_27,In_477,In_52);
or U28 (N_28,In_71,In_46);
nand U29 (N_29,In_109,In_152);
nor U30 (N_30,In_44,In_299);
nor U31 (N_31,In_86,In_343);
nor U32 (N_32,In_51,In_73);
or U33 (N_33,In_266,In_457);
nor U34 (N_34,In_264,In_288);
or U35 (N_35,In_305,In_169);
and U36 (N_36,In_433,In_473);
or U37 (N_37,In_21,In_374);
nor U38 (N_38,In_131,In_291);
nand U39 (N_39,In_446,In_412);
and U40 (N_40,In_156,In_292);
and U41 (N_41,In_101,In_407);
nor U42 (N_42,In_234,In_206);
or U43 (N_43,In_197,In_115);
or U44 (N_44,In_431,In_176);
or U45 (N_45,In_259,In_373);
or U46 (N_46,In_201,In_348);
and U47 (N_47,In_455,In_239);
nor U48 (N_48,In_36,In_123);
nand U49 (N_49,In_2,In_163);
nand U50 (N_50,In_49,In_443);
nand U51 (N_51,In_187,In_145);
nor U52 (N_52,In_483,In_434);
nor U53 (N_53,In_278,In_66);
nand U54 (N_54,In_214,In_405);
or U55 (N_55,In_54,In_141);
nand U56 (N_56,In_360,In_312);
and U57 (N_57,In_50,In_254);
and U58 (N_58,In_361,In_193);
nor U59 (N_59,In_463,In_487);
nor U60 (N_60,In_130,In_415);
nand U61 (N_61,In_68,In_230);
and U62 (N_62,In_350,In_318);
or U63 (N_63,In_236,In_242);
or U64 (N_64,In_280,In_353);
nor U65 (N_65,In_317,N_57);
or U66 (N_66,In_398,In_268);
or U67 (N_67,In_355,In_249);
xnor U68 (N_68,In_413,N_30);
nor U69 (N_69,In_128,In_428);
nor U70 (N_70,In_388,In_41);
xor U71 (N_71,In_231,In_253);
or U72 (N_72,In_26,In_330);
nand U73 (N_73,In_263,In_127);
and U74 (N_74,In_6,In_246);
nand U75 (N_75,In_250,In_306);
nand U76 (N_76,In_351,In_94);
and U77 (N_77,In_30,In_45);
and U78 (N_78,N_41,In_470);
and U79 (N_79,In_186,N_45);
or U80 (N_80,In_209,In_224);
or U81 (N_81,In_14,In_283);
and U82 (N_82,In_76,In_314);
nor U83 (N_83,In_89,In_233);
nand U84 (N_84,N_51,In_339);
or U85 (N_85,In_174,In_498);
nand U86 (N_86,In_142,In_418);
and U87 (N_87,N_1,In_400);
or U88 (N_88,N_11,In_19);
nand U89 (N_89,In_84,In_401);
nor U90 (N_90,In_437,In_110);
or U91 (N_91,In_358,In_223);
nor U92 (N_92,In_274,In_432);
xor U93 (N_93,N_49,In_311);
xnor U94 (N_94,In_345,In_265);
and U95 (N_95,N_22,N_50);
nor U96 (N_96,In_35,In_448);
nor U97 (N_97,In_425,In_55);
xor U98 (N_98,In_341,In_245);
or U99 (N_99,In_474,In_328);
xnor U100 (N_100,N_58,In_116);
and U101 (N_101,In_33,N_14);
nor U102 (N_102,In_177,In_155);
nor U103 (N_103,N_35,In_436);
nor U104 (N_104,N_2,In_380);
nor U105 (N_105,In_347,In_298);
and U106 (N_106,In_248,In_64);
nor U107 (N_107,In_414,In_327);
and U108 (N_108,In_423,In_261);
nand U109 (N_109,In_281,In_365);
or U110 (N_110,In_173,N_56);
nor U111 (N_111,In_424,In_464);
nand U112 (N_112,N_28,N_4);
nand U113 (N_113,In_93,In_12);
nand U114 (N_114,N_20,In_332);
nand U115 (N_115,N_6,In_378);
or U116 (N_116,In_149,In_24);
or U117 (N_117,In_408,In_402);
nand U118 (N_118,N_59,In_22);
nor U119 (N_119,In_167,In_217);
nor U120 (N_120,In_421,In_48);
nor U121 (N_121,In_475,N_89);
nor U122 (N_122,In_32,In_178);
nor U123 (N_123,In_366,In_17);
and U124 (N_124,In_183,In_168);
or U125 (N_125,In_300,N_0);
nor U126 (N_126,In_229,N_86);
nor U127 (N_127,In_106,N_13);
nor U128 (N_128,In_137,In_257);
or U129 (N_129,In_375,N_82);
nand U130 (N_130,In_212,N_10);
nand U131 (N_131,N_5,N_109);
and U132 (N_132,N_66,In_83);
or U133 (N_133,In_385,In_336);
nor U134 (N_134,In_112,N_116);
nor U135 (N_135,N_12,In_42);
nand U136 (N_136,In_1,In_387);
and U137 (N_137,In_286,In_16);
and U138 (N_138,In_139,In_309);
nand U139 (N_139,In_135,In_335);
and U140 (N_140,In_485,In_235);
nor U141 (N_141,In_452,N_80);
nor U142 (N_142,N_19,In_31);
and U143 (N_143,In_62,In_99);
and U144 (N_144,In_60,In_331);
nor U145 (N_145,In_107,In_469);
and U146 (N_146,In_490,N_107);
and U147 (N_147,In_85,In_471);
nor U148 (N_148,In_454,In_252);
and U149 (N_149,N_75,In_482);
nor U150 (N_150,In_100,In_491);
nand U151 (N_151,In_170,In_496);
or U152 (N_152,N_24,In_480);
or U153 (N_153,N_96,In_409);
nor U154 (N_154,In_466,In_256);
or U155 (N_155,N_36,In_467);
nand U156 (N_156,In_308,N_84);
and U157 (N_157,In_435,In_29);
and U158 (N_158,In_329,In_95);
and U159 (N_159,In_427,N_110);
nor U160 (N_160,In_13,In_322);
or U161 (N_161,N_97,In_481);
nor U162 (N_162,In_53,In_164);
and U163 (N_163,N_29,N_53);
nor U164 (N_164,N_98,In_476);
nand U165 (N_165,In_450,In_119);
and U166 (N_166,In_90,In_494);
or U167 (N_167,In_392,In_129);
or U168 (N_168,In_395,N_104);
and U169 (N_169,N_119,In_180);
nand U170 (N_170,In_211,N_67);
nand U171 (N_171,N_61,N_25);
and U172 (N_172,In_205,N_112);
or U173 (N_173,N_46,In_10);
and U174 (N_174,N_81,In_9);
nor U175 (N_175,In_63,In_97);
or U176 (N_176,In_357,In_293);
or U177 (N_177,In_303,In_382);
and U178 (N_178,In_228,In_153);
xnor U179 (N_179,In_190,In_441);
nand U180 (N_180,In_404,In_182);
nand U181 (N_181,N_123,In_126);
nor U182 (N_182,N_37,In_389);
nor U183 (N_183,In_104,N_134);
nor U184 (N_184,N_160,In_3);
nand U185 (N_185,N_111,In_376);
and U186 (N_186,N_74,N_64);
nand U187 (N_187,N_43,In_354);
or U188 (N_188,In_323,N_161);
nor U189 (N_189,N_85,In_27);
and U190 (N_190,In_226,N_172);
nor U191 (N_191,In_121,N_140);
and U192 (N_192,N_105,In_105);
nand U193 (N_193,In_195,In_67);
and U194 (N_194,N_124,In_459);
nor U195 (N_195,N_32,In_227);
and U196 (N_196,N_142,In_478);
nor U197 (N_197,In_296,N_152);
nor U198 (N_198,N_102,N_145);
nand U199 (N_199,N_179,N_168);
and U200 (N_200,In_43,N_108);
and U201 (N_201,N_147,N_166);
nand U202 (N_202,In_319,In_411);
or U203 (N_203,In_200,In_77);
nand U204 (N_204,In_262,In_181);
nand U205 (N_205,In_460,In_316);
nor U206 (N_206,In_136,In_222);
nand U207 (N_207,N_90,N_83);
or U208 (N_208,N_158,N_7);
nand U209 (N_209,In_244,In_241);
nand U210 (N_210,In_18,In_218);
or U211 (N_211,N_103,In_194);
nand U212 (N_212,N_77,In_438);
nor U213 (N_213,N_33,N_164);
nand U214 (N_214,N_165,N_131);
or U215 (N_215,In_451,N_169);
or U216 (N_216,In_0,In_210);
nand U217 (N_217,In_162,In_80);
or U218 (N_218,In_157,N_17);
nand U219 (N_219,In_220,N_156);
nand U220 (N_220,In_406,In_240);
or U221 (N_221,In_290,In_82);
nor U222 (N_222,In_426,In_301);
nor U223 (N_223,N_143,In_47);
nor U224 (N_224,In_237,N_146);
or U225 (N_225,In_189,N_76);
nor U226 (N_226,N_170,N_106);
nor U227 (N_227,N_31,N_63);
nor U228 (N_228,In_488,In_271);
nand U229 (N_229,In_65,In_208);
nand U230 (N_230,In_117,N_71);
nor U231 (N_231,N_157,In_108);
nor U232 (N_232,N_155,In_364);
and U233 (N_233,N_129,In_92);
and U234 (N_234,In_166,N_92);
or U235 (N_235,N_162,N_173);
nor U236 (N_236,N_144,N_137);
and U237 (N_237,In_165,N_69);
nor U238 (N_238,N_148,In_258);
nand U239 (N_239,In_196,In_381);
and U240 (N_240,N_65,N_88);
nor U241 (N_241,In_315,N_122);
nor U242 (N_242,In_161,In_140);
or U243 (N_243,In_295,In_171);
nand U244 (N_244,In_184,N_235);
and U245 (N_245,In_356,N_115);
nor U246 (N_246,N_95,N_177);
and U247 (N_247,N_68,N_47);
nand U248 (N_248,N_21,N_231);
or U249 (N_249,N_159,N_127);
nor U250 (N_250,N_54,N_132);
or U251 (N_251,In_87,N_15);
or U252 (N_252,In_461,N_100);
and U253 (N_253,In_445,In_260);
or U254 (N_254,In_216,In_272);
and U255 (N_255,In_103,N_222);
or U256 (N_256,N_113,In_144);
nor U257 (N_257,N_23,In_377);
or U258 (N_258,In_185,N_99);
nor U259 (N_259,N_151,N_154);
nand U260 (N_260,N_194,N_220);
and U261 (N_261,In_453,In_304);
or U262 (N_262,N_228,In_72);
nor U263 (N_263,In_337,N_171);
nand U264 (N_264,In_133,N_167);
xnor U265 (N_265,In_192,N_87);
and U266 (N_266,In_399,In_279);
and U267 (N_267,In_390,N_125);
or U268 (N_268,In_199,In_338);
nand U269 (N_269,In_148,In_371);
and U270 (N_270,In_98,N_175);
nor U271 (N_271,In_172,In_134);
and U272 (N_272,N_199,In_120);
xor U273 (N_273,In_160,In_4);
nand U274 (N_274,N_16,In_232);
nor U275 (N_275,In_363,In_270);
nor U276 (N_276,N_153,N_239);
nor U277 (N_277,N_193,N_187);
or U278 (N_278,In_150,In_58);
or U279 (N_279,N_196,In_215);
and U280 (N_280,In_277,N_120);
or U281 (N_281,N_9,In_440);
nand U282 (N_282,In_386,N_188);
xnor U283 (N_283,N_73,N_211);
nand U284 (N_284,N_236,In_34);
nor U285 (N_285,In_267,N_206);
nor U286 (N_286,In_61,N_208);
or U287 (N_287,In_403,In_251);
nor U288 (N_288,In_458,In_489);
and U289 (N_289,In_359,N_27);
and U290 (N_290,N_198,N_136);
nand U291 (N_291,N_118,N_52);
nor U292 (N_292,N_221,N_121);
nor U293 (N_293,In_368,N_163);
nor U294 (N_294,In_282,In_307);
or U295 (N_295,In_203,In_154);
nand U296 (N_296,N_212,In_102);
and U297 (N_297,N_210,N_192);
and U298 (N_298,N_191,N_218);
xnor U299 (N_299,In_497,N_216);
xnor U300 (N_300,N_60,In_158);
or U301 (N_301,N_72,N_291);
nor U302 (N_302,N_270,N_185);
and U303 (N_303,In_255,N_44);
and U304 (N_304,N_117,In_479);
and U305 (N_305,N_254,N_261);
nor U306 (N_306,N_255,N_243);
or U307 (N_307,In_143,N_201);
and U308 (N_308,N_260,N_256);
nor U309 (N_309,In_342,N_289);
or U310 (N_310,N_287,In_147);
and U311 (N_311,N_280,In_369);
or U312 (N_312,N_259,In_238);
or U313 (N_313,N_18,N_246);
or U314 (N_314,N_79,In_75);
nand U315 (N_315,N_180,In_340);
nand U316 (N_316,N_268,N_264);
nand U317 (N_317,In_159,In_333);
nor U318 (N_318,In_297,In_396);
nor U319 (N_319,N_138,N_62);
or U320 (N_320,In_204,N_42);
nand U321 (N_321,In_37,N_233);
nand U322 (N_322,N_141,N_269);
nand U323 (N_323,In_15,N_181);
and U324 (N_324,N_213,N_288);
and U325 (N_325,N_176,N_265);
and U326 (N_326,N_258,N_273);
nor U327 (N_327,N_217,N_240);
and U328 (N_328,In_419,In_146);
nand U329 (N_329,In_56,N_214);
and U330 (N_330,N_128,N_223);
nand U331 (N_331,N_133,In_472);
nor U332 (N_332,N_227,In_334);
and U333 (N_333,N_241,In_384);
nand U334 (N_334,N_285,In_40);
and U335 (N_335,N_224,N_101);
or U336 (N_336,N_182,N_245);
and U337 (N_337,N_279,N_209);
or U338 (N_338,N_135,In_379);
or U339 (N_339,N_174,In_96);
nor U340 (N_340,In_91,N_93);
or U341 (N_341,In_410,N_48);
xnor U342 (N_342,N_225,In_430);
nand U343 (N_343,N_149,N_40);
and U344 (N_344,N_250,N_232);
or U345 (N_345,In_422,N_200);
nand U346 (N_346,N_282,N_70);
nand U347 (N_347,In_74,N_203);
or U348 (N_348,N_294,In_493);
and U349 (N_349,N_94,N_26);
or U350 (N_350,In_465,N_299);
or U351 (N_351,In_321,N_130);
or U352 (N_352,N_219,In_462);
and U353 (N_353,N_230,N_266);
nor U354 (N_354,N_284,N_114);
xor U355 (N_355,In_370,N_286);
and U356 (N_356,N_3,N_139);
or U357 (N_357,N_226,N_38);
nor U358 (N_358,In_11,N_234);
and U359 (N_359,In_362,N_278);
nor U360 (N_360,N_207,In_284);
and U361 (N_361,N_237,N_150);
and U362 (N_362,N_305,N_39);
and U363 (N_363,N_263,N_307);
nand U364 (N_364,N_186,N_281);
or U365 (N_365,N_356,N_331);
and U366 (N_366,N_300,N_197);
or U367 (N_367,In_70,N_296);
or U368 (N_368,N_78,N_251);
xnor U369 (N_369,N_178,N_336);
or U370 (N_370,N_349,N_276);
and U371 (N_371,N_253,N_342);
or U372 (N_372,N_252,N_272);
or U373 (N_373,N_351,N_340);
or U374 (N_374,N_229,N_326);
nor U375 (N_375,N_323,In_113);
nor U376 (N_376,In_28,N_347);
or U377 (N_377,N_277,N_184);
or U378 (N_378,In_225,N_249);
or U379 (N_379,N_310,In_287);
nand U380 (N_380,N_344,N_55);
nand U381 (N_381,N_298,N_244);
or U382 (N_382,N_91,In_320);
and U383 (N_383,N_315,N_334);
nor U384 (N_384,N_327,N_357);
nand U385 (N_385,N_348,N_332);
xor U386 (N_386,In_273,N_353);
nor U387 (N_387,In_394,N_328);
and U388 (N_388,In_5,N_303);
nand U389 (N_389,In_449,In_179);
nand U390 (N_390,N_358,N_304);
nand U391 (N_391,N_346,N_335);
or U392 (N_392,N_34,N_195);
nor U393 (N_393,N_262,In_302);
or U394 (N_394,N_316,N_295);
and U395 (N_395,N_350,N_333);
nor U396 (N_396,N_267,N_204);
and U397 (N_397,N_343,N_242);
and U398 (N_398,In_417,N_8);
and U399 (N_399,N_317,N_271);
or U400 (N_400,N_306,In_349);
nor U401 (N_401,In_202,N_248);
nor U402 (N_402,N_359,N_283);
or U403 (N_403,N_309,N_352);
or U404 (N_404,N_301,N_302);
nand U405 (N_405,N_313,N_290);
nor U406 (N_406,N_311,In_468);
nor U407 (N_407,N_314,In_81);
and U408 (N_408,N_354,N_183);
and U409 (N_409,N_318,N_322);
nor U410 (N_410,N_190,N_324);
nand U411 (N_411,N_321,N_247);
or U412 (N_412,N_189,In_420);
or U413 (N_413,N_319,In_122);
nor U414 (N_414,In_429,N_275);
or U415 (N_415,N_297,N_345);
nor U416 (N_416,N_338,In_456);
or U417 (N_417,N_308,N_126);
nand U418 (N_418,N_274,N_325);
nor U419 (N_419,In_294,N_337);
or U420 (N_420,N_373,N_389);
nand U421 (N_421,N_378,N_388);
nor U422 (N_422,N_384,N_408);
nor U423 (N_423,In_352,N_416);
or U424 (N_424,N_404,N_257);
and U425 (N_425,N_205,N_368);
and U426 (N_426,N_366,N_406);
nor U427 (N_427,N_329,N_375);
nand U428 (N_428,N_369,N_409);
xor U429 (N_429,N_382,N_341);
nor U430 (N_430,N_412,N_370);
or U431 (N_431,N_377,N_405);
nand U432 (N_432,N_396,N_293);
or U433 (N_433,N_320,N_398);
nor U434 (N_434,In_59,N_312);
nand U435 (N_435,N_376,In_383);
or U436 (N_436,N_363,N_215);
nor U437 (N_437,N_360,N_397);
nand U438 (N_438,N_390,N_371);
and U439 (N_439,N_387,N_383);
nor U440 (N_440,N_380,N_367);
and U441 (N_441,N_364,N_400);
nand U442 (N_442,N_407,N_238);
nor U443 (N_443,N_374,N_413);
xnor U444 (N_444,N_391,N_392);
and U445 (N_445,N_402,N_394);
or U446 (N_446,N_393,N_292);
nor U447 (N_447,N_361,N_202);
and U448 (N_448,N_419,N_401);
nand U449 (N_449,In_138,N_399);
nor U450 (N_450,N_386,N_362);
and U451 (N_451,N_339,N_385);
or U452 (N_452,N_330,N_381);
or U453 (N_453,N_395,N_415);
or U454 (N_454,N_410,N_418);
nand U455 (N_455,In_397,N_365);
and U456 (N_456,N_379,In_247);
nand U457 (N_457,N_417,N_355);
or U458 (N_458,N_372,N_411);
or U459 (N_459,N_414,N_403);
nor U460 (N_460,N_383,N_399);
nor U461 (N_461,N_418,N_391);
nor U462 (N_462,N_402,In_397);
and U463 (N_463,N_238,N_413);
nor U464 (N_464,N_397,N_395);
nor U465 (N_465,N_376,N_361);
nand U466 (N_466,In_397,In_352);
or U467 (N_467,N_341,N_385);
and U468 (N_468,N_363,N_369);
or U469 (N_469,N_390,N_392);
nor U470 (N_470,N_398,N_385);
or U471 (N_471,N_390,N_418);
nor U472 (N_472,N_398,N_379);
or U473 (N_473,N_382,N_396);
and U474 (N_474,N_341,N_360);
nand U475 (N_475,N_320,N_361);
nor U476 (N_476,N_373,In_59);
and U477 (N_477,N_320,N_368);
nand U478 (N_478,N_410,N_381);
nand U479 (N_479,N_339,N_376);
nand U480 (N_480,N_470,N_426);
nor U481 (N_481,N_461,N_451);
nand U482 (N_482,N_457,N_458);
nor U483 (N_483,N_432,N_428);
nor U484 (N_484,N_423,N_476);
nand U485 (N_485,N_427,N_455);
or U486 (N_486,N_473,N_436);
or U487 (N_487,N_429,N_456);
nor U488 (N_488,N_462,N_475);
nand U489 (N_489,N_454,N_464);
nand U490 (N_490,N_441,N_438);
or U491 (N_491,N_422,N_437);
nand U492 (N_492,N_468,N_425);
or U493 (N_493,N_420,N_474);
nand U494 (N_494,N_446,N_469);
nand U495 (N_495,N_450,N_421);
nor U496 (N_496,N_433,N_449);
or U497 (N_497,N_445,N_448);
or U498 (N_498,N_440,N_471);
nor U499 (N_499,N_472,N_443);
and U500 (N_500,N_435,N_452);
or U501 (N_501,N_453,N_460);
nand U502 (N_502,N_431,N_424);
and U503 (N_503,N_467,N_444);
nor U504 (N_504,N_463,N_466);
nand U505 (N_505,N_478,N_442);
and U506 (N_506,N_477,N_465);
nand U507 (N_507,N_479,N_434);
nor U508 (N_508,N_430,N_459);
nor U509 (N_509,N_447,N_439);
and U510 (N_510,N_459,N_470);
or U511 (N_511,N_477,N_429);
nor U512 (N_512,N_447,N_471);
or U513 (N_513,N_450,N_472);
and U514 (N_514,N_475,N_474);
or U515 (N_515,N_432,N_463);
or U516 (N_516,N_449,N_456);
nand U517 (N_517,N_452,N_465);
nand U518 (N_518,N_463,N_446);
nand U519 (N_519,N_449,N_455);
or U520 (N_520,N_434,N_421);
or U521 (N_521,N_448,N_465);
or U522 (N_522,N_447,N_450);
or U523 (N_523,N_442,N_446);
nand U524 (N_524,N_478,N_464);
or U525 (N_525,N_432,N_434);
nand U526 (N_526,N_450,N_469);
or U527 (N_527,N_477,N_470);
nand U528 (N_528,N_432,N_445);
or U529 (N_529,N_432,N_436);
nand U530 (N_530,N_469,N_459);
and U531 (N_531,N_449,N_468);
and U532 (N_532,N_429,N_438);
nor U533 (N_533,N_455,N_442);
nor U534 (N_534,N_450,N_431);
nand U535 (N_535,N_421,N_459);
nor U536 (N_536,N_422,N_474);
or U537 (N_537,N_477,N_427);
and U538 (N_538,N_446,N_422);
or U539 (N_539,N_473,N_460);
nor U540 (N_540,N_533,N_524);
or U541 (N_541,N_519,N_498);
or U542 (N_542,N_532,N_517);
nor U543 (N_543,N_534,N_530);
or U544 (N_544,N_480,N_504);
nand U545 (N_545,N_535,N_529);
nand U546 (N_546,N_490,N_483);
and U547 (N_547,N_503,N_481);
or U548 (N_548,N_489,N_523);
nor U549 (N_549,N_501,N_518);
and U550 (N_550,N_496,N_510);
nor U551 (N_551,N_515,N_506);
nand U552 (N_552,N_497,N_485);
or U553 (N_553,N_486,N_484);
or U554 (N_554,N_538,N_507);
or U555 (N_555,N_493,N_495);
or U556 (N_556,N_525,N_491);
and U557 (N_557,N_521,N_531);
nor U558 (N_558,N_488,N_487);
nor U559 (N_559,N_494,N_537);
or U560 (N_560,N_508,N_499);
nand U561 (N_561,N_528,N_539);
xor U562 (N_562,N_505,N_513);
and U563 (N_563,N_511,N_522);
nand U564 (N_564,N_516,N_512);
and U565 (N_565,N_482,N_520);
nor U566 (N_566,N_509,N_536);
and U567 (N_567,N_527,N_492);
nand U568 (N_568,N_500,N_502);
and U569 (N_569,N_526,N_514);
and U570 (N_570,N_483,N_524);
nor U571 (N_571,N_527,N_501);
nor U572 (N_572,N_519,N_510);
nor U573 (N_573,N_509,N_526);
and U574 (N_574,N_528,N_501);
nand U575 (N_575,N_514,N_507);
nand U576 (N_576,N_490,N_500);
nand U577 (N_577,N_526,N_515);
nor U578 (N_578,N_531,N_517);
nand U579 (N_579,N_503,N_518);
or U580 (N_580,N_512,N_525);
nand U581 (N_581,N_503,N_502);
and U582 (N_582,N_495,N_506);
or U583 (N_583,N_539,N_494);
nand U584 (N_584,N_484,N_537);
nor U585 (N_585,N_509,N_508);
nand U586 (N_586,N_527,N_526);
or U587 (N_587,N_528,N_493);
or U588 (N_588,N_526,N_489);
nand U589 (N_589,N_535,N_490);
nor U590 (N_590,N_515,N_516);
and U591 (N_591,N_492,N_519);
nand U592 (N_592,N_502,N_539);
nand U593 (N_593,N_482,N_536);
and U594 (N_594,N_512,N_508);
nand U595 (N_595,N_536,N_503);
nor U596 (N_596,N_509,N_483);
or U597 (N_597,N_489,N_511);
and U598 (N_598,N_536,N_499);
nand U599 (N_599,N_515,N_480);
or U600 (N_600,N_552,N_565);
and U601 (N_601,N_581,N_562);
and U602 (N_602,N_572,N_574);
nor U603 (N_603,N_585,N_564);
nand U604 (N_604,N_557,N_556);
and U605 (N_605,N_577,N_599);
or U606 (N_606,N_570,N_590);
xnor U607 (N_607,N_593,N_549);
and U608 (N_608,N_547,N_584);
or U609 (N_609,N_586,N_580);
nor U610 (N_610,N_553,N_567);
nor U611 (N_611,N_595,N_558);
xor U612 (N_612,N_540,N_555);
nor U613 (N_613,N_550,N_598);
and U614 (N_614,N_541,N_578);
or U615 (N_615,N_592,N_583);
or U616 (N_616,N_576,N_566);
nor U617 (N_617,N_559,N_596);
and U618 (N_618,N_594,N_569);
or U619 (N_619,N_573,N_543);
and U620 (N_620,N_563,N_545);
or U621 (N_621,N_571,N_548);
nand U622 (N_622,N_589,N_591);
nand U623 (N_623,N_582,N_597);
nand U624 (N_624,N_544,N_561);
nor U625 (N_625,N_551,N_560);
and U626 (N_626,N_568,N_579);
nor U627 (N_627,N_587,N_575);
or U628 (N_628,N_554,N_546);
and U629 (N_629,N_588,N_542);
and U630 (N_630,N_596,N_550);
nand U631 (N_631,N_554,N_544);
or U632 (N_632,N_568,N_573);
nand U633 (N_633,N_550,N_557);
xor U634 (N_634,N_568,N_577);
nand U635 (N_635,N_549,N_579);
or U636 (N_636,N_549,N_585);
or U637 (N_637,N_584,N_574);
and U638 (N_638,N_547,N_563);
or U639 (N_639,N_561,N_545);
nand U640 (N_640,N_546,N_563);
and U641 (N_641,N_596,N_591);
or U642 (N_642,N_567,N_582);
nand U643 (N_643,N_572,N_577);
nor U644 (N_644,N_582,N_596);
or U645 (N_645,N_588,N_595);
or U646 (N_646,N_543,N_563);
nor U647 (N_647,N_567,N_591);
and U648 (N_648,N_585,N_575);
and U649 (N_649,N_560,N_582);
or U650 (N_650,N_542,N_545);
xnor U651 (N_651,N_554,N_589);
nand U652 (N_652,N_574,N_569);
nand U653 (N_653,N_581,N_595);
nor U654 (N_654,N_583,N_587);
and U655 (N_655,N_542,N_578);
or U656 (N_656,N_551,N_554);
nor U657 (N_657,N_555,N_592);
nor U658 (N_658,N_568,N_576);
xor U659 (N_659,N_577,N_578);
nor U660 (N_660,N_625,N_647);
nand U661 (N_661,N_614,N_601);
nand U662 (N_662,N_621,N_659);
nor U663 (N_663,N_613,N_654);
or U664 (N_664,N_610,N_623);
nand U665 (N_665,N_608,N_615);
and U666 (N_666,N_635,N_600);
or U667 (N_667,N_620,N_633);
or U668 (N_668,N_637,N_656);
nor U669 (N_669,N_611,N_616);
or U670 (N_670,N_602,N_642);
nor U671 (N_671,N_624,N_639);
nor U672 (N_672,N_630,N_612);
and U673 (N_673,N_652,N_646);
nor U674 (N_674,N_653,N_629);
and U675 (N_675,N_607,N_632);
nor U676 (N_676,N_657,N_618);
and U677 (N_677,N_605,N_655);
xor U678 (N_678,N_617,N_658);
nand U679 (N_679,N_627,N_638);
and U680 (N_680,N_645,N_644);
and U681 (N_681,N_619,N_606);
nand U682 (N_682,N_636,N_643);
and U683 (N_683,N_604,N_634);
and U684 (N_684,N_603,N_648);
nor U685 (N_685,N_641,N_649);
and U686 (N_686,N_640,N_628);
nor U687 (N_687,N_609,N_651);
nand U688 (N_688,N_626,N_631);
nand U689 (N_689,N_622,N_650);
and U690 (N_690,N_655,N_606);
nand U691 (N_691,N_652,N_634);
and U692 (N_692,N_627,N_637);
nand U693 (N_693,N_658,N_631);
nor U694 (N_694,N_606,N_612);
and U695 (N_695,N_619,N_617);
nand U696 (N_696,N_640,N_652);
nor U697 (N_697,N_618,N_623);
nor U698 (N_698,N_646,N_614);
nand U699 (N_699,N_644,N_646);
and U700 (N_700,N_612,N_641);
xnor U701 (N_701,N_609,N_656);
or U702 (N_702,N_623,N_615);
nor U703 (N_703,N_606,N_638);
and U704 (N_704,N_643,N_651);
nor U705 (N_705,N_607,N_640);
nor U706 (N_706,N_629,N_656);
nor U707 (N_707,N_610,N_647);
xnor U708 (N_708,N_610,N_656);
nor U709 (N_709,N_645,N_603);
or U710 (N_710,N_644,N_603);
and U711 (N_711,N_629,N_631);
or U712 (N_712,N_632,N_619);
nor U713 (N_713,N_631,N_646);
and U714 (N_714,N_640,N_617);
nor U715 (N_715,N_611,N_659);
or U716 (N_716,N_620,N_639);
or U717 (N_717,N_650,N_636);
and U718 (N_718,N_657,N_624);
nor U719 (N_719,N_617,N_643);
and U720 (N_720,N_669,N_689);
nand U721 (N_721,N_680,N_701);
xnor U722 (N_722,N_672,N_714);
or U723 (N_723,N_700,N_718);
or U724 (N_724,N_682,N_707);
and U725 (N_725,N_691,N_719);
nand U726 (N_726,N_661,N_702);
nor U727 (N_727,N_710,N_686);
nor U728 (N_728,N_666,N_681);
nand U729 (N_729,N_676,N_664);
or U730 (N_730,N_693,N_692);
nor U731 (N_731,N_683,N_663);
or U732 (N_732,N_705,N_685);
nand U733 (N_733,N_698,N_668);
and U734 (N_734,N_674,N_688);
and U735 (N_735,N_716,N_704);
nand U736 (N_736,N_695,N_667);
and U737 (N_737,N_709,N_665);
and U738 (N_738,N_673,N_671);
or U739 (N_739,N_694,N_675);
nor U740 (N_740,N_706,N_715);
nor U741 (N_741,N_708,N_699);
nand U742 (N_742,N_670,N_703);
nand U743 (N_743,N_687,N_677);
and U744 (N_744,N_717,N_696);
or U745 (N_745,N_678,N_712);
or U746 (N_746,N_684,N_713);
nand U747 (N_747,N_697,N_690);
or U748 (N_748,N_711,N_660);
nand U749 (N_749,N_662,N_679);
or U750 (N_750,N_711,N_668);
or U751 (N_751,N_713,N_678);
or U752 (N_752,N_690,N_710);
or U753 (N_753,N_701,N_660);
or U754 (N_754,N_672,N_687);
and U755 (N_755,N_680,N_668);
and U756 (N_756,N_681,N_707);
and U757 (N_757,N_708,N_702);
or U758 (N_758,N_691,N_677);
or U759 (N_759,N_718,N_715);
or U760 (N_760,N_664,N_689);
nand U761 (N_761,N_713,N_702);
or U762 (N_762,N_702,N_706);
or U763 (N_763,N_692,N_663);
nor U764 (N_764,N_666,N_680);
and U765 (N_765,N_679,N_663);
xor U766 (N_766,N_691,N_707);
nor U767 (N_767,N_696,N_708);
or U768 (N_768,N_675,N_712);
nand U769 (N_769,N_680,N_713);
and U770 (N_770,N_702,N_660);
or U771 (N_771,N_705,N_662);
and U772 (N_772,N_719,N_675);
nand U773 (N_773,N_663,N_699);
nand U774 (N_774,N_671,N_691);
and U775 (N_775,N_681,N_682);
or U776 (N_776,N_710,N_680);
nand U777 (N_777,N_710,N_698);
and U778 (N_778,N_685,N_661);
and U779 (N_779,N_696,N_697);
and U780 (N_780,N_737,N_768);
nand U781 (N_781,N_749,N_729);
nor U782 (N_782,N_745,N_765);
nand U783 (N_783,N_753,N_735);
or U784 (N_784,N_770,N_726);
nor U785 (N_785,N_747,N_752);
and U786 (N_786,N_762,N_734);
or U787 (N_787,N_778,N_777);
nand U788 (N_788,N_739,N_721);
nand U789 (N_789,N_766,N_733);
or U790 (N_790,N_748,N_776);
or U791 (N_791,N_722,N_757);
and U792 (N_792,N_756,N_724);
xnor U793 (N_793,N_723,N_758);
nor U794 (N_794,N_754,N_744);
and U795 (N_795,N_741,N_727);
or U796 (N_796,N_779,N_743);
nand U797 (N_797,N_769,N_736);
and U798 (N_798,N_771,N_761);
or U799 (N_799,N_773,N_742);
nor U800 (N_800,N_730,N_746);
or U801 (N_801,N_764,N_772);
nor U802 (N_802,N_740,N_751);
and U803 (N_803,N_728,N_760);
or U804 (N_804,N_755,N_725);
nand U805 (N_805,N_767,N_759);
or U806 (N_806,N_732,N_731);
nor U807 (N_807,N_775,N_720);
nor U808 (N_808,N_738,N_750);
and U809 (N_809,N_763,N_774);
nor U810 (N_810,N_771,N_748);
nand U811 (N_811,N_749,N_762);
or U812 (N_812,N_765,N_761);
nor U813 (N_813,N_723,N_736);
nor U814 (N_814,N_772,N_768);
or U815 (N_815,N_759,N_726);
nand U816 (N_816,N_728,N_772);
and U817 (N_817,N_745,N_740);
or U818 (N_818,N_745,N_752);
and U819 (N_819,N_720,N_769);
and U820 (N_820,N_767,N_723);
nor U821 (N_821,N_763,N_730);
nor U822 (N_822,N_728,N_745);
nand U823 (N_823,N_762,N_733);
and U824 (N_824,N_760,N_747);
nand U825 (N_825,N_728,N_749);
nor U826 (N_826,N_778,N_779);
nand U827 (N_827,N_772,N_761);
nor U828 (N_828,N_769,N_748);
and U829 (N_829,N_763,N_743);
or U830 (N_830,N_768,N_732);
nor U831 (N_831,N_747,N_761);
or U832 (N_832,N_746,N_739);
or U833 (N_833,N_748,N_772);
nand U834 (N_834,N_754,N_741);
or U835 (N_835,N_729,N_739);
nand U836 (N_836,N_767,N_753);
nor U837 (N_837,N_729,N_761);
nor U838 (N_838,N_745,N_771);
or U839 (N_839,N_762,N_772);
nand U840 (N_840,N_795,N_837);
and U841 (N_841,N_796,N_785);
and U842 (N_842,N_836,N_833);
or U843 (N_843,N_780,N_814);
nand U844 (N_844,N_812,N_827);
nor U845 (N_845,N_790,N_800);
and U846 (N_846,N_803,N_788);
nor U847 (N_847,N_817,N_807);
and U848 (N_848,N_808,N_825);
nor U849 (N_849,N_799,N_835);
or U850 (N_850,N_810,N_828);
nand U851 (N_851,N_793,N_782);
and U852 (N_852,N_809,N_820);
and U853 (N_853,N_829,N_816);
nand U854 (N_854,N_826,N_813);
nand U855 (N_855,N_834,N_818);
and U856 (N_856,N_821,N_783);
nor U857 (N_857,N_786,N_791);
and U858 (N_858,N_797,N_804);
nand U859 (N_859,N_831,N_794);
or U860 (N_860,N_838,N_801);
nand U861 (N_861,N_805,N_822);
or U862 (N_862,N_830,N_781);
and U863 (N_863,N_823,N_802);
and U864 (N_864,N_824,N_789);
and U865 (N_865,N_787,N_806);
or U866 (N_866,N_839,N_798);
nor U867 (N_867,N_832,N_792);
nor U868 (N_868,N_811,N_815);
nand U869 (N_869,N_784,N_819);
and U870 (N_870,N_796,N_784);
and U871 (N_871,N_780,N_837);
nand U872 (N_872,N_829,N_795);
and U873 (N_873,N_781,N_818);
nand U874 (N_874,N_838,N_810);
and U875 (N_875,N_821,N_798);
or U876 (N_876,N_789,N_832);
and U877 (N_877,N_816,N_814);
nand U878 (N_878,N_796,N_810);
and U879 (N_879,N_829,N_805);
nor U880 (N_880,N_811,N_798);
or U881 (N_881,N_820,N_826);
nand U882 (N_882,N_830,N_829);
or U883 (N_883,N_817,N_820);
or U884 (N_884,N_837,N_792);
nor U885 (N_885,N_788,N_796);
nor U886 (N_886,N_827,N_796);
or U887 (N_887,N_819,N_832);
xnor U888 (N_888,N_828,N_820);
and U889 (N_889,N_824,N_814);
and U890 (N_890,N_820,N_812);
nand U891 (N_891,N_831,N_838);
and U892 (N_892,N_811,N_791);
nor U893 (N_893,N_824,N_828);
or U894 (N_894,N_820,N_785);
nor U895 (N_895,N_783,N_781);
xnor U896 (N_896,N_819,N_825);
and U897 (N_897,N_824,N_781);
nor U898 (N_898,N_812,N_794);
nand U899 (N_899,N_803,N_821);
or U900 (N_900,N_887,N_853);
nand U901 (N_901,N_876,N_842);
nor U902 (N_902,N_873,N_878);
and U903 (N_903,N_857,N_883);
nand U904 (N_904,N_863,N_865);
nor U905 (N_905,N_874,N_858);
nor U906 (N_906,N_880,N_862);
xor U907 (N_907,N_893,N_879);
nor U908 (N_908,N_871,N_840);
or U909 (N_909,N_864,N_895);
nor U910 (N_910,N_866,N_892);
nand U911 (N_911,N_891,N_847);
xnor U912 (N_912,N_899,N_872);
or U913 (N_913,N_884,N_861);
or U914 (N_914,N_885,N_867);
nand U915 (N_915,N_849,N_881);
nand U916 (N_916,N_869,N_888);
or U917 (N_917,N_841,N_886);
and U918 (N_918,N_868,N_894);
nand U919 (N_919,N_852,N_877);
and U920 (N_920,N_846,N_845);
and U921 (N_921,N_855,N_889);
or U922 (N_922,N_897,N_860);
nor U923 (N_923,N_859,N_870);
or U924 (N_924,N_875,N_890);
xor U925 (N_925,N_856,N_854);
and U926 (N_926,N_850,N_898);
nor U927 (N_927,N_843,N_882);
xnor U928 (N_928,N_844,N_851);
nor U929 (N_929,N_848,N_896);
nor U930 (N_930,N_899,N_840);
nor U931 (N_931,N_892,N_859);
nor U932 (N_932,N_881,N_850);
nor U933 (N_933,N_874,N_852);
and U934 (N_934,N_888,N_858);
and U935 (N_935,N_864,N_855);
and U936 (N_936,N_869,N_850);
nor U937 (N_937,N_888,N_879);
and U938 (N_938,N_856,N_867);
and U939 (N_939,N_856,N_863);
and U940 (N_940,N_857,N_873);
nand U941 (N_941,N_885,N_855);
and U942 (N_942,N_841,N_877);
and U943 (N_943,N_883,N_899);
and U944 (N_944,N_881,N_857);
and U945 (N_945,N_870,N_848);
nor U946 (N_946,N_878,N_895);
and U947 (N_947,N_891,N_850);
and U948 (N_948,N_843,N_850);
and U949 (N_949,N_864,N_840);
or U950 (N_950,N_868,N_864);
nor U951 (N_951,N_851,N_861);
nor U952 (N_952,N_893,N_844);
and U953 (N_953,N_892,N_860);
or U954 (N_954,N_894,N_856);
or U955 (N_955,N_879,N_873);
nor U956 (N_956,N_868,N_874);
and U957 (N_957,N_847,N_892);
and U958 (N_958,N_894,N_851);
nor U959 (N_959,N_862,N_853);
nor U960 (N_960,N_903,N_949);
nor U961 (N_961,N_942,N_909);
or U962 (N_962,N_901,N_951);
nor U963 (N_963,N_953,N_956);
or U964 (N_964,N_917,N_957);
nand U965 (N_965,N_950,N_954);
nand U966 (N_966,N_922,N_932);
and U967 (N_967,N_928,N_945);
or U968 (N_968,N_925,N_934);
nor U969 (N_969,N_952,N_938);
and U970 (N_970,N_923,N_924);
nand U971 (N_971,N_930,N_908);
nand U972 (N_972,N_937,N_955);
or U973 (N_973,N_931,N_905);
nand U974 (N_974,N_902,N_913);
or U975 (N_975,N_916,N_941);
or U976 (N_976,N_918,N_912);
or U977 (N_977,N_936,N_959);
and U978 (N_978,N_948,N_929);
or U979 (N_979,N_904,N_935);
or U980 (N_980,N_919,N_907);
nor U981 (N_981,N_944,N_927);
nand U982 (N_982,N_958,N_947);
nand U983 (N_983,N_933,N_911);
nor U984 (N_984,N_940,N_900);
nor U985 (N_985,N_926,N_943);
and U986 (N_986,N_910,N_921);
or U987 (N_987,N_906,N_939);
nor U988 (N_988,N_946,N_915);
and U989 (N_989,N_920,N_914);
nor U990 (N_990,N_956,N_957);
and U991 (N_991,N_935,N_903);
nand U992 (N_992,N_930,N_944);
nor U993 (N_993,N_906,N_920);
nand U994 (N_994,N_951,N_935);
nand U995 (N_995,N_912,N_944);
nor U996 (N_996,N_923,N_958);
nand U997 (N_997,N_912,N_940);
and U998 (N_998,N_934,N_900);
or U999 (N_999,N_912,N_956);
nor U1000 (N_1000,N_930,N_921);
nand U1001 (N_1001,N_901,N_932);
xor U1002 (N_1002,N_921,N_918);
or U1003 (N_1003,N_915,N_942);
nand U1004 (N_1004,N_949,N_931);
and U1005 (N_1005,N_926,N_923);
or U1006 (N_1006,N_912,N_929);
or U1007 (N_1007,N_955,N_951);
nand U1008 (N_1008,N_944,N_911);
or U1009 (N_1009,N_925,N_906);
nor U1010 (N_1010,N_914,N_952);
or U1011 (N_1011,N_934,N_930);
nor U1012 (N_1012,N_927,N_936);
and U1013 (N_1013,N_911,N_907);
and U1014 (N_1014,N_933,N_958);
nor U1015 (N_1015,N_933,N_922);
or U1016 (N_1016,N_914,N_911);
and U1017 (N_1017,N_948,N_928);
or U1018 (N_1018,N_934,N_931);
or U1019 (N_1019,N_935,N_953);
or U1020 (N_1020,N_1006,N_969);
nand U1021 (N_1021,N_978,N_961);
or U1022 (N_1022,N_963,N_967);
nand U1023 (N_1023,N_1015,N_987);
nor U1024 (N_1024,N_1014,N_995);
nor U1025 (N_1025,N_968,N_986);
nor U1026 (N_1026,N_996,N_984);
nor U1027 (N_1027,N_990,N_998);
nand U1028 (N_1028,N_1004,N_1000);
nand U1029 (N_1029,N_965,N_966);
and U1030 (N_1030,N_993,N_1008);
or U1031 (N_1031,N_962,N_988);
nand U1032 (N_1032,N_1007,N_1002);
and U1033 (N_1033,N_973,N_994);
and U1034 (N_1034,N_991,N_997);
nor U1035 (N_1035,N_989,N_999);
nor U1036 (N_1036,N_1019,N_1010);
nor U1037 (N_1037,N_1003,N_985);
nand U1038 (N_1038,N_983,N_976);
and U1039 (N_1039,N_1013,N_1011);
nand U1040 (N_1040,N_964,N_970);
and U1041 (N_1041,N_982,N_971);
nand U1042 (N_1042,N_1009,N_1005);
or U1043 (N_1043,N_979,N_975);
or U1044 (N_1044,N_960,N_992);
or U1045 (N_1045,N_1012,N_1016);
or U1046 (N_1046,N_1018,N_981);
and U1047 (N_1047,N_980,N_977);
nand U1048 (N_1048,N_1017,N_972);
and U1049 (N_1049,N_1001,N_974);
and U1050 (N_1050,N_1018,N_969);
nor U1051 (N_1051,N_984,N_973);
nand U1052 (N_1052,N_1017,N_961);
or U1053 (N_1053,N_976,N_1004);
nor U1054 (N_1054,N_1007,N_1005);
and U1055 (N_1055,N_979,N_973);
nand U1056 (N_1056,N_971,N_1015);
xnor U1057 (N_1057,N_991,N_990);
or U1058 (N_1058,N_1001,N_963);
xor U1059 (N_1059,N_993,N_982);
and U1060 (N_1060,N_998,N_972);
nor U1061 (N_1061,N_1011,N_996);
nor U1062 (N_1062,N_1017,N_969);
nand U1063 (N_1063,N_986,N_984);
and U1064 (N_1064,N_1017,N_1009);
and U1065 (N_1065,N_1014,N_1003);
nor U1066 (N_1066,N_1008,N_975);
nor U1067 (N_1067,N_985,N_976);
nor U1068 (N_1068,N_980,N_963);
and U1069 (N_1069,N_990,N_974);
nor U1070 (N_1070,N_961,N_1010);
nand U1071 (N_1071,N_986,N_973);
nand U1072 (N_1072,N_1019,N_986);
nand U1073 (N_1073,N_976,N_1018);
or U1074 (N_1074,N_1015,N_1005);
and U1075 (N_1075,N_991,N_994);
nand U1076 (N_1076,N_998,N_1007);
xor U1077 (N_1077,N_1013,N_1012);
and U1078 (N_1078,N_994,N_992);
nand U1079 (N_1079,N_985,N_961);
or U1080 (N_1080,N_1035,N_1056);
or U1081 (N_1081,N_1076,N_1025);
nor U1082 (N_1082,N_1052,N_1037);
nor U1083 (N_1083,N_1022,N_1078);
nor U1084 (N_1084,N_1040,N_1049);
and U1085 (N_1085,N_1079,N_1069);
and U1086 (N_1086,N_1026,N_1021);
nor U1087 (N_1087,N_1059,N_1030);
or U1088 (N_1088,N_1073,N_1039);
nand U1089 (N_1089,N_1067,N_1033);
nand U1090 (N_1090,N_1054,N_1042);
or U1091 (N_1091,N_1023,N_1058);
and U1092 (N_1092,N_1055,N_1072);
or U1093 (N_1093,N_1068,N_1050);
and U1094 (N_1094,N_1065,N_1028);
nor U1095 (N_1095,N_1074,N_1041);
nor U1096 (N_1096,N_1043,N_1044);
nand U1097 (N_1097,N_1057,N_1064);
nand U1098 (N_1098,N_1034,N_1046);
nand U1099 (N_1099,N_1047,N_1031);
and U1100 (N_1100,N_1071,N_1066);
and U1101 (N_1101,N_1048,N_1038);
and U1102 (N_1102,N_1036,N_1062);
nand U1103 (N_1103,N_1060,N_1027);
xnor U1104 (N_1104,N_1061,N_1063);
nor U1105 (N_1105,N_1024,N_1045);
nor U1106 (N_1106,N_1020,N_1053);
nand U1107 (N_1107,N_1077,N_1075);
nor U1108 (N_1108,N_1032,N_1070);
or U1109 (N_1109,N_1051,N_1029);
and U1110 (N_1110,N_1059,N_1036);
nor U1111 (N_1111,N_1070,N_1023);
nor U1112 (N_1112,N_1045,N_1074);
nor U1113 (N_1113,N_1075,N_1071);
nor U1114 (N_1114,N_1046,N_1030);
nor U1115 (N_1115,N_1020,N_1047);
nand U1116 (N_1116,N_1066,N_1074);
or U1117 (N_1117,N_1070,N_1046);
nand U1118 (N_1118,N_1037,N_1056);
nand U1119 (N_1119,N_1034,N_1075);
and U1120 (N_1120,N_1032,N_1021);
or U1121 (N_1121,N_1030,N_1073);
nor U1122 (N_1122,N_1061,N_1022);
nand U1123 (N_1123,N_1068,N_1070);
nand U1124 (N_1124,N_1059,N_1061);
or U1125 (N_1125,N_1048,N_1075);
nor U1126 (N_1126,N_1038,N_1058);
and U1127 (N_1127,N_1061,N_1070);
nand U1128 (N_1128,N_1075,N_1046);
or U1129 (N_1129,N_1044,N_1063);
or U1130 (N_1130,N_1044,N_1054);
nand U1131 (N_1131,N_1058,N_1071);
nand U1132 (N_1132,N_1031,N_1030);
xor U1133 (N_1133,N_1063,N_1055);
nand U1134 (N_1134,N_1022,N_1040);
nand U1135 (N_1135,N_1069,N_1058);
and U1136 (N_1136,N_1044,N_1069);
nand U1137 (N_1137,N_1067,N_1040);
and U1138 (N_1138,N_1035,N_1045);
nor U1139 (N_1139,N_1042,N_1035);
nand U1140 (N_1140,N_1087,N_1127);
nor U1141 (N_1141,N_1119,N_1106);
or U1142 (N_1142,N_1089,N_1086);
or U1143 (N_1143,N_1108,N_1082);
and U1144 (N_1144,N_1133,N_1107);
and U1145 (N_1145,N_1081,N_1088);
nand U1146 (N_1146,N_1115,N_1116);
or U1147 (N_1147,N_1137,N_1094);
or U1148 (N_1148,N_1105,N_1136);
nand U1149 (N_1149,N_1113,N_1126);
nor U1150 (N_1150,N_1124,N_1093);
and U1151 (N_1151,N_1128,N_1132);
nor U1152 (N_1152,N_1109,N_1090);
or U1153 (N_1153,N_1102,N_1125);
nor U1154 (N_1154,N_1117,N_1092);
and U1155 (N_1155,N_1123,N_1096);
and U1156 (N_1156,N_1091,N_1122);
or U1157 (N_1157,N_1111,N_1098);
and U1158 (N_1158,N_1100,N_1121);
or U1159 (N_1159,N_1112,N_1131);
nand U1160 (N_1160,N_1080,N_1101);
or U1161 (N_1161,N_1130,N_1099);
nor U1162 (N_1162,N_1104,N_1103);
or U1163 (N_1163,N_1095,N_1135);
nand U1164 (N_1164,N_1083,N_1139);
nand U1165 (N_1165,N_1114,N_1110);
nor U1166 (N_1166,N_1084,N_1118);
or U1167 (N_1167,N_1134,N_1097);
or U1168 (N_1168,N_1138,N_1120);
nand U1169 (N_1169,N_1129,N_1085);
nand U1170 (N_1170,N_1124,N_1122);
nand U1171 (N_1171,N_1128,N_1126);
nor U1172 (N_1172,N_1110,N_1129);
nor U1173 (N_1173,N_1109,N_1088);
nand U1174 (N_1174,N_1125,N_1138);
and U1175 (N_1175,N_1101,N_1117);
and U1176 (N_1176,N_1123,N_1116);
nor U1177 (N_1177,N_1124,N_1101);
nor U1178 (N_1178,N_1080,N_1120);
nor U1179 (N_1179,N_1132,N_1112);
or U1180 (N_1180,N_1082,N_1086);
or U1181 (N_1181,N_1122,N_1088);
nand U1182 (N_1182,N_1089,N_1084);
and U1183 (N_1183,N_1107,N_1116);
and U1184 (N_1184,N_1102,N_1124);
and U1185 (N_1185,N_1115,N_1127);
nand U1186 (N_1186,N_1125,N_1090);
or U1187 (N_1187,N_1138,N_1113);
or U1188 (N_1188,N_1099,N_1119);
or U1189 (N_1189,N_1110,N_1105);
nor U1190 (N_1190,N_1096,N_1132);
nand U1191 (N_1191,N_1099,N_1136);
and U1192 (N_1192,N_1124,N_1092);
and U1193 (N_1193,N_1090,N_1089);
and U1194 (N_1194,N_1117,N_1102);
and U1195 (N_1195,N_1088,N_1121);
nand U1196 (N_1196,N_1116,N_1102);
nand U1197 (N_1197,N_1137,N_1122);
and U1198 (N_1198,N_1129,N_1086);
or U1199 (N_1199,N_1121,N_1135);
nor U1200 (N_1200,N_1186,N_1174);
nor U1201 (N_1201,N_1184,N_1185);
and U1202 (N_1202,N_1154,N_1146);
nor U1203 (N_1203,N_1178,N_1198);
or U1204 (N_1204,N_1153,N_1147);
nand U1205 (N_1205,N_1199,N_1144);
nand U1206 (N_1206,N_1192,N_1163);
nor U1207 (N_1207,N_1169,N_1183);
nor U1208 (N_1208,N_1190,N_1143);
nor U1209 (N_1209,N_1181,N_1177);
or U1210 (N_1210,N_1191,N_1155);
or U1211 (N_1211,N_1149,N_1172);
nor U1212 (N_1212,N_1179,N_1170);
nand U1213 (N_1213,N_1193,N_1189);
nor U1214 (N_1214,N_1156,N_1194);
and U1215 (N_1215,N_1162,N_1188);
nor U1216 (N_1216,N_1159,N_1141);
nor U1217 (N_1217,N_1187,N_1161);
xnor U1218 (N_1218,N_1160,N_1166);
and U1219 (N_1219,N_1168,N_1175);
and U1220 (N_1220,N_1182,N_1197);
nor U1221 (N_1221,N_1195,N_1173);
and U1222 (N_1222,N_1171,N_1148);
nor U1223 (N_1223,N_1152,N_1158);
nor U1224 (N_1224,N_1164,N_1157);
and U1225 (N_1225,N_1150,N_1165);
nand U1226 (N_1226,N_1167,N_1176);
nand U1227 (N_1227,N_1180,N_1196);
nor U1228 (N_1228,N_1140,N_1151);
or U1229 (N_1229,N_1142,N_1145);
and U1230 (N_1230,N_1191,N_1185);
nand U1231 (N_1231,N_1146,N_1192);
nand U1232 (N_1232,N_1143,N_1180);
nand U1233 (N_1233,N_1159,N_1176);
nand U1234 (N_1234,N_1143,N_1185);
or U1235 (N_1235,N_1191,N_1159);
nor U1236 (N_1236,N_1192,N_1157);
and U1237 (N_1237,N_1166,N_1161);
nor U1238 (N_1238,N_1147,N_1191);
or U1239 (N_1239,N_1174,N_1192);
nor U1240 (N_1240,N_1158,N_1147);
nand U1241 (N_1241,N_1141,N_1153);
or U1242 (N_1242,N_1152,N_1151);
nand U1243 (N_1243,N_1179,N_1181);
nand U1244 (N_1244,N_1158,N_1142);
nor U1245 (N_1245,N_1194,N_1140);
xor U1246 (N_1246,N_1153,N_1183);
and U1247 (N_1247,N_1160,N_1187);
and U1248 (N_1248,N_1160,N_1155);
or U1249 (N_1249,N_1144,N_1179);
nand U1250 (N_1250,N_1147,N_1187);
nand U1251 (N_1251,N_1171,N_1152);
nor U1252 (N_1252,N_1144,N_1140);
and U1253 (N_1253,N_1152,N_1199);
nand U1254 (N_1254,N_1174,N_1158);
nand U1255 (N_1255,N_1195,N_1199);
nand U1256 (N_1256,N_1142,N_1185);
or U1257 (N_1257,N_1198,N_1183);
and U1258 (N_1258,N_1195,N_1140);
or U1259 (N_1259,N_1157,N_1176);
nor U1260 (N_1260,N_1247,N_1242);
nor U1261 (N_1261,N_1225,N_1251);
and U1262 (N_1262,N_1210,N_1214);
nor U1263 (N_1263,N_1218,N_1206);
or U1264 (N_1264,N_1259,N_1241);
and U1265 (N_1265,N_1211,N_1212);
nand U1266 (N_1266,N_1237,N_1256);
nor U1267 (N_1267,N_1230,N_1227);
nand U1268 (N_1268,N_1207,N_1213);
and U1269 (N_1269,N_1231,N_1228);
nand U1270 (N_1270,N_1201,N_1222);
or U1271 (N_1271,N_1229,N_1217);
nand U1272 (N_1272,N_1203,N_1252);
xor U1273 (N_1273,N_1253,N_1238);
nor U1274 (N_1274,N_1245,N_1255);
nand U1275 (N_1275,N_1220,N_1205);
nor U1276 (N_1276,N_1258,N_1243);
and U1277 (N_1277,N_1254,N_1209);
nand U1278 (N_1278,N_1257,N_1226);
and U1279 (N_1279,N_1219,N_1204);
and U1280 (N_1280,N_1244,N_1248);
nor U1281 (N_1281,N_1235,N_1240);
nand U1282 (N_1282,N_1233,N_1223);
and U1283 (N_1283,N_1232,N_1224);
or U1284 (N_1284,N_1239,N_1202);
or U1285 (N_1285,N_1234,N_1250);
and U1286 (N_1286,N_1200,N_1246);
and U1287 (N_1287,N_1215,N_1208);
nor U1288 (N_1288,N_1236,N_1216);
or U1289 (N_1289,N_1221,N_1249);
nor U1290 (N_1290,N_1242,N_1238);
and U1291 (N_1291,N_1249,N_1219);
or U1292 (N_1292,N_1247,N_1238);
nor U1293 (N_1293,N_1247,N_1237);
and U1294 (N_1294,N_1252,N_1204);
nand U1295 (N_1295,N_1203,N_1213);
or U1296 (N_1296,N_1250,N_1239);
and U1297 (N_1297,N_1243,N_1241);
and U1298 (N_1298,N_1228,N_1222);
or U1299 (N_1299,N_1246,N_1224);
and U1300 (N_1300,N_1223,N_1243);
and U1301 (N_1301,N_1257,N_1216);
nand U1302 (N_1302,N_1240,N_1231);
nor U1303 (N_1303,N_1228,N_1201);
nand U1304 (N_1304,N_1216,N_1210);
and U1305 (N_1305,N_1254,N_1208);
nand U1306 (N_1306,N_1247,N_1209);
or U1307 (N_1307,N_1200,N_1215);
nor U1308 (N_1308,N_1202,N_1241);
nand U1309 (N_1309,N_1213,N_1243);
and U1310 (N_1310,N_1205,N_1212);
or U1311 (N_1311,N_1215,N_1213);
xnor U1312 (N_1312,N_1253,N_1202);
nand U1313 (N_1313,N_1234,N_1205);
or U1314 (N_1314,N_1242,N_1224);
nor U1315 (N_1315,N_1239,N_1235);
or U1316 (N_1316,N_1207,N_1254);
and U1317 (N_1317,N_1243,N_1239);
nand U1318 (N_1318,N_1257,N_1211);
nor U1319 (N_1319,N_1236,N_1214);
nor U1320 (N_1320,N_1306,N_1279);
or U1321 (N_1321,N_1318,N_1268);
or U1322 (N_1322,N_1276,N_1269);
and U1323 (N_1323,N_1287,N_1282);
nor U1324 (N_1324,N_1304,N_1274);
nand U1325 (N_1325,N_1280,N_1281);
or U1326 (N_1326,N_1292,N_1295);
nor U1327 (N_1327,N_1308,N_1266);
nor U1328 (N_1328,N_1293,N_1310);
or U1329 (N_1329,N_1264,N_1315);
and U1330 (N_1330,N_1297,N_1296);
and U1331 (N_1331,N_1286,N_1262);
and U1332 (N_1332,N_1271,N_1275);
nand U1333 (N_1333,N_1288,N_1284);
or U1334 (N_1334,N_1290,N_1300);
nor U1335 (N_1335,N_1313,N_1314);
nand U1336 (N_1336,N_1302,N_1311);
nor U1337 (N_1337,N_1270,N_1307);
or U1338 (N_1338,N_1283,N_1317);
nand U1339 (N_1339,N_1278,N_1265);
and U1340 (N_1340,N_1272,N_1298);
or U1341 (N_1341,N_1273,N_1291);
nor U1342 (N_1342,N_1299,N_1277);
and U1343 (N_1343,N_1316,N_1261);
nor U1344 (N_1344,N_1285,N_1305);
nor U1345 (N_1345,N_1263,N_1267);
or U1346 (N_1346,N_1312,N_1301);
nand U1347 (N_1347,N_1309,N_1260);
and U1348 (N_1348,N_1303,N_1289);
and U1349 (N_1349,N_1294,N_1319);
nand U1350 (N_1350,N_1281,N_1301);
xor U1351 (N_1351,N_1307,N_1263);
or U1352 (N_1352,N_1289,N_1319);
or U1353 (N_1353,N_1295,N_1310);
nor U1354 (N_1354,N_1294,N_1310);
and U1355 (N_1355,N_1316,N_1305);
or U1356 (N_1356,N_1288,N_1274);
nor U1357 (N_1357,N_1313,N_1289);
nor U1358 (N_1358,N_1278,N_1268);
or U1359 (N_1359,N_1280,N_1296);
xor U1360 (N_1360,N_1282,N_1264);
nand U1361 (N_1361,N_1278,N_1281);
or U1362 (N_1362,N_1288,N_1295);
or U1363 (N_1363,N_1261,N_1317);
and U1364 (N_1364,N_1262,N_1317);
nor U1365 (N_1365,N_1307,N_1261);
nor U1366 (N_1366,N_1270,N_1298);
nand U1367 (N_1367,N_1263,N_1275);
nor U1368 (N_1368,N_1274,N_1281);
nor U1369 (N_1369,N_1273,N_1299);
nand U1370 (N_1370,N_1276,N_1264);
or U1371 (N_1371,N_1299,N_1275);
xnor U1372 (N_1372,N_1310,N_1315);
or U1373 (N_1373,N_1282,N_1296);
or U1374 (N_1374,N_1260,N_1276);
nor U1375 (N_1375,N_1280,N_1287);
nor U1376 (N_1376,N_1264,N_1297);
and U1377 (N_1377,N_1267,N_1266);
and U1378 (N_1378,N_1295,N_1273);
nor U1379 (N_1379,N_1290,N_1263);
nand U1380 (N_1380,N_1331,N_1378);
and U1381 (N_1381,N_1348,N_1374);
nor U1382 (N_1382,N_1367,N_1340);
xnor U1383 (N_1383,N_1350,N_1328);
and U1384 (N_1384,N_1372,N_1351);
and U1385 (N_1385,N_1332,N_1342);
nand U1386 (N_1386,N_1346,N_1352);
or U1387 (N_1387,N_1344,N_1361);
or U1388 (N_1388,N_1324,N_1338);
nand U1389 (N_1389,N_1377,N_1336);
nand U1390 (N_1390,N_1371,N_1327);
nand U1391 (N_1391,N_1323,N_1376);
nand U1392 (N_1392,N_1356,N_1357);
or U1393 (N_1393,N_1370,N_1373);
and U1394 (N_1394,N_1362,N_1363);
and U1395 (N_1395,N_1321,N_1349);
and U1396 (N_1396,N_1320,N_1353);
nor U1397 (N_1397,N_1359,N_1347);
nand U1398 (N_1398,N_1379,N_1368);
nor U1399 (N_1399,N_1355,N_1341);
or U1400 (N_1400,N_1354,N_1358);
or U1401 (N_1401,N_1345,N_1329);
and U1402 (N_1402,N_1334,N_1337);
or U1403 (N_1403,N_1369,N_1326);
nand U1404 (N_1404,N_1325,N_1343);
or U1405 (N_1405,N_1360,N_1322);
and U1406 (N_1406,N_1364,N_1366);
nor U1407 (N_1407,N_1330,N_1365);
nand U1408 (N_1408,N_1339,N_1335);
nor U1409 (N_1409,N_1333,N_1375);
nand U1410 (N_1410,N_1342,N_1358);
and U1411 (N_1411,N_1350,N_1347);
and U1412 (N_1412,N_1338,N_1343);
or U1413 (N_1413,N_1368,N_1367);
nor U1414 (N_1414,N_1376,N_1343);
and U1415 (N_1415,N_1328,N_1359);
nor U1416 (N_1416,N_1343,N_1346);
nand U1417 (N_1417,N_1336,N_1320);
nand U1418 (N_1418,N_1326,N_1375);
nand U1419 (N_1419,N_1352,N_1323);
or U1420 (N_1420,N_1338,N_1327);
or U1421 (N_1421,N_1350,N_1353);
or U1422 (N_1422,N_1377,N_1362);
nor U1423 (N_1423,N_1324,N_1350);
or U1424 (N_1424,N_1332,N_1377);
or U1425 (N_1425,N_1356,N_1330);
and U1426 (N_1426,N_1326,N_1360);
nand U1427 (N_1427,N_1327,N_1322);
or U1428 (N_1428,N_1363,N_1342);
or U1429 (N_1429,N_1333,N_1378);
and U1430 (N_1430,N_1322,N_1338);
or U1431 (N_1431,N_1330,N_1354);
or U1432 (N_1432,N_1375,N_1360);
and U1433 (N_1433,N_1324,N_1374);
nor U1434 (N_1434,N_1343,N_1353);
nor U1435 (N_1435,N_1378,N_1347);
and U1436 (N_1436,N_1333,N_1328);
nor U1437 (N_1437,N_1352,N_1349);
nor U1438 (N_1438,N_1368,N_1365);
nand U1439 (N_1439,N_1356,N_1368);
or U1440 (N_1440,N_1415,N_1424);
nand U1441 (N_1441,N_1402,N_1388);
or U1442 (N_1442,N_1407,N_1417);
nand U1443 (N_1443,N_1389,N_1382);
nand U1444 (N_1444,N_1429,N_1400);
and U1445 (N_1445,N_1380,N_1408);
nand U1446 (N_1446,N_1398,N_1381);
or U1447 (N_1447,N_1426,N_1401);
nor U1448 (N_1448,N_1396,N_1385);
nor U1449 (N_1449,N_1437,N_1394);
nor U1450 (N_1450,N_1423,N_1416);
or U1451 (N_1451,N_1386,N_1436);
or U1452 (N_1452,N_1420,N_1390);
nor U1453 (N_1453,N_1410,N_1397);
nand U1454 (N_1454,N_1432,N_1418);
or U1455 (N_1455,N_1419,N_1431);
nor U1456 (N_1456,N_1412,N_1383);
and U1457 (N_1457,N_1406,N_1439);
nor U1458 (N_1458,N_1427,N_1422);
or U1459 (N_1459,N_1414,N_1399);
or U1460 (N_1460,N_1428,N_1413);
nor U1461 (N_1461,N_1404,N_1409);
nor U1462 (N_1462,N_1387,N_1430);
and U1463 (N_1463,N_1434,N_1435);
nor U1464 (N_1464,N_1392,N_1405);
nor U1465 (N_1465,N_1393,N_1403);
or U1466 (N_1466,N_1425,N_1391);
or U1467 (N_1467,N_1433,N_1395);
nand U1468 (N_1468,N_1411,N_1421);
nand U1469 (N_1469,N_1438,N_1384);
and U1470 (N_1470,N_1384,N_1404);
nand U1471 (N_1471,N_1407,N_1405);
or U1472 (N_1472,N_1431,N_1380);
nand U1473 (N_1473,N_1383,N_1416);
nor U1474 (N_1474,N_1435,N_1436);
nor U1475 (N_1475,N_1403,N_1386);
and U1476 (N_1476,N_1418,N_1388);
nor U1477 (N_1477,N_1435,N_1439);
or U1478 (N_1478,N_1413,N_1427);
nor U1479 (N_1479,N_1428,N_1430);
and U1480 (N_1480,N_1410,N_1382);
and U1481 (N_1481,N_1398,N_1394);
and U1482 (N_1482,N_1413,N_1439);
and U1483 (N_1483,N_1425,N_1436);
and U1484 (N_1484,N_1398,N_1401);
or U1485 (N_1485,N_1404,N_1433);
or U1486 (N_1486,N_1430,N_1424);
and U1487 (N_1487,N_1402,N_1430);
and U1488 (N_1488,N_1430,N_1434);
nand U1489 (N_1489,N_1417,N_1411);
nor U1490 (N_1490,N_1382,N_1438);
nand U1491 (N_1491,N_1385,N_1410);
nand U1492 (N_1492,N_1430,N_1410);
nand U1493 (N_1493,N_1425,N_1430);
nor U1494 (N_1494,N_1387,N_1417);
nor U1495 (N_1495,N_1396,N_1439);
nand U1496 (N_1496,N_1415,N_1418);
nand U1497 (N_1497,N_1433,N_1428);
or U1498 (N_1498,N_1408,N_1417);
or U1499 (N_1499,N_1426,N_1381);
and U1500 (N_1500,N_1480,N_1464);
and U1501 (N_1501,N_1499,N_1466);
or U1502 (N_1502,N_1484,N_1474);
nor U1503 (N_1503,N_1476,N_1463);
and U1504 (N_1504,N_1483,N_1446);
nand U1505 (N_1505,N_1485,N_1482);
xor U1506 (N_1506,N_1455,N_1481);
nor U1507 (N_1507,N_1487,N_1465);
nand U1508 (N_1508,N_1447,N_1461);
and U1509 (N_1509,N_1498,N_1450);
or U1510 (N_1510,N_1469,N_1452);
and U1511 (N_1511,N_1453,N_1468);
or U1512 (N_1512,N_1492,N_1491);
and U1513 (N_1513,N_1462,N_1471);
nand U1514 (N_1514,N_1490,N_1449);
and U1515 (N_1515,N_1493,N_1445);
nand U1516 (N_1516,N_1470,N_1472);
nand U1517 (N_1517,N_1495,N_1460);
or U1518 (N_1518,N_1441,N_1497);
xor U1519 (N_1519,N_1458,N_1477);
nor U1520 (N_1520,N_1475,N_1486);
or U1521 (N_1521,N_1440,N_1454);
nor U1522 (N_1522,N_1448,N_1473);
and U1523 (N_1523,N_1459,N_1479);
and U1524 (N_1524,N_1457,N_1443);
nor U1525 (N_1525,N_1456,N_1488);
nor U1526 (N_1526,N_1451,N_1478);
and U1527 (N_1527,N_1467,N_1496);
and U1528 (N_1528,N_1442,N_1489);
and U1529 (N_1529,N_1444,N_1494);
or U1530 (N_1530,N_1495,N_1494);
xor U1531 (N_1531,N_1485,N_1478);
or U1532 (N_1532,N_1495,N_1483);
and U1533 (N_1533,N_1490,N_1494);
nand U1534 (N_1534,N_1489,N_1460);
nor U1535 (N_1535,N_1461,N_1457);
nand U1536 (N_1536,N_1481,N_1471);
and U1537 (N_1537,N_1495,N_1453);
nor U1538 (N_1538,N_1478,N_1459);
or U1539 (N_1539,N_1495,N_1496);
nor U1540 (N_1540,N_1444,N_1465);
nand U1541 (N_1541,N_1497,N_1464);
or U1542 (N_1542,N_1487,N_1490);
and U1543 (N_1543,N_1484,N_1490);
or U1544 (N_1544,N_1474,N_1448);
nor U1545 (N_1545,N_1473,N_1440);
and U1546 (N_1546,N_1464,N_1481);
nand U1547 (N_1547,N_1445,N_1466);
and U1548 (N_1548,N_1471,N_1465);
or U1549 (N_1549,N_1492,N_1495);
nor U1550 (N_1550,N_1460,N_1496);
or U1551 (N_1551,N_1467,N_1492);
nand U1552 (N_1552,N_1456,N_1458);
or U1553 (N_1553,N_1459,N_1462);
and U1554 (N_1554,N_1491,N_1460);
or U1555 (N_1555,N_1485,N_1446);
and U1556 (N_1556,N_1447,N_1471);
nand U1557 (N_1557,N_1492,N_1446);
and U1558 (N_1558,N_1492,N_1472);
nand U1559 (N_1559,N_1456,N_1485);
and U1560 (N_1560,N_1523,N_1509);
nand U1561 (N_1561,N_1506,N_1557);
or U1562 (N_1562,N_1501,N_1518);
nand U1563 (N_1563,N_1548,N_1526);
and U1564 (N_1564,N_1534,N_1515);
or U1565 (N_1565,N_1552,N_1539);
and U1566 (N_1566,N_1528,N_1524);
or U1567 (N_1567,N_1502,N_1549);
or U1568 (N_1568,N_1540,N_1541);
nor U1569 (N_1569,N_1503,N_1521);
or U1570 (N_1570,N_1520,N_1538);
nand U1571 (N_1571,N_1510,N_1508);
and U1572 (N_1572,N_1533,N_1514);
nand U1573 (N_1573,N_1543,N_1529);
and U1574 (N_1574,N_1554,N_1542);
and U1575 (N_1575,N_1504,N_1556);
nand U1576 (N_1576,N_1550,N_1530);
and U1577 (N_1577,N_1559,N_1525);
and U1578 (N_1578,N_1507,N_1537);
or U1579 (N_1579,N_1546,N_1531);
nand U1580 (N_1580,N_1512,N_1536);
or U1581 (N_1581,N_1553,N_1547);
nor U1582 (N_1582,N_1517,N_1544);
and U1583 (N_1583,N_1500,N_1551);
nand U1584 (N_1584,N_1555,N_1545);
or U1585 (N_1585,N_1519,N_1513);
and U1586 (N_1586,N_1535,N_1522);
xor U1587 (N_1587,N_1516,N_1511);
or U1588 (N_1588,N_1527,N_1532);
nor U1589 (N_1589,N_1505,N_1558);
or U1590 (N_1590,N_1557,N_1544);
nor U1591 (N_1591,N_1531,N_1513);
nand U1592 (N_1592,N_1514,N_1515);
nand U1593 (N_1593,N_1556,N_1544);
nor U1594 (N_1594,N_1523,N_1535);
nor U1595 (N_1595,N_1538,N_1541);
or U1596 (N_1596,N_1557,N_1508);
and U1597 (N_1597,N_1518,N_1529);
nor U1598 (N_1598,N_1516,N_1536);
nor U1599 (N_1599,N_1541,N_1504);
and U1600 (N_1600,N_1537,N_1544);
nor U1601 (N_1601,N_1524,N_1536);
or U1602 (N_1602,N_1510,N_1542);
and U1603 (N_1603,N_1557,N_1547);
nor U1604 (N_1604,N_1525,N_1540);
xnor U1605 (N_1605,N_1539,N_1529);
or U1606 (N_1606,N_1520,N_1550);
and U1607 (N_1607,N_1546,N_1513);
or U1608 (N_1608,N_1506,N_1522);
or U1609 (N_1609,N_1532,N_1526);
and U1610 (N_1610,N_1532,N_1503);
and U1611 (N_1611,N_1528,N_1550);
or U1612 (N_1612,N_1529,N_1514);
and U1613 (N_1613,N_1557,N_1509);
xor U1614 (N_1614,N_1503,N_1543);
nand U1615 (N_1615,N_1543,N_1545);
nor U1616 (N_1616,N_1525,N_1531);
nor U1617 (N_1617,N_1545,N_1539);
or U1618 (N_1618,N_1516,N_1529);
nor U1619 (N_1619,N_1538,N_1546);
and U1620 (N_1620,N_1565,N_1568);
xnor U1621 (N_1621,N_1580,N_1594);
nand U1622 (N_1622,N_1613,N_1563);
nand U1623 (N_1623,N_1569,N_1598);
or U1624 (N_1624,N_1561,N_1618);
or U1625 (N_1625,N_1592,N_1577);
nand U1626 (N_1626,N_1583,N_1574);
nand U1627 (N_1627,N_1591,N_1570);
and U1628 (N_1628,N_1612,N_1560);
xor U1629 (N_1629,N_1584,N_1603);
and U1630 (N_1630,N_1599,N_1575);
nor U1631 (N_1631,N_1571,N_1595);
nand U1632 (N_1632,N_1601,N_1610);
and U1633 (N_1633,N_1578,N_1616);
nand U1634 (N_1634,N_1586,N_1576);
nand U1635 (N_1635,N_1581,N_1589);
or U1636 (N_1636,N_1608,N_1573);
and U1637 (N_1637,N_1604,N_1579);
and U1638 (N_1638,N_1602,N_1597);
nor U1639 (N_1639,N_1619,N_1572);
xor U1640 (N_1640,N_1611,N_1606);
nand U1641 (N_1641,N_1596,N_1587);
xor U1642 (N_1642,N_1590,N_1588);
nand U1643 (N_1643,N_1564,N_1605);
nor U1644 (N_1644,N_1607,N_1600);
and U1645 (N_1645,N_1566,N_1582);
nor U1646 (N_1646,N_1615,N_1585);
xnor U1647 (N_1647,N_1614,N_1562);
nand U1648 (N_1648,N_1617,N_1567);
nand U1649 (N_1649,N_1593,N_1609);
nand U1650 (N_1650,N_1600,N_1596);
or U1651 (N_1651,N_1594,N_1618);
nand U1652 (N_1652,N_1569,N_1603);
nor U1653 (N_1653,N_1604,N_1581);
and U1654 (N_1654,N_1578,N_1603);
or U1655 (N_1655,N_1589,N_1596);
nor U1656 (N_1656,N_1609,N_1570);
nand U1657 (N_1657,N_1563,N_1566);
and U1658 (N_1658,N_1597,N_1589);
or U1659 (N_1659,N_1575,N_1595);
or U1660 (N_1660,N_1608,N_1598);
nand U1661 (N_1661,N_1607,N_1580);
and U1662 (N_1662,N_1577,N_1609);
nand U1663 (N_1663,N_1615,N_1571);
nor U1664 (N_1664,N_1569,N_1571);
nor U1665 (N_1665,N_1595,N_1600);
nand U1666 (N_1666,N_1575,N_1571);
and U1667 (N_1667,N_1573,N_1565);
nand U1668 (N_1668,N_1596,N_1608);
and U1669 (N_1669,N_1602,N_1603);
or U1670 (N_1670,N_1598,N_1592);
or U1671 (N_1671,N_1563,N_1579);
nor U1672 (N_1672,N_1605,N_1603);
nand U1673 (N_1673,N_1572,N_1585);
and U1674 (N_1674,N_1613,N_1584);
nor U1675 (N_1675,N_1599,N_1582);
or U1676 (N_1676,N_1591,N_1585);
and U1677 (N_1677,N_1612,N_1583);
nor U1678 (N_1678,N_1597,N_1596);
or U1679 (N_1679,N_1608,N_1592);
or U1680 (N_1680,N_1658,N_1634);
or U1681 (N_1681,N_1676,N_1630);
nor U1682 (N_1682,N_1672,N_1649);
xnor U1683 (N_1683,N_1660,N_1663);
or U1684 (N_1684,N_1656,N_1640);
nor U1685 (N_1685,N_1670,N_1641);
and U1686 (N_1686,N_1645,N_1621);
nand U1687 (N_1687,N_1624,N_1625);
and U1688 (N_1688,N_1642,N_1638);
nor U1689 (N_1689,N_1647,N_1654);
and U1690 (N_1690,N_1653,N_1666);
or U1691 (N_1691,N_1651,N_1655);
nand U1692 (N_1692,N_1673,N_1678);
and U1693 (N_1693,N_1648,N_1644);
nor U1694 (N_1694,N_1646,N_1629);
nor U1695 (N_1695,N_1677,N_1620);
or U1696 (N_1696,N_1650,N_1659);
and U1697 (N_1697,N_1633,N_1665);
or U1698 (N_1698,N_1622,N_1662);
or U1699 (N_1699,N_1628,N_1632);
nor U1700 (N_1700,N_1627,N_1679);
and U1701 (N_1701,N_1635,N_1664);
or U1702 (N_1702,N_1675,N_1626);
and U1703 (N_1703,N_1668,N_1639);
nand U1704 (N_1704,N_1657,N_1669);
nand U1705 (N_1705,N_1623,N_1652);
nor U1706 (N_1706,N_1636,N_1674);
nor U1707 (N_1707,N_1667,N_1637);
nand U1708 (N_1708,N_1631,N_1643);
nor U1709 (N_1709,N_1671,N_1661);
and U1710 (N_1710,N_1660,N_1652);
nor U1711 (N_1711,N_1642,N_1678);
nor U1712 (N_1712,N_1632,N_1642);
nor U1713 (N_1713,N_1674,N_1655);
nor U1714 (N_1714,N_1670,N_1629);
and U1715 (N_1715,N_1645,N_1663);
and U1716 (N_1716,N_1673,N_1665);
nand U1717 (N_1717,N_1631,N_1627);
nor U1718 (N_1718,N_1651,N_1654);
nor U1719 (N_1719,N_1631,N_1678);
or U1720 (N_1720,N_1658,N_1672);
or U1721 (N_1721,N_1653,N_1672);
nor U1722 (N_1722,N_1625,N_1627);
nor U1723 (N_1723,N_1641,N_1647);
or U1724 (N_1724,N_1634,N_1674);
and U1725 (N_1725,N_1665,N_1635);
nor U1726 (N_1726,N_1643,N_1646);
nand U1727 (N_1727,N_1649,N_1630);
or U1728 (N_1728,N_1636,N_1651);
nor U1729 (N_1729,N_1626,N_1673);
and U1730 (N_1730,N_1678,N_1647);
or U1731 (N_1731,N_1669,N_1651);
and U1732 (N_1732,N_1672,N_1648);
nand U1733 (N_1733,N_1630,N_1635);
xor U1734 (N_1734,N_1652,N_1653);
nor U1735 (N_1735,N_1649,N_1636);
nand U1736 (N_1736,N_1661,N_1627);
xor U1737 (N_1737,N_1655,N_1633);
nand U1738 (N_1738,N_1621,N_1649);
nand U1739 (N_1739,N_1671,N_1626);
nor U1740 (N_1740,N_1719,N_1709);
or U1741 (N_1741,N_1701,N_1697);
or U1742 (N_1742,N_1703,N_1689);
or U1743 (N_1743,N_1708,N_1711);
or U1744 (N_1744,N_1698,N_1684);
nand U1745 (N_1745,N_1725,N_1715);
nor U1746 (N_1746,N_1736,N_1735);
nor U1747 (N_1747,N_1718,N_1724);
nand U1748 (N_1748,N_1693,N_1681);
or U1749 (N_1749,N_1702,N_1730);
nor U1750 (N_1750,N_1721,N_1717);
or U1751 (N_1751,N_1733,N_1731);
or U1752 (N_1752,N_1699,N_1696);
nand U1753 (N_1753,N_1683,N_1707);
nor U1754 (N_1754,N_1704,N_1714);
nor U1755 (N_1755,N_1726,N_1706);
nand U1756 (N_1756,N_1720,N_1738);
or U1757 (N_1757,N_1685,N_1692);
nand U1758 (N_1758,N_1729,N_1728);
nand U1759 (N_1759,N_1710,N_1727);
nand U1760 (N_1760,N_1737,N_1687);
nand U1761 (N_1761,N_1680,N_1723);
or U1762 (N_1762,N_1688,N_1734);
and U1763 (N_1763,N_1722,N_1691);
or U1764 (N_1764,N_1712,N_1739);
and U1765 (N_1765,N_1690,N_1716);
nand U1766 (N_1766,N_1694,N_1686);
nor U1767 (N_1767,N_1695,N_1700);
and U1768 (N_1768,N_1732,N_1713);
nand U1769 (N_1769,N_1682,N_1705);
nor U1770 (N_1770,N_1709,N_1731);
nand U1771 (N_1771,N_1711,N_1687);
xor U1772 (N_1772,N_1703,N_1714);
or U1773 (N_1773,N_1715,N_1686);
nand U1774 (N_1774,N_1685,N_1693);
or U1775 (N_1775,N_1713,N_1705);
nor U1776 (N_1776,N_1719,N_1698);
and U1777 (N_1777,N_1704,N_1683);
nand U1778 (N_1778,N_1726,N_1725);
or U1779 (N_1779,N_1735,N_1680);
and U1780 (N_1780,N_1712,N_1711);
or U1781 (N_1781,N_1682,N_1700);
or U1782 (N_1782,N_1721,N_1735);
xnor U1783 (N_1783,N_1736,N_1730);
nand U1784 (N_1784,N_1703,N_1736);
or U1785 (N_1785,N_1693,N_1691);
nand U1786 (N_1786,N_1682,N_1707);
or U1787 (N_1787,N_1729,N_1730);
and U1788 (N_1788,N_1700,N_1722);
nor U1789 (N_1789,N_1738,N_1703);
or U1790 (N_1790,N_1705,N_1703);
nand U1791 (N_1791,N_1680,N_1703);
nand U1792 (N_1792,N_1694,N_1681);
nand U1793 (N_1793,N_1714,N_1686);
and U1794 (N_1794,N_1727,N_1720);
nor U1795 (N_1795,N_1715,N_1731);
nor U1796 (N_1796,N_1719,N_1728);
and U1797 (N_1797,N_1711,N_1709);
or U1798 (N_1798,N_1738,N_1704);
nor U1799 (N_1799,N_1727,N_1738);
nor U1800 (N_1800,N_1771,N_1795);
or U1801 (N_1801,N_1749,N_1748);
or U1802 (N_1802,N_1783,N_1785);
nor U1803 (N_1803,N_1753,N_1798);
nor U1804 (N_1804,N_1769,N_1786);
or U1805 (N_1805,N_1752,N_1767);
and U1806 (N_1806,N_1746,N_1772);
nand U1807 (N_1807,N_1778,N_1759);
nor U1808 (N_1808,N_1776,N_1747);
and U1809 (N_1809,N_1773,N_1763);
and U1810 (N_1810,N_1794,N_1789);
or U1811 (N_1811,N_1770,N_1775);
and U1812 (N_1812,N_1788,N_1755);
nand U1813 (N_1813,N_1741,N_1762);
and U1814 (N_1814,N_1782,N_1745);
nand U1815 (N_1815,N_1779,N_1796);
nor U1816 (N_1816,N_1765,N_1781);
nand U1817 (N_1817,N_1792,N_1784);
nand U1818 (N_1818,N_1761,N_1757);
or U1819 (N_1819,N_1793,N_1768);
nor U1820 (N_1820,N_1780,N_1787);
nor U1821 (N_1821,N_1742,N_1774);
nand U1822 (N_1822,N_1766,N_1799);
nor U1823 (N_1823,N_1743,N_1764);
nor U1824 (N_1824,N_1754,N_1740);
or U1825 (N_1825,N_1744,N_1777);
and U1826 (N_1826,N_1751,N_1791);
nor U1827 (N_1827,N_1756,N_1760);
nor U1828 (N_1828,N_1797,N_1750);
nor U1829 (N_1829,N_1790,N_1758);
nor U1830 (N_1830,N_1799,N_1748);
nor U1831 (N_1831,N_1796,N_1751);
and U1832 (N_1832,N_1751,N_1785);
nor U1833 (N_1833,N_1748,N_1774);
or U1834 (N_1834,N_1781,N_1746);
nand U1835 (N_1835,N_1790,N_1757);
nand U1836 (N_1836,N_1761,N_1785);
nand U1837 (N_1837,N_1756,N_1787);
nand U1838 (N_1838,N_1760,N_1753);
and U1839 (N_1839,N_1753,N_1774);
nand U1840 (N_1840,N_1787,N_1786);
or U1841 (N_1841,N_1763,N_1749);
and U1842 (N_1842,N_1784,N_1766);
nor U1843 (N_1843,N_1754,N_1771);
nand U1844 (N_1844,N_1753,N_1746);
and U1845 (N_1845,N_1752,N_1749);
or U1846 (N_1846,N_1767,N_1759);
or U1847 (N_1847,N_1793,N_1752);
nand U1848 (N_1848,N_1757,N_1760);
or U1849 (N_1849,N_1756,N_1789);
and U1850 (N_1850,N_1792,N_1775);
nand U1851 (N_1851,N_1799,N_1765);
and U1852 (N_1852,N_1749,N_1742);
nor U1853 (N_1853,N_1749,N_1751);
and U1854 (N_1854,N_1776,N_1785);
or U1855 (N_1855,N_1768,N_1745);
or U1856 (N_1856,N_1754,N_1784);
nand U1857 (N_1857,N_1771,N_1748);
nor U1858 (N_1858,N_1745,N_1793);
nor U1859 (N_1859,N_1740,N_1798);
and U1860 (N_1860,N_1842,N_1804);
or U1861 (N_1861,N_1809,N_1845);
and U1862 (N_1862,N_1846,N_1822);
and U1863 (N_1863,N_1813,N_1853);
and U1864 (N_1864,N_1816,N_1837);
or U1865 (N_1865,N_1856,N_1851);
xnor U1866 (N_1866,N_1859,N_1818);
xor U1867 (N_1867,N_1811,N_1849);
nand U1868 (N_1868,N_1828,N_1805);
nand U1869 (N_1869,N_1826,N_1810);
nor U1870 (N_1870,N_1802,N_1834);
nor U1871 (N_1871,N_1807,N_1850);
or U1872 (N_1872,N_1835,N_1803);
and U1873 (N_1873,N_1825,N_1857);
xnor U1874 (N_1874,N_1824,N_1831);
nand U1875 (N_1875,N_1847,N_1823);
and U1876 (N_1876,N_1821,N_1800);
nor U1877 (N_1877,N_1830,N_1815);
and U1878 (N_1878,N_1836,N_1801);
nand U1879 (N_1879,N_1827,N_1812);
nor U1880 (N_1880,N_1817,N_1841);
and U1881 (N_1881,N_1852,N_1839);
nor U1882 (N_1882,N_1858,N_1848);
or U1883 (N_1883,N_1854,N_1806);
nand U1884 (N_1884,N_1838,N_1829);
nor U1885 (N_1885,N_1808,N_1840);
and U1886 (N_1886,N_1814,N_1844);
nor U1887 (N_1887,N_1820,N_1833);
or U1888 (N_1888,N_1832,N_1855);
nor U1889 (N_1889,N_1843,N_1819);
nor U1890 (N_1890,N_1817,N_1819);
or U1891 (N_1891,N_1856,N_1850);
or U1892 (N_1892,N_1800,N_1811);
nand U1893 (N_1893,N_1812,N_1845);
nand U1894 (N_1894,N_1807,N_1840);
nand U1895 (N_1895,N_1824,N_1812);
and U1896 (N_1896,N_1831,N_1828);
nor U1897 (N_1897,N_1813,N_1802);
nand U1898 (N_1898,N_1830,N_1808);
or U1899 (N_1899,N_1814,N_1843);
and U1900 (N_1900,N_1816,N_1850);
nor U1901 (N_1901,N_1844,N_1832);
nand U1902 (N_1902,N_1834,N_1852);
nand U1903 (N_1903,N_1853,N_1828);
nor U1904 (N_1904,N_1813,N_1846);
nand U1905 (N_1905,N_1800,N_1803);
nand U1906 (N_1906,N_1837,N_1826);
nor U1907 (N_1907,N_1856,N_1811);
nand U1908 (N_1908,N_1858,N_1841);
or U1909 (N_1909,N_1801,N_1826);
nor U1910 (N_1910,N_1818,N_1819);
and U1911 (N_1911,N_1855,N_1851);
nor U1912 (N_1912,N_1848,N_1856);
nand U1913 (N_1913,N_1810,N_1815);
nor U1914 (N_1914,N_1806,N_1819);
nor U1915 (N_1915,N_1851,N_1827);
or U1916 (N_1916,N_1846,N_1845);
nor U1917 (N_1917,N_1809,N_1847);
or U1918 (N_1918,N_1808,N_1805);
nor U1919 (N_1919,N_1803,N_1852);
xnor U1920 (N_1920,N_1891,N_1910);
and U1921 (N_1921,N_1879,N_1900);
or U1922 (N_1922,N_1911,N_1897);
and U1923 (N_1923,N_1861,N_1906);
nor U1924 (N_1924,N_1881,N_1864);
nand U1925 (N_1925,N_1901,N_1874);
or U1926 (N_1926,N_1903,N_1880);
and U1927 (N_1927,N_1902,N_1894);
nand U1928 (N_1928,N_1913,N_1918);
and U1929 (N_1929,N_1919,N_1865);
nand U1930 (N_1930,N_1871,N_1899);
and U1931 (N_1931,N_1863,N_1895);
and U1932 (N_1932,N_1883,N_1915);
nor U1933 (N_1933,N_1905,N_1917);
nand U1934 (N_1934,N_1892,N_1882);
nor U1935 (N_1935,N_1870,N_1908);
nor U1936 (N_1936,N_1878,N_1896);
nor U1937 (N_1937,N_1890,N_1862);
and U1938 (N_1938,N_1886,N_1914);
and U1939 (N_1939,N_1909,N_1876);
and U1940 (N_1940,N_1887,N_1867);
and U1941 (N_1941,N_1866,N_1868);
and U1942 (N_1942,N_1872,N_1873);
or U1943 (N_1943,N_1898,N_1875);
nor U1944 (N_1944,N_1904,N_1884);
nand U1945 (N_1945,N_1885,N_1907);
and U1946 (N_1946,N_1860,N_1912);
xnor U1947 (N_1947,N_1877,N_1888);
and U1948 (N_1948,N_1893,N_1889);
and U1949 (N_1949,N_1916,N_1869);
nand U1950 (N_1950,N_1908,N_1901);
or U1951 (N_1951,N_1904,N_1877);
nor U1952 (N_1952,N_1873,N_1880);
nand U1953 (N_1953,N_1900,N_1902);
and U1954 (N_1954,N_1887,N_1912);
and U1955 (N_1955,N_1874,N_1897);
or U1956 (N_1956,N_1910,N_1906);
nor U1957 (N_1957,N_1892,N_1897);
and U1958 (N_1958,N_1900,N_1880);
nor U1959 (N_1959,N_1870,N_1873);
or U1960 (N_1960,N_1899,N_1917);
or U1961 (N_1961,N_1876,N_1880);
and U1962 (N_1962,N_1904,N_1882);
and U1963 (N_1963,N_1865,N_1862);
nand U1964 (N_1964,N_1898,N_1895);
or U1965 (N_1965,N_1897,N_1888);
nor U1966 (N_1966,N_1888,N_1913);
and U1967 (N_1967,N_1861,N_1895);
nor U1968 (N_1968,N_1903,N_1889);
xnor U1969 (N_1969,N_1884,N_1911);
nand U1970 (N_1970,N_1902,N_1896);
nand U1971 (N_1971,N_1907,N_1883);
nor U1972 (N_1972,N_1917,N_1864);
and U1973 (N_1973,N_1913,N_1861);
or U1974 (N_1974,N_1863,N_1881);
and U1975 (N_1975,N_1907,N_1910);
or U1976 (N_1976,N_1875,N_1887);
or U1977 (N_1977,N_1894,N_1868);
nor U1978 (N_1978,N_1892,N_1910);
and U1979 (N_1979,N_1885,N_1891);
or U1980 (N_1980,N_1941,N_1961);
nor U1981 (N_1981,N_1956,N_1959);
nor U1982 (N_1982,N_1923,N_1927);
and U1983 (N_1983,N_1924,N_1973);
and U1984 (N_1984,N_1943,N_1975);
nand U1985 (N_1985,N_1921,N_1949);
and U1986 (N_1986,N_1979,N_1965);
nor U1987 (N_1987,N_1969,N_1958);
xnor U1988 (N_1988,N_1948,N_1942);
nand U1989 (N_1989,N_1955,N_1947);
or U1990 (N_1990,N_1929,N_1944);
or U1991 (N_1991,N_1954,N_1926);
nor U1992 (N_1992,N_1936,N_1974);
nor U1993 (N_1993,N_1930,N_1952);
nor U1994 (N_1994,N_1967,N_1968);
and U1995 (N_1995,N_1938,N_1920);
and U1996 (N_1996,N_1957,N_1928);
and U1997 (N_1997,N_1922,N_1951);
nor U1998 (N_1998,N_1953,N_1939);
or U1999 (N_1999,N_1972,N_1925);
nor U2000 (N_2000,N_1978,N_1962);
nor U2001 (N_2001,N_1937,N_1977);
nor U2002 (N_2002,N_1960,N_1950);
or U2003 (N_2003,N_1976,N_1940);
and U2004 (N_2004,N_1964,N_1933);
nor U2005 (N_2005,N_1932,N_1963);
nand U2006 (N_2006,N_1934,N_1945);
and U2007 (N_2007,N_1946,N_1966);
nor U2008 (N_2008,N_1935,N_1970);
or U2009 (N_2009,N_1931,N_1971);
nand U2010 (N_2010,N_1960,N_1929);
nor U2011 (N_2011,N_1958,N_1967);
and U2012 (N_2012,N_1960,N_1976);
nor U2013 (N_2013,N_1923,N_1968);
or U2014 (N_2014,N_1940,N_1920);
and U2015 (N_2015,N_1940,N_1954);
or U2016 (N_2016,N_1949,N_1939);
nand U2017 (N_2017,N_1961,N_1950);
nor U2018 (N_2018,N_1937,N_1951);
or U2019 (N_2019,N_1948,N_1952);
and U2020 (N_2020,N_1975,N_1963);
nor U2021 (N_2021,N_1927,N_1955);
and U2022 (N_2022,N_1927,N_1924);
and U2023 (N_2023,N_1957,N_1923);
and U2024 (N_2024,N_1932,N_1943);
nor U2025 (N_2025,N_1971,N_1936);
and U2026 (N_2026,N_1935,N_1943);
nand U2027 (N_2027,N_1924,N_1955);
and U2028 (N_2028,N_1959,N_1941);
and U2029 (N_2029,N_1932,N_1927);
or U2030 (N_2030,N_1925,N_1927);
and U2031 (N_2031,N_1942,N_1960);
or U2032 (N_2032,N_1975,N_1922);
nand U2033 (N_2033,N_1976,N_1945);
or U2034 (N_2034,N_1930,N_1924);
nor U2035 (N_2035,N_1965,N_1936);
or U2036 (N_2036,N_1970,N_1965);
nor U2037 (N_2037,N_1926,N_1956);
and U2038 (N_2038,N_1943,N_1956);
and U2039 (N_2039,N_1934,N_1972);
nand U2040 (N_2040,N_2015,N_1985);
and U2041 (N_2041,N_2035,N_2033);
or U2042 (N_2042,N_2001,N_2012);
or U2043 (N_2043,N_2026,N_2021);
and U2044 (N_2044,N_2027,N_2007);
nor U2045 (N_2045,N_2011,N_2023);
or U2046 (N_2046,N_2019,N_2022);
and U2047 (N_2047,N_2031,N_2002);
nor U2048 (N_2048,N_2013,N_2030);
and U2049 (N_2049,N_2024,N_1989);
nand U2050 (N_2050,N_2032,N_1983);
nor U2051 (N_2051,N_1994,N_1984);
nand U2052 (N_2052,N_2034,N_2008);
nand U2053 (N_2053,N_2004,N_2039);
nor U2054 (N_2054,N_2028,N_2006);
or U2055 (N_2055,N_2005,N_2017);
nand U2056 (N_2056,N_2009,N_1995);
nor U2057 (N_2057,N_1997,N_1993);
nor U2058 (N_2058,N_1999,N_2016);
or U2059 (N_2059,N_1986,N_1980);
or U2060 (N_2060,N_1996,N_1987);
nor U2061 (N_2061,N_2020,N_2000);
nor U2062 (N_2062,N_2018,N_1990);
nand U2063 (N_2063,N_1998,N_1988);
and U2064 (N_2064,N_2036,N_2037);
nor U2065 (N_2065,N_2014,N_2029);
nand U2066 (N_2066,N_2003,N_2025);
nor U2067 (N_2067,N_1992,N_1982);
nand U2068 (N_2068,N_1981,N_1991);
or U2069 (N_2069,N_2010,N_2038);
and U2070 (N_2070,N_2004,N_2029);
nor U2071 (N_2071,N_1993,N_2010);
and U2072 (N_2072,N_1982,N_2017);
or U2073 (N_2073,N_2004,N_1998);
nand U2074 (N_2074,N_2022,N_2030);
and U2075 (N_2075,N_2022,N_2029);
nand U2076 (N_2076,N_2001,N_2011);
and U2077 (N_2077,N_2009,N_2037);
xnor U2078 (N_2078,N_1989,N_1984);
nor U2079 (N_2079,N_2013,N_1989);
or U2080 (N_2080,N_2002,N_2020);
nand U2081 (N_2081,N_2009,N_2031);
nand U2082 (N_2082,N_2015,N_2023);
nor U2083 (N_2083,N_2016,N_2015);
and U2084 (N_2084,N_1998,N_1987);
nand U2085 (N_2085,N_2025,N_2024);
and U2086 (N_2086,N_2008,N_2002);
nand U2087 (N_2087,N_2020,N_2027);
nor U2088 (N_2088,N_2026,N_2038);
or U2089 (N_2089,N_1989,N_1996);
and U2090 (N_2090,N_1991,N_2036);
or U2091 (N_2091,N_1989,N_1998);
nor U2092 (N_2092,N_2001,N_2029);
nand U2093 (N_2093,N_2027,N_1997);
nand U2094 (N_2094,N_1992,N_2021);
nor U2095 (N_2095,N_2034,N_2004);
nor U2096 (N_2096,N_2036,N_2025);
or U2097 (N_2097,N_2033,N_2034);
and U2098 (N_2098,N_1980,N_2038);
or U2099 (N_2099,N_2038,N_2005);
xnor U2100 (N_2100,N_2047,N_2096);
nand U2101 (N_2101,N_2046,N_2055);
or U2102 (N_2102,N_2050,N_2075);
and U2103 (N_2103,N_2097,N_2071);
or U2104 (N_2104,N_2056,N_2092);
nand U2105 (N_2105,N_2067,N_2044);
and U2106 (N_2106,N_2090,N_2041);
or U2107 (N_2107,N_2085,N_2065);
or U2108 (N_2108,N_2070,N_2045);
nor U2109 (N_2109,N_2077,N_2066);
or U2110 (N_2110,N_2072,N_2087);
nand U2111 (N_2111,N_2080,N_2076);
and U2112 (N_2112,N_2063,N_2064);
nand U2113 (N_2113,N_2051,N_2083);
or U2114 (N_2114,N_2082,N_2068);
and U2115 (N_2115,N_2089,N_2052);
or U2116 (N_2116,N_2048,N_2084);
nand U2117 (N_2117,N_2078,N_2074);
nor U2118 (N_2118,N_2053,N_2093);
or U2119 (N_2119,N_2086,N_2054);
nand U2120 (N_2120,N_2091,N_2094);
and U2121 (N_2121,N_2057,N_2060);
nor U2122 (N_2122,N_2040,N_2058);
and U2123 (N_2123,N_2098,N_2059);
nand U2124 (N_2124,N_2099,N_2073);
nand U2125 (N_2125,N_2079,N_2043);
or U2126 (N_2126,N_2081,N_2061);
or U2127 (N_2127,N_2042,N_2088);
and U2128 (N_2128,N_2049,N_2062);
nor U2129 (N_2129,N_2069,N_2095);
nor U2130 (N_2130,N_2097,N_2057);
and U2131 (N_2131,N_2088,N_2044);
or U2132 (N_2132,N_2054,N_2050);
nand U2133 (N_2133,N_2069,N_2055);
nor U2134 (N_2134,N_2089,N_2079);
nand U2135 (N_2135,N_2053,N_2083);
and U2136 (N_2136,N_2045,N_2091);
nand U2137 (N_2137,N_2093,N_2076);
nor U2138 (N_2138,N_2088,N_2043);
nor U2139 (N_2139,N_2074,N_2097);
nor U2140 (N_2140,N_2092,N_2040);
nand U2141 (N_2141,N_2060,N_2096);
or U2142 (N_2142,N_2068,N_2044);
nor U2143 (N_2143,N_2074,N_2073);
nand U2144 (N_2144,N_2062,N_2084);
nand U2145 (N_2145,N_2082,N_2089);
nor U2146 (N_2146,N_2073,N_2055);
or U2147 (N_2147,N_2041,N_2042);
or U2148 (N_2148,N_2066,N_2060);
nor U2149 (N_2149,N_2079,N_2047);
or U2150 (N_2150,N_2041,N_2070);
and U2151 (N_2151,N_2054,N_2078);
nor U2152 (N_2152,N_2087,N_2044);
nand U2153 (N_2153,N_2069,N_2056);
nand U2154 (N_2154,N_2052,N_2057);
nor U2155 (N_2155,N_2060,N_2043);
nand U2156 (N_2156,N_2088,N_2053);
nor U2157 (N_2157,N_2069,N_2099);
nand U2158 (N_2158,N_2071,N_2079);
nor U2159 (N_2159,N_2071,N_2083);
nor U2160 (N_2160,N_2123,N_2113);
nand U2161 (N_2161,N_2150,N_2153);
or U2162 (N_2162,N_2151,N_2116);
nor U2163 (N_2163,N_2112,N_2146);
nand U2164 (N_2164,N_2125,N_2136);
nor U2165 (N_2165,N_2140,N_2114);
nor U2166 (N_2166,N_2156,N_2159);
nor U2167 (N_2167,N_2120,N_2135);
or U2168 (N_2168,N_2128,N_2148);
nor U2169 (N_2169,N_2131,N_2122);
nor U2170 (N_2170,N_2115,N_2145);
and U2171 (N_2171,N_2105,N_2100);
and U2172 (N_2172,N_2138,N_2134);
nand U2173 (N_2173,N_2139,N_2101);
nor U2174 (N_2174,N_2118,N_2137);
or U2175 (N_2175,N_2152,N_2154);
nor U2176 (N_2176,N_2132,N_2109);
and U2177 (N_2177,N_2157,N_2144);
nand U2178 (N_2178,N_2141,N_2127);
nand U2179 (N_2179,N_2158,N_2133);
and U2180 (N_2180,N_2119,N_2155);
and U2181 (N_2181,N_2111,N_2129);
and U2182 (N_2182,N_2126,N_2142);
nor U2183 (N_2183,N_2147,N_2143);
nor U2184 (N_2184,N_2117,N_2130);
or U2185 (N_2185,N_2102,N_2121);
and U2186 (N_2186,N_2108,N_2103);
or U2187 (N_2187,N_2104,N_2110);
nor U2188 (N_2188,N_2107,N_2124);
nand U2189 (N_2189,N_2106,N_2149);
and U2190 (N_2190,N_2113,N_2101);
nand U2191 (N_2191,N_2128,N_2103);
nor U2192 (N_2192,N_2103,N_2141);
nand U2193 (N_2193,N_2128,N_2121);
or U2194 (N_2194,N_2142,N_2146);
nand U2195 (N_2195,N_2152,N_2141);
and U2196 (N_2196,N_2124,N_2125);
and U2197 (N_2197,N_2137,N_2112);
nand U2198 (N_2198,N_2159,N_2106);
xnor U2199 (N_2199,N_2157,N_2107);
nand U2200 (N_2200,N_2111,N_2105);
nor U2201 (N_2201,N_2146,N_2133);
and U2202 (N_2202,N_2104,N_2148);
or U2203 (N_2203,N_2121,N_2110);
or U2204 (N_2204,N_2101,N_2151);
nor U2205 (N_2205,N_2138,N_2104);
xor U2206 (N_2206,N_2153,N_2154);
nor U2207 (N_2207,N_2114,N_2144);
nand U2208 (N_2208,N_2145,N_2125);
nand U2209 (N_2209,N_2110,N_2126);
nand U2210 (N_2210,N_2101,N_2100);
and U2211 (N_2211,N_2109,N_2103);
nor U2212 (N_2212,N_2155,N_2124);
nor U2213 (N_2213,N_2115,N_2148);
nor U2214 (N_2214,N_2126,N_2146);
nand U2215 (N_2215,N_2140,N_2135);
or U2216 (N_2216,N_2101,N_2153);
nor U2217 (N_2217,N_2130,N_2147);
and U2218 (N_2218,N_2102,N_2142);
and U2219 (N_2219,N_2127,N_2136);
and U2220 (N_2220,N_2210,N_2161);
nand U2221 (N_2221,N_2182,N_2201);
nand U2222 (N_2222,N_2217,N_2171);
or U2223 (N_2223,N_2183,N_2199);
and U2224 (N_2224,N_2191,N_2186);
and U2225 (N_2225,N_2170,N_2196);
nand U2226 (N_2226,N_2185,N_2179);
and U2227 (N_2227,N_2180,N_2169);
and U2228 (N_2228,N_2218,N_2193);
or U2229 (N_2229,N_2187,N_2173);
or U2230 (N_2230,N_2176,N_2162);
and U2231 (N_2231,N_2163,N_2197);
nand U2232 (N_2232,N_2211,N_2209);
nand U2233 (N_2233,N_2160,N_2216);
nand U2234 (N_2234,N_2204,N_2203);
or U2235 (N_2235,N_2181,N_2190);
nand U2236 (N_2236,N_2166,N_2205);
nor U2237 (N_2237,N_2215,N_2178);
or U2238 (N_2238,N_2172,N_2206);
nor U2239 (N_2239,N_2207,N_2189);
nand U2240 (N_2240,N_2200,N_2175);
or U2241 (N_2241,N_2164,N_2192);
nor U2242 (N_2242,N_2202,N_2184);
xnor U2243 (N_2243,N_2167,N_2213);
nand U2244 (N_2244,N_2195,N_2165);
and U2245 (N_2245,N_2212,N_2188);
nand U2246 (N_2246,N_2174,N_2208);
nand U2247 (N_2247,N_2198,N_2168);
nand U2248 (N_2248,N_2219,N_2177);
and U2249 (N_2249,N_2194,N_2214);
nand U2250 (N_2250,N_2176,N_2182);
or U2251 (N_2251,N_2218,N_2179);
or U2252 (N_2252,N_2169,N_2200);
nor U2253 (N_2253,N_2196,N_2193);
nor U2254 (N_2254,N_2188,N_2192);
or U2255 (N_2255,N_2197,N_2170);
nor U2256 (N_2256,N_2197,N_2191);
nor U2257 (N_2257,N_2217,N_2191);
nor U2258 (N_2258,N_2183,N_2204);
nor U2259 (N_2259,N_2192,N_2219);
nor U2260 (N_2260,N_2200,N_2201);
nand U2261 (N_2261,N_2213,N_2207);
or U2262 (N_2262,N_2176,N_2202);
and U2263 (N_2263,N_2185,N_2181);
and U2264 (N_2264,N_2197,N_2171);
nand U2265 (N_2265,N_2184,N_2218);
nand U2266 (N_2266,N_2163,N_2194);
nor U2267 (N_2267,N_2193,N_2177);
xnor U2268 (N_2268,N_2209,N_2207);
and U2269 (N_2269,N_2195,N_2188);
nor U2270 (N_2270,N_2211,N_2180);
nor U2271 (N_2271,N_2197,N_2211);
and U2272 (N_2272,N_2162,N_2214);
nor U2273 (N_2273,N_2199,N_2193);
or U2274 (N_2274,N_2184,N_2193);
or U2275 (N_2275,N_2164,N_2211);
and U2276 (N_2276,N_2161,N_2180);
xnor U2277 (N_2277,N_2213,N_2160);
or U2278 (N_2278,N_2204,N_2191);
and U2279 (N_2279,N_2170,N_2212);
nand U2280 (N_2280,N_2241,N_2221);
and U2281 (N_2281,N_2250,N_2260);
nand U2282 (N_2282,N_2230,N_2234);
and U2283 (N_2283,N_2277,N_2273);
nor U2284 (N_2284,N_2238,N_2236);
nand U2285 (N_2285,N_2247,N_2252);
or U2286 (N_2286,N_2267,N_2239);
nor U2287 (N_2287,N_2220,N_2256);
nor U2288 (N_2288,N_2246,N_2253);
nand U2289 (N_2289,N_2264,N_2271);
nand U2290 (N_2290,N_2278,N_2257);
and U2291 (N_2291,N_2225,N_2233);
and U2292 (N_2292,N_2274,N_2272);
nand U2293 (N_2293,N_2262,N_2227);
nor U2294 (N_2294,N_2240,N_2259);
or U2295 (N_2295,N_2266,N_2245);
or U2296 (N_2296,N_2251,N_2255);
or U2297 (N_2297,N_2224,N_2265);
and U2298 (N_2298,N_2276,N_2229);
xor U2299 (N_2299,N_2242,N_2244);
nand U2300 (N_2300,N_2237,N_2263);
nor U2301 (N_2301,N_2226,N_2248);
and U2302 (N_2302,N_2232,N_2235);
nor U2303 (N_2303,N_2261,N_2275);
or U2304 (N_2304,N_2268,N_2254);
nor U2305 (N_2305,N_2279,N_2223);
or U2306 (N_2306,N_2228,N_2269);
nor U2307 (N_2307,N_2243,N_2249);
nand U2308 (N_2308,N_2258,N_2270);
or U2309 (N_2309,N_2222,N_2231);
and U2310 (N_2310,N_2277,N_2251);
nand U2311 (N_2311,N_2236,N_2247);
or U2312 (N_2312,N_2239,N_2238);
nand U2313 (N_2313,N_2242,N_2252);
nor U2314 (N_2314,N_2259,N_2266);
and U2315 (N_2315,N_2258,N_2252);
nor U2316 (N_2316,N_2271,N_2278);
nand U2317 (N_2317,N_2231,N_2240);
or U2318 (N_2318,N_2271,N_2236);
nand U2319 (N_2319,N_2222,N_2263);
nor U2320 (N_2320,N_2247,N_2237);
nand U2321 (N_2321,N_2223,N_2268);
nand U2322 (N_2322,N_2272,N_2270);
nor U2323 (N_2323,N_2261,N_2269);
or U2324 (N_2324,N_2275,N_2227);
nor U2325 (N_2325,N_2239,N_2263);
nand U2326 (N_2326,N_2237,N_2277);
or U2327 (N_2327,N_2236,N_2234);
xor U2328 (N_2328,N_2237,N_2248);
nor U2329 (N_2329,N_2255,N_2245);
nor U2330 (N_2330,N_2255,N_2257);
and U2331 (N_2331,N_2276,N_2250);
nor U2332 (N_2332,N_2224,N_2237);
nor U2333 (N_2333,N_2249,N_2235);
and U2334 (N_2334,N_2268,N_2237);
nand U2335 (N_2335,N_2222,N_2262);
and U2336 (N_2336,N_2250,N_2263);
or U2337 (N_2337,N_2253,N_2226);
nor U2338 (N_2338,N_2266,N_2244);
and U2339 (N_2339,N_2237,N_2227);
and U2340 (N_2340,N_2327,N_2291);
and U2341 (N_2341,N_2317,N_2331);
or U2342 (N_2342,N_2281,N_2313);
nand U2343 (N_2343,N_2314,N_2323);
nand U2344 (N_2344,N_2336,N_2297);
and U2345 (N_2345,N_2283,N_2318);
or U2346 (N_2346,N_2294,N_2311);
nand U2347 (N_2347,N_2302,N_2339);
or U2348 (N_2348,N_2310,N_2285);
nor U2349 (N_2349,N_2290,N_2284);
and U2350 (N_2350,N_2319,N_2335);
or U2351 (N_2351,N_2322,N_2312);
nor U2352 (N_2352,N_2328,N_2300);
or U2353 (N_2353,N_2309,N_2295);
xor U2354 (N_2354,N_2301,N_2303);
nand U2355 (N_2355,N_2324,N_2296);
nor U2356 (N_2356,N_2315,N_2286);
or U2357 (N_2357,N_2337,N_2304);
or U2358 (N_2358,N_2293,N_2316);
nand U2359 (N_2359,N_2298,N_2292);
nand U2360 (N_2360,N_2338,N_2326);
or U2361 (N_2361,N_2334,N_2320);
or U2362 (N_2362,N_2305,N_2330);
nand U2363 (N_2363,N_2325,N_2282);
nand U2364 (N_2364,N_2308,N_2306);
nor U2365 (N_2365,N_2321,N_2287);
or U2366 (N_2366,N_2288,N_2299);
and U2367 (N_2367,N_2333,N_2289);
nor U2368 (N_2368,N_2329,N_2280);
or U2369 (N_2369,N_2307,N_2332);
xor U2370 (N_2370,N_2305,N_2287);
nor U2371 (N_2371,N_2320,N_2325);
nor U2372 (N_2372,N_2330,N_2304);
nand U2373 (N_2373,N_2285,N_2283);
nor U2374 (N_2374,N_2332,N_2321);
and U2375 (N_2375,N_2310,N_2330);
nor U2376 (N_2376,N_2338,N_2336);
or U2377 (N_2377,N_2324,N_2297);
nor U2378 (N_2378,N_2314,N_2311);
nor U2379 (N_2379,N_2288,N_2307);
and U2380 (N_2380,N_2306,N_2317);
nand U2381 (N_2381,N_2305,N_2290);
nand U2382 (N_2382,N_2330,N_2286);
nand U2383 (N_2383,N_2326,N_2329);
and U2384 (N_2384,N_2310,N_2280);
or U2385 (N_2385,N_2295,N_2284);
and U2386 (N_2386,N_2300,N_2281);
nor U2387 (N_2387,N_2303,N_2316);
nand U2388 (N_2388,N_2296,N_2292);
nor U2389 (N_2389,N_2329,N_2312);
nor U2390 (N_2390,N_2328,N_2281);
nor U2391 (N_2391,N_2338,N_2307);
and U2392 (N_2392,N_2293,N_2322);
or U2393 (N_2393,N_2303,N_2281);
nand U2394 (N_2394,N_2310,N_2333);
or U2395 (N_2395,N_2280,N_2323);
or U2396 (N_2396,N_2337,N_2322);
and U2397 (N_2397,N_2296,N_2328);
nand U2398 (N_2398,N_2328,N_2332);
nand U2399 (N_2399,N_2320,N_2310);
nand U2400 (N_2400,N_2384,N_2359);
or U2401 (N_2401,N_2390,N_2386);
or U2402 (N_2402,N_2389,N_2355);
nor U2403 (N_2403,N_2373,N_2376);
nand U2404 (N_2404,N_2382,N_2363);
nor U2405 (N_2405,N_2361,N_2349);
or U2406 (N_2406,N_2396,N_2371);
nor U2407 (N_2407,N_2365,N_2368);
or U2408 (N_2408,N_2340,N_2375);
nor U2409 (N_2409,N_2399,N_2378);
nand U2410 (N_2410,N_2350,N_2362);
and U2411 (N_2411,N_2345,N_2381);
nand U2412 (N_2412,N_2351,N_2357);
nand U2413 (N_2413,N_2356,N_2385);
xor U2414 (N_2414,N_2377,N_2379);
and U2415 (N_2415,N_2344,N_2391);
xnor U2416 (N_2416,N_2360,N_2342);
nor U2417 (N_2417,N_2353,N_2374);
and U2418 (N_2418,N_2364,N_2372);
or U2419 (N_2419,N_2347,N_2348);
and U2420 (N_2420,N_2366,N_2367);
xnor U2421 (N_2421,N_2358,N_2352);
nor U2422 (N_2422,N_2394,N_2354);
nand U2423 (N_2423,N_2343,N_2369);
and U2424 (N_2424,N_2370,N_2383);
and U2425 (N_2425,N_2398,N_2395);
or U2426 (N_2426,N_2393,N_2380);
nor U2427 (N_2427,N_2346,N_2392);
and U2428 (N_2428,N_2397,N_2387);
nor U2429 (N_2429,N_2341,N_2388);
nor U2430 (N_2430,N_2386,N_2351);
nand U2431 (N_2431,N_2387,N_2390);
and U2432 (N_2432,N_2397,N_2395);
nand U2433 (N_2433,N_2376,N_2399);
and U2434 (N_2434,N_2383,N_2389);
nand U2435 (N_2435,N_2370,N_2397);
nand U2436 (N_2436,N_2373,N_2378);
nor U2437 (N_2437,N_2385,N_2391);
and U2438 (N_2438,N_2365,N_2399);
or U2439 (N_2439,N_2377,N_2348);
nand U2440 (N_2440,N_2346,N_2382);
or U2441 (N_2441,N_2366,N_2371);
or U2442 (N_2442,N_2376,N_2360);
and U2443 (N_2443,N_2383,N_2368);
nor U2444 (N_2444,N_2372,N_2367);
nand U2445 (N_2445,N_2344,N_2364);
or U2446 (N_2446,N_2371,N_2389);
and U2447 (N_2447,N_2385,N_2399);
nand U2448 (N_2448,N_2372,N_2344);
or U2449 (N_2449,N_2355,N_2341);
or U2450 (N_2450,N_2385,N_2376);
nand U2451 (N_2451,N_2368,N_2366);
or U2452 (N_2452,N_2373,N_2367);
nand U2453 (N_2453,N_2378,N_2367);
nand U2454 (N_2454,N_2369,N_2358);
nor U2455 (N_2455,N_2341,N_2358);
or U2456 (N_2456,N_2393,N_2364);
or U2457 (N_2457,N_2391,N_2372);
nand U2458 (N_2458,N_2349,N_2374);
nand U2459 (N_2459,N_2368,N_2382);
or U2460 (N_2460,N_2450,N_2453);
nor U2461 (N_2461,N_2444,N_2406);
xor U2462 (N_2462,N_2452,N_2412);
nor U2463 (N_2463,N_2410,N_2446);
nor U2464 (N_2464,N_2403,N_2424);
nand U2465 (N_2465,N_2442,N_2405);
and U2466 (N_2466,N_2449,N_2459);
nor U2467 (N_2467,N_2404,N_2416);
xnor U2468 (N_2468,N_2438,N_2420);
and U2469 (N_2469,N_2425,N_2423);
nand U2470 (N_2470,N_2428,N_2440);
xor U2471 (N_2471,N_2445,N_2419);
nor U2472 (N_2472,N_2431,N_2417);
or U2473 (N_2473,N_2421,N_2436);
nor U2474 (N_2474,N_2454,N_2407);
and U2475 (N_2475,N_2447,N_2401);
or U2476 (N_2476,N_2448,N_2455);
nor U2477 (N_2477,N_2433,N_2429);
nor U2478 (N_2478,N_2408,N_2458);
nand U2479 (N_2479,N_2435,N_2418);
and U2480 (N_2480,N_2427,N_2443);
nand U2481 (N_2481,N_2413,N_2441);
nor U2482 (N_2482,N_2414,N_2422);
nand U2483 (N_2483,N_2415,N_2457);
and U2484 (N_2484,N_2411,N_2400);
or U2485 (N_2485,N_2426,N_2432);
or U2486 (N_2486,N_2434,N_2402);
xor U2487 (N_2487,N_2456,N_2439);
or U2488 (N_2488,N_2437,N_2409);
or U2489 (N_2489,N_2451,N_2430);
or U2490 (N_2490,N_2448,N_2418);
and U2491 (N_2491,N_2434,N_2413);
and U2492 (N_2492,N_2424,N_2405);
or U2493 (N_2493,N_2404,N_2401);
or U2494 (N_2494,N_2413,N_2444);
or U2495 (N_2495,N_2436,N_2400);
and U2496 (N_2496,N_2445,N_2434);
nand U2497 (N_2497,N_2439,N_2402);
nor U2498 (N_2498,N_2452,N_2434);
and U2499 (N_2499,N_2447,N_2424);
nor U2500 (N_2500,N_2448,N_2446);
nor U2501 (N_2501,N_2414,N_2454);
nor U2502 (N_2502,N_2423,N_2406);
and U2503 (N_2503,N_2442,N_2409);
nand U2504 (N_2504,N_2441,N_2422);
nand U2505 (N_2505,N_2409,N_2419);
nand U2506 (N_2506,N_2411,N_2451);
nor U2507 (N_2507,N_2458,N_2402);
nand U2508 (N_2508,N_2415,N_2447);
nor U2509 (N_2509,N_2426,N_2429);
and U2510 (N_2510,N_2454,N_2434);
nand U2511 (N_2511,N_2408,N_2422);
and U2512 (N_2512,N_2416,N_2450);
nor U2513 (N_2513,N_2408,N_2451);
nor U2514 (N_2514,N_2415,N_2451);
or U2515 (N_2515,N_2429,N_2449);
and U2516 (N_2516,N_2400,N_2416);
or U2517 (N_2517,N_2457,N_2433);
nor U2518 (N_2518,N_2434,N_2409);
or U2519 (N_2519,N_2402,N_2442);
nand U2520 (N_2520,N_2508,N_2507);
nand U2521 (N_2521,N_2519,N_2500);
nor U2522 (N_2522,N_2476,N_2517);
or U2523 (N_2523,N_2475,N_2467);
nor U2524 (N_2524,N_2463,N_2481);
nand U2525 (N_2525,N_2472,N_2461);
nand U2526 (N_2526,N_2460,N_2502);
and U2527 (N_2527,N_2496,N_2491);
or U2528 (N_2528,N_2513,N_2487);
nand U2529 (N_2529,N_2480,N_2469);
or U2530 (N_2530,N_2510,N_2489);
nand U2531 (N_2531,N_2468,N_2465);
nor U2532 (N_2532,N_2515,N_2494);
nand U2533 (N_2533,N_2490,N_2504);
and U2534 (N_2534,N_2477,N_2514);
or U2535 (N_2535,N_2486,N_2493);
xnor U2536 (N_2536,N_2512,N_2485);
and U2537 (N_2537,N_2505,N_2518);
nand U2538 (N_2538,N_2473,N_2488);
nand U2539 (N_2539,N_2506,N_2474);
and U2540 (N_2540,N_2501,N_2462);
nand U2541 (N_2541,N_2483,N_2503);
xnor U2542 (N_2542,N_2471,N_2466);
nor U2543 (N_2543,N_2470,N_2509);
nor U2544 (N_2544,N_2516,N_2499);
nor U2545 (N_2545,N_2479,N_2478);
nor U2546 (N_2546,N_2498,N_2495);
and U2547 (N_2547,N_2497,N_2464);
nand U2548 (N_2548,N_2484,N_2482);
and U2549 (N_2549,N_2511,N_2492);
nand U2550 (N_2550,N_2471,N_2484);
nand U2551 (N_2551,N_2497,N_2483);
or U2552 (N_2552,N_2484,N_2506);
and U2553 (N_2553,N_2502,N_2498);
and U2554 (N_2554,N_2513,N_2509);
or U2555 (N_2555,N_2477,N_2490);
nor U2556 (N_2556,N_2473,N_2508);
nor U2557 (N_2557,N_2509,N_2506);
and U2558 (N_2558,N_2497,N_2506);
nand U2559 (N_2559,N_2466,N_2515);
or U2560 (N_2560,N_2501,N_2465);
nand U2561 (N_2561,N_2501,N_2505);
nand U2562 (N_2562,N_2501,N_2488);
nand U2563 (N_2563,N_2510,N_2513);
nor U2564 (N_2564,N_2479,N_2514);
and U2565 (N_2565,N_2488,N_2495);
and U2566 (N_2566,N_2498,N_2509);
nor U2567 (N_2567,N_2506,N_2517);
or U2568 (N_2568,N_2480,N_2466);
and U2569 (N_2569,N_2480,N_2502);
nor U2570 (N_2570,N_2461,N_2497);
nor U2571 (N_2571,N_2461,N_2498);
and U2572 (N_2572,N_2489,N_2509);
xnor U2573 (N_2573,N_2470,N_2497);
xnor U2574 (N_2574,N_2475,N_2478);
and U2575 (N_2575,N_2511,N_2508);
and U2576 (N_2576,N_2485,N_2472);
or U2577 (N_2577,N_2519,N_2478);
or U2578 (N_2578,N_2479,N_2488);
xor U2579 (N_2579,N_2463,N_2480);
and U2580 (N_2580,N_2567,N_2530);
nand U2581 (N_2581,N_2561,N_2548);
or U2582 (N_2582,N_2542,N_2539);
and U2583 (N_2583,N_2556,N_2570);
or U2584 (N_2584,N_2524,N_2577);
and U2585 (N_2585,N_2560,N_2523);
and U2586 (N_2586,N_2564,N_2576);
or U2587 (N_2587,N_2563,N_2536);
nand U2588 (N_2588,N_2573,N_2545);
nor U2589 (N_2589,N_2557,N_2575);
or U2590 (N_2590,N_2553,N_2551);
or U2591 (N_2591,N_2525,N_2546);
xnor U2592 (N_2592,N_2558,N_2574);
nor U2593 (N_2593,N_2527,N_2543);
nand U2594 (N_2594,N_2522,N_2544);
nand U2595 (N_2595,N_2538,N_2559);
and U2596 (N_2596,N_2521,N_2520);
nand U2597 (N_2597,N_2529,N_2534);
nor U2598 (N_2598,N_2572,N_2569);
or U2599 (N_2599,N_2537,N_2540);
and U2600 (N_2600,N_2555,N_2526);
nor U2601 (N_2601,N_2533,N_2550);
nand U2602 (N_2602,N_2532,N_2535);
or U2603 (N_2603,N_2566,N_2552);
nor U2604 (N_2604,N_2565,N_2579);
and U2605 (N_2605,N_2531,N_2541);
nor U2606 (N_2606,N_2528,N_2562);
and U2607 (N_2607,N_2554,N_2578);
or U2608 (N_2608,N_2568,N_2549);
xor U2609 (N_2609,N_2547,N_2571);
and U2610 (N_2610,N_2545,N_2557);
nand U2611 (N_2611,N_2571,N_2539);
or U2612 (N_2612,N_2572,N_2532);
xnor U2613 (N_2613,N_2525,N_2522);
nand U2614 (N_2614,N_2547,N_2540);
and U2615 (N_2615,N_2572,N_2561);
or U2616 (N_2616,N_2520,N_2548);
nor U2617 (N_2617,N_2548,N_2524);
and U2618 (N_2618,N_2544,N_2521);
and U2619 (N_2619,N_2521,N_2571);
nand U2620 (N_2620,N_2567,N_2547);
or U2621 (N_2621,N_2539,N_2533);
or U2622 (N_2622,N_2532,N_2576);
and U2623 (N_2623,N_2579,N_2561);
nand U2624 (N_2624,N_2527,N_2576);
nor U2625 (N_2625,N_2552,N_2576);
nor U2626 (N_2626,N_2531,N_2560);
nor U2627 (N_2627,N_2528,N_2577);
nor U2628 (N_2628,N_2578,N_2551);
or U2629 (N_2629,N_2574,N_2530);
and U2630 (N_2630,N_2573,N_2575);
nand U2631 (N_2631,N_2550,N_2548);
nor U2632 (N_2632,N_2523,N_2566);
and U2633 (N_2633,N_2567,N_2550);
or U2634 (N_2634,N_2524,N_2568);
nor U2635 (N_2635,N_2574,N_2571);
and U2636 (N_2636,N_2571,N_2541);
nor U2637 (N_2637,N_2579,N_2576);
xor U2638 (N_2638,N_2541,N_2547);
and U2639 (N_2639,N_2526,N_2531);
nand U2640 (N_2640,N_2626,N_2584);
nor U2641 (N_2641,N_2594,N_2617);
or U2642 (N_2642,N_2625,N_2611);
or U2643 (N_2643,N_2614,N_2605);
and U2644 (N_2644,N_2635,N_2629);
or U2645 (N_2645,N_2608,N_2633);
xor U2646 (N_2646,N_2609,N_2613);
and U2647 (N_2647,N_2589,N_2619);
and U2648 (N_2648,N_2598,N_2639);
nor U2649 (N_2649,N_2600,N_2583);
and U2650 (N_2650,N_2585,N_2631);
or U2651 (N_2651,N_2616,N_2622);
or U2652 (N_2652,N_2628,N_2607);
xor U2653 (N_2653,N_2630,N_2615);
nand U2654 (N_2654,N_2618,N_2581);
nor U2655 (N_2655,N_2597,N_2582);
nor U2656 (N_2656,N_2620,N_2596);
nor U2657 (N_2657,N_2624,N_2593);
nor U2658 (N_2658,N_2636,N_2602);
and U2659 (N_2659,N_2634,N_2588);
or U2660 (N_2660,N_2612,N_2592);
nor U2661 (N_2661,N_2599,N_2621);
and U2662 (N_2662,N_2632,N_2601);
nor U2663 (N_2663,N_2627,N_2595);
nor U2664 (N_2664,N_2590,N_2587);
nand U2665 (N_2665,N_2610,N_2638);
xor U2666 (N_2666,N_2580,N_2623);
and U2667 (N_2667,N_2606,N_2586);
or U2668 (N_2668,N_2604,N_2591);
nand U2669 (N_2669,N_2637,N_2603);
and U2670 (N_2670,N_2625,N_2618);
or U2671 (N_2671,N_2600,N_2610);
and U2672 (N_2672,N_2612,N_2625);
nor U2673 (N_2673,N_2585,N_2627);
nand U2674 (N_2674,N_2611,N_2603);
nor U2675 (N_2675,N_2597,N_2594);
nor U2676 (N_2676,N_2612,N_2583);
or U2677 (N_2677,N_2627,N_2613);
and U2678 (N_2678,N_2588,N_2624);
and U2679 (N_2679,N_2631,N_2601);
and U2680 (N_2680,N_2602,N_2603);
or U2681 (N_2681,N_2625,N_2617);
nor U2682 (N_2682,N_2639,N_2637);
xor U2683 (N_2683,N_2624,N_2616);
and U2684 (N_2684,N_2624,N_2629);
xnor U2685 (N_2685,N_2619,N_2628);
nor U2686 (N_2686,N_2625,N_2616);
nand U2687 (N_2687,N_2591,N_2583);
or U2688 (N_2688,N_2600,N_2636);
nand U2689 (N_2689,N_2618,N_2633);
and U2690 (N_2690,N_2599,N_2603);
or U2691 (N_2691,N_2616,N_2605);
nand U2692 (N_2692,N_2637,N_2633);
and U2693 (N_2693,N_2624,N_2631);
and U2694 (N_2694,N_2603,N_2584);
nand U2695 (N_2695,N_2627,N_2631);
and U2696 (N_2696,N_2638,N_2604);
nand U2697 (N_2697,N_2590,N_2623);
xnor U2698 (N_2698,N_2590,N_2609);
or U2699 (N_2699,N_2623,N_2627);
nor U2700 (N_2700,N_2655,N_2643);
and U2701 (N_2701,N_2648,N_2665);
or U2702 (N_2702,N_2682,N_2645);
nor U2703 (N_2703,N_2649,N_2659);
nor U2704 (N_2704,N_2647,N_2667);
nand U2705 (N_2705,N_2677,N_2686);
nand U2706 (N_2706,N_2652,N_2694);
or U2707 (N_2707,N_2660,N_2685);
and U2708 (N_2708,N_2671,N_2693);
nor U2709 (N_2709,N_2668,N_2669);
and U2710 (N_2710,N_2662,N_2661);
nor U2711 (N_2711,N_2666,N_2684);
or U2712 (N_2712,N_2650,N_2688);
and U2713 (N_2713,N_2675,N_2644);
nand U2714 (N_2714,N_2680,N_2698);
or U2715 (N_2715,N_2654,N_2687);
nand U2716 (N_2716,N_2663,N_2656);
nor U2717 (N_2717,N_2699,N_2690);
or U2718 (N_2718,N_2679,N_2692);
nand U2719 (N_2719,N_2683,N_2657);
nor U2720 (N_2720,N_2695,N_2642);
and U2721 (N_2721,N_2640,N_2651);
and U2722 (N_2722,N_2678,N_2641);
nand U2723 (N_2723,N_2674,N_2670);
and U2724 (N_2724,N_2658,N_2664);
or U2725 (N_2725,N_2681,N_2676);
nor U2726 (N_2726,N_2691,N_2653);
nand U2727 (N_2727,N_2646,N_2672);
nor U2728 (N_2728,N_2673,N_2696);
or U2729 (N_2729,N_2697,N_2689);
nand U2730 (N_2730,N_2662,N_2697);
or U2731 (N_2731,N_2664,N_2650);
nand U2732 (N_2732,N_2643,N_2646);
or U2733 (N_2733,N_2695,N_2657);
nor U2734 (N_2734,N_2670,N_2679);
or U2735 (N_2735,N_2690,N_2695);
or U2736 (N_2736,N_2669,N_2645);
and U2737 (N_2737,N_2682,N_2673);
or U2738 (N_2738,N_2664,N_2667);
or U2739 (N_2739,N_2689,N_2667);
or U2740 (N_2740,N_2695,N_2655);
or U2741 (N_2741,N_2657,N_2661);
and U2742 (N_2742,N_2659,N_2684);
or U2743 (N_2743,N_2686,N_2688);
nand U2744 (N_2744,N_2642,N_2653);
nor U2745 (N_2745,N_2697,N_2665);
and U2746 (N_2746,N_2661,N_2695);
or U2747 (N_2747,N_2672,N_2696);
nand U2748 (N_2748,N_2661,N_2664);
or U2749 (N_2749,N_2643,N_2676);
or U2750 (N_2750,N_2645,N_2661);
nor U2751 (N_2751,N_2648,N_2682);
and U2752 (N_2752,N_2643,N_2668);
nor U2753 (N_2753,N_2659,N_2655);
nor U2754 (N_2754,N_2668,N_2652);
nor U2755 (N_2755,N_2643,N_2640);
nor U2756 (N_2756,N_2680,N_2658);
or U2757 (N_2757,N_2656,N_2689);
and U2758 (N_2758,N_2691,N_2664);
or U2759 (N_2759,N_2652,N_2660);
and U2760 (N_2760,N_2759,N_2724);
and U2761 (N_2761,N_2719,N_2737);
and U2762 (N_2762,N_2743,N_2753);
xor U2763 (N_2763,N_2731,N_2733);
nand U2764 (N_2764,N_2745,N_2751);
and U2765 (N_2765,N_2716,N_2711);
nor U2766 (N_2766,N_2707,N_2755);
nand U2767 (N_2767,N_2723,N_2727);
nand U2768 (N_2768,N_2756,N_2700);
and U2769 (N_2769,N_2747,N_2757);
and U2770 (N_2770,N_2721,N_2718);
or U2771 (N_2771,N_2744,N_2705);
xor U2772 (N_2772,N_2750,N_2736);
and U2773 (N_2773,N_2730,N_2735);
nand U2774 (N_2774,N_2701,N_2706);
or U2775 (N_2775,N_2752,N_2739);
or U2776 (N_2776,N_2715,N_2710);
and U2777 (N_2777,N_2740,N_2702);
or U2778 (N_2778,N_2742,N_2734);
or U2779 (N_2779,N_2712,N_2709);
or U2780 (N_2780,N_2704,N_2738);
and U2781 (N_2781,N_2726,N_2729);
or U2782 (N_2782,N_2714,N_2754);
or U2783 (N_2783,N_2703,N_2708);
or U2784 (N_2784,N_2758,N_2749);
or U2785 (N_2785,N_2748,N_2725);
or U2786 (N_2786,N_2713,N_2722);
and U2787 (N_2787,N_2746,N_2720);
nor U2788 (N_2788,N_2732,N_2717);
nor U2789 (N_2789,N_2741,N_2728);
nand U2790 (N_2790,N_2739,N_2702);
nor U2791 (N_2791,N_2731,N_2746);
nor U2792 (N_2792,N_2738,N_2705);
and U2793 (N_2793,N_2718,N_2749);
nand U2794 (N_2794,N_2729,N_2724);
nor U2795 (N_2795,N_2717,N_2738);
and U2796 (N_2796,N_2723,N_2747);
and U2797 (N_2797,N_2725,N_2756);
and U2798 (N_2798,N_2711,N_2723);
or U2799 (N_2799,N_2749,N_2716);
xnor U2800 (N_2800,N_2714,N_2734);
nor U2801 (N_2801,N_2715,N_2712);
nand U2802 (N_2802,N_2704,N_2733);
nor U2803 (N_2803,N_2730,N_2747);
nor U2804 (N_2804,N_2721,N_2714);
or U2805 (N_2805,N_2756,N_2709);
nand U2806 (N_2806,N_2739,N_2736);
and U2807 (N_2807,N_2738,N_2730);
nand U2808 (N_2808,N_2745,N_2717);
nand U2809 (N_2809,N_2755,N_2731);
nand U2810 (N_2810,N_2736,N_2735);
nor U2811 (N_2811,N_2746,N_2735);
or U2812 (N_2812,N_2755,N_2746);
nor U2813 (N_2813,N_2745,N_2752);
nor U2814 (N_2814,N_2726,N_2750);
nor U2815 (N_2815,N_2741,N_2713);
nor U2816 (N_2816,N_2718,N_2722);
xor U2817 (N_2817,N_2700,N_2712);
nand U2818 (N_2818,N_2715,N_2702);
or U2819 (N_2819,N_2724,N_2749);
nand U2820 (N_2820,N_2804,N_2816);
nor U2821 (N_2821,N_2780,N_2774);
nor U2822 (N_2822,N_2806,N_2801);
and U2823 (N_2823,N_2815,N_2772);
nand U2824 (N_2824,N_2764,N_2776);
or U2825 (N_2825,N_2788,N_2791);
nand U2826 (N_2826,N_2773,N_2799);
nand U2827 (N_2827,N_2818,N_2771);
nand U2828 (N_2828,N_2813,N_2808);
nor U2829 (N_2829,N_2777,N_2761);
and U2830 (N_2830,N_2807,N_2785);
nand U2831 (N_2831,N_2770,N_2809);
nand U2832 (N_2832,N_2817,N_2798);
nand U2833 (N_2833,N_2819,N_2767);
xor U2834 (N_2834,N_2763,N_2779);
nor U2835 (N_2835,N_2793,N_2795);
nor U2836 (N_2836,N_2796,N_2814);
nand U2837 (N_2837,N_2794,N_2800);
or U2838 (N_2838,N_2762,N_2768);
and U2839 (N_2839,N_2805,N_2790);
nor U2840 (N_2840,N_2760,N_2769);
and U2841 (N_2841,N_2802,N_2778);
or U2842 (N_2842,N_2792,N_2789);
and U2843 (N_2843,N_2782,N_2783);
nand U2844 (N_2844,N_2811,N_2812);
nor U2845 (N_2845,N_2766,N_2784);
and U2846 (N_2846,N_2781,N_2797);
or U2847 (N_2847,N_2765,N_2786);
nand U2848 (N_2848,N_2803,N_2775);
or U2849 (N_2849,N_2787,N_2810);
or U2850 (N_2850,N_2780,N_2792);
xor U2851 (N_2851,N_2813,N_2775);
and U2852 (N_2852,N_2773,N_2760);
nor U2853 (N_2853,N_2774,N_2788);
or U2854 (N_2854,N_2801,N_2790);
nand U2855 (N_2855,N_2761,N_2784);
xnor U2856 (N_2856,N_2796,N_2785);
and U2857 (N_2857,N_2779,N_2772);
and U2858 (N_2858,N_2796,N_2807);
or U2859 (N_2859,N_2805,N_2804);
nor U2860 (N_2860,N_2772,N_2812);
nand U2861 (N_2861,N_2772,N_2777);
nand U2862 (N_2862,N_2763,N_2798);
nand U2863 (N_2863,N_2763,N_2799);
nor U2864 (N_2864,N_2818,N_2766);
or U2865 (N_2865,N_2771,N_2813);
and U2866 (N_2866,N_2771,N_2814);
and U2867 (N_2867,N_2802,N_2794);
xnor U2868 (N_2868,N_2783,N_2789);
nand U2869 (N_2869,N_2811,N_2762);
nor U2870 (N_2870,N_2792,N_2777);
nand U2871 (N_2871,N_2764,N_2795);
or U2872 (N_2872,N_2791,N_2778);
nor U2873 (N_2873,N_2787,N_2782);
nor U2874 (N_2874,N_2811,N_2763);
nor U2875 (N_2875,N_2809,N_2819);
nand U2876 (N_2876,N_2782,N_2802);
nor U2877 (N_2877,N_2786,N_2789);
and U2878 (N_2878,N_2812,N_2762);
or U2879 (N_2879,N_2795,N_2805);
or U2880 (N_2880,N_2869,N_2848);
or U2881 (N_2881,N_2859,N_2879);
nor U2882 (N_2882,N_2853,N_2873);
or U2883 (N_2883,N_2862,N_2833);
and U2884 (N_2884,N_2826,N_2877);
or U2885 (N_2885,N_2874,N_2829);
nand U2886 (N_2886,N_2823,N_2825);
and U2887 (N_2887,N_2855,N_2864);
or U2888 (N_2888,N_2842,N_2820);
or U2889 (N_2889,N_2821,N_2841);
nor U2890 (N_2890,N_2846,N_2844);
nor U2891 (N_2891,N_2871,N_2827);
or U2892 (N_2892,N_2838,N_2872);
nand U2893 (N_2893,N_2832,N_2824);
and U2894 (N_2894,N_2851,N_2868);
or U2895 (N_2895,N_2878,N_2836);
and U2896 (N_2896,N_2852,N_2843);
nor U2897 (N_2897,N_2828,N_2865);
xnor U2898 (N_2898,N_2856,N_2861);
nand U2899 (N_2899,N_2857,N_2875);
nor U2900 (N_2900,N_2866,N_2845);
nor U2901 (N_2901,N_2863,N_2830);
or U2902 (N_2902,N_2831,N_2835);
and U2903 (N_2903,N_2870,N_2867);
and U2904 (N_2904,N_2834,N_2837);
nor U2905 (N_2905,N_2858,N_2849);
or U2906 (N_2906,N_2839,N_2840);
and U2907 (N_2907,N_2847,N_2876);
and U2908 (N_2908,N_2822,N_2850);
and U2909 (N_2909,N_2854,N_2860);
or U2910 (N_2910,N_2876,N_2863);
nand U2911 (N_2911,N_2865,N_2837);
and U2912 (N_2912,N_2857,N_2848);
or U2913 (N_2913,N_2820,N_2870);
xnor U2914 (N_2914,N_2858,N_2830);
or U2915 (N_2915,N_2842,N_2832);
nor U2916 (N_2916,N_2847,N_2820);
xor U2917 (N_2917,N_2822,N_2823);
nand U2918 (N_2918,N_2828,N_2851);
or U2919 (N_2919,N_2858,N_2862);
nand U2920 (N_2920,N_2857,N_2878);
nand U2921 (N_2921,N_2823,N_2872);
nor U2922 (N_2922,N_2829,N_2850);
and U2923 (N_2923,N_2845,N_2831);
nand U2924 (N_2924,N_2833,N_2829);
and U2925 (N_2925,N_2855,N_2852);
nand U2926 (N_2926,N_2847,N_2834);
xor U2927 (N_2927,N_2832,N_2876);
and U2928 (N_2928,N_2829,N_2842);
nor U2929 (N_2929,N_2825,N_2839);
nand U2930 (N_2930,N_2822,N_2847);
nand U2931 (N_2931,N_2848,N_2853);
nor U2932 (N_2932,N_2829,N_2827);
and U2933 (N_2933,N_2840,N_2824);
nand U2934 (N_2934,N_2858,N_2865);
nand U2935 (N_2935,N_2835,N_2848);
nor U2936 (N_2936,N_2852,N_2860);
and U2937 (N_2937,N_2853,N_2867);
nor U2938 (N_2938,N_2821,N_2827);
nor U2939 (N_2939,N_2825,N_2833);
and U2940 (N_2940,N_2918,N_2890);
nand U2941 (N_2941,N_2911,N_2932);
or U2942 (N_2942,N_2920,N_2883);
or U2943 (N_2943,N_2902,N_2905);
and U2944 (N_2944,N_2916,N_2894);
and U2945 (N_2945,N_2899,N_2935);
or U2946 (N_2946,N_2912,N_2939);
and U2947 (N_2947,N_2930,N_2910);
or U2948 (N_2948,N_2887,N_2927);
nand U2949 (N_2949,N_2908,N_2934);
nor U2950 (N_2950,N_2917,N_2938);
or U2951 (N_2951,N_2892,N_2888);
or U2952 (N_2952,N_2931,N_2897);
and U2953 (N_2953,N_2923,N_2881);
or U2954 (N_2954,N_2919,N_2909);
nand U2955 (N_2955,N_2903,N_2900);
nand U2956 (N_2956,N_2884,N_2913);
nand U2957 (N_2957,N_2898,N_2922);
or U2958 (N_2958,N_2882,N_2924);
nor U2959 (N_2959,N_2914,N_2891);
and U2960 (N_2960,N_2936,N_2937);
or U2961 (N_2961,N_2906,N_2926);
and U2962 (N_2962,N_2907,N_2895);
and U2963 (N_2963,N_2915,N_2886);
nand U2964 (N_2964,N_2904,N_2929);
and U2965 (N_2965,N_2889,N_2896);
xor U2966 (N_2966,N_2928,N_2901);
and U2967 (N_2967,N_2893,N_2925);
nand U2968 (N_2968,N_2933,N_2885);
nor U2969 (N_2969,N_2880,N_2921);
or U2970 (N_2970,N_2927,N_2920);
nor U2971 (N_2971,N_2903,N_2924);
or U2972 (N_2972,N_2894,N_2897);
and U2973 (N_2973,N_2919,N_2897);
and U2974 (N_2974,N_2918,N_2903);
nand U2975 (N_2975,N_2888,N_2891);
and U2976 (N_2976,N_2897,N_2892);
and U2977 (N_2977,N_2934,N_2883);
nand U2978 (N_2978,N_2935,N_2918);
xnor U2979 (N_2979,N_2928,N_2930);
and U2980 (N_2980,N_2895,N_2887);
or U2981 (N_2981,N_2914,N_2905);
or U2982 (N_2982,N_2911,N_2884);
or U2983 (N_2983,N_2927,N_2910);
and U2984 (N_2984,N_2927,N_2936);
and U2985 (N_2985,N_2882,N_2885);
nor U2986 (N_2986,N_2920,N_2891);
nand U2987 (N_2987,N_2904,N_2906);
nor U2988 (N_2988,N_2938,N_2909);
and U2989 (N_2989,N_2936,N_2926);
and U2990 (N_2990,N_2888,N_2925);
nor U2991 (N_2991,N_2898,N_2927);
nand U2992 (N_2992,N_2923,N_2910);
and U2993 (N_2993,N_2883,N_2899);
or U2994 (N_2994,N_2913,N_2931);
or U2995 (N_2995,N_2918,N_2926);
xor U2996 (N_2996,N_2937,N_2935);
nor U2997 (N_2997,N_2902,N_2915);
and U2998 (N_2998,N_2916,N_2936);
nor U2999 (N_2999,N_2919,N_2920);
nor UO_0 (O_0,N_2978,N_2999);
nand UO_1 (O_1,N_2969,N_2994);
and UO_2 (O_2,N_2990,N_2943);
nand UO_3 (O_3,N_2997,N_2959);
or UO_4 (O_4,N_2940,N_2965);
nand UO_5 (O_5,N_2974,N_2961);
or UO_6 (O_6,N_2995,N_2964);
nor UO_7 (O_7,N_2991,N_2973);
or UO_8 (O_8,N_2976,N_2942);
nand UO_9 (O_9,N_2984,N_2968);
nor UO_10 (O_10,N_2947,N_2963);
nor UO_11 (O_11,N_2966,N_2958);
nand UO_12 (O_12,N_2987,N_2989);
nor UO_13 (O_13,N_2950,N_2988);
or UO_14 (O_14,N_2941,N_2944);
or UO_15 (O_15,N_2983,N_2962);
nor UO_16 (O_16,N_2954,N_2993);
nor UO_17 (O_17,N_2967,N_2951);
nand UO_18 (O_18,N_2971,N_2981);
or UO_19 (O_19,N_2956,N_2957);
or UO_20 (O_20,N_2980,N_2985);
nor UO_21 (O_21,N_2946,N_2953);
or UO_22 (O_22,N_2952,N_2998);
nand UO_23 (O_23,N_2948,N_2945);
and UO_24 (O_24,N_2970,N_2955);
nand UO_25 (O_25,N_2975,N_2972);
nand UO_26 (O_26,N_2996,N_2992);
and UO_27 (O_27,N_2949,N_2979);
or UO_28 (O_28,N_2977,N_2986);
and UO_29 (O_29,N_2960,N_2982);
and UO_30 (O_30,N_2948,N_2941);
or UO_31 (O_31,N_2985,N_2963);
nor UO_32 (O_32,N_2985,N_2975);
nor UO_33 (O_33,N_2963,N_2984);
nand UO_34 (O_34,N_2997,N_2991);
nor UO_35 (O_35,N_2948,N_2947);
nand UO_36 (O_36,N_2974,N_2981);
nand UO_37 (O_37,N_2947,N_2944);
nand UO_38 (O_38,N_2963,N_2983);
nand UO_39 (O_39,N_2973,N_2954);
nand UO_40 (O_40,N_2983,N_2976);
or UO_41 (O_41,N_2941,N_2953);
nor UO_42 (O_42,N_2955,N_2957);
nor UO_43 (O_43,N_2966,N_2977);
nand UO_44 (O_44,N_2991,N_2940);
or UO_45 (O_45,N_2971,N_2969);
or UO_46 (O_46,N_2998,N_2976);
nor UO_47 (O_47,N_2974,N_2956);
or UO_48 (O_48,N_2981,N_2997);
or UO_49 (O_49,N_2953,N_2973);
and UO_50 (O_50,N_2954,N_2981);
and UO_51 (O_51,N_2978,N_2977);
and UO_52 (O_52,N_2970,N_2967);
nor UO_53 (O_53,N_2947,N_2964);
and UO_54 (O_54,N_2955,N_2971);
and UO_55 (O_55,N_2985,N_2944);
or UO_56 (O_56,N_2997,N_2949);
nor UO_57 (O_57,N_2946,N_2982);
nand UO_58 (O_58,N_2967,N_2966);
nor UO_59 (O_59,N_2951,N_2979);
nand UO_60 (O_60,N_2952,N_2967);
nand UO_61 (O_61,N_2946,N_2947);
and UO_62 (O_62,N_2950,N_2983);
and UO_63 (O_63,N_2948,N_2993);
or UO_64 (O_64,N_2981,N_2996);
or UO_65 (O_65,N_2997,N_2958);
and UO_66 (O_66,N_2948,N_2942);
nand UO_67 (O_67,N_2990,N_2952);
or UO_68 (O_68,N_2984,N_2989);
and UO_69 (O_69,N_2991,N_2954);
and UO_70 (O_70,N_2983,N_2966);
and UO_71 (O_71,N_2980,N_2947);
nand UO_72 (O_72,N_2960,N_2951);
nand UO_73 (O_73,N_2963,N_2943);
and UO_74 (O_74,N_2950,N_2955);
nor UO_75 (O_75,N_2970,N_2951);
nand UO_76 (O_76,N_2997,N_2985);
nor UO_77 (O_77,N_2958,N_2969);
nand UO_78 (O_78,N_2963,N_2999);
nor UO_79 (O_79,N_2950,N_2959);
or UO_80 (O_80,N_2979,N_2968);
or UO_81 (O_81,N_2985,N_2996);
nand UO_82 (O_82,N_2983,N_2965);
or UO_83 (O_83,N_2965,N_2958);
nor UO_84 (O_84,N_2975,N_2943);
and UO_85 (O_85,N_2946,N_2958);
and UO_86 (O_86,N_2975,N_2994);
or UO_87 (O_87,N_2983,N_2953);
or UO_88 (O_88,N_2994,N_2953);
nand UO_89 (O_89,N_2994,N_2944);
and UO_90 (O_90,N_2999,N_2957);
or UO_91 (O_91,N_2964,N_2955);
or UO_92 (O_92,N_2942,N_2958);
and UO_93 (O_93,N_2950,N_2999);
nand UO_94 (O_94,N_2948,N_2962);
or UO_95 (O_95,N_2946,N_2979);
or UO_96 (O_96,N_2988,N_2999);
nand UO_97 (O_97,N_2996,N_2965);
and UO_98 (O_98,N_2963,N_2949);
nor UO_99 (O_99,N_2991,N_2975);
nor UO_100 (O_100,N_2998,N_2946);
or UO_101 (O_101,N_2942,N_2941);
and UO_102 (O_102,N_2992,N_2980);
and UO_103 (O_103,N_2952,N_2997);
nand UO_104 (O_104,N_2996,N_2999);
and UO_105 (O_105,N_2964,N_2994);
or UO_106 (O_106,N_2998,N_2965);
and UO_107 (O_107,N_2952,N_2947);
nand UO_108 (O_108,N_2954,N_2969);
or UO_109 (O_109,N_2957,N_2977);
and UO_110 (O_110,N_2947,N_2992);
or UO_111 (O_111,N_2948,N_2951);
and UO_112 (O_112,N_2984,N_2967);
nand UO_113 (O_113,N_2985,N_2961);
and UO_114 (O_114,N_2973,N_2979);
or UO_115 (O_115,N_2964,N_2946);
nand UO_116 (O_116,N_2948,N_2981);
or UO_117 (O_117,N_2959,N_2961);
nand UO_118 (O_118,N_2956,N_2977);
nor UO_119 (O_119,N_2945,N_2950);
nand UO_120 (O_120,N_2978,N_2972);
nand UO_121 (O_121,N_2974,N_2982);
nand UO_122 (O_122,N_2961,N_2958);
and UO_123 (O_123,N_2990,N_2988);
nor UO_124 (O_124,N_2942,N_2994);
and UO_125 (O_125,N_2981,N_2990);
and UO_126 (O_126,N_2976,N_2973);
nand UO_127 (O_127,N_2982,N_2958);
nand UO_128 (O_128,N_2948,N_2989);
xor UO_129 (O_129,N_2961,N_2972);
or UO_130 (O_130,N_2955,N_2991);
nor UO_131 (O_131,N_2955,N_2943);
nor UO_132 (O_132,N_2989,N_2970);
or UO_133 (O_133,N_2993,N_2953);
nor UO_134 (O_134,N_2998,N_2999);
and UO_135 (O_135,N_2967,N_2971);
nor UO_136 (O_136,N_2949,N_2981);
and UO_137 (O_137,N_2968,N_2993);
and UO_138 (O_138,N_2995,N_2958);
nor UO_139 (O_139,N_2967,N_2978);
nand UO_140 (O_140,N_2953,N_2972);
or UO_141 (O_141,N_2999,N_2993);
or UO_142 (O_142,N_2946,N_2960);
nor UO_143 (O_143,N_2997,N_2988);
nand UO_144 (O_144,N_2955,N_2986);
nor UO_145 (O_145,N_2950,N_2962);
and UO_146 (O_146,N_2983,N_2994);
or UO_147 (O_147,N_2957,N_2987);
or UO_148 (O_148,N_2971,N_2942);
nor UO_149 (O_149,N_2972,N_2976);
nor UO_150 (O_150,N_2991,N_2947);
or UO_151 (O_151,N_2942,N_2977);
nand UO_152 (O_152,N_2940,N_2967);
or UO_153 (O_153,N_2970,N_2961);
or UO_154 (O_154,N_2995,N_2982);
nand UO_155 (O_155,N_2966,N_2944);
nor UO_156 (O_156,N_2941,N_2956);
xnor UO_157 (O_157,N_2972,N_2995);
nand UO_158 (O_158,N_2989,N_2977);
nand UO_159 (O_159,N_2982,N_2984);
and UO_160 (O_160,N_2966,N_2994);
or UO_161 (O_161,N_2967,N_2989);
and UO_162 (O_162,N_2945,N_2963);
nor UO_163 (O_163,N_2943,N_2976);
or UO_164 (O_164,N_2983,N_2967);
nand UO_165 (O_165,N_2951,N_2999);
and UO_166 (O_166,N_2942,N_2988);
and UO_167 (O_167,N_2970,N_2962);
or UO_168 (O_168,N_2992,N_2961);
nand UO_169 (O_169,N_2949,N_2945);
nor UO_170 (O_170,N_2988,N_2989);
nand UO_171 (O_171,N_2966,N_2995);
nand UO_172 (O_172,N_2979,N_2957);
xor UO_173 (O_173,N_2962,N_2995);
and UO_174 (O_174,N_2975,N_2945);
nor UO_175 (O_175,N_2953,N_2990);
nand UO_176 (O_176,N_2985,N_2994);
and UO_177 (O_177,N_2959,N_2954);
and UO_178 (O_178,N_2984,N_2978);
nor UO_179 (O_179,N_2961,N_2987);
or UO_180 (O_180,N_2988,N_2973);
and UO_181 (O_181,N_2999,N_2966);
nor UO_182 (O_182,N_2973,N_2985);
nand UO_183 (O_183,N_2984,N_2953);
xor UO_184 (O_184,N_2949,N_2966);
nor UO_185 (O_185,N_2976,N_2958);
or UO_186 (O_186,N_2977,N_2951);
or UO_187 (O_187,N_2976,N_2981);
xor UO_188 (O_188,N_2979,N_2998);
or UO_189 (O_189,N_2975,N_2955);
and UO_190 (O_190,N_2971,N_2941);
nand UO_191 (O_191,N_2991,N_2943);
nand UO_192 (O_192,N_2949,N_2955);
or UO_193 (O_193,N_2980,N_2962);
nand UO_194 (O_194,N_2967,N_2975);
or UO_195 (O_195,N_2986,N_2943);
nor UO_196 (O_196,N_2959,N_2971);
nand UO_197 (O_197,N_2971,N_2947);
and UO_198 (O_198,N_2950,N_2964);
and UO_199 (O_199,N_2978,N_2961);
nand UO_200 (O_200,N_2943,N_2946);
nor UO_201 (O_201,N_2949,N_2994);
and UO_202 (O_202,N_2970,N_2982);
nor UO_203 (O_203,N_2977,N_2965);
or UO_204 (O_204,N_2947,N_2956);
and UO_205 (O_205,N_2987,N_2959);
nor UO_206 (O_206,N_2948,N_2965);
or UO_207 (O_207,N_2958,N_2943);
and UO_208 (O_208,N_2941,N_2986);
nor UO_209 (O_209,N_2987,N_2990);
nand UO_210 (O_210,N_2946,N_2948);
nand UO_211 (O_211,N_2998,N_2971);
or UO_212 (O_212,N_2982,N_2942);
and UO_213 (O_213,N_2979,N_2963);
or UO_214 (O_214,N_2996,N_2993);
nand UO_215 (O_215,N_2956,N_2971);
or UO_216 (O_216,N_2974,N_2973);
or UO_217 (O_217,N_2990,N_2968);
or UO_218 (O_218,N_2969,N_2957);
nor UO_219 (O_219,N_2975,N_2988);
or UO_220 (O_220,N_2983,N_2957);
or UO_221 (O_221,N_2994,N_2998);
and UO_222 (O_222,N_2993,N_2967);
or UO_223 (O_223,N_2978,N_2947);
or UO_224 (O_224,N_2981,N_2984);
nor UO_225 (O_225,N_2985,N_2995);
and UO_226 (O_226,N_2963,N_2989);
nand UO_227 (O_227,N_2977,N_2970);
nor UO_228 (O_228,N_2956,N_2946);
and UO_229 (O_229,N_2993,N_2983);
or UO_230 (O_230,N_2953,N_2979);
nand UO_231 (O_231,N_2960,N_2947);
and UO_232 (O_232,N_2973,N_2963);
and UO_233 (O_233,N_2995,N_2944);
nand UO_234 (O_234,N_2966,N_2954);
nand UO_235 (O_235,N_2948,N_2940);
and UO_236 (O_236,N_2953,N_2981);
nor UO_237 (O_237,N_2962,N_2988);
and UO_238 (O_238,N_2989,N_2999);
nor UO_239 (O_239,N_2942,N_2956);
or UO_240 (O_240,N_2981,N_2942);
nor UO_241 (O_241,N_2945,N_2990);
and UO_242 (O_242,N_2974,N_2983);
and UO_243 (O_243,N_2993,N_2975);
or UO_244 (O_244,N_2996,N_2988);
nor UO_245 (O_245,N_2964,N_2944);
and UO_246 (O_246,N_2960,N_2986);
nand UO_247 (O_247,N_2966,N_2991);
nand UO_248 (O_248,N_2973,N_2977);
or UO_249 (O_249,N_2988,N_2992);
nand UO_250 (O_250,N_2944,N_2949);
nor UO_251 (O_251,N_2968,N_2950);
nor UO_252 (O_252,N_2982,N_2943);
nor UO_253 (O_253,N_2954,N_2950);
and UO_254 (O_254,N_2961,N_2963);
nand UO_255 (O_255,N_2959,N_2980);
or UO_256 (O_256,N_2999,N_2949);
or UO_257 (O_257,N_2945,N_2946);
nor UO_258 (O_258,N_2989,N_2995);
nor UO_259 (O_259,N_2944,N_2981);
nand UO_260 (O_260,N_2950,N_2948);
or UO_261 (O_261,N_2942,N_2992);
nand UO_262 (O_262,N_2942,N_2950);
and UO_263 (O_263,N_2941,N_2989);
xor UO_264 (O_264,N_2970,N_2944);
and UO_265 (O_265,N_2942,N_2975);
nand UO_266 (O_266,N_2959,N_2949);
nand UO_267 (O_267,N_2954,N_2995);
or UO_268 (O_268,N_2989,N_2954);
and UO_269 (O_269,N_2980,N_2969);
nand UO_270 (O_270,N_2966,N_2957);
or UO_271 (O_271,N_2962,N_2951);
nor UO_272 (O_272,N_2960,N_2956);
and UO_273 (O_273,N_2951,N_2992);
and UO_274 (O_274,N_2994,N_2956);
nor UO_275 (O_275,N_2969,N_2997);
nor UO_276 (O_276,N_2967,N_2948);
nand UO_277 (O_277,N_2995,N_2945);
nand UO_278 (O_278,N_2965,N_2956);
and UO_279 (O_279,N_2995,N_2977);
nand UO_280 (O_280,N_2990,N_2986);
nand UO_281 (O_281,N_2949,N_2998);
nand UO_282 (O_282,N_2998,N_2995);
nand UO_283 (O_283,N_2945,N_2966);
and UO_284 (O_284,N_2974,N_2953);
nor UO_285 (O_285,N_2963,N_2965);
nor UO_286 (O_286,N_2943,N_2969);
xor UO_287 (O_287,N_2960,N_2954);
nand UO_288 (O_288,N_2949,N_2961);
nand UO_289 (O_289,N_2944,N_2971);
or UO_290 (O_290,N_2972,N_2941);
nor UO_291 (O_291,N_2949,N_2952);
nand UO_292 (O_292,N_2945,N_2993);
nor UO_293 (O_293,N_2950,N_2965);
and UO_294 (O_294,N_2973,N_2957);
nand UO_295 (O_295,N_2940,N_2944);
or UO_296 (O_296,N_2952,N_2976);
nor UO_297 (O_297,N_2972,N_2984);
or UO_298 (O_298,N_2955,N_2940);
nor UO_299 (O_299,N_2973,N_2959);
or UO_300 (O_300,N_2967,N_2946);
nor UO_301 (O_301,N_2964,N_2972);
and UO_302 (O_302,N_2977,N_2954);
nand UO_303 (O_303,N_2957,N_2953);
or UO_304 (O_304,N_2985,N_2945);
nand UO_305 (O_305,N_2974,N_2969);
xor UO_306 (O_306,N_2954,N_2996);
and UO_307 (O_307,N_2977,N_2997);
nand UO_308 (O_308,N_2949,N_2962);
xor UO_309 (O_309,N_2990,N_2963);
and UO_310 (O_310,N_2973,N_2997);
nand UO_311 (O_311,N_2976,N_2997);
nor UO_312 (O_312,N_2991,N_2944);
and UO_313 (O_313,N_2964,N_2981);
and UO_314 (O_314,N_2968,N_2958);
and UO_315 (O_315,N_2958,N_2998);
nand UO_316 (O_316,N_2968,N_2967);
nand UO_317 (O_317,N_2950,N_2951);
and UO_318 (O_318,N_2958,N_2996);
or UO_319 (O_319,N_2970,N_2969);
nand UO_320 (O_320,N_2961,N_2984);
nor UO_321 (O_321,N_2989,N_2960);
nand UO_322 (O_322,N_2960,N_2993);
nor UO_323 (O_323,N_2985,N_2979);
nor UO_324 (O_324,N_2964,N_2973);
nor UO_325 (O_325,N_2971,N_2982);
and UO_326 (O_326,N_2947,N_2961);
or UO_327 (O_327,N_2984,N_2945);
nor UO_328 (O_328,N_2973,N_2995);
nand UO_329 (O_329,N_2955,N_2963);
nor UO_330 (O_330,N_2956,N_2954);
nor UO_331 (O_331,N_2975,N_2960);
and UO_332 (O_332,N_2959,N_2945);
and UO_333 (O_333,N_2960,N_2987);
nand UO_334 (O_334,N_2960,N_2999);
and UO_335 (O_335,N_2983,N_2971);
or UO_336 (O_336,N_2953,N_2940);
nand UO_337 (O_337,N_2988,N_2986);
nor UO_338 (O_338,N_2953,N_2950);
or UO_339 (O_339,N_2998,N_2972);
nand UO_340 (O_340,N_2975,N_2963);
or UO_341 (O_341,N_2999,N_2958);
nor UO_342 (O_342,N_2942,N_2954);
nand UO_343 (O_343,N_2992,N_2965);
nor UO_344 (O_344,N_2984,N_2946);
and UO_345 (O_345,N_2952,N_2960);
nor UO_346 (O_346,N_2962,N_2994);
nand UO_347 (O_347,N_2943,N_2950);
or UO_348 (O_348,N_2972,N_2962);
nor UO_349 (O_349,N_2963,N_2982);
nor UO_350 (O_350,N_2954,N_2958);
and UO_351 (O_351,N_2973,N_2969);
nand UO_352 (O_352,N_2987,N_2969);
or UO_353 (O_353,N_2989,N_2955);
nand UO_354 (O_354,N_2998,N_2962);
and UO_355 (O_355,N_2985,N_2941);
or UO_356 (O_356,N_2971,N_2950);
or UO_357 (O_357,N_2950,N_2975);
and UO_358 (O_358,N_2948,N_2999);
nor UO_359 (O_359,N_2957,N_2961);
and UO_360 (O_360,N_2945,N_2955);
nand UO_361 (O_361,N_2989,N_2961);
nand UO_362 (O_362,N_2972,N_2996);
nor UO_363 (O_363,N_2949,N_2970);
nand UO_364 (O_364,N_2990,N_2959);
nor UO_365 (O_365,N_2996,N_2957);
nor UO_366 (O_366,N_2963,N_2974);
xor UO_367 (O_367,N_2954,N_2944);
and UO_368 (O_368,N_2976,N_2989);
nand UO_369 (O_369,N_2971,N_2963);
or UO_370 (O_370,N_2992,N_2940);
and UO_371 (O_371,N_2963,N_2967);
nor UO_372 (O_372,N_2990,N_2944);
nand UO_373 (O_373,N_2950,N_2941);
and UO_374 (O_374,N_2952,N_2965);
nor UO_375 (O_375,N_2942,N_2978);
nand UO_376 (O_376,N_2964,N_2970);
nor UO_377 (O_377,N_2955,N_2941);
xnor UO_378 (O_378,N_2948,N_2983);
or UO_379 (O_379,N_2985,N_2974);
or UO_380 (O_380,N_2943,N_2959);
or UO_381 (O_381,N_2964,N_2976);
or UO_382 (O_382,N_2947,N_2994);
nor UO_383 (O_383,N_2953,N_2959);
xor UO_384 (O_384,N_2997,N_2956);
xnor UO_385 (O_385,N_2941,N_2978);
and UO_386 (O_386,N_2948,N_2966);
or UO_387 (O_387,N_2973,N_2942);
nand UO_388 (O_388,N_2955,N_2994);
and UO_389 (O_389,N_2945,N_2947);
or UO_390 (O_390,N_2992,N_2995);
nand UO_391 (O_391,N_2957,N_2971);
or UO_392 (O_392,N_2985,N_2965);
or UO_393 (O_393,N_2976,N_2969);
and UO_394 (O_394,N_2964,N_2960);
nand UO_395 (O_395,N_2958,N_2993);
nor UO_396 (O_396,N_2982,N_2986);
nand UO_397 (O_397,N_2971,N_2953);
nand UO_398 (O_398,N_2976,N_2970);
and UO_399 (O_399,N_2967,N_2977);
nor UO_400 (O_400,N_2976,N_2999);
nor UO_401 (O_401,N_2959,N_2952);
nor UO_402 (O_402,N_2998,N_2977);
nand UO_403 (O_403,N_2944,N_2989);
or UO_404 (O_404,N_2943,N_2970);
nor UO_405 (O_405,N_2965,N_2973);
and UO_406 (O_406,N_2968,N_2987);
or UO_407 (O_407,N_2977,N_2944);
and UO_408 (O_408,N_2986,N_2947);
or UO_409 (O_409,N_2957,N_2997);
nor UO_410 (O_410,N_2991,N_2959);
nor UO_411 (O_411,N_2961,N_2950);
xor UO_412 (O_412,N_2979,N_2987);
nand UO_413 (O_413,N_2992,N_2974);
and UO_414 (O_414,N_2949,N_2958);
and UO_415 (O_415,N_2954,N_2976);
nor UO_416 (O_416,N_2945,N_2941);
or UO_417 (O_417,N_2958,N_2967);
or UO_418 (O_418,N_2976,N_2962);
or UO_419 (O_419,N_2999,N_2992);
nand UO_420 (O_420,N_2947,N_2943);
xor UO_421 (O_421,N_2973,N_2972);
nand UO_422 (O_422,N_2972,N_2958);
or UO_423 (O_423,N_2962,N_2946);
nor UO_424 (O_424,N_2973,N_2984);
or UO_425 (O_425,N_2969,N_2944);
or UO_426 (O_426,N_2986,N_2958);
and UO_427 (O_427,N_2942,N_2974);
and UO_428 (O_428,N_2980,N_2976);
nand UO_429 (O_429,N_2955,N_2978);
and UO_430 (O_430,N_2982,N_2968);
nand UO_431 (O_431,N_2969,N_2985);
nand UO_432 (O_432,N_2942,N_2967);
or UO_433 (O_433,N_2958,N_2945);
or UO_434 (O_434,N_2954,N_2987);
nand UO_435 (O_435,N_2982,N_2959);
or UO_436 (O_436,N_2967,N_2945);
and UO_437 (O_437,N_2974,N_2995);
nand UO_438 (O_438,N_2998,N_2988);
nor UO_439 (O_439,N_2994,N_2990);
nand UO_440 (O_440,N_2979,N_2999);
and UO_441 (O_441,N_2975,N_2959);
xnor UO_442 (O_442,N_2996,N_2998);
and UO_443 (O_443,N_2951,N_2959);
and UO_444 (O_444,N_2962,N_2990);
nand UO_445 (O_445,N_2945,N_2965);
or UO_446 (O_446,N_2990,N_2946);
and UO_447 (O_447,N_2984,N_2954);
nor UO_448 (O_448,N_2964,N_2958);
nor UO_449 (O_449,N_2957,N_2940);
nand UO_450 (O_450,N_2968,N_2946);
nand UO_451 (O_451,N_2979,N_2986);
nand UO_452 (O_452,N_2960,N_2963);
nand UO_453 (O_453,N_2990,N_2999);
or UO_454 (O_454,N_2996,N_2953);
or UO_455 (O_455,N_2982,N_2990);
nand UO_456 (O_456,N_2995,N_2952);
xor UO_457 (O_457,N_2969,N_2984);
nand UO_458 (O_458,N_2968,N_2985);
and UO_459 (O_459,N_2962,N_2984);
and UO_460 (O_460,N_2978,N_2995);
or UO_461 (O_461,N_2971,N_2975);
and UO_462 (O_462,N_2972,N_2986);
and UO_463 (O_463,N_2983,N_2998);
nor UO_464 (O_464,N_2980,N_2987);
or UO_465 (O_465,N_2963,N_2941);
nand UO_466 (O_466,N_2985,N_2940);
or UO_467 (O_467,N_2997,N_2995);
and UO_468 (O_468,N_2943,N_2983);
and UO_469 (O_469,N_2998,N_2968);
and UO_470 (O_470,N_2978,N_2989);
and UO_471 (O_471,N_2946,N_2987);
nor UO_472 (O_472,N_2949,N_2996);
nand UO_473 (O_473,N_2963,N_2992);
nor UO_474 (O_474,N_2968,N_2942);
or UO_475 (O_475,N_2942,N_2961);
and UO_476 (O_476,N_2973,N_2992);
nor UO_477 (O_477,N_2966,N_2984);
nor UO_478 (O_478,N_2967,N_2961);
nand UO_479 (O_479,N_2947,N_2987);
nor UO_480 (O_480,N_2954,N_2946);
nand UO_481 (O_481,N_2967,N_2994);
nor UO_482 (O_482,N_2989,N_2953);
or UO_483 (O_483,N_2981,N_2987);
or UO_484 (O_484,N_2941,N_2977);
or UO_485 (O_485,N_2957,N_2989);
nor UO_486 (O_486,N_2978,N_2976);
nor UO_487 (O_487,N_2948,N_2954);
or UO_488 (O_488,N_2960,N_2958);
nand UO_489 (O_489,N_2942,N_2970);
nand UO_490 (O_490,N_2973,N_2986);
nand UO_491 (O_491,N_2963,N_2970);
nor UO_492 (O_492,N_2995,N_2943);
nand UO_493 (O_493,N_2995,N_2986);
and UO_494 (O_494,N_2992,N_2966);
nand UO_495 (O_495,N_2983,N_2980);
nor UO_496 (O_496,N_2971,N_2987);
and UO_497 (O_497,N_2959,N_2964);
or UO_498 (O_498,N_2977,N_2984);
nand UO_499 (O_499,N_2985,N_2960);
endmodule