module basic_500_3000_500_5_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_287,In_164);
or U1 (N_1,In_68,In_418);
and U2 (N_2,In_489,In_170);
or U3 (N_3,In_254,In_342);
nand U4 (N_4,In_422,In_35);
nand U5 (N_5,In_497,In_385);
or U6 (N_6,In_340,In_33);
or U7 (N_7,In_350,In_114);
nand U8 (N_8,In_207,In_21);
nand U9 (N_9,In_144,In_393);
nor U10 (N_10,In_488,In_433);
and U11 (N_11,In_466,In_80);
nor U12 (N_12,In_183,In_267);
and U13 (N_13,In_362,In_237);
xor U14 (N_14,In_384,In_136);
and U15 (N_15,In_224,In_367);
or U16 (N_16,In_440,In_389);
and U17 (N_17,In_27,In_477);
and U18 (N_18,In_391,In_451);
or U19 (N_19,In_218,In_223);
xnor U20 (N_20,In_143,In_19);
xor U21 (N_21,In_409,In_402);
and U22 (N_22,In_438,In_354);
nor U23 (N_23,In_308,In_177);
nor U24 (N_24,In_394,In_448);
nor U25 (N_25,In_172,In_372);
and U26 (N_26,In_8,In_423);
or U27 (N_27,In_375,In_84);
xor U28 (N_28,In_386,In_127);
nand U29 (N_29,In_148,In_395);
or U30 (N_30,In_399,In_26);
nand U31 (N_31,In_61,In_91);
or U32 (N_32,In_62,In_307);
nor U33 (N_33,In_412,In_234);
and U34 (N_34,In_64,In_443);
xnor U35 (N_35,In_428,In_481);
or U36 (N_36,In_496,In_94);
or U37 (N_37,In_392,In_141);
and U38 (N_38,In_301,In_9);
and U39 (N_39,In_447,In_309);
xor U40 (N_40,In_231,In_12);
nand U41 (N_41,In_346,In_187);
nor U42 (N_42,In_321,In_390);
nand U43 (N_43,In_37,In_209);
or U44 (N_44,In_408,In_159);
xnor U45 (N_45,In_155,In_171);
and U46 (N_46,In_17,In_400);
or U47 (N_47,In_365,In_67);
xnor U48 (N_48,In_225,In_230);
or U49 (N_49,In_473,In_229);
xnor U50 (N_50,In_344,In_135);
and U51 (N_51,In_429,In_279);
nand U52 (N_52,In_458,In_405);
or U53 (N_53,In_269,In_194);
nand U54 (N_54,In_154,In_425);
and U55 (N_55,In_305,In_197);
nand U56 (N_56,In_388,In_191);
and U57 (N_57,In_174,In_180);
nor U58 (N_58,In_205,In_470);
xnor U59 (N_59,In_368,In_14);
or U60 (N_60,In_36,In_338);
or U61 (N_61,In_160,In_216);
or U62 (N_62,In_288,In_247);
or U63 (N_63,In_427,In_20);
xnor U64 (N_64,In_450,In_480);
xor U65 (N_65,In_414,In_461);
or U66 (N_66,In_168,In_292);
xnor U67 (N_67,In_356,In_485);
xor U68 (N_68,In_378,In_352);
nand U69 (N_69,In_252,In_289);
or U70 (N_70,In_30,In_283);
nand U71 (N_71,In_266,In_233);
nand U72 (N_72,In_272,In_7);
or U73 (N_73,In_430,In_286);
nand U74 (N_74,In_364,In_52);
or U75 (N_75,In_97,In_326);
or U76 (N_76,In_341,In_432);
nand U77 (N_77,In_472,In_157);
xnor U78 (N_78,In_436,In_328);
xor U79 (N_79,In_10,In_92);
or U80 (N_80,In_111,In_156);
and U81 (N_81,In_6,In_370);
nand U82 (N_82,In_398,In_406);
nand U83 (N_83,In_220,In_121);
xor U84 (N_84,In_351,In_208);
or U85 (N_85,In_163,In_119);
xor U86 (N_86,In_323,In_206);
and U87 (N_87,In_39,In_312);
or U88 (N_88,In_242,In_420);
or U89 (N_89,In_465,In_210);
xor U90 (N_90,In_235,In_474);
nor U91 (N_91,In_445,In_437);
nor U92 (N_92,In_484,In_302);
nand U93 (N_93,In_217,In_335);
xor U94 (N_94,In_416,In_181);
nand U95 (N_95,In_204,In_463);
nor U96 (N_96,In_34,In_349);
and U97 (N_97,In_81,In_322);
and U98 (N_98,In_40,In_494);
nand U99 (N_99,In_23,In_245);
nand U100 (N_100,In_435,In_101);
nor U101 (N_101,In_4,In_296);
nand U102 (N_102,In_401,In_357);
and U103 (N_103,In_125,In_250);
nor U104 (N_104,In_16,In_377);
xnor U105 (N_105,In_479,In_263);
nor U106 (N_106,In_31,In_417);
nand U107 (N_107,In_89,In_59);
nand U108 (N_108,In_201,In_434);
nand U109 (N_109,In_366,In_330);
or U110 (N_110,In_228,In_18);
xor U111 (N_111,In_293,In_495);
or U112 (N_112,In_1,In_190);
nor U113 (N_113,In_280,In_153);
xnor U114 (N_114,In_139,In_424);
xor U115 (N_115,In_345,In_32);
nor U116 (N_116,In_256,In_83);
nor U117 (N_117,In_195,In_70);
nor U118 (N_118,In_109,In_348);
xor U119 (N_119,In_277,In_469);
nor U120 (N_120,In_117,In_99);
nor U121 (N_121,In_215,In_452);
or U122 (N_122,In_490,In_358);
or U123 (N_123,In_100,In_381);
xnor U124 (N_124,In_306,In_442);
and U125 (N_125,In_145,In_189);
nand U126 (N_126,In_86,In_421);
nor U127 (N_127,In_222,In_66);
and U128 (N_128,In_123,In_238);
nor U129 (N_129,In_282,In_491);
nor U130 (N_130,In_53,In_161);
or U131 (N_131,In_38,In_104);
nand U132 (N_132,In_300,In_290);
and U133 (N_133,In_102,In_343);
or U134 (N_134,In_456,In_167);
or U135 (N_135,In_498,In_260);
and U136 (N_136,In_107,In_76);
or U137 (N_137,In_314,In_128);
xnor U138 (N_138,In_198,In_152);
xor U139 (N_139,In_98,In_446);
nor U140 (N_140,In_58,In_332);
nand U141 (N_141,In_202,In_82);
xor U142 (N_142,In_142,In_146);
or U143 (N_143,In_95,In_459);
and U144 (N_144,In_407,In_476);
nor U145 (N_145,In_15,In_361);
and U146 (N_146,In_151,In_2);
nor U147 (N_147,In_371,In_410);
or U148 (N_148,In_25,In_244);
and U149 (N_149,In_51,In_44);
or U150 (N_150,In_72,In_29);
or U151 (N_151,In_212,In_77);
or U152 (N_152,In_103,In_69);
nor U153 (N_153,In_105,In_298);
xor U154 (N_154,In_178,In_297);
nand U155 (N_155,In_96,In_219);
xor U156 (N_156,In_131,In_487);
or U157 (N_157,In_379,In_294);
or U158 (N_158,In_257,In_255);
xnor U159 (N_159,In_110,In_106);
xor U160 (N_160,In_325,In_24);
xnor U161 (N_161,In_65,In_457);
nand U162 (N_162,In_60,In_173);
or U163 (N_163,In_275,In_493);
and U164 (N_164,In_129,In_55);
and U165 (N_165,In_130,In_274);
or U166 (N_166,In_449,In_48);
nand U167 (N_167,In_241,In_134);
and U168 (N_168,In_45,In_369);
nand U169 (N_169,In_374,In_57);
or U170 (N_170,In_259,In_133);
nor U171 (N_171,In_382,In_320);
nand U172 (N_172,In_175,In_120);
or U173 (N_173,In_49,In_41);
xor U174 (N_174,In_213,In_108);
nand U175 (N_175,In_336,In_334);
nand U176 (N_176,In_380,In_486);
and U177 (N_177,In_79,In_415);
xnor U178 (N_178,In_196,In_192);
xor U179 (N_179,In_426,In_243);
xor U180 (N_180,In_471,In_253);
xor U181 (N_181,In_54,In_363);
nor U182 (N_182,In_87,In_271);
xnor U183 (N_183,In_453,In_179);
and U184 (N_184,In_132,In_310);
nand U185 (N_185,In_13,In_455);
nand U186 (N_186,In_158,In_124);
xnor U187 (N_187,In_118,In_295);
and U188 (N_188,In_318,In_444);
nand U189 (N_189,In_88,In_285);
xnor U190 (N_190,In_47,In_90);
and U191 (N_191,In_126,In_278);
xor U192 (N_192,In_193,In_147);
nor U193 (N_193,In_339,In_284);
or U194 (N_194,In_116,In_137);
or U195 (N_195,In_276,In_214);
xor U196 (N_196,In_478,In_211);
and U197 (N_197,In_93,In_236);
or U198 (N_198,In_258,In_387);
nand U199 (N_199,In_176,In_63);
and U200 (N_200,In_397,In_200);
xor U201 (N_201,In_264,In_475);
nor U202 (N_202,In_431,In_316);
xor U203 (N_203,In_28,In_22);
or U204 (N_204,In_221,In_439);
and U205 (N_205,In_319,In_186);
xor U206 (N_206,In_5,In_311);
nand U207 (N_207,In_337,In_331);
nor U208 (N_208,In_467,In_317);
xor U209 (N_209,In_0,In_75);
nand U210 (N_210,In_50,In_329);
nor U211 (N_211,In_441,In_246);
nor U212 (N_212,In_166,In_324);
nand U213 (N_213,In_71,In_138);
xnor U214 (N_214,In_268,In_383);
and U215 (N_215,In_353,In_199);
xor U216 (N_216,In_454,In_203);
and U217 (N_217,In_73,In_122);
xnor U218 (N_218,In_304,In_3);
xnor U219 (N_219,In_149,In_232);
nand U220 (N_220,In_227,In_419);
and U221 (N_221,In_468,In_376);
nand U222 (N_222,In_162,In_460);
nor U223 (N_223,In_413,In_403);
nand U224 (N_224,In_270,In_239);
nand U225 (N_225,In_188,In_373);
nand U226 (N_226,In_291,In_184);
or U227 (N_227,In_251,In_315);
and U228 (N_228,In_150,In_482);
nor U229 (N_229,In_85,In_273);
xor U230 (N_230,In_404,In_185);
nand U231 (N_231,In_43,In_226);
and U232 (N_232,In_140,In_299);
xnor U233 (N_233,In_281,In_56);
or U234 (N_234,In_262,In_359);
or U235 (N_235,In_78,In_333);
and U236 (N_236,In_360,In_115);
or U237 (N_237,In_492,In_303);
xnor U238 (N_238,In_248,In_499);
or U239 (N_239,In_313,In_42);
and U240 (N_240,In_240,In_327);
or U241 (N_241,In_11,In_464);
xor U242 (N_242,In_462,In_74);
or U243 (N_243,In_355,In_46);
nor U244 (N_244,In_396,In_483);
nor U245 (N_245,In_169,In_249);
nand U246 (N_246,In_261,In_182);
or U247 (N_247,In_265,In_112);
nor U248 (N_248,In_411,In_165);
nand U249 (N_249,In_113,In_347);
xor U250 (N_250,In_54,In_268);
and U251 (N_251,In_74,In_267);
or U252 (N_252,In_400,In_316);
and U253 (N_253,In_181,In_495);
nor U254 (N_254,In_19,In_351);
and U255 (N_255,In_428,In_376);
or U256 (N_256,In_322,In_142);
nor U257 (N_257,In_66,In_423);
or U258 (N_258,In_254,In_31);
and U259 (N_259,In_99,In_467);
xor U260 (N_260,In_165,In_281);
nand U261 (N_261,In_436,In_163);
xnor U262 (N_262,In_212,In_308);
nor U263 (N_263,In_0,In_387);
xnor U264 (N_264,In_246,In_216);
nand U265 (N_265,In_273,In_477);
xor U266 (N_266,In_99,In_296);
and U267 (N_267,In_352,In_143);
nor U268 (N_268,In_298,In_18);
xnor U269 (N_269,In_49,In_214);
nand U270 (N_270,In_245,In_330);
and U271 (N_271,In_487,In_483);
nand U272 (N_272,In_101,In_491);
and U273 (N_273,In_21,In_445);
xnor U274 (N_274,In_109,In_290);
or U275 (N_275,In_196,In_470);
or U276 (N_276,In_7,In_43);
and U277 (N_277,In_104,In_253);
nand U278 (N_278,In_447,In_16);
or U279 (N_279,In_80,In_114);
and U280 (N_280,In_138,In_385);
nor U281 (N_281,In_178,In_100);
or U282 (N_282,In_233,In_64);
xnor U283 (N_283,In_124,In_473);
xnor U284 (N_284,In_355,In_384);
and U285 (N_285,In_64,In_278);
or U286 (N_286,In_292,In_44);
nand U287 (N_287,In_390,In_447);
nand U288 (N_288,In_293,In_230);
nand U289 (N_289,In_369,In_481);
and U290 (N_290,In_146,In_246);
nor U291 (N_291,In_353,In_98);
xor U292 (N_292,In_181,In_178);
xnor U293 (N_293,In_228,In_134);
nand U294 (N_294,In_132,In_24);
xor U295 (N_295,In_98,In_141);
and U296 (N_296,In_494,In_193);
nor U297 (N_297,In_139,In_30);
or U298 (N_298,In_181,In_146);
and U299 (N_299,In_254,In_34);
xor U300 (N_300,In_439,In_241);
nand U301 (N_301,In_386,In_173);
nor U302 (N_302,In_133,In_160);
and U303 (N_303,In_165,In_481);
or U304 (N_304,In_476,In_227);
xor U305 (N_305,In_301,In_216);
or U306 (N_306,In_396,In_126);
or U307 (N_307,In_226,In_298);
or U308 (N_308,In_444,In_109);
and U309 (N_309,In_395,In_290);
nand U310 (N_310,In_96,In_439);
nor U311 (N_311,In_426,In_336);
nand U312 (N_312,In_451,In_240);
xnor U313 (N_313,In_8,In_100);
xor U314 (N_314,In_139,In_57);
or U315 (N_315,In_211,In_347);
and U316 (N_316,In_378,In_491);
xor U317 (N_317,In_416,In_98);
or U318 (N_318,In_450,In_255);
and U319 (N_319,In_361,In_124);
nor U320 (N_320,In_475,In_206);
or U321 (N_321,In_374,In_425);
nor U322 (N_322,In_103,In_239);
nand U323 (N_323,In_23,In_3);
nor U324 (N_324,In_302,In_94);
or U325 (N_325,In_52,In_233);
or U326 (N_326,In_52,In_193);
xnor U327 (N_327,In_391,In_253);
xnor U328 (N_328,In_138,In_369);
nor U329 (N_329,In_495,In_386);
nor U330 (N_330,In_67,In_465);
nor U331 (N_331,In_46,In_142);
nor U332 (N_332,In_83,In_308);
xor U333 (N_333,In_484,In_147);
xor U334 (N_334,In_286,In_314);
and U335 (N_335,In_386,In_359);
or U336 (N_336,In_20,In_493);
nand U337 (N_337,In_52,In_195);
xor U338 (N_338,In_136,In_367);
nor U339 (N_339,In_338,In_189);
nor U340 (N_340,In_140,In_417);
or U341 (N_341,In_210,In_437);
xnor U342 (N_342,In_10,In_474);
or U343 (N_343,In_104,In_131);
or U344 (N_344,In_311,In_473);
nand U345 (N_345,In_419,In_449);
and U346 (N_346,In_16,In_374);
and U347 (N_347,In_492,In_399);
nand U348 (N_348,In_62,In_301);
xnor U349 (N_349,In_60,In_420);
nor U350 (N_350,In_312,In_455);
or U351 (N_351,In_35,In_202);
or U352 (N_352,In_260,In_208);
xor U353 (N_353,In_166,In_258);
or U354 (N_354,In_379,In_104);
nor U355 (N_355,In_304,In_218);
or U356 (N_356,In_150,In_127);
nor U357 (N_357,In_29,In_82);
or U358 (N_358,In_320,In_175);
nand U359 (N_359,In_360,In_489);
xnor U360 (N_360,In_368,In_198);
or U361 (N_361,In_375,In_377);
or U362 (N_362,In_280,In_441);
and U363 (N_363,In_441,In_466);
or U364 (N_364,In_364,In_419);
or U365 (N_365,In_459,In_1);
nand U366 (N_366,In_52,In_455);
nor U367 (N_367,In_383,In_203);
nor U368 (N_368,In_157,In_455);
and U369 (N_369,In_198,In_267);
nor U370 (N_370,In_88,In_280);
nor U371 (N_371,In_375,In_63);
xnor U372 (N_372,In_433,In_109);
nor U373 (N_373,In_149,In_413);
nor U374 (N_374,In_368,In_173);
xnor U375 (N_375,In_496,In_60);
and U376 (N_376,In_374,In_402);
nor U377 (N_377,In_204,In_88);
xnor U378 (N_378,In_103,In_10);
and U379 (N_379,In_489,In_240);
xor U380 (N_380,In_412,In_119);
and U381 (N_381,In_381,In_40);
or U382 (N_382,In_304,In_277);
nor U383 (N_383,In_363,In_200);
nand U384 (N_384,In_263,In_495);
xnor U385 (N_385,In_108,In_39);
or U386 (N_386,In_115,In_287);
nand U387 (N_387,In_38,In_31);
or U388 (N_388,In_481,In_310);
nand U389 (N_389,In_314,In_130);
or U390 (N_390,In_143,In_139);
and U391 (N_391,In_372,In_279);
nor U392 (N_392,In_141,In_410);
or U393 (N_393,In_44,In_305);
and U394 (N_394,In_224,In_5);
or U395 (N_395,In_387,In_116);
nor U396 (N_396,In_5,In_317);
xor U397 (N_397,In_16,In_211);
or U398 (N_398,In_211,In_440);
and U399 (N_399,In_484,In_476);
xnor U400 (N_400,In_60,In_213);
nor U401 (N_401,In_209,In_283);
nor U402 (N_402,In_321,In_211);
and U403 (N_403,In_399,In_383);
or U404 (N_404,In_215,In_484);
xor U405 (N_405,In_167,In_352);
xor U406 (N_406,In_213,In_390);
xor U407 (N_407,In_66,In_296);
or U408 (N_408,In_284,In_244);
and U409 (N_409,In_243,In_432);
and U410 (N_410,In_133,In_263);
nor U411 (N_411,In_400,In_158);
nor U412 (N_412,In_233,In_326);
and U413 (N_413,In_76,In_1);
nand U414 (N_414,In_121,In_7);
nand U415 (N_415,In_200,In_469);
and U416 (N_416,In_127,In_279);
nor U417 (N_417,In_150,In_490);
nand U418 (N_418,In_122,In_346);
nand U419 (N_419,In_281,In_136);
nor U420 (N_420,In_334,In_245);
and U421 (N_421,In_356,In_495);
xnor U422 (N_422,In_450,In_193);
and U423 (N_423,In_100,In_270);
nor U424 (N_424,In_132,In_116);
nor U425 (N_425,In_477,In_479);
or U426 (N_426,In_294,In_263);
or U427 (N_427,In_475,In_305);
nor U428 (N_428,In_449,In_301);
and U429 (N_429,In_281,In_324);
xor U430 (N_430,In_443,In_50);
and U431 (N_431,In_170,In_313);
and U432 (N_432,In_135,In_36);
nand U433 (N_433,In_395,In_411);
or U434 (N_434,In_369,In_86);
and U435 (N_435,In_481,In_84);
or U436 (N_436,In_24,In_422);
and U437 (N_437,In_239,In_218);
xor U438 (N_438,In_28,In_307);
or U439 (N_439,In_402,In_460);
xnor U440 (N_440,In_183,In_260);
and U441 (N_441,In_182,In_429);
nand U442 (N_442,In_243,In_106);
or U443 (N_443,In_123,In_232);
nand U444 (N_444,In_334,In_322);
nand U445 (N_445,In_265,In_31);
or U446 (N_446,In_173,In_0);
and U447 (N_447,In_478,In_97);
nor U448 (N_448,In_13,In_495);
nand U449 (N_449,In_327,In_354);
xnor U450 (N_450,In_479,In_329);
xor U451 (N_451,In_458,In_189);
nor U452 (N_452,In_54,In_200);
nand U453 (N_453,In_328,In_207);
nor U454 (N_454,In_370,In_402);
and U455 (N_455,In_250,In_423);
xnor U456 (N_456,In_237,In_413);
nor U457 (N_457,In_342,In_115);
nor U458 (N_458,In_428,In_463);
nor U459 (N_459,In_467,In_447);
and U460 (N_460,In_68,In_232);
xor U461 (N_461,In_487,In_106);
nand U462 (N_462,In_23,In_458);
or U463 (N_463,In_300,In_77);
and U464 (N_464,In_281,In_300);
nor U465 (N_465,In_493,In_403);
nor U466 (N_466,In_423,In_248);
and U467 (N_467,In_204,In_170);
nor U468 (N_468,In_442,In_468);
nand U469 (N_469,In_240,In_257);
and U470 (N_470,In_296,In_409);
nand U471 (N_471,In_445,In_284);
or U472 (N_472,In_82,In_60);
and U473 (N_473,In_185,In_490);
or U474 (N_474,In_277,In_284);
xnor U475 (N_475,In_173,In_306);
or U476 (N_476,In_79,In_485);
and U477 (N_477,In_351,In_469);
or U478 (N_478,In_416,In_372);
and U479 (N_479,In_259,In_141);
or U480 (N_480,In_426,In_492);
and U481 (N_481,In_353,In_466);
nand U482 (N_482,In_229,In_421);
and U483 (N_483,In_468,In_361);
or U484 (N_484,In_110,In_166);
nor U485 (N_485,In_425,In_98);
nor U486 (N_486,In_239,In_363);
nor U487 (N_487,In_262,In_207);
or U488 (N_488,In_47,In_365);
or U489 (N_489,In_411,In_148);
and U490 (N_490,In_341,In_191);
nand U491 (N_491,In_16,In_194);
nand U492 (N_492,In_80,In_264);
and U493 (N_493,In_182,In_165);
and U494 (N_494,In_31,In_10);
or U495 (N_495,In_258,In_366);
and U496 (N_496,In_496,In_106);
or U497 (N_497,In_157,In_467);
and U498 (N_498,In_71,In_494);
and U499 (N_499,In_68,In_429);
nor U500 (N_500,In_356,In_354);
and U501 (N_501,In_198,In_178);
or U502 (N_502,In_40,In_193);
nor U503 (N_503,In_109,In_436);
nand U504 (N_504,In_378,In_69);
or U505 (N_505,In_156,In_398);
or U506 (N_506,In_380,In_438);
xor U507 (N_507,In_168,In_76);
nand U508 (N_508,In_399,In_250);
xor U509 (N_509,In_226,In_200);
or U510 (N_510,In_430,In_94);
xnor U511 (N_511,In_366,In_114);
or U512 (N_512,In_425,In_169);
xnor U513 (N_513,In_437,In_243);
nand U514 (N_514,In_49,In_121);
nand U515 (N_515,In_27,In_270);
and U516 (N_516,In_407,In_43);
or U517 (N_517,In_142,In_84);
nand U518 (N_518,In_158,In_157);
nor U519 (N_519,In_463,In_64);
or U520 (N_520,In_471,In_360);
nor U521 (N_521,In_407,In_131);
nor U522 (N_522,In_164,In_172);
or U523 (N_523,In_312,In_113);
xor U524 (N_524,In_273,In_150);
or U525 (N_525,In_283,In_438);
nand U526 (N_526,In_106,In_399);
or U527 (N_527,In_111,In_217);
and U528 (N_528,In_437,In_254);
nand U529 (N_529,In_83,In_341);
and U530 (N_530,In_221,In_405);
and U531 (N_531,In_30,In_289);
and U532 (N_532,In_282,In_107);
nor U533 (N_533,In_220,In_328);
nand U534 (N_534,In_185,In_402);
and U535 (N_535,In_198,In_223);
or U536 (N_536,In_489,In_322);
xor U537 (N_537,In_103,In_268);
nor U538 (N_538,In_57,In_280);
nor U539 (N_539,In_187,In_447);
nand U540 (N_540,In_427,In_243);
and U541 (N_541,In_98,In_308);
or U542 (N_542,In_171,In_247);
or U543 (N_543,In_466,In_112);
nor U544 (N_544,In_364,In_149);
nor U545 (N_545,In_368,In_109);
xor U546 (N_546,In_46,In_164);
xnor U547 (N_547,In_229,In_148);
nor U548 (N_548,In_289,In_350);
nor U549 (N_549,In_220,In_332);
nand U550 (N_550,In_148,In_172);
nor U551 (N_551,In_310,In_206);
or U552 (N_552,In_484,In_120);
nor U553 (N_553,In_139,In_487);
nor U554 (N_554,In_7,In_497);
nand U555 (N_555,In_234,In_0);
or U556 (N_556,In_395,In_297);
nor U557 (N_557,In_184,In_417);
nor U558 (N_558,In_495,In_73);
nand U559 (N_559,In_477,In_183);
nor U560 (N_560,In_102,In_119);
xnor U561 (N_561,In_9,In_65);
nand U562 (N_562,In_63,In_29);
and U563 (N_563,In_60,In_230);
xor U564 (N_564,In_384,In_420);
nor U565 (N_565,In_360,In_261);
and U566 (N_566,In_423,In_245);
nor U567 (N_567,In_146,In_251);
and U568 (N_568,In_224,In_50);
and U569 (N_569,In_288,In_128);
nand U570 (N_570,In_207,In_195);
nor U571 (N_571,In_186,In_57);
or U572 (N_572,In_172,In_316);
xor U573 (N_573,In_294,In_449);
nand U574 (N_574,In_382,In_431);
nor U575 (N_575,In_390,In_193);
nand U576 (N_576,In_80,In_423);
and U577 (N_577,In_265,In_206);
xor U578 (N_578,In_389,In_447);
xnor U579 (N_579,In_352,In_304);
xnor U580 (N_580,In_344,In_487);
xor U581 (N_581,In_374,In_111);
or U582 (N_582,In_186,In_182);
and U583 (N_583,In_74,In_327);
and U584 (N_584,In_126,In_168);
nand U585 (N_585,In_247,In_59);
or U586 (N_586,In_295,In_388);
xnor U587 (N_587,In_10,In_486);
xnor U588 (N_588,In_432,In_197);
or U589 (N_589,In_480,In_231);
nor U590 (N_590,In_188,In_436);
and U591 (N_591,In_490,In_459);
and U592 (N_592,In_280,In_497);
xnor U593 (N_593,In_429,In_358);
or U594 (N_594,In_187,In_62);
nor U595 (N_595,In_38,In_197);
nor U596 (N_596,In_30,In_457);
and U597 (N_597,In_199,In_160);
nand U598 (N_598,In_311,In_343);
xnor U599 (N_599,In_386,In_465);
and U600 (N_600,N_65,N_462);
and U601 (N_601,N_72,N_475);
nand U602 (N_602,N_530,N_409);
xor U603 (N_603,N_471,N_46);
xor U604 (N_604,N_196,N_287);
nand U605 (N_605,N_386,N_436);
xor U606 (N_606,N_33,N_428);
xor U607 (N_607,N_396,N_402);
and U608 (N_608,N_239,N_414);
xor U609 (N_609,N_96,N_417);
nor U610 (N_610,N_551,N_218);
nor U611 (N_611,N_264,N_518);
or U612 (N_612,N_511,N_103);
or U613 (N_613,N_464,N_589);
nand U614 (N_614,N_17,N_482);
or U615 (N_615,N_419,N_274);
nand U616 (N_616,N_582,N_523);
nor U617 (N_617,N_398,N_435);
or U618 (N_618,N_496,N_517);
nand U619 (N_619,N_459,N_413);
xnor U620 (N_620,N_294,N_463);
nor U621 (N_621,N_584,N_217);
and U622 (N_622,N_32,N_19);
nor U623 (N_623,N_83,N_315);
nand U624 (N_624,N_240,N_524);
or U625 (N_625,N_140,N_451);
nor U626 (N_626,N_539,N_429);
or U627 (N_627,N_534,N_44);
xor U628 (N_628,N_380,N_10);
nand U629 (N_629,N_59,N_329);
nor U630 (N_630,N_228,N_452);
nand U631 (N_631,N_8,N_61);
nand U632 (N_632,N_559,N_194);
nor U633 (N_633,N_123,N_467);
nor U634 (N_634,N_245,N_576);
and U635 (N_635,N_260,N_591);
xnor U636 (N_636,N_388,N_62);
nor U637 (N_637,N_1,N_349);
or U638 (N_638,N_331,N_531);
nand U639 (N_639,N_420,N_197);
and U640 (N_640,N_312,N_105);
xor U641 (N_641,N_495,N_49);
xor U642 (N_642,N_535,N_439);
and U643 (N_643,N_195,N_512);
nor U644 (N_644,N_509,N_7);
xnor U645 (N_645,N_401,N_204);
nand U646 (N_646,N_433,N_290);
or U647 (N_647,N_541,N_16);
nor U648 (N_648,N_53,N_106);
and U649 (N_649,N_416,N_492);
nor U650 (N_650,N_11,N_24);
xor U651 (N_651,N_514,N_368);
and U652 (N_652,N_100,N_599);
or U653 (N_653,N_48,N_30);
xor U654 (N_654,N_18,N_596);
or U655 (N_655,N_45,N_389);
nor U656 (N_656,N_552,N_441);
and U657 (N_657,N_450,N_164);
and U658 (N_658,N_126,N_288);
xnor U659 (N_659,N_366,N_483);
or U660 (N_660,N_200,N_494);
nor U661 (N_661,N_285,N_157);
xnor U662 (N_662,N_47,N_281);
nand U663 (N_663,N_387,N_493);
nor U664 (N_664,N_359,N_58);
xor U665 (N_665,N_588,N_360);
xor U666 (N_666,N_491,N_310);
or U667 (N_667,N_77,N_379);
nand U668 (N_668,N_256,N_15);
and U669 (N_669,N_51,N_305);
or U670 (N_670,N_567,N_598);
nand U671 (N_671,N_585,N_262);
nor U672 (N_672,N_527,N_333);
nand U673 (N_673,N_469,N_258);
nand U674 (N_674,N_377,N_532);
or U675 (N_675,N_302,N_374);
xor U676 (N_676,N_298,N_4);
nand U677 (N_677,N_587,N_507);
xor U678 (N_678,N_460,N_533);
and U679 (N_679,N_201,N_519);
xnor U680 (N_680,N_313,N_537);
and U681 (N_681,N_23,N_131);
xnor U682 (N_682,N_210,N_267);
and U683 (N_683,N_146,N_573);
xnor U684 (N_684,N_253,N_306);
and U685 (N_685,N_373,N_248);
or U686 (N_686,N_352,N_52);
nor U687 (N_687,N_521,N_251);
and U688 (N_688,N_544,N_309);
or U689 (N_689,N_138,N_236);
or U690 (N_690,N_406,N_390);
xnor U691 (N_691,N_430,N_74);
nand U692 (N_692,N_297,N_391);
and U693 (N_693,N_299,N_508);
xnor U694 (N_694,N_6,N_479);
or U695 (N_695,N_27,N_367);
and U696 (N_696,N_487,N_295);
or U697 (N_697,N_14,N_421);
xor U698 (N_698,N_89,N_37);
and U699 (N_699,N_142,N_229);
nor U700 (N_700,N_209,N_80);
nand U701 (N_701,N_449,N_415);
xor U702 (N_702,N_453,N_268);
nand U703 (N_703,N_246,N_81);
xnor U704 (N_704,N_120,N_163);
nor U705 (N_705,N_199,N_43);
nor U706 (N_706,N_597,N_321);
nand U707 (N_707,N_147,N_92);
nor U708 (N_708,N_124,N_443);
or U709 (N_709,N_226,N_590);
xnor U710 (N_710,N_134,N_404);
nand U711 (N_711,N_102,N_350);
xor U712 (N_712,N_176,N_444);
or U713 (N_713,N_474,N_136);
nand U714 (N_714,N_500,N_456);
nand U715 (N_715,N_183,N_91);
xor U716 (N_716,N_107,N_108);
xor U717 (N_717,N_580,N_446);
nand U718 (N_718,N_381,N_98);
nand U719 (N_719,N_113,N_568);
and U720 (N_720,N_562,N_181);
nor U721 (N_721,N_144,N_238);
nand U722 (N_722,N_411,N_31);
and U723 (N_723,N_277,N_270);
nand U724 (N_724,N_498,N_472);
or U725 (N_725,N_93,N_161);
nor U726 (N_726,N_426,N_536);
nand U727 (N_727,N_528,N_520);
and U728 (N_728,N_340,N_121);
nor U729 (N_729,N_154,N_9);
or U730 (N_730,N_445,N_280);
xor U731 (N_731,N_3,N_114);
or U732 (N_732,N_431,N_484);
or U733 (N_733,N_579,N_364);
and U734 (N_734,N_328,N_110);
and U735 (N_735,N_5,N_119);
xnor U736 (N_736,N_334,N_137);
nand U737 (N_737,N_75,N_455);
and U738 (N_738,N_82,N_88);
nand U739 (N_739,N_526,N_499);
nor U740 (N_740,N_172,N_221);
nor U741 (N_741,N_68,N_203);
nand U742 (N_742,N_595,N_90);
or U743 (N_743,N_423,N_546);
nor U744 (N_744,N_447,N_322);
and U745 (N_745,N_87,N_501);
nor U746 (N_746,N_362,N_506);
nor U747 (N_747,N_12,N_545);
xor U748 (N_748,N_522,N_156);
nand U749 (N_749,N_178,N_357);
or U750 (N_750,N_468,N_189);
or U751 (N_751,N_242,N_99);
nor U752 (N_752,N_291,N_224);
or U753 (N_753,N_454,N_478);
and U754 (N_754,N_410,N_515);
nand U755 (N_755,N_529,N_177);
and U756 (N_756,N_564,N_561);
and U757 (N_757,N_345,N_505);
nand U758 (N_758,N_132,N_319);
nor U759 (N_759,N_572,N_35);
nand U760 (N_760,N_66,N_489);
or U761 (N_761,N_307,N_555);
nor U762 (N_762,N_158,N_198);
nand U763 (N_763,N_525,N_21);
xor U764 (N_764,N_570,N_97);
and U765 (N_765,N_205,N_293);
and U766 (N_766,N_575,N_351);
and U767 (N_767,N_143,N_41);
nor U768 (N_768,N_42,N_261);
and U769 (N_769,N_438,N_314);
or U770 (N_770,N_193,N_278);
xnor U771 (N_771,N_399,N_392);
xnor U772 (N_772,N_407,N_286);
or U773 (N_773,N_141,N_273);
or U774 (N_774,N_272,N_67);
or U775 (N_775,N_13,N_486);
and U776 (N_776,N_271,N_202);
xnor U777 (N_777,N_481,N_540);
or U778 (N_778,N_332,N_64);
nor U779 (N_779,N_466,N_227);
nand U780 (N_780,N_476,N_342);
nor U781 (N_781,N_384,N_40);
or U782 (N_782,N_247,N_234);
nand U783 (N_783,N_289,N_275);
and U784 (N_784,N_583,N_369);
or U785 (N_785,N_155,N_29);
and U786 (N_786,N_382,N_422);
nand U787 (N_787,N_71,N_465);
and U788 (N_788,N_424,N_578);
nor U789 (N_789,N_324,N_111);
nand U790 (N_790,N_112,N_296);
or U791 (N_791,N_300,N_152);
and U792 (N_792,N_173,N_383);
nor U793 (N_793,N_337,N_554);
or U794 (N_794,N_222,N_473);
nor U795 (N_795,N_361,N_316);
xnor U796 (N_796,N_346,N_115);
nor U797 (N_797,N_581,N_553);
nor U798 (N_798,N_403,N_513);
nand U799 (N_799,N_393,N_57);
nand U800 (N_800,N_348,N_243);
and U801 (N_801,N_254,N_263);
and U802 (N_802,N_442,N_510);
or U803 (N_803,N_470,N_214);
and U804 (N_804,N_212,N_179);
or U805 (N_805,N_170,N_558);
or U806 (N_806,N_418,N_569);
nand U807 (N_807,N_125,N_25);
xor U808 (N_808,N_38,N_215);
xnor U809 (N_809,N_353,N_265);
or U810 (N_810,N_548,N_320);
nor U811 (N_811,N_405,N_190);
nor U812 (N_812,N_542,N_150);
nand U813 (N_813,N_175,N_192);
xor U814 (N_814,N_184,N_394);
nor U815 (N_815,N_358,N_104);
xor U816 (N_816,N_148,N_437);
nor U817 (N_817,N_308,N_412);
xnor U818 (N_818,N_318,N_371);
nor U819 (N_819,N_376,N_76);
and U820 (N_820,N_84,N_241);
or U821 (N_821,N_237,N_266);
or U822 (N_822,N_169,N_344);
xnor U823 (N_823,N_211,N_127);
nor U824 (N_824,N_168,N_182);
nor U825 (N_825,N_480,N_165);
or U826 (N_826,N_327,N_325);
xor U827 (N_827,N_118,N_69);
nor U828 (N_828,N_26,N_223);
nand U829 (N_829,N_370,N_504);
xor U830 (N_830,N_355,N_130);
nor U831 (N_831,N_101,N_180);
nand U832 (N_832,N_220,N_216);
nand U833 (N_833,N_94,N_341);
xnor U834 (N_834,N_28,N_231);
and U835 (N_835,N_206,N_70);
or U836 (N_836,N_135,N_86);
xor U837 (N_837,N_55,N_257);
nor U838 (N_838,N_60,N_339);
xnor U839 (N_839,N_282,N_503);
xnor U840 (N_840,N_485,N_365);
nand U841 (N_841,N_385,N_276);
nand U842 (N_842,N_160,N_249);
or U843 (N_843,N_593,N_188);
nand U844 (N_844,N_162,N_39);
nor U845 (N_845,N_284,N_232);
and U846 (N_846,N_149,N_85);
xnor U847 (N_847,N_372,N_323);
and U848 (N_848,N_233,N_303);
nand U849 (N_849,N_2,N_255);
or U850 (N_850,N_252,N_129);
or U851 (N_851,N_457,N_95);
and U852 (N_852,N_317,N_347);
and U853 (N_853,N_538,N_434);
xnor U854 (N_854,N_448,N_171);
nand U855 (N_855,N_283,N_574);
xor U856 (N_856,N_225,N_54);
and U857 (N_857,N_34,N_311);
or U858 (N_858,N_36,N_207);
or U859 (N_859,N_326,N_185);
xor U860 (N_860,N_73,N_354);
or U861 (N_861,N_244,N_556);
and U862 (N_862,N_79,N_56);
nor U863 (N_863,N_139,N_116);
and U864 (N_864,N_269,N_235);
and U865 (N_865,N_477,N_490);
nor U866 (N_866,N_378,N_565);
xor U867 (N_867,N_458,N_63);
or U868 (N_868,N_336,N_547);
nor U869 (N_869,N_122,N_586);
or U870 (N_870,N_167,N_400);
nand U871 (N_871,N_592,N_128);
or U872 (N_872,N_440,N_166);
and U873 (N_873,N_488,N_549);
or U874 (N_874,N_566,N_50);
nand U875 (N_875,N_159,N_230);
and U876 (N_876,N_153,N_279);
nand U877 (N_877,N_594,N_151);
xnor U878 (N_878,N_117,N_497);
and U879 (N_879,N_408,N_109);
nor U880 (N_880,N_145,N_375);
xor U881 (N_881,N_250,N_577);
nand U882 (N_882,N_550,N_343);
xnor U883 (N_883,N_461,N_427);
or U884 (N_884,N_191,N_363);
and U885 (N_885,N_356,N_571);
nand U886 (N_886,N_208,N_395);
or U887 (N_887,N_304,N_335);
xnor U888 (N_888,N_133,N_219);
nor U889 (N_889,N_563,N_557);
nor U890 (N_890,N_174,N_543);
and U891 (N_891,N_0,N_432);
nor U892 (N_892,N_397,N_425);
nand U893 (N_893,N_516,N_502);
nand U894 (N_894,N_292,N_22);
and U895 (N_895,N_186,N_187);
xor U896 (N_896,N_213,N_259);
nand U897 (N_897,N_560,N_338);
nor U898 (N_898,N_330,N_78);
nor U899 (N_899,N_301,N_20);
or U900 (N_900,N_68,N_401);
xor U901 (N_901,N_514,N_546);
nor U902 (N_902,N_511,N_149);
and U903 (N_903,N_121,N_384);
xor U904 (N_904,N_376,N_398);
or U905 (N_905,N_265,N_317);
and U906 (N_906,N_439,N_576);
xor U907 (N_907,N_560,N_308);
nand U908 (N_908,N_422,N_171);
nor U909 (N_909,N_592,N_166);
nand U910 (N_910,N_363,N_494);
nand U911 (N_911,N_583,N_353);
nand U912 (N_912,N_334,N_325);
nor U913 (N_913,N_543,N_166);
xnor U914 (N_914,N_379,N_576);
or U915 (N_915,N_285,N_458);
or U916 (N_916,N_276,N_201);
nor U917 (N_917,N_326,N_496);
nand U918 (N_918,N_19,N_183);
xnor U919 (N_919,N_147,N_126);
xor U920 (N_920,N_8,N_11);
nor U921 (N_921,N_531,N_44);
or U922 (N_922,N_299,N_323);
nor U923 (N_923,N_11,N_386);
and U924 (N_924,N_331,N_248);
nand U925 (N_925,N_434,N_420);
xor U926 (N_926,N_114,N_39);
nand U927 (N_927,N_227,N_307);
xor U928 (N_928,N_134,N_587);
or U929 (N_929,N_458,N_517);
xnor U930 (N_930,N_305,N_162);
nor U931 (N_931,N_427,N_107);
nand U932 (N_932,N_96,N_200);
or U933 (N_933,N_58,N_332);
and U934 (N_934,N_258,N_248);
nor U935 (N_935,N_494,N_463);
nand U936 (N_936,N_180,N_146);
nor U937 (N_937,N_87,N_404);
nor U938 (N_938,N_517,N_167);
and U939 (N_939,N_61,N_29);
nor U940 (N_940,N_582,N_592);
nand U941 (N_941,N_102,N_485);
xnor U942 (N_942,N_363,N_435);
nor U943 (N_943,N_452,N_20);
xnor U944 (N_944,N_319,N_34);
xnor U945 (N_945,N_131,N_508);
and U946 (N_946,N_286,N_564);
or U947 (N_947,N_317,N_597);
and U948 (N_948,N_313,N_440);
nor U949 (N_949,N_182,N_23);
nor U950 (N_950,N_272,N_119);
xnor U951 (N_951,N_181,N_168);
xnor U952 (N_952,N_80,N_334);
xor U953 (N_953,N_493,N_146);
xnor U954 (N_954,N_526,N_283);
nand U955 (N_955,N_307,N_396);
or U956 (N_956,N_502,N_216);
or U957 (N_957,N_312,N_129);
or U958 (N_958,N_29,N_469);
nor U959 (N_959,N_506,N_234);
or U960 (N_960,N_464,N_415);
and U961 (N_961,N_72,N_441);
xor U962 (N_962,N_147,N_355);
nand U963 (N_963,N_339,N_18);
and U964 (N_964,N_341,N_517);
and U965 (N_965,N_214,N_541);
nor U966 (N_966,N_547,N_576);
or U967 (N_967,N_241,N_8);
or U968 (N_968,N_239,N_39);
xor U969 (N_969,N_44,N_325);
xnor U970 (N_970,N_86,N_478);
xor U971 (N_971,N_301,N_103);
and U972 (N_972,N_541,N_121);
xor U973 (N_973,N_424,N_313);
nor U974 (N_974,N_490,N_273);
nor U975 (N_975,N_163,N_562);
xnor U976 (N_976,N_119,N_327);
and U977 (N_977,N_568,N_571);
nor U978 (N_978,N_478,N_140);
xor U979 (N_979,N_404,N_591);
or U980 (N_980,N_304,N_546);
xnor U981 (N_981,N_412,N_49);
nand U982 (N_982,N_501,N_34);
nor U983 (N_983,N_317,N_480);
xor U984 (N_984,N_509,N_519);
nand U985 (N_985,N_363,N_226);
and U986 (N_986,N_203,N_250);
nand U987 (N_987,N_379,N_409);
nor U988 (N_988,N_558,N_166);
and U989 (N_989,N_65,N_253);
and U990 (N_990,N_18,N_279);
nand U991 (N_991,N_538,N_457);
xor U992 (N_992,N_448,N_235);
and U993 (N_993,N_82,N_192);
nand U994 (N_994,N_17,N_228);
xnor U995 (N_995,N_553,N_141);
and U996 (N_996,N_138,N_35);
nand U997 (N_997,N_128,N_499);
and U998 (N_998,N_179,N_348);
nand U999 (N_999,N_345,N_555);
nor U1000 (N_1000,N_468,N_5);
or U1001 (N_1001,N_64,N_194);
xor U1002 (N_1002,N_184,N_294);
nor U1003 (N_1003,N_403,N_494);
or U1004 (N_1004,N_375,N_265);
or U1005 (N_1005,N_513,N_223);
and U1006 (N_1006,N_271,N_181);
or U1007 (N_1007,N_194,N_510);
nor U1008 (N_1008,N_545,N_289);
xor U1009 (N_1009,N_348,N_214);
xnor U1010 (N_1010,N_181,N_374);
nor U1011 (N_1011,N_309,N_530);
and U1012 (N_1012,N_219,N_123);
and U1013 (N_1013,N_35,N_33);
and U1014 (N_1014,N_473,N_42);
nor U1015 (N_1015,N_583,N_211);
xnor U1016 (N_1016,N_418,N_200);
nor U1017 (N_1017,N_325,N_443);
nand U1018 (N_1018,N_202,N_5);
nand U1019 (N_1019,N_153,N_518);
xor U1020 (N_1020,N_202,N_424);
and U1021 (N_1021,N_138,N_25);
xnor U1022 (N_1022,N_484,N_243);
nor U1023 (N_1023,N_198,N_543);
nand U1024 (N_1024,N_70,N_469);
xnor U1025 (N_1025,N_497,N_538);
nand U1026 (N_1026,N_18,N_449);
nor U1027 (N_1027,N_80,N_397);
or U1028 (N_1028,N_40,N_12);
and U1029 (N_1029,N_321,N_401);
xor U1030 (N_1030,N_92,N_223);
nor U1031 (N_1031,N_309,N_406);
and U1032 (N_1032,N_52,N_360);
nor U1033 (N_1033,N_328,N_180);
xor U1034 (N_1034,N_140,N_27);
xnor U1035 (N_1035,N_385,N_467);
nor U1036 (N_1036,N_358,N_318);
nor U1037 (N_1037,N_262,N_47);
nor U1038 (N_1038,N_66,N_250);
nand U1039 (N_1039,N_210,N_216);
nor U1040 (N_1040,N_542,N_133);
and U1041 (N_1041,N_214,N_443);
and U1042 (N_1042,N_275,N_422);
nor U1043 (N_1043,N_233,N_271);
or U1044 (N_1044,N_551,N_538);
nand U1045 (N_1045,N_166,N_544);
xor U1046 (N_1046,N_187,N_129);
nand U1047 (N_1047,N_88,N_33);
nor U1048 (N_1048,N_377,N_479);
xor U1049 (N_1049,N_179,N_214);
xnor U1050 (N_1050,N_178,N_503);
and U1051 (N_1051,N_223,N_393);
and U1052 (N_1052,N_419,N_598);
and U1053 (N_1053,N_18,N_282);
nand U1054 (N_1054,N_56,N_500);
or U1055 (N_1055,N_244,N_557);
and U1056 (N_1056,N_382,N_194);
or U1057 (N_1057,N_168,N_34);
nand U1058 (N_1058,N_16,N_366);
or U1059 (N_1059,N_48,N_378);
nand U1060 (N_1060,N_201,N_526);
or U1061 (N_1061,N_151,N_292);
or U1062 (N_1062,N_355,N_597);
nand U1063 (N_1063,N_445,N_540);
xnor U1064 (N_1064,N_345,N_224);
xor U1065 (N_1065,N_559,N_491);
nand U1066 (N_1066,N_28,N_286);
nor U1067 (N_1067,N_126,N_343);
or U1068 (N_1068,N_18,N_437);
xor U1069 (N_1069,N_379,N_16);
nand U1070 (N_1070,N_82,N_400);
nand U1071 (N_1071,N_273,N_103);
nand U1072 (N_1072,N_518,N_297);
nor U1073 (N_1073,N_173,N_585);
nand U1074 (N_1074,N_72,N_208);
and U1075 (N_1075,N_20,N_575);
nand U1076 (N_1076,N_150,N_496);
or U1077 (N_1077,N_128,N_278);
nor U1078 (N_1078,N_60,N_587);
xor U1079 (N_1079,N_371,N_224);
and U1080 (N_1080,N_467,N_489);
and U1081 (N_1081,N_467,N_484);
and U1082 (N_1082,N_294,N_304);
nand U1083 (N_1083,N_185,N_315);
or U1084 (N_1084,N_449,N_359);
nor U1085 (N_1085,N_540,N_287);
nor U1086 (N_1086,N_180,N_197);
nand U1087 (N_1087,N_448,N_450);
and U1088 (N_1088,N_303,N_507);
nor U1089 (N_1089,N_28,N_288);
xor U1090 (N_1090,N_487,N_483);
xor U1091 (N_1091,N_395,N_94);
nor U1092 (N_1092,N_524,N_587);
nand U1093 (N_1093,N_240,N_62);
nand U1094 (N_1094,N_510,N_390);
and U1095 (N_1095,N_572,N_177);
xnor U1096 (N_1096,N_373,N_579);
nor U1097 (N_1097,N_229,N_517);
or U1098 (N_1098,N_290,N_143);
nor U1099 (N_1099,N_32,N_483);
nor U1100 (N_1100,N_233,N_510);
nor U1101 (N_1101,N_35,N_225);
nand U1102 (N_1102,N_342,N_44);
and U1103 (N_1103,N_243,N_397);
xnor U1104 (N_1104,N_598,N_560);
nand U1105 (N_1105,N_496,N_555);
xor U1106 (N_1106,N_225,N_489);
nand U1107 (N_1107,N_187,N_154);
xnor U1108 (N_1108,N_518,N_599);
or U1109 (N_1109,N_502,N_583);
and U1110 (N_1110,N_482,N_450);
nand U1111 (N_1111,N_344,N_1);
nor U1112 (N_1112,N_519,N_27);
xnor U1113 (N_1113,N_468,N_238);
xor U1114 (N_1114,N_306,N_4);
and U1115 (N_1115,N_478,N_414);
and U1116 (N_1116,N_379,N_64);
nor U1117 (N_1117,N_362,N_190);
xor U1118 (N_1118,N_458,N_475);
nand U1119 (N_1119,N_320,N_569);
nor U1120 (N_1120,N_291,N_335);
and U1121 (N_1121,N_28,N_479);
nor U1122 (N_1122,N_593,N_89);
nor U1123 (N_1123,N_60,N_407);
or U1124 (N_1124,N_451,N_410);
xnor U1125 (N_1125,N_127,N_117);
nand U1126 (N_1126,N_265,N_333);
nor U1127 (N_1127,N_159,N_148);
or U1128 (N_1128,N_231,N_159);
or U1129 (N_1129,N_215,N_166);
xor U1130 (N_1130,N_59,N_461);
nor U1131 (N_1131,N_403,N_566);
or U1132 (N_1132,N_259,N_242);
and U1133 (N_1133,N_232,N_570);
nand U1134 (N_1134,N_216,N_81);
nor U1135 (N_1135,N_169,N_279);
and U1136 (N_1136,N_38,N_156);
nor U1137 (N_1137,N_429,N_244);
or U1138 (N_1138,N_258,N_70);
nor U1139 (N_1139,N_217,N_331);
xnor U1140 (N_1140,N_509,N_261);
nand U1141 (N_1141,N_555,N_329);
nand U1142 (N_1142,N_564,N_81);
xor U1143 (N_1143,N_329,N_35);
nor U1144 (N_1144,N_110,N_342);
nor U1145 (N_1145,N_420,N_383);
xnor U1146 (N_1146,N_180,N_112);
and U1147 (N_1147,N_288,N_157);
or U1148 (N_1148,N_505,N_176);
or U1149 (N_1149,N_216,N_589);
and U1150 (N_1150,N_578,N_465);
and U1151 (N_1151,N_395,N_16);
nand U1152 (N_1152,N_200,N_53);
nand U1153 (N_1153,N_45,N_348);
and U1154 (N_1154,N_179,N_591);
or U1155 (N_1155,N_1,N_555);
or U1156 (N_1156,N_301,N_230);
or U1157 (N_1157,N_328,N_69);
xnor U1158 (N_1158,N_351,N_564);
xor U1159 (N_1159,N_229,N_256);
nand U1160 (N_1160,N_352,N_119);
xor U1161 (N_1161,N_20,N_230);
xnor U1162 (N_1162,N_10,N_438);
nor U1163 (N_1163,N_428,N_78);
nor U1164 (N_1164,N_56,N_466);
xnor U1165 (N_1165,N_308,N_337);
or U1166 (N_1166,N_259,N_65);
xor U1167 (N_1167,N_434,N_414);
xnor U1168 (N_1168,N_528,N_479);
or U1169 (N_1169,N_550,N_206);
xnor U1170 (N_1170,N_582,N_451);
nand U1171 (N_1171,N_96,N_454);
or U1172 (N_1172,N_562,N_504);
nand U1173 (N_1173,N_422,N_567);
and U1174 (N_1174,N_358,N_73);
or U1175 (N_1175,N_472,N_284);
xnor U1176 (N_1176,N_571,N_67);
xor U1177 (N_1177,N_514,N_369);
or U1178 (N_1178,N_432,N_435);
xnor U1179 (N_1179,N_545,N_468);
nor U1180 (N_1180,N_117,N_222);
nand U1181 (N_1181,N_143,N_286);
nand U1182 (N_1182,N_347,N_412);
or U1183 (N_1183,N_397,N_484);
nand U1184 (N_1184,N_329,N_598);
and U1185 (N_1185,N_494,N_108);
nor U1186 (N_1186,N_433,N_223);
and U1187 (N_1187,N_273,N_261);
and U1188 (N_1188,N_187,N_114);
and U1189 (N_1189,N_50,N_413);
nor U1190 (N_1190,N_452,N_64);
or U1191 (N_1191,N_342,N_122);
nand U1192 (N_1192,N_173,N_240);
and U1193 (N_1193,N_554,N_338);
xor U1194 (N_1194,N_301,N_65);
or U1195 (N_1195,N_277,N_250);
nand U1196 (N_1196,N_40,N_422);
or U1197 (N_1197,N_292,N_148);
and U1198 (N_1198,N_369,N_444);
nand U1199 (N_1199,N_20,N_386);
and U1200 (N_1200,N_680,N_684);
and U1201 (N_1201,N_886,N_999);
nand U1202 (N_1202,N_1122,N_1039);
nand U1203 (N_1203,N_957,N_965);
or U1204 (N_1204,N_1141,N_784);
xnor U1205 (N_1205,N_880,N_1045);
nor U1206 (N_1206,N_1005,N_1065);
nand U1207 (N_1207,N_725,N_668);
nor U1208 (N_1208,N_788,N_777);
and U1209 (N_1209,N_620,N_612);
nand U1210 (N_1210,N_915,N_653);
nor U1211 (N_1211,N_933,N_702);
nor U1212 (N_1212,N_1073,N_1074);
xor U1213 (N_1213,N_786,N_610);
nand U1214 (N_1214,N_1159,N_736);
nor U1215 (N_1215,N_940,N_616);
and U1216 (N_1216,N_1067,N_969);
and U1217 (N_1217,N_604,N_1058);
or U1218 (N_1218,N_663,N_879);
and U1219 (N_1219,N_1018,N_1127);
xor U1220 (N_1220,N_895,N_1196);
nor U1221 (N_1221,N_1164,N_1042);
nor U1222 (N_1222,N_693,N_919);
and U1223 (N_1223,N_623,N_1170);
or U1224 (N_1224,N_681,N_1143);
xor U1225 (N_1225,N_722,N_639);
nand U1226 (N_1226,N_821,N_1036);
or U1227 (N_1227,N_1043,N_1081);
and U1228 (N_1228,N_660,N_1025);
xor U1229 (N_1229,N_1140,N_1101);
xor U1230 (N_1230,N_982,N_968);
or U1231 (N_1231,N_923,N_988);
or U1232 (N_1232,N_689,N_629);
xnor U1233 (N_1233,N_905,N_666);
nand U1234 (N_1234,N_892,N_954);
xnor U1235 (N_1235,N_1031,N_749);
or U1236 (N_1236,N_914,N_832);
xor U1237 (N_1237,N_964,N_1047);
and U1238 (N_1238,N_995,N_1168);
and U1239 (N_1239,N_1151,N_1169);
xor U1240 (N_1240,N_730,N_1097);
xor U1241 (N_1241,N_643,N_1082);
nor U1242 (N_1242,N_978,N_973);
or U1243 (N_1243,N_753,N_633);
nand U1244 (N_1244,N_641,N_1048);
and U1245 (N_1245,N_761,N_1112);
and U1246 (N_1246,N_671,N_697);
or U1247 (N_1247,N_764,N_1075);
or U1248 (N_1248,N_757,N_867);
nand U1249 (N_1249,N_1123,N_841);
nand U1250 (N_1250,N_1152,N_854);
nor U1251 (N_1251,N_1035,N_834);
xor U1252 (N_1252,N_876,N_719);
xnor U1253 (N_1253,N_951,N_600);
nor U1254 (N_1254,N_1120,N_714);
nor U1255 (N_1255,N_760,N_618);
nand U1256 (N_1256,N_1165,N_1109);
or U1257 (N_1257,N_1024,N_744);
and U1258 (N_1258,N_601,N_648);
and U1259 (N_1259,N_898,N_657);
nor U1260 (N_1260,N_903,N_930);
xnor U1261 (N_1261,N_955,N_1193);
and U1262 (N_1262,N_864,N_1192);
nor U1263 (N_1263,N_750,N_1153);
nand U1264 (N_1264,N_1029,N_613);
and U1265 (N_1265,N_1080,N_781);
nand U1266 (N_1266,N_1040,N_806);
and U1267 (N_1267,N_796,N_920);
or U1268 (N_1268,N_927,N_826);
nand U1269 (N_1269,N_908,N_807);
xor U1270 (N_1270,N_603,N_1055);
nor U1271 (N_1271,N_1066,N_887);
xor U1272 (N_1272,N_823,N_634);
and U1273 (N_1273,N_789,N_1077);
or U1274 (N_1274,N_1136,N_651);
or U1275 (N_1275,N_983,N_907);
or U1276 (N_1276,N_1102,N_1034);
nand U1277 (N_1277,N_607,N_893);
xnor U1278 (N_1278,N_659,N_683);
or U1279 (N_1279,N_1117,N_961);
nand U1280 (N_1280,N_669,N_738);
or U1281 (N_1281,N_809,N_1100);
nand U1282 (N_1282,N_705,N_677);
xnor U1283 (N_1283,N_992,N_1172);
xnor U1284 (N_1284,N_791,N_1147);
xnor U1285 (N_1285,N_1161,N_828);
nor U1286 (N_1286,N_850,N_1114);
or U1287 (N_1287,N_863,N_1162);
nand U1288 (N_1288,N_870,N_743);
or U1289 (N_1289,N_942,N_1020);
nor U1290 (N_1290,N_696,N_793);
nor U1291 (N_1291,N_716,N_859);
or U1292 (N_1292,N_820,N_773);
or U1293 (N_1293,N_765,N_759);
xnor U1294 (N_1294,N_993,N_990);
nor U1295 (N_1295,N_687,N_1017);
and U1296 (N_1296,N_1022,N_852);
or U1297 (N_1297,N_718,N_1190);
xor U1298 (N_1298,N_1076,N_1186);
and U1299 (N_1299,N_658,N_924);
nand U1300 (N_1300,N_721,N_937);
nor U1301 (N_1301,N_1188,N_906);
and U1302 (N_1302,N_873,N_966);
nor U1303 (N_1303,N_1057,N_1146);
nand U1304 (N_1304,N_824,N_679);
nor U1305 (N_1305,N_934,N_799);
nand U1306 (N_1306,N_742,N_912);
nor U1307 (N_1307,N_960,N_1134);
nand U1308 (N_1308,N_900,N_896);
xnor U1309 (N_1309,N_814,N_1090);
nor U1310 (N_1310,N_1012,N_655);
nor U1311 (N_1311,N_808,N_1118);
nand U1312 (N_1312,N_1108,N_1062);
and U1313 (N_1313,N_1079,N_916);
xor U1314 (N_1314,N_813,N_747);
or U1315 (N_1315,N_728,N_953);
and U1316 (N_1316,N_1160,N_812);
or U1317 (N_1317,N_1156,N_897);
nand U1318 (N_1318,N_994,N_614);
xor U1319 (N_1319,N_1011,N_1054);
xor U1320 (N_1320,N_845,N_611);
and U1321 (N_1321,N_1182,N_706);
or U1322 (N_1322,N_1126,N_1111);
nor U1323 (N_1323,N_1183,N_805);
xnor U1324 (N_1324,N_678,N_856);
xnor U1325 (N_1325,N_1178,N_727);
nor U1326 (N_1326,N_810,N_1091);
nand U1327 (N_1327,N_1105,N_630);
or U1328 (N_1328,N_1032,N_710);
and U1329 (N_1329,N_875,N_1095);
and U1330 (N_1330,N_1119,N_804);
nand U1331 (N_1331,N_976,N_979);
and U1332 (N_1332,N_956,N_825);
xor U1333 (N_1333,N_617,N_1155);
or U1334 (N_1334,N_1157,N_1015);
nand U1335 (N_1335,N_688,N_936);
xor U1336 (N_1336,N_1129,N_817);
or U1337 (N_1337,N_741,N_962);
nor U1338 (N_1338,N_762,N_1027);
xor U1339 (N_1339,N_866,N_846);
nor U1340 (N_1340,N_944,N_1049);
xor U1341 (N_1341,N_709,N_1007);
and U1342 (N_1342,N_798,N_874);
nand U1343 (N_1343,N_700,N_1026);
and U1344 (N_1344,N_783,N_989);
nand U1345 (N_1345,N_1063,N_949);
or U1346 (N_1346,N_1071,N_682);
and U1347 (N_1347,N_608,N_885);
and U1348 (N_1348,N_827,N_918);
xor U1349 (N_1349,N_1056,N_667);
and U1350 (N_1350,N_1130,N_1115);
nand U1351 (N_1351,N_977,N_1059);
and U1352 (N_1352,N_890,N_844);
nand U1353 (N_1353,N_769,N_1093);
nand U1354 (N_1354,N_981,N_627);
and U1355 (N_1355,N_837,N_819);
or U1356 (N_1356,N_899,N_642);
and U1357 (N_1357,N_654,N_763);
nor U1358 (N_1358,N_686,N_779);
and U1359 (N_1359,N_1008,N_1016);
or U1360 (N_1360,N_996,N_662);
xor U1361 (N_1361,N_647,N_665);
or U1362 (N_1362,N_921,N_1124);
and U1363 (N_1363,N_800,N_1089);
and U1364 (N_1364,N_1087,N_902);
xnor U1365 (N_1365,N_815,N_843);
nand U1366 (N_1366,N_913,N_928);
nand U1367 (N_1367,N_1158,N_871);
xor U1368 (N_1368,N_755,N_778);
xor U1369 (N_1369,N_1006,N_615);
or U1370 (N_1370,N_987,N_1171);
and U1371 (N_1371,N_1173,N_782);
xnor U1372 (N_1372,N_605,N_652);
xor U1373 (N_1373,N_676,N_766);
or U1374 (N_1374,N_858,N_790);
and U1375 (N_1375,N_768,N_882);
nor U1376 (N_1376,N_947,N_1154);
or U1377 (N_1377,N_1070,N_860);
nor U1378 (N_1378,N_664,N_831);
xnor U1379 (N_1379,N_963,N_708);
nand U1380 (N_1380,N_904,N_1191);
nor U1381 (N_1381,N_938,N_1103);
and U1382 (N_1382,N_646,N_1104);
nor U1383 (N_1383,N_967,N_816);
and U1384 (N_1384,N_707,N_1085);
nand U1385 (N_1385,N_948,N_717);
or U1386 (N_1386,N_1096,N_830);
nand U1387 (N_1387,N_1002,N_980);
nand U1388 (N_1388,N_1083,N_1060);
nand U1389 (N_1389,N_929,N_649);
nor U1390 (N_1390,N_1133,N_839);
or U1391 (N_1391,N_1116,N_1013);
or U1392 (N_1392,N_1189,N_853);
nand U1393 (N_1393,N_704,N_1144);
xnor U1394 (N_1394,N_1199,N_703);
xnor U1395 (N_1395,N_1181,N_661);
and U1396 (N_1396,N_1064,N_803);
nor U1397 (N_1397,N_884,N_1028);
and U1398 (N_1398,N_1180,N_971);
nand U1399 (N_1399,N_1044,N_972);
or U1400 (N_1400,N_986,N_1110);
and U1401 (N_1401,N_731,N_776);
nand U1402 (N_1402,N_1125,N_1021);
nor U1403 (N_1403,N_970,N_732);
nand U1404 (N_1404,N_619,N_720);
and U1405 (N_1405,N_606,N_1038);
or U1406 (N_1406,N_801,N_640);
nor U1407 (N_1407,N_1037,N_984);
and U1408 (N_1408,N_701,N_881);
and U1409 (N_1409,N_950,N_1184);
nand U1410 (N_1410,N_739,N_877);
xnor U1411 (N_1411,N_1174,N_670);
and U1412 (N_1412,N_746,N_822);
xnor U1413 (N_1413,N_1092,N_811);
and U1414 (N_1414,N_626,N_998);
nor U1415 (N_1415,N_855,N_997);
and U1416 (N_1416,N_775,N_770);
nor U1417 (N_1417,N_1142,N_723);
nor U1418 (N_1418,N_637,N_1072);
nor U1419 (N_1419,N_932,N_935);
nor U1420 (N_1420,N_835,N_926);
or U1421 (N_1421,N_985,N_868);
nand U1422 (N_1422,N_780,N_840);
xnor U1423 (N_1423,N_851,N_1084);
nand U1424 (N_1424,N_712,N_636);
nand U1425 (N_1425,N_645,N_925);
nor U1426 (N_1426,N_748,N_958);
nor U1427 (N_1427,N_901,N_1001);
nor U1428 (N_1428,N_733,N_838);
nor U1429 (N_1429,N_1010,N_847);
nor U1430 (N_1430,N_959,N_889);
and U1431 (N_1431,N_910,N_865);
or U1432 (N_1432,N_1198,N_772);
nand U1433 (N_1433,N_656,N_735);
nor U1434 (N_1434,N_1138,N_1053);
and U1435 (N_1435,N_609,N_695);
nand U1436 (N_1436,N_1150,N_861);
nand U1437 (N_1437,N_690,N_692);
or U1438 (N_1438,N_1061,N_1113);
and U1439 (N_1439,N_767,N_726);
and U1440 (N_1440,N_891,N_917);
and U1441 (N_1441,N_795,N_740);
nand U1442 (N_1442,N_931,N_1023);
xnor U1443 (N_1443,N_1088,N_1166);
nor U1444 (N_1444,N_1078,N_751);
xnor U1445 (N_1445,N_1187,N_1009);
nand U1446 (N_1446,N_713,N_1195);
nor U1447 (N_1447,N_1137,N_797);
nand U1448 (N_1448,N_715,N_632);
xnor U1449 (N_1449,N_1149,N_602);
or U1450 (N_1450,N_1177,N_974);
and U1451 (N_1451,N_1176,N_675);
nor U1452 (N_1452,N_754,N_939);
nor U1453 (N_1453,N_758,N_1197);
nor U1454 (N_1454,N_1106,N_941);
xnor U1455 (N_1455,N_638,N_699);
or U1456 (N_1456,N_1019,N_1046);
nor U1457 (N_1457,N_1014,N_1163);
nand U1458 (N_1458,N_878,N_894);
and U1459 (N_1459,N_1132,N_787);
and U1460 (N_1460,N_631,N_1068);
xnor U1461 (N_1461,N_922,N_737);
and U1462 (N_1462,N_1069,N_622);
or U1463 (N_1463,N_673,N_624);
nand U1464 (N_1464,N_946,N_991);
and U1465 (N_1465,N_1131,N_945);
nor U1466 (N_1466,N_952,N_883);
and U1467 (N_1467,N_729,N_818);
nand U1468 (N_1468,N_848,N_1175);
or U1469 (N_1469,N_1128,N_711);
nand U1470 (N_1470,N_857,N_911);
nand U1471 (N_1471,N_694,N_650);
nand U1472 (N_1472,N_1145,N_1139);
nor U1473 (N_1473,N_836,N_685);
nor U1474 (N_1474,N_909,N_1033);
and U1475 (N_1475,N_745,N_829);
nor U1476 (N_1476,N_625,N_1094);
or U1477 (N_1477,N_1107,N_635);
nand U1478 (N_1478,N_792,N_1041);
or U1479 (N_1479,N_621,N_842);
and U1480 (N_1480,N_888,N_774);
nand U1481 (N_1481,N_833,N_1003);
xor U1482 (N_1482,N_1000,N_1099);
and U1483 (N_1483,N_1050,N_1004);
and U1484 (N_1484,N_1098,N_794);
nor U1485 (N_1485,N_1135,N_1167);
nor U1486 (N_1486,N_975,N_1086);
nand U1487 (N_1487,N_1185,N_752);
and U1488 (N_1488,N_869,N_862);
xor U1489 (N_1489,N_1051,N_771);
and U1490 (N_1490,N_1194,N_644);
nor U1491 (N_1491,N_1121,N_672);
and U1492 (N_1492,N_802,N_1052);
xor U1493 (N_1493,N_674,N_785);
and U1494 (N_1494,N_628,N_734);
nand U1495 (N_1495,N_872,N_1179);
xor U1496 (N_1496,N_691,N_943);
nor U1497 (N_1497,N_698,N_1030);
nand U1498 (N_1498,N_724,N_756);
and U1499 (N_1499,N_1148,N_849);
or U1500 (N_1500,N_1076,N_1185);
nor U1501 (N_1501,N_1063,N_652);
nor U1502 (N_1502,N_838,N_1023);
nand U1503 (N_1503,N_615,N_1011);
xor U1504 (N_1504,N_723,N_887);
xnor U1505 (N_1505,N_799,N_824);
nand U1506 (N_1506,N_1146,N_668);
xnor U1507 (N_1507,N_956,N_697);
xor U1508 (N_1508,N_957,N_900);
or U1509 (N_1509,N_711,N_830);
xnor U1510 (N_1510,N_725,N_944);
nand U1511 (N_1511,N_1144,N_728);
nor U1512 (N_1512,N_787,N_898);
nor U1513 (N_1513,N_1141,N_1126);
nor U1514 (N_1514,N_891,N_973);
nor U1515 (N_1515,N_1126,N_1001);
nor U1516 (N_1516,N_864,N_649);
xor U1517 (N_1517,N_912,N_922);
nand U1518 (N_1518,N_1043,N_722);
and U1519 (N_1519,N_753,N_1140);
and U1520 (N_1520,N_1172,N_738);
xor U1521 (N_1521,N_935,N_1018);
nand U1522 (N_1522,N_1164,N_1098);
and U1523 (N_1523,N_658,N_739);
or U1524 (N_1524,N_623,N_1115);
nand U1525 (N_1525,N_1183,N_820);
xnor U1526 (N_1526,N_1138,N_1042);
nor U1527 (N_1527,N_738,N_1134);
or U1528 (N_1528,N_658,N_857);
or U1529 (N_1529,N_988,N_925);
nand U1530 (N_1530,N_1159,N_658);
nor U1531 (N_1531,N_1096,N_721);
nor U1532 (N_1532,N_610,N_811);
nor U1533 (N_1533,N_937,N_1101);
and U1534 (N_1534,N_798,N_1014);
nor U1535 (N_1535,N_633,N_1098);
nand U1536 (N_1536,N_707,N_961);
nand U1537 (N_1537,N_1172,N_1167);
nand U1538 (N_1538,N_1180,N_999);
nand U1539 (N_1539,N_1139,N_675);
nand U1540 (N_1540,N_1176,N_1088);
or U1541 (N_1541,N_1042,N_1126);
or U1542 (N_1542,N_903,N_999);
xnor U1543 (N_1543,N_730,N_639);
nor U1544 (N_1544,N_998,N_949);
or U1545 (N_1545,N_771,N_754);
xnor U1546 (N_1546,N_740,N_703);
nor U1547 (N_1547,N_671,N_970);
xor U1548 (N_1548,N_870,N_893);
nor U1549 (N_1549,N_963,N_1115);
xnor U1550 (N_1550,N_628,N_774);
nor U1551 (N_1551,N_719,N_958);
nand U1552 (N_1552,N_799,N_919);
xor U1553 (N_1553,N_821,N_858);
xnor U1554 (N_1554,N_887,N_655);
nor U1555 (N_1555,N_707,N_948);
or U1556 (N_1556,N_1098,N_652);
xnor U1557 (N_1557,N_1156,N_975);
xnor U1558 (N_1558,N_776,N_913);
or U1559 (N_1559,N_657,N_930);
xor U1560 (N_1560,N_819,N_620);
xnor U1561 (N_1561,N_639,N_1199);
nor U1562 (N_1562,N_611,N_1038);
and U1563 (N_1563,N_709,N_1189);
xnor U1564 (N_1564,N_991,N_1050);
or U1565 (N_1565,N_848,N_855);
or U1566 (N_1566,N_1040,N_953);
xor U1567 (N_1567,N_1043,N_713);
and U1568 (N_1568,N_1115,N_916);
and U1569 (N_1569,N_988,N_1167);
xnor U1570 (N_1570,N_852,N_779);
or U1571 (N_1571,N_644,N_1029);
or U1572 (N_1572,N_852,N_863);
xor U1573 (N_1573,N_1073,N_1091);
and U1574 (N_1574,N_1119,N_895);
or U1575 (N_1575,N_1057,N_1052);
nand U1576 (N_1576,N_960,N_993);
nor U1577 (N_1577,N_634,N_1138);
or U1578 (N_1578,N_681,N_1122);
nand U1579 (N_1579,N_948,N_669);
nand U1580 (N_1580,N_749,N_830);
xor U1581 (N_1581,N_1094,N_878);
xnor U1582 (N_1582,N_1195,N_753);
xnor U1583 (N_1583,N_1148,N_1146);
nor U1584 (N_1584,N_952,N_1083);
and U1585 (N_1585,N_1042,N_702);
xnor U1586 (N_1586,N_746,N_756);
nand U1587 (N_1587,N_830,N_807);
xor U1588 (N_1588,N_770,N_1132);
or U1589 (N_1589,N_692,N_802);
xor U1590 (N_1590,N_979,N_988);
xor U1591 (N_1591,N_646,N_816);
nand U1592 (N_1592,N_883,N_735);
and U1593 (N_1593,N_842,N_608);
or U1594 (N_1594,N_949,N_1113);
nand U1595 (N_1595,N_915,N_1100);
xnor U1596 (N_1596,N_795,N_904);
or U1597 (N_1597,N_833,N_1176);
or U1598 (N_1598,N_772,N_792);
nor U1599 (N_1599,N_1037,N_1069);
or U1600 (N_1600,N_633,N_788);
xor U1601 (N_1601,N_859,N_1107);
nand U1602 (N_1602,N_1168,N_839);
and U1603 (N_1603,N_1039,N_1045);
and U1604 (N_1604,N_668,N_682);
nor U1605 (N_1605,N_784,N_670);
nand U1606 (N_1606,N_802,N_634);
nand U1607 (N_1607,N_1113,N_765);
and U1608 (N_1608,N_845,N_1032);
and U1609 (N_1609,N_1039,N_772);
xnor U1610 (N_1610,N_1077,N_1005);
xor U1611 (N_1611,N_1165,N_1153);
nand U1612 (N_1612,N_880,N_1163);
xor U1613 (N_1613,N_1133,N_780);
or U1614 (N_1614,N_794,N_675);
and U1615 (N_1615,N_1059,N_939);
or U1616 (N_1616,N_764,N_1015);
and U1617 (N_1617,N_860,N_698);
nor U1618 (N_1618,N_787,N_1010);
nand U1619 (N_1619,N_1172,N_1044);
nand U1620 (N_1620,N_1145,N_1179);
or U1621 (N_1621,N_680,N_715);
or U1622 (N_1622,N_863,N_817);
nand U1623 (N_1623,N_1114,N_667);
nor U1624 (N_1624,N_839,N_781);
and U1625 (N_1625,N_1176,N_709);
nand U1626 (N_1626,N_617,N_1010);
xnor U1627 (N_1627,N_982,N_779);
nor U1628 (N_1628,N_861,N_898);
or U1629 (N_1629,N_811,N_700);
nand U1630 (N_1630,N_794,N_1097);
or U1631 (N_1631,N_943,N_647);
nand U1632 (N_1632,N_704,N_987);
or U1633 (N_1633,N_611,N_1042);
nor U1634 (N_1634,N_809,N_1118);
xor U1635 (N_1635,N_857,N_628);
nand U1636 (N_1636,N_765,N_1119);
or U1637 (N_1637,N_784,N_1116);
and U1638 (N_1638,N_971,N_669);
nand U1639 (N_1639,N_703,N_1088);
nor U1640 (N_1640,N_650,N_1158);
nand U1641 (N_1641,N_1081,N_775);
nor U1642 (N_1642,N_776,N_948);
nor U1643 (N_1643,N_736,N_1199);
nor U1644 (N_1644,N_1198,N_946);
or U1645 (N_1645,N_693,N_1179);
xor U1646 (N_1646,N_694,N_1138);
nand U1647 (N_1647,N_819,N_671);
and U1648 (N_1648,N_1194,N_914);
nor U1649 (N_1649,N_1043,N_810);
and U1650 (N_1650,N_1016,N_716);
nor U1651 (N_1651,N_828,N_1140);
xnor U1652 (N_1652,N_1064,N_671);
or U1653 (N_1653,N_750,N_982);
or U1654 (N_1654,N_955,N_917);
xor U1655 (N_1655,N_1080,N_676);
or U1656 (N_1656,N_602,N_808);
or U1657 (N_1657,N_720,N_925);
and U1658 (N_1658,N_1124,N_816);
and U1659 (N_1659,N_1104,N_783);
or U1660 (N_1660,N_721,N_1164);
and U1661 (N_1661,N_979,N_1179);
nor U1662 (N_1662,N_678,N_607);
xor U1663 (N_1663,N_1024,N_814);
xnor U1664 (N_1664,N_1075,N_748);
and U1665 (N_1665,N_1103,N_1109);
and U1666 (N_1666,N_1107,N_840);
nand U1667 (N_1667,N_850,N_841);
or U1668 (N_1668,N_1173,N_945);
xor U1669 (N_1669,N_1142,N_756);
and U1670 (N_1670,N_855,N_725);
nand U1671 (N_1671,N_896,N_1085);
nor U1672 (N_1672,N_877,N_737);
xor U1673 (N_1673,N_718,N_872);
or U1674 (N_1674,N_812,N_938);
nand U1675 (N_1675,N_1127,N_699);
and U1676 (N_1676,N_1161,N_902);
xor U1677 (N_1677,N_765,N_737);
and U1678 (N_1678,N_1180,N_908);
nand U1679 (N_1679,N_962,N_802);
or U1680 (N_1680,N_768,N_1012);
or U1681 (N_1681,N_883,N_1166);
or U1682 (N_1682,N_722,N_1033);
xnor U1683 (N_1683,N_667,N_913);
nand U1684 (N_1684,N_1178,N_660);
nor U1685 (N_1685,N_926,N_1020);
xor U1686 (N_1686,N_754,N_1173);
nor U1687 (N_1687,N_699,N_1117);
and U1688 (N_1688,N_669,N_993);
nor U1689 (N_1689,N_994,N_800);
nand U1690 (N_1690,N_792,N_1106);
or U1691 (N_1691,N_778,N_1159);
xor U1692 (N_1692,N_644,N_1080);
and U1693 (N_1693,N_787,N_781);
or U1694 (N_1694,N_1140,N_966);
xnor U1695 (N_1695,N_760,N_816);
or U1696 (N_1696,N_992,N_640);
or U1697 (N_1697,N_937,N_1014);
nor U1698 (N_1698,N_1080,N_855);
nor U1699 (N_1699,N_920,N_1011);
nand U1700 (N_1700,N_844,N_911);
xor U1701 (N_1701,N_1060,N_771);
xor U1702 (N_1702,N_1101,N_1159);
nand U1703 (N_1703,N_967,N_1002);
nor U1704 (N_1704,N_981,N_691);
xor U1705 (N_1705,N_1157,N_904);
nand U1706 (N_1706,N_1009,N_903);
nor U1707 (N_1707,N_1044,N_887);
nand U1708 (N_1708,N_629,N_832);
nor U1709 (N_1709,N_672,N_643);
nand U1710 (N_1710,N_912,N_1033);
nor U1711 (N_1711,N_691,N_900);
and U1712 (N_1712,N_634,N_749);
nand U1713 (N_1713,N_683,N_901);
nand U1714 (N_1714,N_643,N_967);
or U1715 (N_1715,N_1011,N_737);
nor U1716 (N_1716,N_984,N_766);
nor U1717 (N_1717,N_883,N_1022);
nand U1718 (N_1718,N_837,N_675);
nand U1719 (N_1719,N_901,N_1147);
xor U1720 (N_1720,N_1126,N_783);
and U1721 (N_1721,N_679,N_956);
or U1722 (N_1722,N_1082,N_1036);
and U1723 (N_1723,N_890,N_984);
and U1724 (N_1724,N_1100,N_1091);
or U1725 (N_1725,N_1038,N_914);
nand U1726 (N_1726,N_1170,N_793);
and U1727 (N_1727,N_1081,N_998);
nor U1728 (N_1728,N_649,N_918);
nor U1729 (N_1729,N_1066,N_1048);
or U1730 (N_1730,N_705,N_980);
xnor U1731 (N_1731,N_821,N_1135);
and U1732 (N_1732,N_650,N_958);
or U1733 (N_1733,N_855,N_1165);
nor U1734 (N_1734,N_1038,N_781);
and U1735 (N_1735,N_1047,N_1057);
nor U1736 (N_1736,N_931,N_789);
or U1737 (N_1737,N_698,N_1146);
xnor U1738 (N_1738,N_665,N_1085);
xnor U1739 (N_1739,N_634,N_1042);
xnor U1740 (N_1740,N_1070,N_842);
and U1741 (N_1741,N_1039,N_908);
nand U1742 (N_1742,N_876,N_1113);
and U1743 (N_1743,N_1062,N_824);
or U1744 (N_1744,N_719,N_986);
and U1745 (N_1745,N_1146,N_1082);
xor U1746 (N_1746,N_629,N_942);
nand U1747 (N_1747,N_916,N_851);
nand U1748 (N_1748,N_1118,N_814);
and U1749 (N_1749,N_927,N_880);
nand U1750 (N_1750,N_614,N_1014);
xnor U1751 (N_1751,N_1031,N_1117);
or U1752 (N_1752,N_1180,N_989);
or U1753 (N_1753,N_1171,N_670);
or U1754 (N_1754,N_1066,N_1018);
nor U1755 (N_1755,N_849,N_717);
and U1756 (N_1756,N_1178,N_724);
or U1757 (N_1757,N_962,N_914);
nand U1758 (N_1758,N_1002,N_946);
nand U1759 (N_1759,N_1112,N_842);
xnor U1760 (N_1760,N_779,N_1181);
xnor U1761 (N_1761,N_670,N_1018);
and U1762 (N_1762,N_910,N_1109);
and U1763 (N_1763,N_938,N_774);
and U1764 (N_1764,N_763,N_693);
nor U1765 (N_1765,N_1133,N_825);
and U1766 (N_1766,N_920,N_720);
or U1767 (N_1767,N_956,N_817);
nor U1768 (N_1768,N_621,N_672);
nor U1769 (N_1769,N_609,N_725);
nor U1770 (N_1770,N_1107,N_650);
nand U1771 (N_1771,N_975,N_1190);
and U1772 (N_1772,N_1143,N_732);
nor U1773 (N_1773,N_630,N_1182);
and U1774 (N_1774,N_1134,N_703);
and U1775 (N_1775,N_627,N_966);
nor U1776 (N_1776,N_767,N_700);
or U1777 (N_1777,N_1134,N_1070);
nor U1778 (N_1778,N_729,N_1122);
or U1779 (N_1779,N_1078,N_1134);
nor U1780 (N_1780,N_815,N_878);
nand U1781 (N_1781,N_837,N_934);
xnor U1782 (N_1782,N_819,N_829);
and U1783 (N_1783,N_798,N_1145);
nor U1784 (N_1784,N_626,N_940);
xnor U1785 (N_1785,N_1030,N_877);
nand U1786 (N_1786,N_845,N_669);
nand U1787 (N_1787,N_686,N_1117);
nor U1788 (N_1788,N_932,N_766);
xnor U1789 (N_1789,N_865,N_723);
nand U1790 (N_1790,N_641,N_710);
or U1791 (N_1791,N_603,N_630);
and U1792 (N_1792,N_811,N_999);
xnor U1793 (N_1793,N_1109,N_666);
nor U1794 (N_1794,N_629,N_665);
xnor U1795 (N_1795,N_864,N_675);
xnor U1796 (N_1796,N_1056,N_883);
xor U1797 (N_1797,N_1070,N_939);
or U1798 (N_1798,N_916,N_782);
or U1799 (N_1799,N_923,N_835);
xnor U1800 (N_1800,N_1649,N_1203);
nor U1801 (N_1801,N_1664,N_1469);
nor U1802 (N_1802,N_1316,N_1650);
or U1803 (N_1803,N_1769,N_1459);
xnor U1804 (N_1804,N_1416,N_1578);
and U1805 (N_1805,N_1538,N_1251);
and U1806 (N_1806,N_1645,N_1663);
or U1807 (N_1807,N_1750,N_1308);
xor U1808 (N_1808,N_1736,N_1660);
xor U1809 (N_1809,N_1684,N_1255);
xor U1810 (N_1810,N_1572,N_1345);
nand U1811 (N_1811,N_1247,N_1629);
and U1812 (N_1812,N_1365,N_1404);
xor U1813 (N_1813,N_1363,N_1519);
and U1814 (N_1814,N_1794,N_1682);
nand U1815 (N_1815,N_1557,N_1334);
xor U1816 (N_1816,N_1237,N_1597);
nand U1817 (N_1817,N_1554,N_1398);
and U1818 (N_1818,N_1479,N_1333);
and U1819 (N_1819,N_1386,N_1689);
or U1820 (N_1820,N_1435,N_1327);
nand U1821 (N_1821,N_1499,N_1558);
or U1822 (N_1822,N_1394,N_1244);
nor U1823 (N_1823,N_1235,N_1708);
nand U1824 (N_1824,N_1477,N_1523);
xor U1825 (N_1825,N_1662,N_1419);
or U1826 (N_1826,N_1376,N_1261);
or U1827 (N_1827,N_1711,N_1298);
xnor U1828 (N_1828,N_1757,N_1322);
nand U1829 (N_1829,N_1588,N_1290);
and U1830 (N_1830,N_1269,N_1521);
xor U1831 (N_1831,N_1569,N_1200);
and U1832 (N_1832,N_1699,N_1703);
nor U1833 (N_1833,N_1691,N_1604);
nor U1834 (N_1834,N_1696,N_1370);
xor U1835 (N_1835,N_1674,N_1591);
and U1836 (N_1836,N_1665,N_1391);
nand U1837 (N_1837,N_1389,N_1765);
or U1838 (N_1838,N_1671,N_1344);
and U1839 (N_1839,N_1752,N_1722);
or U1840 (N_1840,N_1229,N_1314);
nor U1841 (N_1841,N_1202,N_1762);
xnor U1842 (N_1842,N_1677,N_1718);
xnor U1843 (N_1843,N_1568,N_1458);
nor U1844 (N_1844,N_1421,N_1425);
nor U1845 (N_1845,N_1481,N_1328);
nor U1846 (N_1846,N_1501,N_1434);
xnor U1847 (N_1847,N_1346,N_1270);
nand U1848 (N_1848,N_1271,N_1473);
nand U1849 (N_1849,N_1624,N_1442);
or U1850 (N_1850,N_1617,N_1369);
or U1851 (N_1851,N_1413,N_1599);
and U1852 (N_1852,N_1697,N_1304);
nor U1853 (N_1853,N_1594,N_1383);
nor U1854 (N_1854,N_1508,N_1709);
and U1855 (N_1855,N_1209,N_1638);
or U1856 (N_1856,N_1563,N_1751);
nor U1857 (N_1857,N_1758,N_1549);
nand U1858 (N_1858,N_1786,N_1770);
nand U1859 (N_1859,N_1492,N_1301);
and U1860 (N_1860,N_1385,N_1755);
and U1861 (N_1861,N_1518,N_1546);
xor U1862 (N_1862,N_1215,N_1742);
or U1863 (N_1863,N_1252,N_1222);
nand U1864 (N_1864,N_1302,N_1631);
or U1865 (N_1865,N_1616,N_1228);
nor U1866 (N_1866,N_1676,N_1651);
and U1867 (N_1867,N_1330,N_1586);
nor U1868 (N_1868,N_1720,N_1497);
or U1869 (N_1869,N_1642,N_1507);
nand U1870 (N_1870,N_1207,N_1342);
nand U1871 (N_1871,N_1289,N_1489);
and U1872 (N_1872,N_1254,N_1509);
nand U1873 (N_1873,N_1547,N_1279);
or U1874 (N_1874,N_1657,N_1653);
and U1875 (N_1875,N_1749,N_1500);
and U1876 (N_1876,N_1233,N_1799);
xnor U1877 (N_1877,N_1582,N_1743);
nand U1878 (N_1878,N_1777,N_1730);
nor U1879 (N_1879,N_1789,N_1715);
or U1880 (N_1880,N_1319,N_1357);
nor U1881 (N_1881,N_1323,N_1293);
nand U1882 (N_1882,N_1717,N_1451);
and U1883 (N_1883,N_1428,N_1223);
or U1884 (N_1884,N_1351,N_1764);
nor U1885 (N_1885,N_1714,N_1600);
or U1886 (N_1886,N_1362,N_1669);
or U1887 (N_1887,N_1213,N_1384);
nand U1888 (N_1888,N_1338,N_1763);
nor U1889 (N_1889,N_1679,N_1352);
nand U1890 (N_1890,N_1273,N_1598);
nor U1891 (N_1891,N_1639,N_1776);
nand U1892 (N_1892,N_1388,N_1297);
or U1893 (N_1893,N_1392,N_1567);
or U1894 (N_1894,N_1529,N_1545);
nor U1895 (N_1895,N_1414,N_1461);
nor U1896 (N_1896,N_1221,N_1748);
nand U1897 (N_1897,N_1356,N_1692);
nor U1898 (N_1898,N_1517,N_1723);
nand U1899 (N_1899,N_1373,N_1390);
nor U1900 (N_1900,N_1731,N_1410);
nand U1901 (N_1901,N_1292,N_1454);
or U1902 (N_1902,N_1412,N_1219);
nor U1903 (N_1903,N_1277,N_1329);
nand U1904 (N_1904,N_1475,N_1733);
and U1905 (N_1905,N_1424,N_1490);
xor U1906 (N_1906,N_1609,N_1408);
nor U1907 (N_1907,N_1622,N_1710);
or U1908 (N_1908,N_1779,N_1409);
nand U1909 (N_1909,N_1628,N_1283);
and U1910 (N_1910,N_1349,N_1258);
nor U1911 (N_1911,N_1612,N_1713);
nor U1912 (N_1912,N_1212,N_1484);
and U1913 (N_1913,N_1619,N_1401);
or U1914 (N_1914,N_1287,N_1480);
and U1915 (N_1915,N_1584,N_1783);
and U1916 (N_1916,N_1539,N_1487);
or U1917 (N_1917,N_1399,N_1552);
or U1918 (N_1918,N_1672,N_1756);
and U1919 (N_1919,N_1530,N_1433);
xor U1920 (N_1920,N_1732,N_1746);
nor U1921 (N_1921,N_1260,N_1621);
nor U1922 (N_1922,N_1462,N_1526);
xor U1923 (N_1923,N_1635,N_1256);
and U1924 (N_1924,N_1744,N_1214);
nand U1925 (N_1925,N_1627,N_1793);
xnor U1926 (N_1926,N_1513,N_1637);
or U1927 (N_1927,N_1460,N_1647);
xor U1928 (N_1928,N_1358,N_1464);
xnor U1929 (N_1929,N_1375,N_1792);
nand U1930 (N_1930,N_1693,N_1436);
or U1931 (N_1931,N_1550,N_1371);
xnor U1932 (N_1932,N_1551,N_1211);
xor U1933 (N_1933,N_1630,N_1368);
nor U1934 (N_1934,N_1564,N_1361);
nor U1935 (N_1935,N_1537,N_1332);
and U1936 (N_1936,N_1309,N_1378);
and U1937 (N_1937,N_1658,N_1206);
xor U1938 (N_1938,N_1307,N_1680);
xnor U1939 (N_1939,N_1263,N_1575);
nand U1940 (N_1940,N_1686,N_1246);
or U1941 (N_1941,N_1716,N_1753);
nor U1942 (N_1942,N_1522,N_1668);
and U1943 (N_1943,N_1278,N_1589);
and U1944 (N_1944,N_1734,N_1285);
or U1945 (N_1945,N_1326,N_1620);
or U1946 (N_1946,N_1335,N_1601);
and U1947 (N_1947,N_1262,N_1656);
and U1948 (N_1948,N_1667,N_1640);
xor U1949 (N_1949,N_1670,N_1305);
xor U1950 (N_1950,N_1585,N_1313);
nand U1951 (N_1951,N_1700,N_1511);
xnor U1952 (N_1952,N_1347,N_1790);
or U1953 (N_1953,N_1232,N_1341);
and U1954 (N_1954,N_1610,N_1795);
or U1955 (N_1955,N_1320,N_1466);
or U1956 (N_1956,N_1216,N_1259);
or U1957 (N_1957,N_1739,N_1448);
nand U1958 (N_1958,N_1618,N_1415);
or U1959 (N_1959,N_1496,N_1536);
or U1960 (N_1960,N_1471,N_1317);
nand U1961 (N_1961,N_1303,N_1623);
or U1962 (N_1962,N_1245,N_1583);
xor U1963 (N_1963,N_1615,N_1350);
nor U1964 (N_1964,N_1728,N_1535);
xor U1965 (N_1965,N_1774,N_1798);
xor U1966 (N_1966,N_1590,N_1659);
nor U1967 (N_1967,N_1455,N_1236);
nor U1968 (N_1968,N_1655,N_1775);
or U1969 (N_1969,N_1423,N_1275);
and U1970 (N_1970,N_1465,N_1504);
xnor U1971 (N_1971,N_1566,N_1761);
nand U1972 (N_1972,N_1268,N_1544);
nand U1973 (N_1973,N_1422,N_1579);
xnor U1974 (N_1974,N_1791,N_1543);
xnor U1975 (N_1975,N_1485,N_1472);
nand U1976 (N_1976,N_1493,N_1681);
and U1977 (N_1977,N_1272,N_1772);
nor U1978 (N_1978,N_1540,N_1441);
xnor U1979 (N_1979,N_1288,N_1354);
xnor U1980 (N_1980,N_1432,N_1644);
nand U1981 (N_1981,N_1224,N_1311);
or U1982 (N_1982,N_1407,N_1514);
nor U1983 (N_1983,N_1675,N_1754);
or U1984 (N_1984,N_1515,N_1516);
xor U1985 (N_1985,N_1555,N_1463);
nand U1986 (N_1986,N_1225,N_1249);
and U1987 (N_1987,N_1593,N_1318);
xnor U1988 (N_1988,N_1456,N_1737);
xor U1989 (N_1989,N_1698,N_1611);
nand U1990 (N_1990,N_1778,N_1296);
nand U1991 (N_1991,N_1444,N_1524);
and U1992 (N_1992,N_1581,N_1274);
nor U1993 (N_1993,N_1712,N_1607);
or U1994 (N_1994,N_1439,N_1280);
nand U1995 (N_1995,N_1602,N_1577);
nand U1996 (N_1996,N_1661,N_1721);
and U1997 (N_1997,N_1702,N_1380);
and U1998 (N_1998,N_1678,N_1633);
nor U1999 (N_1999,N_1606,N_1706);
nand U2000 (N_2000,N_1427,N_1747);
xnor U2001 (N_2001,N_1695,N_1587);
xnor U2002 (N_2002,N_1553,N_1201);
xor U2003 (N_2003,N_1353,N_1315);
nor U2004 (N_2004,N_1646,N_1542);
xor U2005 (N_2005,N_1701,N_1360);
and U2006 (N_2006,N_1527,N_1241);
nand U2007 (N_2007,N_1411,N_1418);
or U2008 (N_2008,N_1773,N_1438);
and U2009 (N_2009,N_1239,N_1395);
nand U2010 (N_2010,N_1242,N_1210);
nand U2011 (N_2011,N_1760,N_1226);
and U2012 (N_2012,N_1306,N_1687);
and U2013 (N_2013,N_1382,N_1688);
nand U2014 (N_2014,N_1417,N_1406);
nor U2015 (N_2015,N_1768,N_1548);
or U2016 (N_2016,N_1512,N_1488);
nand U2017 (N_2017,N_1781,N_1396);
xor U2018 (N_2018,N_1387,N_1727);
xnor U2019 (N_2019,N_1648,N_1377);
nor U2020 (N_2020,N_1498,N_1788);
nand U2021 (N_2021,N_1367,N_1403);
xnor U2022 (N_2022,N_1420,N_1576);
and U2023 (N_2023,N_1447,N_1603);
or U2024 (N_2024,N_1476,N_1431);
nor U2025 (N_2025,N_1331,N_1295);
and U2026 (N_2026,N_1771,N_1467);
and U2027 (N_2027,N_1528,N_1291);
nor U2028 (N_2028,N_1250,N_1673);
or U2029 (N_2029,N_1457,N_1596);
nor U2030 (N_2030,N_1741,N_1784);
nor U2031 (N_2031,N_1281,N_1220);
or U2032 (N_2032,N_1449,N_1690);
xnor U2033 (N_2033,N_1726,N_1299);
nand U2034 (N_2034,N_1243,N_1453);
nor U2035 (N_2035,N_1379,N_1474);
nor U2036 (N_2036,N_1446,N_1486);
nand U2037 (N_2037,N_1608,N_1312);
or U2038 (N_2038,N_1445,N_1321);
or U2039 (N_2039,N_1257,N_1227);
or U2040 (N_2040,N_1574,N_1300);
or U2041 (N_2041,N_1372,N_1374);
or U2042 (N_2042,N_1533,N_1704);
or U2043 (N_2043,N_1218,N_1759);
and U2044 (N_2044,N_1248,N_1560);
nand U2045 (N_2045,N_1614,N_1234);
xnor U2046 (N_2046,N_1787,N_1452);
nor U2047 (N_2047,N_1208,N_1632);
xor U2048 (N_2048,N_1429,N_1641);
xor U2049 (N_2049,N_1595,N_1561);
and U2050 (N_2050,N_1294,N_1559);
or U2051 (N_2051,N_1740,N_1766);
nor U2052 (N_2052,N_1592,N_1397);
nand U2053 (N_2053,N_1562,N_1336);
xnor U2054 (N_2054,N_1780,N_1468);
and U2055 (N_2055,N_1738,N_1310);
or U2056 (N_2056,N_1405,N_1719);
nor U2057 (N_2057,N_1652,N_1643);
and U2058 (N_2058,N_1525,N_1393);
nor U2059 (N_2059,N_1478,N_1483);
nor U2060 (N_2060,N_1426,N_1541);
nor U2061 (N_2061,N_1654,N_1520);
or U2062 (N_2062,N_1797,N_1694);
nand U2063 (N_2063,N_1324,N_1534);
nor U2064 (N_2064,N_1284,N_1276);
nor U2065 (N_2065,N_1364,N_1556);
nand U2066 (N_2066,N_1286,N_1782);
xnor U2067 (N_2067,N_1724,N_1613);
or U2068 (N_2068,N_1725,N_1400);
and U2069 (N_2069,N_1502,N_1343);
or U2070 (N_2070,N_1217,N_1767);
or U2071 (N_2071,N_1443,N_1339);
or U2072 (N_2072,N_1348,N_1253);
xor U2073 (N_2073,N_1625,N_1626);
and U2074 (N_2074,N_1340,N_1491);
or U2075 (N_2075,N_1231,N_1683);
nand U2076 (N_2076,N_1636,N_1402);
and U2077 (N_2077,N_1510,N_1230);
or U2078 (N_2078,N_1796,N_1440);
nand U2079 (N_2079,N_1573,N_1470);
and U2080 (N_2080,N_1450,N_1531);
nand U2081 (N_2081,N_1240,N_1205);
xnor U2082 (N_2082,N_1532,N_1494);
xor U2083 (N_2083,N_1482,N_1503);
or U2084 (N_2084,N_1437,N_1204);
xor U2085 (N_2085,N_1729,N_1282);
or U2086 (N_2086,N_1565,N_1707);
nor U2087 (N_2087,N_1430,N_1238);
xnor U2088 (N_2088,N_1366,N_1735);
or U2089 (N_2089,N_1265,N_1605);
or U2090 (N_2090,N_1570,N_1266);
and U2091 (N_2091,N_1506,N_1785);
or U2092 (N_2092,N_1495,N_1325);
nand U2093 (N_2093,N_1505,N_1381);
and U2094 (N_2094,N_1666,N_1359);
xnor U2095 (N_2095,N_1685,N_1580);
nor U2096 (N_2096,N_1571,N_1267);
nor U2097 (N_2097,N_1705,N_1264);
nand U2098 (N_2098,N_1634,N_1337);
and U2099 (N_2099,N_1355,N_1745);
nand U2100 (N_2100,N_1677,N_1227);
nand U2101 (N_2101,N_1624,N_1242);
nor U2102 (N_2102,N_1447,N_1491);
nand U2103 (N_2103,N_1658,N_1350);
nor U2104 (N_2104,N_1667,N_1714);
xor U2105 (N_2105,N_1368,N_1470);
nor U2106 (N_2106,N_1606,N_1777);
nand U2107 (N_2107,N_1305,N_1284);
nand U2108 (N_2108,N_1677,N_1519);
nand U2109 (N_2109,N_1340,N_1573);
nor U2110 (N_2110,N_1506,N_1485);
nand U2111 (N_2111,N_1226,N_1669);
or U2112 (N_2112,N_1291,N_1295);
xor U2113 (N_2113,N_1713,N_1737);
or U2114 (N_2114,N_1543,N_1284);
xnor U2115 (N_2115,N_1326,N_1431);
nand U2116 (N_2116,N_1357,N_1504);
nor U2117 (N_2117,N_1715,N_1332);
nand U2118 (N_2118,N_1601,N_1210);
and U2119 (N_2119,N_1243,N_1318);
or U2120 (N_2120,N_1396,N_1318);
or U2121 (N_2121,N_1422,N_1306);
nor U2122 (N_2122,N_1268,N_1690);
xor U2123 (N_2123,N_1287,N_1672);
and U2124 (N_2124,N_1667,N_1210);
and U2125 (N_2125,N_1602,N_1500);
and U2126 (N_2126,N_1614,N_1331);
xnor U2127 (N_2127,N_1445,N_1781);
and U2128 (N_2128,N_1453,N_1416);
nor U2129 (N_2129,N_1503,N_1691);
nand U2130 (N_2130,N_1353,N_1705);
or U2131 (N_2131,N_1520,N_1273);
nor U2132 (N_2132,N_1514,N_1641);
and U2133 (N_2133,N_1213,N_1652);
or U2134 (N_2134,N_1580,N_1409);
or U2135 (N_2135,N_1508,N_1424);
xnor U2136 (N_2136,N_1561,N_1349);
nand U2137 (N_2137,N_1689,N_1383);
or U2138 (N_2138,N_1567,N_1634);
xor U2139 (N_2139,N_1702,N_1299);
xor U2140 (N_2140,N_1528,N_1363);
nand U2141 (N_2141,N_1433,N_1497);
nand U2142 (N_2142,N_1400,N_1337);
and U2143 (N_2143,N_1510,N_1466);
and U2144 (N_2144,N_1544,N_1680);
and U2145 (N_2145,N_1205,N_1680);
nor U2146 (N_2146,N_1609,N_1765);
nand U2147 (N_2147,N_1390,N_1486);
or U2148 (N_2148,N_1372,N_1611);
nand U2149 (N_2149,N_1509,N_1725);
xor U2150 (N_2150,N_1349,N_1790);
or U2151 (N_2151,N_1300,N_1497);
and U2152 (N_2152,N_1287,N_1710);
or U2153 (N_2153,N_1614,N_1368);
xnor U2154 (N_2154,N_1732,N_1241);
nor U2155 (N_2155,N_1383,N_1223);
nand U2156 (N_2156,N_1693,N_1377);
and U2157 (N_2157,N_1246,N_1329);
nand U2158 (N_2158,N_1781,N_1388);
xor U2159 (N_2159,N_1415,N_1506);
and U2160 (N_2160,N_1570,N_1285);
nand U2161 (N_2161,N_1576,N_1287);
xnor U2162 (N_2162,N_1410,N_1399);
xor U2163 (N_2163,N_1454,N_1584);
and U2164 (N_2164,N_1355,N_1270);
and U2165 (N_2165,N_1402,N_1215);
or U2166 (N_2166,N_1433,N_1558);
or U2167 (N_2167,N_1298,N_1202);
nand U2168 (N_2168,N_1253,N_1691);
nor U2169 (N_2169,N_1468,N_1684);
or U2170 (N_2170,N_1539,N_1225);
and U2171 (N_2171,N_1720,N_1346);
nand U2172 (N_2172,N_1228,N_1675);
or U2173 (N_2173,N_1529,N_1458);
and U2174 (N_2174,N_1386,N_1472);
nand U2175 (N_2175,N_1480,N_1671);
and U2176 (N_2176,N_1628,N_1783);
and U2177 (N_2177,N_1646,N_1774);
or U2178 (N_2178,N_1715,N_1686);
and U2179 (N_2179,N_1632,N_1386);
and U2180 (N_2180,N_1477,N_1632);
or U2181 (N_2181,N_1377,N_1643);
or U2182 (N_2182,N_1522,N_1385);
and U2183 (N_2183,N_1332,N_1474);
or U2184 (N_2184,N_1521,N_1213);
nor U2185 (N_2185,N_1334,N_1265);
nand U2186 (N_2186,N_1719,N_1251);
or U2187 (N_2187,N_1299,N_1617);
or U2188 (N_2188,N_1596,N_1284);
or U2189 (N_2189,N_1767,N_1234);
or U2190 (N_2190,N_1533,N_1447);
nand U2191 (N_2191,N_1295,N_1350);
or U2192 (N_2192,N_1763,N_1385);
or U2193 (N_2193,N_1510,N_1468);
nand U2194 (N_2194,N_1498,N_1301);
or U2195 (N_2195,N_1319,N_1719);
nand U2196 (N_2196,N_1374,N_1436);
nor U2197 (N_2197,N_1223,N_1415);
nor U2198 (N_2198,N_1211,N_1640);
nor U2199 (N_2199,N_1296,N_1748);
and U2200 (N_2200,N_1776,N_1409);
or U2201 (N_2201,N_1774,N_1628);
or U2202 (N_2202,N_1281,N_1502);
nand U2203 (N_2203,N_1433,N_1614);
nor U2204 (N_2204,N_1242,N_1533);
nand U2205 (N_2205,N_1539,N_1218);
nand U2206 (N_2206,N_1258,N_1729);
or U2207 (N_2207,N_1622,N_1516);
and U2208 (N_2208,N_1474,N_1584);
nor U2209 (N_2209,N_1643,N_1560);
xnor U2210 (N_2210,N_1643,N_1695);
nor U2211 (N_2211,N_1719,N_1270);
nor U2212 (N_2212,N_1664,N_1224);
and U2213 (N_2213,N_1417,N_1247);
nand U2214 (N_2214,N_1411,N_1659);
nor U2215 (N_2215,N_1692,N_1672);
and U2216 (N_2216,N_1431,N_1203);
and U2217 (N_2217,N_1669,N_1435);
and U2218 (N_2218,N_1528,N_1289);
nand U2219 (N_2219,N_1532,N_1424);
nand U2220 (N_2220,N_1379,N_1546);
and U2221 (N_2221,N_1455,N_1372);
or U2222 (N_2222,N_1290,N_1792);
and U2223 (N_2223,N_1287,N_1435);
xor U2224 (N_2224,N_1208,N_1748);
or U2225 (N_2225,N_1370,N_1435);
nor U2226 (N_2226,N_1332,N_1355);
and U2227 (N_2227,N_1575,N_1777);
xor U2228 (N_2228,N_1624,N_1679);
xor U2229 (N_2229,N_1528,N_1372);
nor U2230 (N_2230,N_1747,N_1746);
and U2231 (N_2231,N_1430,N_1258);
nand U2232 (N_2232,N_1513,N_1315);
nand U2233 (N_2233,N_1211,N_1309);
nor U2234 (N_2234,N_1560,N_1790);
or U2235 (N_2235,N_1226,N_1757);
xor U2236 (N_2236,N_1332,N_1278);
or U2237 (N_2237,N_1339,N_1241);
and U2238 (N_2238,N_1747,N_1285);
and U2239 (N_2239,N_1713,N_1710);
or U2240 (N_2240,N_1680,N_1539);
nor U2241 (N_2241,N_1351,N_1701);
or U2242 (N_2242,N_1744,N_1626);
xor U2243 (N_2243,N_1232,N_1725);
or U2244 (N_2244,N_1694,N_1209);
nand U2245 (N_2245,N_1781,N_1489);
nand U2246 (N_2246,N_1794,N_1642);
xnor U2247 (N_2247,N_1682,N_1297);
and U2248 (N_2248,N_1576,N_1370);
or U2249 (N_2249,N_1366,N_1641);
and U2250 (N_2250,N_1787,N_1542);
xnor U2251 (N_2251,N_1738,N_1702);
xnor U2252 (N_2252,N_1344,N_1255);
nand U2253 (N_2253,N_1627,N_1277);
xnor U2254 (N_2254,N_1585,N_1476);
nor U2255 (N_2255,N_1208,N_1230);
xor U2256 (N_2256,N_1619,N_1510);
xnor U2257 (N_2257,N_1210,N_1352);
xnor U2258 (N_2258,N_1549,N_1403);
or U2259 (N_2259,N_1582,N_1628);
nor U2260 (N_2260,N_1613,N_1579);
and U2261 (N_2261,N_1480,N_1571);
xnor U2262 (N_2262,N_1542,N_1585);
xnor U2263 (N_2263,N_1402,N_1709);
nand U2264 (N_2264,N_1222,N_1560);
and U2265 (N_2265,N_1476,N_1724);
or U2266 (N_2266,N_1533,N_1790);
or U2267 (N_2267,N_1733,N_1367);
nor U2268 (N_2268,N_1692,N_1274);
and U2269 (N_2269,N_1227,N_1692);
or U2270 (N_2270,N_1605,N_1689);
and U2271 (N_2271,N_1715,N_1405);
or U2272 (N_2272,N_1765,N_1351);
nand U2273 (N_2273,N_1237,N_1510);
xor U2274 (N_2274,N_1769,N_1404);
nor U2275 (N_2275,N_1607,N_1610);
xnor U2276 (N_2276,N_1359,N_1421);
or U2277 (N_2277,N_1681,N_1267);
nor U2278 (N_2278,N_1388,N_1482);
and U2279 (N_2279,N_1591,N_1284);
nor U2280 (N_2280,N_1555,N_1467);
or U2281 (N_2281,N_1262,N_1236);
xor U2282 (N_2282,N_1262,N_1695);
xor U2283 (N_2283,N_1232,N_1658);
nor U2284 (N_2284,N_1525,N_1272);
nand U2285 (N_2285,N_1783,N_1726);
and U2286 (N_2286,N_1327,N_1350);
nand U2287 (N_2287,N_1634,N_1422);
and U2288 (N_2288,N_1208,N_1600);
nand U2289 (N_2289,N_1774,N_1246);
and U2290 (N_2290,N_1776,N_1661);
nand U2291 (N_2291,N_1788,N_1345);
nand U2292 (N_2292,N_1369,N_1600);
or U2293 (N_2293,N_1711,N_1702);
or U2294 (N_2294,N_1201,N_1795);
nor U2295 (N_2295,N_1280,N_1394);
nor U2296 (N_2296,N_1664,N_1460);
xor U2297 (N_2297,N_1623,N_1310);
xor U2298 (N_2298,N_1325,N_1613);
nand U2299 (N_2299,N_1451,N_1455);
nor U2300 (N_2300,N_1499,N_1346);
nand U2301 (N_2301,N_1229,N_1556);
nor U2302 (N_2302,N_1793,N_1647);
nor U2303 (N_2303,N_1660,N_1753);
or U2304 (N_2304,N_1298,N_1243);
or U2305 (N_2305,N_1495,N_1419);
xnor U2306 (N_2306,N_1568,N_1421);
xor U2307 (N_2307,N_1608,N_1441);
nand U2308 (N_2308,N_1758,N_1713);
or U2309 (N_2309,N_1295,N_1337);
xnor U2310 (N_2310,N_1501,N_1616);
nor U2311 (N_2311,N_1736,N_1455);
nor U2312 (N_2312,N_1281,N_1641);
or U2313 (N_2313,N_1509,N_1762);
xnor U2314 (N_2314,N_1550,N_1753);
nor U2315 (N_2315,N_1359,N_1643);
and U2316 (N_2316,N_1493,N_1220);
or U2317 (N_2317,N_1341,N_1461);
and U2318 (N_2318,N_1340,N_1456);
and U2319 (N_2319,N_1746,N_1538);
nand U2320 (N_2320,N_1681,N_1711);
xnor U2321 (N_2321,N_1307,N_1782);
xor U2322 (N_2322,N_1798,N_1703);
or U2323 (N_2323,N_1597,N_1519);
xor U2324 (N_2324,N_1642,N_1594);
nand U2325 (N_2325,N_1360,N_1272);
and U2326 (N_2326,N_1587,N_1580);
nand U2327 (N_2327,N_1716,N_1493);
nor U2328 (N_2328,N_1606,N_1575);
nor U2329 (N_2329,N_1641,N_1719);
or U2330 (N_2330,N_1637,N_1444);
xor U2331 (N_2331,N_1595,N_1451);
xnor U2332 (N_2332,N_1639,N_1670);
xor U2333 (N_2333,N_1404,N_1473);
or U2334 (N_2334,N_1690,N_1608);
nor U2335 (N_2335,N_1620,N_1570);
nor U2336 (N_2336,N_1704,N_1424);
nor U2337 (N_2337,N_1495,N_1674);
nand U2338 (N_2338,N_1415,N_1281);
nor U2339 (N_2339,N_1246,N_1511);
and U2340 (N_2340,N_1422,N_1374);
or U2341 (N_2341,N_1734,N_1578);
nor U2342 (N_2342,N_1301,N_1579);
nand U2343 (N_2343,N_1200,N_1417);
nand U2344 (N_2344,N_1585,N_1297);
or U2345 (N_2345,N_1462,N_1622);
xor U2346 (N_2346,N_1486,N_1247);
nand U2347 (N_2347,N_1454,N_1418);
xor U2348 (N_2348,N_1421,N_1785);
or U2349 (N_2349,N_1734,N_1209);
nor U2350 (N_2350,N_1426,N_1338);
or U2351 (N_2351,N_1372,N_1635);
nor U2352 (N_2352,N_1594,N_1314);
or U2353 (N_2353,N_1228,N_1244);
or U2354 (N_2354,N_1612,N_1720);
and U2355 (N_2355,N_1583,N_1693);
nand U2356 (N_2356,N_1423,N_1609);
and U2357 (N_2357,N_1448,N_1466);
nor U2358 (N_2358,N_1309,N_1688);
or U2359 (N_2359,N_1672,N_1427);
nand U2360 (N_2360,N_1737,N_1706);
or U2361 (N_2361,N_1495,N_1617);
and U2362 (N_2362,N_1685,N_1482);
nor U2363 (N_2363,N_1622,N_1442);
or U2364 (N_2364,N_1553,N_1547);
and U2365 (N_2365,N_1664,N_1603);
xnor U2366 (N_2366,N_1403,N_1287);
nand U2367 (N_2367,N_1376,N_1648);
nor U2368 (N_2368,N_1736,N_1422);
xor U2369 (N_2369,N_1309,N_1347);
xnor U2370 (N_2370,N_1276,N_1775);
and U2371 (N_2371,N_1314,N_1554);
xnor U2372 (N_2372,N_1570,N_1618);
nor U2373 (N_2373,N_1597,N_1436);
nand U2374 (N_2374,N_1546,N_1342);
or U2375 (N_2375,N_1690,N_1703);
nand U2376 (N_2376,N_1426,N_1223);
or U2377 (N_2377,N_1704,N_1387);
nand U2378 (N_2378,N_1408,N_1507);
nand U2379 (N_2379,N_1242,N_1387);
xor U2380 (N_2380,N_1456,N_1767);
xor U2381 (N_2381,N_1222,N_1452);
xor U2382 (N_2382,N_1592,N_1256);
xnor U2383 (N_2383,N_1345,N_1324);
xnor U2384 (N_2384,N_1452,N_1479);
nor U2385 (N_2385,N_1536,N_1201);
xnor U2386 (N_2386,N_1252,N_1778);
xnor U2387 (N_2387,N_1507,N_1730);
nand U2388 (N_2388,N_1705,N_1785);
nand U2389 (N_2389,N_1727,N_1689);
or U2390 (N_2390,N_1384,N_1436);
or U2391 (N_2391,N_1262,N_1255);
nor U2392 (N_2392,N_1438,N_1581);
and U2393 (N_2393,N_1418,N_1553);
and U2394 (N_2394,N_1377,N_1761);
or U2395 (N_2395,N_1220,N_1720);
xnor U2396 (N_2396,N_1299,N_1316);
and U2397 (N_2397,N_1491,N_1414);
and U2398 (N_2398,N_1213,N_1423);
or U2399 (N_2399,N_1583,N_1355);
and U2400 (N_2400,N_2151,N_2290);
nor U2401 (N_2401,N_2355,N_2133);
or U2402 (N_2402,N_2018,N_2137);
or U2403 (N_2403,N_2156,N_2313);
and U2404 (N_2404,N_2061,N_1850);
nand U2405 (N_2405,N_2241,N_2307);
or U2406 (N_2406,N_1914,N_2054);
nor U2407 (N_2407,N_2315,N_2078);
xor U2408 (N_2408,N_2038,N_2396);
and U2409 (N_2409,N_2066,N_1805);
nor U2410 (N_2410,N_1870,N_2282);
nand U2411 (N_2411,N_2037,N_2250);
nor U2412 (N_2412,N_2252,N_2164);
xor U2413 (N_2413,N_1866,N_2081);
nor U2414 (N_2414,N_1908,N_2083);
xor U2415 (N_2415,N_1800,N_2311);
xor U2416 (N_2416,N_1835,N_1841);
xnor U2417 (N_2417,N_1912,N_1921);
or U2418 (N_2418,N_2073,N_2016);
and U2419 (N_2419,N_2102,N_1831);
and U2420 (N_2420,N_2035,N_2027);
xor U2421 (N_2421,N_1815,N_2219);
nand U2422 (N_2422,N_2373,N_2058);
nor U2423 (N_2423,N_1966,N_1843);
xnor U2424 (N_2424,N_2295,N_2055);
nor U2425 (N_2425,N_2129,N_2187);
xor U2426 (N_2426,N_1935,N_1829);
nor U2427 (N_2427,N_2049,N_2134);
and U2428 (N_2428,N_2395,N_2214);
nor U2429 (N_2429,N_2003,N_2362);
xor U2430 (N_2430,N_1885,N_2216);
or U2431 (N_2431,N_2240,N_1923);
and U2432 (N_2432,N_2391,N_2008);
nand U2433 (N_2433,N_1849,N_2297);
nor U2434 (N_2434,N_2166,N_2326);
nand U2435 (N_2435,N_2269,N_2077);
nand U2436 (N_2436,N_2284,N_2288);
xor U2437 (N_2437,N_2167,N_1910);
nand U2438 (N_2438,N_1880,N_1937);
or U2439 (N_2439,N_1814,N_2191);
xnor U2440 (N_2440,N_2338,N_1891);
nor U2441 (N_2441,N_1941,N_2186);
xnor U2442 (N_2442,N_2088,N_2000);
or U2443 (N_2443,N_1872,N_2128);
nand U2444 (N_2444,N_2189,N_2169);
xor U2445 (N_2445,N_2356,N_2254);
or U2446 (N_2446,N_1900,N_2063);
nand U2447 (N_2447,N_2152,N_2346);
nor U2448 (N_2448,N_2322,N_2001);
or U2449 (N_2449,N_2183,N_1957);
or U2450 (N_2450,N_1839,N_2217);
or U2451 (N_2451,N_1958,N_2312);
nor U2452 (N_2452,N_1824,N_2354);
or U2453 (N_2453,N_2278,N_2200);
nand U2454 (N_2454,N_2384,N_1960);
nand U2455 (N_2455,N_1931,N_2321);
xnor U2456 (N_2456,N_2230,N_2323);
xor U2457 (N_2457,N_2341,N_2057);
xnor U2458 (N_2458,N_2030,N_2097);
xnor U2459 (N_2459,N_2333,N_2204);
or U2460 (N_2460,N_1846,N_1905);
nor U2461 (N_2461,N_2065,N_1934);
xnor U2462 (N_2462,N_2223,N_1832);
or U2463 (N_2463,N_2387,N_2398);
and U2464 (N_2464,N_2012,N_2122);
and U2465 (N_2465,N_1947,N_1926);
nor U2466 (N_2466,N_2368,N_1907);
and U2467 (N_2467,N_2046,N_2190);
xor U2468 (N_2468,N_1913,N_1946);
or U2469 (N_2469,N_2337,N_1909);
and U2470 (N_2470,N_1896,N_2222);
or U2471 (N_2471,N_2154,N_2064);
xnor U2472 (N_2472,N_2147,N_2267);
nand U2473 (N_2473,N_2013,N_2011);
nand U2474 (N_2474,N_2024,N_2280);
or U2475 (N_2475,N_2221,N_2075);
nand U2476 (N_2476,N_1810,N_2363);
nand U2477 (N_2477,N_2231,N_1901);
or U2478 (N_2478,N_2182,N_2103);
or U2479 (N_2479,N_2386,N_2079);
nor U2480 (N_2480,N_2270,N_2175);
and U2481 (N_2481,N_1970,N_2101);
xor U2482 (N_2482,N_1986,N_2366);
xnor U2483 (N_2483,N_1916,N_2381);
and U2484 (N_2484,N_2388,N_1995);
or U2485 (N_2485,N_1992,N_2379);
nand U2486 (N_2486,N_2143,N_1857);
xor U2487 (N_2487,N_2202,N_2115);
and U2488 (N_2488,N_1959,N_2275);
or U2489 (N_2489,N_1821,N_1886);
nand U2490 (N_2490,N_2328,N_2113);
nor U2491 (N_2491,N_2244,N_2385);
xnor U2492 (N_2492,N_2159,N_2291);
nand U2493 (N_2493,N_2068,N_2043);
and U2494 (N_2494,N_1943,N_2098);
nor U2495 (N_2495,N_2274,N_1884);
nand U2496 (N_2496,N_2324,N_2399);
and U2497 (N_2497,N_1915,N_2005);
nand U2498 (N_2498,N_1848,N_2150);
and U2499 (N_2499,N_2161,N_2339);
nor U2500 (N_2500,N_2148,N_2184);
and U2501 (N_2501,N_1836,N_2076);
and U2502 (N_2502,N_1894,N_1962);
or U2503 (N_2503,N_2237,N_2211);
or U2504 (N_2504,N_1816,N_1989);
nor U2505 (N_2505,N_2041,N_2296);
and U2506 (N_2506,N_1979,N_1906);
nor U2507 (N_2507,N_2380,N_2032);
xnor U2508 (N_2508,N_1889,N_1869);
xnor U2509 (N_2509,N_2091,N_2242);
nand U2510 (N_2510,N_2365,N_2050);
and U2511 (N_2511,N_2198,N_2201);
nand U2512 (N_2512,N_1903,N_2085);
and U2513 (N_2513,N_2162,N_2273);
xnor U2514 (N_2514,N_1855,N_2177);
xnor U2515 (N_2515,N_2114,N_1878);
nand U2516 (N_2516,N_1830,N_1961);
xor U2517 (N_2517,N_2236,N_1871);
nand U2518 (N_2518,N_2149,N_1892);
nor U2519 (N_2519,N_2206,N_1936);
or U2520 (N_2520,N_2144,N_1840);
nor U2521 (N_2521,N_1801,N_1985);
nand U2522 (N_2522,N_2369,N_1822);
xnor U2523 (N_2523,N_2095,N_1924);
or U2524 (N_2524,N_1945,N_2319);
nor U2525 (N_2525,N_2359,N_2263);
nor U2526 (N_2526,N_2262,N_2199);
xor U2527 (N_2527,N_2256,N_1968);
xor U2528 (N_2528,N_2330,N_2364);
nor U2529 (N_2529,N_1953,N_2350);
nor U2530 (N_2530,N_2245,N_2051);
and U2531 (N_2531,N_1873,N_2357);
and U2532 (N_2532,N_2180,N_1833);
nand U2533 (N_2533,N_1991,N_1812);
nor U2534 (N_2534,N_2179,N_2228);
or U2535 (N_2535,N_2220,N_2099);
or U2536 (N_2536,N_2232,N_2303);
and U2537 (N_2537,N_2253,N_1825);
or U2538 (N_2538,N_1838,N_2208);
nand U2539 (N_2539,N_1965,N_2344);
and U2540 (N_2540,N_1852,N_2185);
or U2541 (N_2541,N_1997,N_2142);
nand U2542 (N_2542,N_2139,N_2020);
nand U2543 (N_2543,N_1863,N_2268);
nand U2544 (N_2544,N_2210,N_1851);
nand U2545 (N_2545,N_2358,N_2233);
or U2546 (N_2546,N_1944,N_2304);
xor U2547 (N_2547,N_2209,N_2034);
and U2548 (N_2548,N_2048,N_2308);
nor U2549 (N_2549,N_2004,N_2009);
or U2550 (N_2550,N_1974,N_1955);
or U2551 (N_2551,N_2094,N_1980);
and U2552 (N_2552,N_2314,N_2173);
or U2553 (N_2553,N_2397,N_1802);
nor U2554 (N_2554,N_2255,N_2086);
and U2555 (N_2555,N_1932,N_2195);
nor U2556 (N_2556,N_1879,N_2377);
xnor U2557 (N_2557,N_2383,N_2006);
or U2558 (N_2558,N_2002,N_1925);
nand U2559 (N_2559,N_2272,N_2372);
nand U2560 (N_2560,N_2259,N_1976);
and U2561 (N_2561,N_2170,N_2132);
or U2562 (N_2562,N_2082,N_2203);
nand U2563 (N_2563,N_2087,N_2286);
nand U2564 (N_2564,N_1876,N_1939);
and U2565 (N_2565,N_2021,N_1977);
nand U2566 (N_2566,N_2276,N_1862);
or U2567 (N_2567,N_2136,N_2145);
and U2568 (N_2568,N_1996,N_1809);
xor U2569 (N_2569,N_2243,N_1856);
xnor U2570 (N_2570,N_1823,N_2109);
or U2571 (N_2571,N_1893,N_2026);
nor U2572 (N_2572,N_1881,N_2347);
xor U2573 (N_2573,N_2155,N_2153);
xor U2574 (N_2574,N_2394,N_1911);
nand U2575 (N_2575,N_2335,N_1888);
or U2576 (N_2576,N_2067,N_1868);
or U2577 (N_2577,N_2258,N_2040);
and U2578 (N_2578,N_2092,N_1969);
and U2579 (N_2579,N_2140,N_2205);
or U2580 (N_2580,N_2281,N_2126);
or U2581 (N_2581,N_2053,N_2039);
xnor U2582 (N_2582,N_2014,N_2283);
and U2583 (N_2583,N_2264,N_1883);
nand U2584 (N_2584,N_1983,N_2375);
nand U2585 (N_2585,N_1927,N_2171);
or U2586 (N_2586,N_2289,N_1948);
or U2587 (N_2587,N_2163,N_2285);
nor U2588 (N_2588,N_1972,N_1919);
and U2589 (N_2589,N_2251,N_1949);
nor U2590 (N_2590,N_2160,N_2127);
xnor U2591 (N_2591,N_2349,N_2080);
nand U2592 (N_2592,N_1845,N_2125);
xnor U2593 (N_2593,N_2192,N_2010);
nor U2594 (N_2594,N_2112,N_1820);
nor U2595 (N_2595,N_2023,N_2239);
and U2596 (N_2596,N_2089,N_1973);
xor U2597 (N_2597,N_1950,N_2389);
xnor U2598 (N_2598,N_2279,N_1837);
nor U2599 (N_2599,N_2332,N_1933);
nand U2600 (N_2600,N_2334,N_1867);
xor U2601 (N_2601,N_1864,N_1813);
or U2602 (N_2602,N_1827,N_1828);
xor U2603 (N_2603,N_2271,N_2093);
xor U2604 (N_2604,N_2052,N_1844);
nand U2605 (N_2605,N_1817,N_2360);
nand U2606 (N_2606,N_2056,N_2172);
nand U2607 (N_2607,N_2025,N_1895);
and U2608 (N_2608,N_2292,N_2351);
nor U2609 (N_2609,N_1963,N_2320);
xnor U2610 (N_2610,N_2100,N_2111);
and U2611 (N_2611,N_1865,N_1982);
or U2612 (N_2612,N_1858,N_2188);
xnor U2613 (N_2613,N_2108,N_1806);
nand U2614 (N_2614,N_1808,N_1951);
nand U2615 (N_2615,N_1819,N_2168);
nor U2616 (N_2616,N_2044,N_2331);
nand U2617 (N_2617,N_1918,N_2124);
or U2618 (N_2618,N_2107,N_1842);
or U2619 (N_2619,N_1834,N_2261);
nor U2620 (N_2620,N_2353,N_2022);
nor U2621 (N_2621,N_1930,N_2120);
nor U2622 (N_2622,N_2227,N_1861);
and U2623 (N_2623,N_1887,N_2310);
xnor U2624 (N_2624,N_1818,N_2249);
or U2625 (N_2625,N_2226,N_2352);
xnor U2626 (N_2626,N_2225,N_2104);
or U2627 (N_2627,N_2327,N_2235);
nand U2628 (N_2628,N_2300,N_2135);
xnor U2629 (N_2629,N_2033,N_2309);
nor U2630 (N_2630,N_2141,N_1938);
nor U2631 (N_2631,N_2106,N_2117);
or U2632 (N_2632,N_2130,N_1999);
nor U2633 (N_2633,N_2340,N_2090);
nor U2634 (N_2634,N_2325,N_1890);
nand U2635 (N_2635,N_2116,N_2376);
xnor U2636 (N_2636,N_2007,N_2345);
or U2637 (N_2637,N_2131,N_2302);
or U2638 (N_2638,N_1981,N_1854);
and U2639 (N_2639,N_2301,N_1811);
nand U2640 (N_2640,N_2316,N_2294);
or U2641 (N_2641,N_1994,N_2181);
and U2642 (N_2642,N_1874,N_2390);
nor U2643 (N_2643,N_1803,N_2348);
xnor U2644 (N_2644,N_2146,N_2382);
nand U2645 (N_2645,N_1860,N_2047);
nand U2646 (N_2646,N_2118,N_2028);
or U2647 (N_2647,N_1882,N_1978);
nor U2648 (N_2648,N_1897,N_1804);
or U2649 (N_2649,N_2266,N_1975);
or U2650 (N_2650,N_2277,N_1807);
nor U2651 (N_2651,N_2029,N_2072);
nand U2652 (N_2652,N_2318,N_2196);
xnor U2653 (N_2653,N_1990,N_1859);
xnor U2654 (N_2654,N_2305,N_2306);
and U2655 (N_2655,N_2212,N_2260);
nor U2656 (N_2656,N_2084,N_2343);
and U2657 (N_2657,N_1920,N_2215);
xnor U2658 (N_2658,N_2257,N_2157);
xor U2659 (N_2659,N_2224,N_1998);
and U2660 (N_2660,N_2392,N_2336);
and U2661 (N_2661,N_2207,N_1899);
xor U2662 (N_2662,N_1929,N_2293);
xor U2663 (N_2663,N_2036,N_1956);
nand U2664 (N_2664,N_2017,N_2031);
or U2665 (N_2665,N_2246,N_2062);
and U2666 (N_2666,N_2197,N_1853);
and U2667 (N_2667,N_1988,N_1922);
nor U2668 (N_2668,N_2298,N_1993);
nand U2669 (N_2669,N_1898,N_2238);
and U2670 (N_2670,N_2265,N_1826);
nor U2671 (N_2671,N_2361,N_1847);
nand U2672 (N_2672,N_2248,N_2178);
and U2673 (N_2673,N_2287,N_2234);
and U2674 (N_2674,N_1877,N_2371);
and U2675 (N_2675,N_2158,N_2105);
and U2676 (N_2676,N_2096,N_2194);
xnor U2677 (N_2677,N_2370,N_2299);
nand U2678 (N_2678,N_1940,N_2071);
xor U2679 (N_2679,N_2165,N_2110);
nand U2680 (N_2680,N_1967,N_2123);
nor U2681 (N_2681,N_2138,N_1917);
nand U2682 (N_2682,N_2193,N_2070);
and U2683 (N_2683,N_1952,N_1928);
nor U2684 (N_2684,N_1875,N_1984);
and U2685 (N_2685,N_2074,N_2213);
and U2686 (N_2686,N_2374,N_1904);
or U2687 (N_2687,N_2317,N_1971);
xor U2688 (N_2688,N_1964,N_2329);
or U2689 (N_2689,N_2174,N_2176);
xnor U2690 (N_2690,N_2218,N_2059);
and U2691 (N_2691,N_2393,N_2042);
xor U2692 (N_2692,N_2019,N_2045);
and U2693 (N_2693,N_2069,N_2015);
and U2694 (N_2694,N_2247,N_2342);
nand U2695 (N_2695,N_1954,N_2121);
or U2696 (N_2696,N_2060,N_2378);
xor U2697 (N_2697,N_2119,N_2229);
nand U2698 (N_2698,N_2367,N_1942);
nor U2699 (N_2699,N_1902,N_1987);
nor U2700 (N_2700,N_1928,N_2229);
or U2701 (N_2701,N_2181,N_2073);
nor U2702 (N_2702,N_2398,N_2349);
xor U2703 (N_2703,N_2251,N_2026);
nor U2704 (N_2704,N_2154,N_2327);
xnor U2705 (N_2705,N_2365,N_2163);
and U2706 (N_2706,N_2239,N_2140);
and U2707 (N_2707,N_2297,N_1927);
nand U2708 (N_2708,N_1815,N_1936);
or U2709 (N_2709,N_2129,N_1896);
and U2710 (N_2710,N_1945,N_1848);
or U2711 (N_2711,N_2180,N_2005);
xor U2712 (N_2712,N_1961,N_2252);
nor U2713 (N_2713,N_2341,N_2118);
or U2714 (N_2714,N_1801,N_2064);
nand U2715 (N_2715,N_2373,N_1838);
nand U2716 (N_2716,N_2287,N_1806);
nand U2717 (N_2717,N_1881,N_2019);
or U2718 (N_2718,N_2024,N_1960);
nand U2719 (N_2719,N_1819,N_2197);
or U2720 (N_2720,N_2145,N_1812);
or U2721 (N_2721,N_2186,N_1815);
or U2722 (N_2722,N_2302,N_2355);
nor U2723 (N_2723,N_1996,N_1897);
and U2724 (N_2724,N_1860,N_2357);
xor U2725 (N_2725,N_2179,N_2232);
nand U2726 (N_2726,N_2015,N_2310);
nand U2727 (N_2727,N_2024,N_2167);
xor U2728 (N_2728,N_2145,N_2211);
or U2729 (N_2729,N_2030,N_1986);
or U2730 (N_2730,N_2340,N_2334);
xnor U2731 (N_2731,N_2345,N_2165);
and U2732 (N_2732,N_2326,N_1819);
nand U2733 (N_2733,N_2086,N_2008);
nand U2734 (N_2734,N_1975,N_1981);
and U2735 (N_2735,N_1843,N_2305);
xnor U2736 (N_2736,N_1943,N_2097);
nor U2737 (N_2737,N_1889,N_2041);
and U2738 (N_2738,N_1807,N_1954);
nand U2739 (N_2739,N_2023,N_2301);
nor U2740 (N_2740,N_1942,N_1821);
and U2741 (N_2741,N_2192,N_2166);
xnor U2742 (N_2742,N_2007,N_1854);
xnor U2743 (N_2743,N_2082,N_2257);
xor U2744 (N_2744,N_2234,N_2033);
and U2745 (N_2745,N_2153,N_2352);
nor U2746 (N_2746,N_2213,N_1911);
nor U2747 (N_2747,N_1857,N_2065);
and U2748 (N_2748,N_1941,N_2001);
nand U2749 (N_2749,N_1916,N_2011);
xnor U2750 (N_2750,N_2221,N_2137);
xor U2751 (N_2751,N_2393,N_2011);
or U2752 (N_2752,N_1927,N_2364);
and U2753 (N_2753,N_1808,N_1968);
xnor U2754 (N_2754,N_2031,N_2189);
nand U2755 (N_2755,N_2013,N_1895);
nand U2756 (N_2756,N_2295,N_2272);
nor U2757 (N_2757,N_2020,N_2006);
nand U2758 (N_2758,N_2394,N_1947);
and U2759 (N_2759,N_1987,N_2332);
nor U2760 (N_2760,N_1995,N_2108);
or U2761 (N_2761,N_2398,N_2173);
or U2762 (N_2762,N_1971,N_2332);
nand U2763 (N_2763,N_2215,N_2246);
and U2764 (N_2764,N_2330,N_2177);
and U2765 (N_2765,N_1875,N_1846);
nor U2766 (N_2766,N_2262,N_2137);
or U2767 (N_2767,N_2332,N_1928);
or U2768 (N_2768,N_1837,N_1863);
nand U2769 (N_2769,N_2257,N_1893);
xnor U2770 (N_2770,N_1947,N_2052);
or U2771 (N_2771,N_2142,N_2359);
nor U2772 (N_2772,N_2172,N_1863);
xnor U2773 (N_2773,N_2385,N_2017);
or U2774 (N_2774,N_2379,N_2159);
nand U2775 (N_2775,N_2328,N_2118);
or U2776 (N_2776,N_2185,N_1867);
nor U2777 (N_2777,N_2158,N_2185);
nor U2778 (N_2778,N_1919,N_1815);
and U2779 (N_2779,N_2034,N_2018);
and U2780 (N_2780,N_2345,N_2258);
nand U2781 (N_2781,N_2062,N_2202);
nor U2782 (N_2782,N_2052,N_2068);
xnor U2783 (N_2783,N_2159,N_1809);
or U2784 (N_2784,N_1858,N_1922);
nand U2785 (N_2785,N_2227,N_2195);
and U2786 (N_2786,N_2110,N_2246);
or U2787 (N_2787,N_2213,N_1864);
nor U2788 (N_2788,N_1981,N_2105);
nand U2789 (N_2789,N_2339,N_1880);
nand U2790 (N_2790,N_2276,N_1924);
and U2791 (N_2791,N_1829,N_1821);
nand U2792 (N_2792,N_2022,N_1890);
or U2793 (N_2793,N_2033,N_2379);
and U2794 (N_2794,N_2375,N_2038);
or U2795 (N_2795,N_1965,N_1915);
and U2796 (N_2796,N_2039,N_1954);
nor U2797 (N_2797,N_2361,N_2048);
and U2798 (N_2798,N_2022,N_1952);
and U2799 (N_2799,N_2133,N_2345);
nand U2800 (N_2800,N_2377,N_1901);
and U2801 (N_2801,N_1963,N_2352);
nand U2802 (N_2802,N_1905,N_2233);
xor U2803 (N_2803,N_2033,N_1976);
or U2804 (N_2804,N_1808,N_1929);
nand U2805 (N_2805,N_2360,N_1843);
nand U2806 (N_2806,N_1957,N_1919);
nand U2807 (N_2807,N_2268,N_2233);
or U2808 (N_2808,N_2004,N_1881);
xor U2809 (N_2809,N_2271,N_2312);
nor U2810 (N_2810,N_1940,N_2126);
nand U2811 (N_2811,N_1977,N_2293);
xor U2812 (N_2812,N_2142,N_1922);
xnor U2813 (N_2813,N_2221,N_2293);
or U2814 (N_2814,N_2319,N_2145);
or U2815 (N_2815,N_1963,N_1942);
nor U2816 (N_2816,N_2006,N_2352);
and U2817 (N_2817,N_2207,N_1823);
xor U2818 (N_2818,N_1840,N_2026);
nand U2819 (N_2819,N_2235,N_1859);
nand U2820 (N_2820,N_2240,N_1818);
xor U2821 (N_2821,N_2303,N_1849);
and U2822 (N_2822,N_1860,N_2027);
nor U2823 (N_2823,N_2077,N_2258);
and U2824 (N_2824,N_2224,N_2121);
xor U2825 (N_2825,N_2029,N_1836);
xor U2826 (N_2826,N_2168,N_1977);
nor U2827 (N_2827,N_2289,N_2171);
or U2828 (N_2828,N_2276,N_1825);
nor U2829 (N_2829,N_2066,N_2228);
nor U2830 (N_2830,N_2068,N_2239);
xnor U2831 (N_2831,N_1959,N_1832);
xor U2832 (N_2832,N_1831,N_1930);
or U2833 (N_2833,N_2243,N_2311);
nor U2834 (N_2834,N_1820,N_1935);
nand U2835 (N_2835,N_2281,N_2003);
xnor U2836 (N_2836,N_2094,N_1880);
nand U2837 (N_2837,N_2074,N_1871);
nor U2838 (N_2838,N_1965,N_2252);
nor U2839 (N_2839,N_2285,N_2374);
nor U2840 (N_2840,N_1896,N_2030);
nor U2841 (N_2841,N_1835,N_1870);
and U2842 (N_2842,N_1915,N_1859);
nor U2843 (N_2843,N_2373,N_2180);
xnor U2844 (N_2844,N_2274,N_2317);
xor U2845 (N_2845,N_2241,N_1813);
or U2846 (N_2846,N_2070,N_1865);
xor U2847 (N_2847,N_2380,N_1932);
nor U2848 (N_2848,N_1860,N_2270);
or U2849 (N_2849,N_1820,N_2245);
xnor U2850 (N_2850,N_1948,N_2089);
xnor U2851 (N_2851,N_2200,N_2013);
or U2852 (N_2852,N_2122,N_2356);
or U2853 (N_2853,N_1890,N_2196);
nand U2854 (N_2854,N_1862,N_2060);
nand U2855 (N_2855,N_2079,N_1890);
or U2856 (N_2856,N_2214,N_1883);
xnor U2857 (N_2857,N_2168,N_2084);
and U2858 (N_2858,N_2221,N_1870);
xnor U2859 (N_2859,N_2311,N_1808);
xnor U2860 (N_2860,N_2093,N_1948);
and U2861 (N_2861,N_1806,N_2086);
xnor U2862 (N_2862,N_2029,N_2117);
nand U2863 (N_2863,N_2117,N_2297);
or U2864 (N_2864,N_2395,N_2147);
xnor U2865 (N_2865,N_2179,N_2052);
nor U2866 (N_2866,N_2163,N_2100);
nor U2867 (N_2867,N_1968,N_1944);
nand U2868 (N_2868,N_2292,N_2247);
or U2869 (N_2869,N_1924,N_2064);
and U2870 (N_2870,N_2150,N_2338);
xor U2871 (N_2871,N_2312,N_2178);
or U2872 (N_2872,N_2048,N_2131);
nand U2873 (N_2873,N_1992,N_1901);
xnor U2874 (N_2874,N_2392,N_2073);
xor U2875 (N_2875,N_1933,N_2048);
nand U2876 (N_2876,N_2155,N_2049);
nand U2877 (N_2877,N_2354,N_2231);
xor U2878 (N_2878,N_2111,N_2102);
xnor U2879 (N_2879,N_2352,N_2379);
nand U2880 (N_2880,N_2267,N_1845);
nor U2881 (N_2881,N_2338,N_1940);
or U2882 (N_2882,N_2055,N_2355);
nand U2883 (N_2883,N_2252,N_2057);
xor U2884 (N_2884,N_2026,N_1826);
and U2885 (N_2885,N_2286,N_2098);
xnor U2886 (N_2886,N_2143,N_2304);
xor U2887 (N_2887,N_1966,N_2002);
and U2888 (N_2888,N_2249,N_2281);
nor U2889 (N_2889,N_1866,N_2352);
nor U2890 (N_2890,N_1913,N_2185);
nor U2891 (N_2891,N_1964,N_1824);
and U2892 (N_2892,N_1910,N_1964);
and U2893 (N_2893,N_1899,N_2000);
and U2894 (N_2894,N_1967,N_1915);
nor U2895 (N_2895,N_1958,N_2124);
nor U2896 (N_2896,N_2112,N_1962);
nand U2897 (N_2897,N_2079,N_2100);
xor U2898 (N_2898,N_2229,N_1964);
nand U2899 (N_2899,N_2121,N_2238);
nor U2900 (N_2900,N_1879,N_2138);
and U2901 (N_2901,N_1833,N_1826);
nand U2902 (N_2902,N_2168,N_1997);
or U2903 (N_2903,N_1900,N_1815);
and U2904 (N_2904,N_2215,N_1929);
xnor U2905 (N_2905,N_1845,N_2008);
xnor U2906 (N_2906,N_2126,N_2187);
nand U2907 (N_2907,N_2282,N_1864);
and U2908 (N_2908,N_2244,N_2317);
xnor U2909 (N_2909,N_1952,N_2156);
nand U2910 (N_2910,N_2184,N_2215);
nand U2911 (N_2911,N_2148,N_1884);
nor U2912 (N_2912,N_2013,N_1930);
xor U2913 (N_2913,N_2137,N_2369);
and U2914 (N_2914,N_1990,N_2307);
nand U2915 (N_2915,N_2057,N_2316);
or U2916 (N_2916,N_1943,N_2233);
xor U2917 (N_2917,N_1951,N_2279);
nand U2918 (N_2918,N_2275,N_2328);
nor U2919 (N_2919,N_1983,N_2351);
and U2920 (N_2920,N_2185,N_2129);
and U2921 (N_2921,N_2015,N_1819);
nor U2922 (N_2922,N_2163,N_2043);
nor U2923 (N_2923,N_2147,N_1915);
and U2924 (N_2924,N_1936,N_2237);
nand U2925 (N_2925,N_2252,N_2249);
nor U2926 (N_2926,N_2377,N_1843);
xnor U2927 (N_2927,N_2350,N_1853);
xor U2928 (N_2928,N_1836,N_1912);
and U2929 (N_2929,N_1869,N_2212);
nand U2930 (N_2930,N_1896,N_1814);
and U2931 (N_2931,N_1990,N_2284);
nand U2932 (N_2932,N_2199,N_2271);
or U2933 (N_2933,N_2081,N_2328);
nor U2934 (N_2934,N_2275,N_1863);
nor U2935 (N_2935,N_1821,N_1972);
or U2936 (N_2936,N_1897,N_2052);
xor U2937 (N_2937,N_2174,N_2399);
nand U2938 (N_2938,N_2145,N_1995);
and U2939 (N_2939,N_1822,N_2125);
nor U2940 (N_2940,N_1834,N_1853);
nand U2941 (N_2941,N_1970,N_2276);
or U2942 (N_2942,N_2077,N_2023);
or U2943 (N_2943,N_1848,N_2371);
or U2944 (N_2944,N_1995,N_2168);
or U2945 (N_2945,N_1926,N_2014);
xnor U2946 (N_2946,N_2188,N_1895);
nor U2947 (N_2947,N_1903,N_2173);
nor U2948 (N_2948,N_2339,N_2086);
nand U2949 (N_2949,N_1907,N_2167);
nand U2950 (N_2950,N_1957,N_2060);
nand U2951 (N_2951,N_1882,N_1888);
nand U2952 (N_2952,N_2241,N_2105);
xor U2953 (N_2953,N_2211,N_1813);
nand U2954 (N_2954,N_2194,N_2253);
and U2955 (N_2955,N_2195,N_2049);
or U2956 (N_2956,N_2130,N_2348);
nor U2957 (N_2957,N_2183,N_2178);
and U2958 (N_2958,N_2104,N_2398);
nor U2959 (N_2959,N_2145,N_2168);
nor U2960 (N_2960,N_2135,N_2111);
nand U2961 (N_2961,N_2150,N_2365);
and U2962 (N_2962,N_2156,N_2120);
xor U2963 (N_2963,N_1862,N_2321);
xor U2964 (N_2964,N_1823,N_2155);
or U2965 (N_2965,N_2381,N_1942);
and U2966 (N_2966,N_2158,N_2184);
xor U2967 (N_2967,N_1825,N_2185);
or U2968 (N_2968,N_1832,N_2226);
nand U2969 (N_2969,N_2358,N_1984);
nor U2970 (N_2970,N_2366,N_1806);
nor U2971 (N_2971,N_2204,N_1965);
nor U2972 (N_2972,N_1884,N_2237);
nand U2973 (N_2973,N_1801,N_2233);
nor U2974 (N_2974,N_2066,N_2056);
nor U2975 (N_2975,N_2172,N_1923);
nand U2976 (N_2976,N_2235,N_2313);
or U2977 (N_2977,N_2106,N_1931);
nor U2978 (N_2978,N_2356,N_1916);
nand U2979 (N_2979,N_2383,N_2169);
xor U2980 (N_2980,N_1966,N_2330);
or U2981 (N_2981,N_2125,N_1814);
nand U2982 (N_2982,N_2259,N_2347);
or U2983 (N_2983,N_1911,N_1837);
or U2984 (N_2984,N_2025,N_2061);
nand U2985 (N_2985,N_2177,N_2063);
nand U2986 (N_2986,N_2158,N_2108);
nand U2987 (N_2987,N_1857,N_2384);
nor U2988 (N_2988,N_2201,N_2117);
xor U2989 (N_2989,N_2190,N_2318);
nand U2990 (N_2990,N_2361,N_2103);
and U2991 (N_2991,N_2228,N_2358);
nor U2992 (N_2992,N_1805,N_2370);
nand U2993 (N_2993,N_2223,N_2121);
nor U2994 (N_2994,N_2052,N_2327);
or U2995 (N_2995,N_2099,N_2002);
and U2996 (N_2996,N_1956,N_2267);
nand U2997 (N_2997,N_2390,N_2168);
nand U2998 (N_2998,N_2228,N_1819);
and U2999 (N_2999,N_2247,N_2232);
or UO_0 (O_0,N_2771,N_2543);
xor UO_1 (O_1,N_2868,N_2716);
and UO_2 (O_2,N_2497,N_2709);
nand UO_3 (O_3,N_2563,N_2812);
nor UO_4 (O_4,N_2718,N_2400);
or UO_5 (O_5,N_2846,N_2991);
or UO_6 (O_6,N_2587,N_2545);
and UO_7 (O_7,N_2479,N_2626);
or UO_8 (O_8,N_2411,N_2614);
and UO_9 (O_9,N_2505,N_2737);
xor UO_10 (O_10,N_2770,N_2474);
nand UO_11 (O_11,N_2939,N_2420);
or UO_12 (O_12,N_2921,N_2572);
nand UO_13 (O_13,N_2819,N_2450);
xor UO_14 (O_14,N_2429,N_2795);
and UO_15 (O_15,N_2944,N_2742);
and UO_16 (O_16,N_2451,N_2849);
nor UO_17 (O_17,N_2647,N_2830);
xor UO_18 (O_18,N_2793,N_2492);
xor UO_19 (O_19,N_2711,N_2606);
or UO_20 (O_20,N_2509,N_2974);
nand UO_21 (O_21,N_2458,N_2982);
or UO_22 (O_22,N_2924,N_2408);
nor UO_23 (O_23,N_2558,N_2759);
nand UO_24 (O_24,N_2950,N_2937);
nand UO_25 (O_25,N_2410,N_2555);
or UO_26 (O_26,N_2705,N_2687);
or UO_27 (O_27,N_2903,N_2964);
nand UO_28 (O_28,N_2895,N_2681);
nand UO_29 (O_29,N_2851,N_2685);
nor UO_30 (O_30,N_2869,N_2710);
and UO_31 (O_31,N_2730,N_2844);
nor UO_32 (O_32,N_2817,N_2569);
xnor UO_33 (O_33,N_2960,N_2578);
nor UO_34 (O_34,N_2740,N_2707);
nand UO_35 (O_35,N_2617,N_2440);
nand UO_36 (O_36,N_2531,N_2412);
nor UO_37 (O_37,N_2931,N_2988);
and UO_38 (O_38,N_2453,N_2955);
nor UO_39 (O_39,N_2632,N_2933);
and UO_40 (O_40,N_2713,N_2579);
nor UO_41 (O_41,N_2719,N_2651);
nand UO_42 (O_42,N_2575,N_2884);
xnor UO_43 (O_43,N_2639,N_2979);
xor UO_44 (O_44,N_2467,N_2739);
and UO_45 (O_45,N_2593,N_2783);
and UO_46 (O_46,N_2946,N_2607);
or UO_47 (O_47,N_2432,N_2715);
nand UO_48 (O_48,N_2422,N_2591);
and UO_49 (O_49,N_2627,N_2965);
nand UO_50 (O_50,N_2640,N_2608);
nand UO_51 (O_51,N_2975,N_2938);
nor UO_52 (O_52,N_2684,N_2989);
and UO_53 (O_53,N_2499,N_2637);
nand UO_54 (O_54,N_2805,N_2860);
or UO_55 (O_55,N_2978,N_2533);
and UO_56 (O_56,N_2417,N_2619);
and UO_57 (O_57,N_2910,N_2642);
nor UO_58 (O_58,N_2724,N_2609);
and UO_59 (O_59,N_2468,N_2953);
nand UO_60 (O_60,N_2403,N_2729);
nor UO_61 (O_61,N_2618,N_2503);
nor UO_62 (O_62,N_2813,N_2706);
or UO_63 (O_63,N_2780,N_2874);
nor UO_64 (O_64,N_2992,N_2465);
and UO_65 (O_65,N_2676,N_2631);
nor UO_66 (O_66,N_2772,N_2732);
nor UO_67 (O_67,N_2947,N_2728);
and UO_68 (O_68,N_2688,N_2776);
and UO_69 (O_69,N_2956,N_2925);
nand UO_70 (O_70,N_2802,N_2641);
nor UO_71 (O_71,N_2501,N_2485);
nand UO_72 (O_72,N_2516,N_2866);
xor UO_73 (O_73,N_2644,N_2424);
and UO_74 (O_74,N_2908,N_2500);
nor UO_75 (O_75,N_2746,N_2514);
nand UO_76 (O_76,N_2784,N_2462);
or UO_77 (O_77,N_2515,N_2405);
xor UO_78 (O_78,N_2835,N_2561);
or UO_79 (O_79,N_2690,N_2804);
xor UO_80 (O_80,N_2611,N_2577);
nand UO_81 (O_81,N_2787,N_2547);
xor UO_82 (O_82,N_2599,N_2550);
xnor UO_83 (O_83,N_2657,N_2472);
xor UO_84 (O_84,N_2527,N_2886);
xnor UO_85 (O_85,N_2562,N_2712);
nand UO_86 (O_86,N_2634,N_2464);
or UO_87 (O_87,N_2686,N_2666);
or UO_88 (O_88,N_2714,N_2494);
or UO_89 (O_89,N_2779,N_2442);
and UO_90 (O_90,N_2794,N_2423);
nor UO_91 (O_91,N_2490,N_2876);
xor UO_92 (O_92,N_2643,N_2894);
and UO_93 (O_93,N_2664,N_2798);
xnor UO_94 (O_94,N_2859,N_2892);
nand UO_95 (O_95,N_2919,N_2801);
xnor UO_96 (O_96,N_2409,N_2778);
nor UO_97 (O_97,N_2855,N_2768);
nor UO_98 (O_98,N_2674,N_2466);
and UO_99 (O_99,N_2504,N_2900);
or UO_100 (O_100,N_2963,N_2736);
and UO_101 (O_101,N_2430,N_2489);
or UO_102 (O_102,N_2506,N_2663);
xor UO_103 (O_103,N_2756,N_2603);
nand UO_104 (O_104,N_2875,N_2620);
nand UO_105 (O_105,N_2404,N_2923);
nand UO_106 (O_106,N_2582,N_2987);
and UO_107 (O_107,N_2590,N_2731);
nand UO_108 (O_108,N_2597,N_2535);
nand UO_109 (O_109,N_2613,N_2808);
and UO_110 (O_110,N_2948,N_2872);
nor UO_111 (O_111,N_2757,N_2822);
xnor UO_112 (O_112,N_2762,N_2751);
nand UO_113 (O_113,N_2616,N_2475);
or UO_114 (O_114,N_2564,N_2668);
xnor UO_115 (O_115,N_2839,N_2702);
xor UO_116 (O_116,N_2915,N_2477);
xor UO_117 (O_117,N_2537,N_2559);
nor UO_118 (O_118,N_2600,N_2445);
nor UO_119 (O_119,N_2897,N_2658);
nor UO_120 (O_120,N_2517,N_2694);
nand UO_121 (O_121,N_2864,N_2754);
xor UO_122 (O_122,N_2806,N_2976);
nand UO_123 (O_123,N_2738,N_2496);
xor UO_124 (O_124,N_2704,N_2434);
nand UO_125 (O_125,N_2788,N_2883);
nor UO_126 (O_126,N_2856,N_2630);
nor UO_127 (O_127,N_2863,N_2461);
nand UO_128 (O_128,N_2867,N_2973);
xnor UO_129 (O_129,N_2548,N_2836);
xor UO_130 (O_130,N_2853,N_2748);
and UO_131 (O_131,N_2495,N_2943);
xor UO_132 (O_132,N_2763,N_2928);
xor UO_133 (O_133,N_2920,N_2692);
and UO_134 (O_134,N_2568,N_2511);
or UO_135 (O_135,N_2435,N_2507);
xnor UO_136 (O_136,N_2598,N_2675);
nand UO_137 (O_137,N_2402,N_2954);
xnor UO_138 (O_138,N_2720,N_2922);
or UO_139 (O_139,N_2602,N_2828);
xnor UO_140 (O_140,N_2695,N_2983);
or UO_141 (O_141,N_2967,N_2588);
nor UO_142 (O_142,N_2749,N_2508);
or UO_143 (O_143,N_2673,N_2528);
xor UO_144 (O_144,N_2436,N_2470);
and UO_145 (O_145,N_2810,N_2857);
nor UO_146 (O_146,N_2469,N_2901);
nand UO_147 (O_147,N_2792,N_2951);
nor UO_148 (O_148,N_2999,N_2907);
nand UO_149 (O_149,N_2833,N_2765);
xor UO_150 (O_150,N_2660,N_2437);
or UO_151 (O_151,N_2913,N_2652);
and UO_152 (O_152,N_2502,N_2530);
and UO_153 (O_153,N_2595,N_2510);
and UO_154 (O_154,N_2821,N_2845);
or UO_155 (O_155,N_2814,N_2483);
xnor UO_156 (O_156,N_2858,N_2957);
xor UO_157 (O_157,N_2743,N_2551);
or UO_158 (O_158,N_2961,N_2522);
or UO_159 (O_159,N_2890,N_2576);
or UO_160 (O_160,N_2952,N_2481);
or UO_161 (O_161,N_2850,N_2993);
or UO_162 (O_162,N_2998,N_2542);
nor UO_163 (O_163,N_2678,N_2916);
or UO_164 (O_164,N_2968,N_2760);
or UO_165 (O_165,N_2661,N_2439);
or UO_166 (O_166,N_2513,N_2985);
nor UO_167 (O_167,N_2520,N_2498);
nand UO_168 (O_168,N_2407,N_2534);
and UO_169 (O_169,N_2766,N_2567);
or UO_170 (O_170,N_2820,N_2841);
xor UO_171 (O_171,N_2428,N_2735);
or UO_172 (O_172,N_2459,N_2460);
or UO_173 (O_173,N_2696,N_2592);
nand UO_174 (O_174,N_2917,N_2902);
nand UO_175 (O_175,N_2940,N_2827);
and UO_176 (O_176,N_2701,N_2689);
or UO_177 (O_177,N_2677,N_2521);
and UO_178 (O_178,N_2905,N_2699);
and UO_179 (O_179,N_2906,N_2977);
or UO_180 (O_180,N_2524,N_2656);
xnor UO_181 (O_181,N_2994,N_2727);
nand UO_182 (O_182,N_2837,N_2764);
nor UO_183 (O_183,N_2529,N_2672);
xnor UO_184 (O_184,N_2838,N_2438);
nand UO_185 (O_185,N_2832,N_2747);
or UO_186 (O_186,N_2476,N_2638);
or UO_187 (O_187,N_2809,N_2544);
xnor UO_188 (O_188,N_2826,N_2726);
nand UO_189 (O_189,N_2636,N_2782);
and UO_190 (O_190,N_2873,N_2899);
nand UO_191 (O_191,N_2717,N_2807);
or UO_192 (O_192,N_2554,N_2816);
or UO_193 (O_193,N_2488,N_2557);
nand UO_194 (O_194,N_2446,N_2654);
nor UO_195 (O_195,N_2777,N_2773);
and UO_196 (O_196,N_2406,N_2421);
xor UO_197 (O_197,N_2862,N_2927);
and UO_198 (O_198,N_2635,N_2444);
or UO_199 (O_199,N_2449,N_2413);
xor UO_200 (O_200,N_2698,N_2518);
nor UO_201 (O_201,N_2478,N_2815);
nor UO_202 (O_202,N_2648,N_2818);
xnor UO_203 (O_203,N_2929,N_2888);
nor UO_204 (O_204,N_2942,N_2659);
nand UO_205 (O_205,N_2538,N_2431);
nand UO_206 (O_206,N_2441,N_2799);
or UO_207 (O_207,N_2725,N_2774);
nand UO_208 (O_208,N_2972,N_2761);
and UO_209 (O_209,N_2452,N_2670);
xnor UO_210 (O_210,N_2848,N_2624);
nand UO_211 (O_211,N_2700,N_2532);
or UO_212 (O_212,N_2893,N_2871);
and UO_213 (O_213,N_2455,N_2553);
nor UO_214 (O_214,N_2854,N_2790);
and UO_215 (O_215,N_2679,N_2891);
or UO_216 (O_216,N_2829,N_2889);
xor UO_217 (O_217,N_2623,N_2448);
nor UO_218 (O_218,N_2825,N_2797);
xor UO_219 (O_219,N_2546,N_2840);
or UO_220 (O_220,N_2693,N_2571);
or UO_221 (O_221,N_2586,N_2811);
nor UO_222 (O_222,N_2791,N_2775);
nand UO_223 (O_223,N_2456,N_2691);
nor UO_224 (O_224,N_2482,N_2615);
and UO_225 (O_225,N_2981,N_2491);
or UO_226 (O_226,N_2789,N_2486);
xnor UO_227 (O_227,N_2433,N_2831);
or UO_228 (O_228,N_2877,N_2512);
or UO_229 (O_229,N_2723,N_2852);
nor UO_230 (O_230,N_2996,N_2669);
or UO_231 (O_231,N_2427,N_2930);
nand UO_232 (O_232,N_2750,N_2912);
or UO_233 (O_233,N_2865,N_2655);
nor UO_234 (O_234,N_2941,N_2904);
nor UO_235 (O_235,N_2758,N_2419);
nor UO_236 (O_236,N_2425,N_2604);
xor UO_237 (O_237,N_2628,N_2580);
or UO_238 (O_238,N_2622,N_2560);
and UO_239 (O_239,N_2414,N_2457);
nor UO_240 (O_240,N_2914,N_2565);
xor UO_241 (O_241,N_2480,N_2682);
xnor UO_242 (O_242,N_2721,N_2583);
and UO_243 (O_243,N_2734,N_2653);
xor UO_244 (O_244,N_2471,N_2573);
xnor UO_245 (O_245,N_2949,N_2443);
nor UO_246 (O_246,N_2484,N_2769);
nand UO_247 (O_247,N_2744,N_2697);
and UO_248 (O_248,N_2898,N_2741);
nand UO_249 (O_249,N_2945,N_2541);
nand UO_250 (O_250,N_2605,N_2980);
or UO_251 (O_251,N_2834,N_2786);
and UO_252 (O_252,N_2882,N_2536);
or UO_253 (O_253,N_2671,N_2847);
or UO_254 (O_254,N_2984,N_2473);
nand UO_255 (O_255,N_2645,N_2416);
and UO_256 (O_256,N_2824,N_2625);
or UO_257 (O_257,N_2881,N_2556);
nor UO_258 (O_258,N_2584,N_2936);
nor UO_259 (O_259,N_2708,N_2552);
nand UO_260 (O_260,N_2447,N_2621);
xnor UO_261 (O_261,N_2997,N_2887);
xor UO_262 (O_262,N_2610,N_2629);
nor UO_263 (O_263,N_2970,N_2896);
nand UO_264 (O_264,N_2540,N_2880);
nand UO_265 (O_265,N_2523,N_2990);
and UO_266 (O_266,N_2935,N_2745);
or UO_267 (O_267,N_2722,N_2526);
or UO_268 (O_268,N_2463,N_2426);
xnor UO_269 (O_269,N_2926,N_2932);
or UO_270 (O_270,N_2909,N_2574);
nor UO_271 (O_271,N_2665,N_2581);
xor UO_272 (O_272,N_2878,N_2601);
nand UO_273 (O_273,N_2454,N_2549);
xnor UO_274 (O_274,N_2823,N_2752);
or UO_275 (O_275,N_2861,N_2879);
xnor UO_276 (O_276,N_2918,N_2800);
nand UO_277 (O_277,N_2959,N_2649);
xor UO_278 (O_278,N_2680,N_2418);
or UO_279 (O_279,N_2870,N_2683);
and UO_280 (O_280,N_2570,N_2962);
xor UO_281 (O_281,N_2585,N_2493);
xnor UO_282 (O_282,N_2667,N_2803);
xor UO_283 (O_283,N_2986,N_2995);
nor UO_284 (O_284,N_2911,N_2796);
nor UO_285 (O_285,N_2753,N_2539);
nand UO_286 (O_286,N_2703,N_2767);
and UO_287 (O_287,N_2487,N_2415);
or UO_288 (O_288,N_2971,N_2612);
and UO_289 (O_289,N_2519,N_2525);
or UO_290 (O_290,N_2842,N_2566);
and UO_291 (O_291,N_2733,N_2594);
xnor UO_292 (O_292,N_2969,N_2662);
nor UO_293 (O_293,N_2885,N_2646);
nor UO_294 (O_294,N_2781,N_2401);
or UO_295 (O_295,N_2958,N_2843);
nor UO_296 (O_296,N_2589,N_2755);
nand UO_297 (O_297,N_2966,N_2785);
and UO_298 (O_298,N_2650,N_2934);
nor UO_299 (O_299,N_2633,N_2596);
nand UO_300 (O_300,N_2489,N_2794);
and UO_301 (O_301,N_2630,N_2901);
nand UO_302 (O_302,N_2946,N_2763);
and UO_303 (O_303,N_2472,N_2757);
or UO_304 (O_304,N_2553,N_2702);
nor UO_305 (O_305,N_2559,N_2621);
nor UO_306 (O_306,N_2619,N_2808);
xor UO_307 (O_307,N_2703,N_2585);
nand UO_308 (O_308,N_2684,N_2717);
xnor UO_309 (O_309,N_2703,N_2547);
nor UO_310 (O_310,N_2956,N_2973);
xor UO_311 (O_311,N_2752,N_2811);
nor UO_312 (O_312,N_2801,N_2999);
xnor UO_313 (O_313,N_2930,N_2890);
and UO_314 (O_314,N_2543,N_2471);
and UO_315 (O_315,N_2697,N_2938);
xor UO_316 (O_316,N_2576,N_2706);
or UO_317 (O_317,N_2891,N_2427);
nand UO_318 (O_318,N_2700,N_2711);
nand UO_319 (O_319,N_2693,N_2566);
or UO_320 (O_320,N_2565,N_2500);
or UO_321 (O_321,N_2622,N_2544);
or UO_322 (O_322,N_2655,N_2625);
nand UO_323 (O_323,N_2748,N_2993);
and UO_324 (O_324,N_2958,N_2595);
nor UO_325 (O_325,N_2562,N_2910);
and UO_326 (O_326,N_2840,N_2406);
xor UO_327 (O_327,N_2430,N_2575);
nand UO_328 (O_328,N_2585,N_2752);
xor UO_329 (O_329,N_2990,N_2503);
nand UO_330 (O_330,N_2410,N_2771);
nand UO_331 (O_331,N_2566,N_2969);
nand UO_332 (O_332,N_2445,N_2674);
nor UO_333 (O_333,N_2862,N_2826);
nand UO_334 (O_334,N_2466,N_2653);
nor UO_335 (O_335,N_2760,N_2836);
or UO_336 (O_336,N_2610,N_2899);
nand UO_337 (O_337,N_2687,N_2589);
or UO_338 (O_338,N_2694,N_2662);
nor UO_339 (O_339,N_2996,N_2667);
nand UO_340 (O_340,N_2409,N_2413);
and UO_341 (O_341,N_2783,N_2868);
nand UO_342 (O_342,N_2455,N_2687);
xnor UO_343 (O_343,N_2530,N_2831);
xor UO_344 (O_344,N_2624,N_2807);
nor UO_345 (O_345,N_2748,N_2528);
or UO_346 (O_346,N_2567,N_2526);
nor UO_347 (O_347,N_2885,N_2655);
or UO_348 (O_348,N_2421,N_2885);
nand UO_349 (O_349,N_2521,N_2740);
nor UO_350 (O_350,N_2521,N_2510);
xnor UO_351 (O_351,N_2723,N_2722);
and UO_352 (O_352,N_2864,N_2952);
nor UO_353 (O_353,N_2483,N_2591);
and UO_354 (O_354,N_2947,N_2767);
or UO_355 (O_355,N_2900,N_2809);
nand UO_356 (O_356,N_2621,N_2969);
nor UO_357 (O_357,N_2542,N_2577);
nor UO_358 (O_358,N_2649,N_2757);
and UO_359 (O_359,N_2768,N_2542);
xor UO_360 (O_360,N_2441,N_2783);
nand UO_361 (O_361,N_2554,N_2866);
or UO_362 (O_362,N_2908,N_2539);
and UO_363 (O_363,N_2796,N_2644);
xor UO_364 (O_364,N_2869,N_2424);
xnor UO_365 (O_365,N_2787,N_2457);
nor UO_366 (O_366,N_2615,N_2913);
xnor UO_367 (O_367,N_2903,N_2715);
nor UO_368 (O_368,N_2856,N_2436);
xnor UO_369 (O_369,N_2621,N_2457);
or UO_370 (O_370,N_2953,N_2665);
or UO_371 (O_371,N_2892,N_2638);
or UO_372 (O_372,N_2863,N_2949);
nand UO_373 (O_373,N_2402,N_2482);
xnor UO_374 (O_374,N_2463,N_2553);
xor UO_375 (O_375,N_2565,N_2862);
nand UO_376 (O_376,N_2897,N_2809);
nand UO_377 (O_377,N_2963,N_2590);
nand UO_378 (O_378,N_2585,N_2490);
nand UO_379 (O_379,N_2712,N_2601);
nor UO_380 (O_380,N_2421,N_2822);
and UO_381 (O_381,N_2961,N_2826);
xnor UO_382 (O_382,N_2948,N_2551);
and UO_383 (O_383,N_2726,N_2601);
xor UO_384 (O_384,N_2971,N_2769);
and UO_385 (O_385,N_2667,N_2973);
xnor UO_386 (O_386,N_2502,N_2454);
nand UO_387 (O_387,N_2447,N_2516);
or UO_388 (O_388,N_2616,N_2902);
nor UO_389 (O_389,N_2593,N_2664);
xnor UO_390 (O_390,N_2436,N_2930);
or UO_391 (O_391,N_2611,N_2489);
nor UO_392 (O_392,N_2743,N_2690);
nor UO_393 (O_393,N_2732,N_2959);
or UO_394 (O_394,N_2942,N_2959);
or UO_395 (O_395,N_2750,N_2467);
xor UO_396 (O_396,N_2488,N_2837);
nor UO_397 (O_397,N_2478,N_2952);
and UO_398 (O_398,N_2789,N_2931);
xor UO_399 (O_399,N_2586,N_2413);
nor UO_400 (O_400,N_2589,N_2469);
nor UO_401 (O_401,N_2943,N_2536);
or UO_402 (O_402,N_2955,N_2740);
and UO_403 (O_403,N_2635,N_2532);
nand UO_404 (O_404,N_2787,N_2919);
nor UO_405 (O_405,N_2410,N_2929);
and UO_406 (O_406,N_2555,N_2716);
nand UO_407 (O_407,N_2422,N_2681);
nor UO_408 (O_408,N_2511,N_2705);
and UO_409 (O_409,N_2767,N_2411);
nor UO_410 (O_410,N_2847,N_2774);
nor UO_411 (O_411,N_2634,N_2570);
nand UO_412 (O_412,N_2739,N_2577);
xnor UO_413 (O_413,N_2599,N_2892);
xor UO_414 (O_414,N_2569,N_2482);
nor UO_415 (O_415,N_2637,N_2957);
nor UO_416 (O_416,N_2730,N_2987);
nand UO_417 (O_417,N_2625,N_2639);
nor UO_418 (O_418,N_2898,N_2417);
nor UO_419 (O_419,N_2468,N_2880);
or UO_420 (O_420,N_2626,N_2464);
nand UO_421 (O_421,N_2632,N_2512);
xor UO_422 (O_422,N_2804,N_2925);
xor UO_423 (O_423,N_2528,N_2715);
nor UO_424 (O_424,N_2552,N_2520);
or UO_425 (O_425,N_2714,N_2688);
xnor UO_426 (O_426,N_2488,N_2468);
nand UO_427 (O_427,N_2442,N_2445);
nand UO_428 (O_428,N_2878,N_2978);
nor UO_429 (O_429,N_2488,N_2578);
or UO_430 (O_430,N_2620,N_2973);
nand UO_431 (O_431,N_2474,N_2707);
nand UO_432 (O_432,N_2508,N_2864);
nand UO_433 (O_433,N_2462,N_2727);
xnor UO_434 (O_434,N_2400,N_2829);
xor UO_435 (O_435,N_2798,N_2888);
and UO_436 (O_436,N_2977,N_2542);
and UO_437 (O_437,N_2571,N_2797);
nand UO_438 (O_438,N_2609,N_2538);
and UO_439 (O_439,N_2789,N_2601);
nand UO_440 (O_440,N_2470,N_2691);
nand UO_441 (O_441,N_2433,N_2887);
or UO_442 (O_442,N_2677,N_2505);
xnor UO_443 (O_443,N_2929,N_2569);
nor UO_444 (O_444,N_2903,N_2409);
nor UO_445 (O_445,N_2660,N_2495);
nand UO_446 (O_446,N_2587,N_2505);
and UO_447 (O_447,N_2555,N_2798);
and UO_448 (O_448,N_2547,N_2693);
xor UO_449 (O_449,N_2674,N_2745);
nand UO_450 (O_450,N_2800,N_2820);
xnor UO_451 (O_451,N_2727,N_2965);
and UO_452 (O_452,N_2549,N_2460);
nand UO_453 (O_453,N_2880,N_2750);
nand UO_454 (O_454,N_2870,N_2886);
nand UO_455 (O_455,N_2452,N_2908);
or UO_456 (O_456,N_2616,N_2909);
nand UO_457 (O_457,N_2949,N_2541);
and UO_458 (O_458,N_2989,N_2651);
nand UO_459 (O_459,N_2571,N_2462);
xor UO_460 (O_460,N_2612,N_2672);
nand UO_461 (O_461,N_2931,N_2419);
nor UO_462 (O_462,N_2660,N_2904);
or UO_463 (O_463,N_2979,N_2795);
xor UO_464 (O_464,N_2435,N_2486);
xnor UO_465 (O_465,N_2651,N_2415);
or UO_466 (O_466,N_2676,N_2661);
or UO_467 (O_467,N_2960,N_2538);
nand UO_468 (O_468,N_2801,N_2456);
nor UO_469 (O_469,N_2949,N_2557);
or UO_470 (O_470,N_2945,N_2927);
or UO_471 (O_471,N_2861,N_2407);
xor UO_472 (O_472,N_2571,N_2803);
or UO_473 (O_473,N_2941,N_2624);
or UO_474 (O_474,N_2452,N_2699);
and UO_475 (O_475,N_2532,N_2406);
nor UO_476 (O_476,N_2734,N_2680);
nand UO_477 (O_477,N_2554,N_2432);
nand UO_478 (O_478,N_2525,N_2729);
xnor UO_479 (O_479,N_2632,N_2580);
nor UO_480 (O_480,N_2685,N_2597);
or UO_481 (O_481,N_2458,N_2732);
or UO_482 (O_482,N_2510,N_2502);
nor UO_483 (O_483,N_2750,N_2642);
or UO_484 (O_484,N_2964,N_2774);
nand UO_485 (O_485,N_2509,N_2432);
or UO_486 (O_486,N_2900,N_2782);
or UO_487 (O_487,N_2683,N_2904);
and UO_488 (O_488,N_2832,N_2534);
xor UO_489 (O_489,N_2756,N_2624);
and UO_490 (O_490,N_2816,N_2483);
xor UO_491 (O_491,N_2638,N_2755);
and UO_492 (O_492,N_2561,N_2761);
nor UO_493 (O_493,N_2610,N_2564);
nand UO_494 (O_494,N_2638,N_2777);
and UO_495 (O_495,N_2790,N_2418);
nand UO_496 (O_496,N_2855,N_2578);
xor UO_497 (O_497,N_2607,N_2778);
xnor UO_498 (O_498,N_2916,N_2851);
xnor UO_499 (O_499,N_2480,N_2434);
endmodule