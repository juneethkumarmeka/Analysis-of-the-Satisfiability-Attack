module basic_750_5000_1000_25_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_613,In_488);
or U1 (N_1,In_691,In_414);
and U2 (N_2,In_26,In_449);
nor U3 (N_3,In_350,In_31);
and U4 (N_4,In_525,In_423);
nand U5 (N_5,In_621,In_33);
and U6 (N_6,In_651,In_61);
nand U7 (N_7,In_85,In_87);
nand U8 (N_8,In_129,In_642);
or U9 (N_9,In_529,In_729);
nand U10 (N_10,In_665,In_552);
or U11 (N_11,In_340,In_40);
nand U12 (N_12,In_275,In_213);
and U13 (N_13,In_479,In_634);
or U14 (N_14,In_27,In_695);
and U15 (N_15,In_468,In_355);
and U16 (N_16,In_491,In_682);
nor U17 (N_17,In_57,In_389);
or U18 (N_18,In_462,In_317);
and U19 (N_19,In_254,In_186);
and U20 (N_20,In_219,In_240);
or U21 (N_21,In_84,In_282);
or U22 (N_22,In_679,In_56);
nor U23 (N_23,In_302,In_636);
and U24 (N_24,In_654,In_161);
and U25 (N_25,In_615,In_232);
or U26 (N_26,In_141,In_579);
nor U27 (N_27,In_432,In_490);
nand U28 (N_28,In_670,In_363);
and U29 (N_29,In_346,In_660);
nand U30 (N_30,In_256,In_481);
and U31 (N_31,In_405,In_110);
nand U32 (N_32,In_703,In_439);
nor U33 (N_33,In_498,In_699);
or U34 (N_34,In_419,In_473);
nor U35 (N_35,In_112,In_319);
and U36 (N_36,In_569,In_381);
and U37 (N_37,In_179,In_404);
nand U38 (N_38,In_560,In_192);
or U39 (N_39,In_524,In_3);
nor U40 (N_40,In_280,In_140);
nor U41 (N_41,In_215,In_693);
and U42 (N_42,In_422,In_217);
nand U43 (N_43,In_399,In_152);
nor U44 (N_44,In_218,In_597);
nand U45 (N_45,In_290,In_148);
nand U46 (N_46,In_690,In_207);
nor U47 (N_47,In_24,In_721);
or U48 (N_48,In_149,In_630);
nand U49 (N_49,In_644,In_180);
or U50 (N_50,In_728,In_410);
and U51 (N_51,In_611,In_706);
nand U52 (N_52,In_203,In_387);
and U53 (N_53,In_584,In_168);
and U54 (N_54,In_64,In_65);
nand U55 (N_55,In_343,In_132);
nor U56 (N_56,In_412,In_45);
nand U57 (N_57,In_322,In_441);
nor U58 (N_58,In_748,In_133);
nor U59 (N_59,In_469,In_115);
nand U60 (N_60,In_216,In_637);
or U61 (N_61,In_633,In_277);
or U62 (N_62,In_445,In_631);
nor U63 (N_63,In_353,In_22);
nand U64 (N_64,In_80,In_554);
nor U65 (N_65,In_749,In_478);
and U66 (N_66,In_7,In_177);
nand U67 (N_67,In_378,In_538);
and U68 (N_68,In_50,In_233);
or U69 (N_69,In_184,In_106);
or U70 (N_70,In_592,In_204);
nor U71 (N_71,In_402,In_181);
nor U72 (N_72,In_540,In_567);
nor U73 (N_73,In_53,In_513);
nor U74 (N_74,In_361,In_640);
or U75 (N_75,In_608,In_570);
or U76 (N_76,In_362,In_74);
nor U77 (N_77,In_261,In_12);
and U78 (N_78,In_21,In_537);
nand U79 (N_79,In_519,In_121);
or U80 (N_80,In_650,In_542);
or U81 (N_81,In_200,In_103);
and U82 (N_82,In_612,In_398);
or U83 (N_83,In_162,In_551);
or U84 (N_84,In_606,In_20);
nor U85 (N_85,In_167,In_413);
nor U86 (N_86,In_674,In_546);
nor U87 (N_87,In_420,In_466);
nor U88 (N_88,In_616,In_734);
nor U89 (N_89,In_9,In_174);
nand U90 (N_90,In_109,In_298);
and U91 (N_91,In_743,In_605);
nor U92 (N_92,In_197,In_659);
and U93 (N_93,In_514,In_238);
nor U94 (N_94,In_223,In_113);
and U95 (N_95,In_36,In_533);
nand U96 (N_96,In_742,In_212);
or U97 (N_97,In_664,In_658);
and U98 (N_98,In_508,In_723);
and U99 (N_99,In_648,In_484);
or U100 (N_100,In_173,In_596);
nand U101 (N_101,In_672,In_522);
nor U102 (N_102,In_497,In_208);
and U103 (N_103,In_435,In_5);
nand U104 (N_104,In_122,In_252);
or U105 (N_105,In_474,In_334);
nand U106 (N_106,In_75,In_312);
or U107 (N_107,In_725,In_495);
and U108 (N_108,In_158,In_736);
nand U109 (N_109,In_98,In_700);
nor U110 (N_110,In_125,In_507);
or U111 (N_111,In_209,In_194);
and U112 (N_112,In_58,In_460);
nand U113 (N_113,In_726,In_117);
and U114 (N_114,In_587,In_499);
nand U115 (N_115,In_15,In_349);
and U116 (N_116,In_688,In_643);
or U117 (N_117,In_292,In_339);
and U118 (N_118,In_747,In_451);
nand U119 (N_119,In_150,In_684);
or U120 (N_120,In_509,In_573);
nand U121 (N_121,In_701,In_599);
and U122 (N_122,In_702,In_321);
nor U123 (N_123,In_196,In_11);
or U124 (N_124,In_281,In_436);
nand U125 (N_125,In_354,In_301);
nand U126 (N_126,In_520,In_687);
xor U127 (N_127,In_718,In_136);
or U128 (N_128,In_458,In_526);
nand U129 (N_129,In_523,In_234);
and U130 (N_130,In_485,In_467);
or U131 (N_131,In_429,In_376);
and U132 (N_132,In_25,In_308);
nor U133 (N_133,In_328,In_2);
nand U134 (N_134,In_244,In_377);
or U135 (N_135,In_105,In_386);
nand U136 (N_136,In_86,In_257);
nor U137 (N_137,In_144,In_590);
nand U138 (N_138,In_696,In_663);
and U139 (N_139,In_126,In_512);
nor U140 (N_140,In_400,In_657);
and U141 (N_141,In_16,In_323);
or U142 (N_142,In_617,In_395);
nand U143 (N_143,In_639,In_374);
and U144 (N_144,In_543,In_297);
and U145 (N_145,In_245,In_265);
nor U146 (N_146,In_268,In_170);
nor U147 (N_147,In_258,In_190);
and U148 (N_148,In_448,In_0);
nor U149 (N_149,In_384,In_511);
or U150 (N_150,In_37,In_236);
nor U151 (N_151,In_368,In_313);
and U152 (N_152,In_198,In_147);
nand U153 (N_153,In_284,In_171);
or U154 (N_154,In_666,In_437);
nor U155 (N_155,In_576,In_409);
and U156 (N_156,In_250,In_243);
nor U157 (N_157,In_685,In_314);
or U158 (N_158,In_226,In_146);
or U159 (N_159,In_375,In_735);
and U160 (N_160,In_686,In_202);
or U161 (N_161,In_502,In_388);
and U162 (N_162,In_505,In_135);
nand U163 (N_163,In_591,In_273);
or U164 (N_164,In_571,In_553);
and U165 (N_165,In_371,In_338);
nand U166 (N_166,In_272,In_516);
nand U167 (N_167,In_673,In_418);
and U168 (N_168,In_330,In_730);
and U169 (N_169,In_521,In_549);
and U170 (N_170,In_119,In_28);
or U171 (N_171,In_416,In_360);
nor U172 (N_172,In_4,In_506);
nand U173 (N_173,In_626,In_283);
nand U174 (N_174,In_47,In_698);
nand U175 (N_175,In_34,In_603);
nor U176 (N_176,In_607,In_32);
or U177 (N_177,In_391,In_139);
or U178 (N_178,In_475,In_694);
and U179 (N_179,In_138,In_396);
or U180 (N_180,In_310,In_54);
and U181 (N_181,In_604,In_638);
nor U182 (N_182,In_731,In_300);
nand U183 (N_183,In_737,In_421);
nor U184 (N_184,In_348,In_276);
and U185 (N_185,In_18,In_248);
nand U186 (N_186,In_357,In_496);
and U187 (N_187,In_93,In_225);
nor U188 (N_188,In_427,In_438);
nor U189 (N_189,In_30,In_434);
nand U190 (N_190,In_267,In_531);
nor U191 (N_191,In_500,In_46);
nor U192 (N_192,In_588,In_678);
and U193 (N_193,In_189,In_424);
nand U194 (N_194,In_131,In_296);
nor U195 (N_195,In_35,In_315);
nor U196 (N_196,In_380,In_455);
and U197 (N_197,In_707,In_331);
nor U198 (N_198,In_600,In_733);
or U199 (N_199,In_528,In_337);
nor U200 (N_200,In_77,In_137);
or U201 (N_201,N_79,N_172);
and U202 (N_202,N_0,N_186);
nand U203 (N_203,In_14,In_251);
or U204 (N_204,In_403,N_64);
and U205 (N_205,In_622,In_266);
nor U206 (N_206,In_114,In_545);
nor U207 (N_207,In_23,In_714);
or U208 (N_208,In_715,N_101);
or U209 (N_209,N_30,In_472);
or U210 (N_210,N_107,In_394);
nor U211 (N_211,In_536,In_235);
nor U212 (N_212,N_151,N_185);
nand U213 (N_213,N_84,N_118);
nor U214 (N_214,N_10,In_453);
and U215 (N_215,In_556,N_168);
nor U216 (N_216,In_352,In_483);
nor U217 (N_217,In_365,In_704);
or U218 (N_218,In_359,N_35);
xor U219 (N_219,N_182,In_72);
and U220 (N_220,N_193,In_333);
nor U221 (N_221,N_6,In_653);
nand U222 (N_222,In_153,N_98);
or U223 (N_223,In_185,N_125);
or U224 (N_224,In_351,N_160);
or U225 (N_225,In_29,N_12);
nor U226 (N_226,In_318,N_110);
nand U227 (N_227,N_133,In_629);
and U228 (N_228,In_425,In_614);
and U229 (N_229,N_69,N_159);
xor U230 (N_230,In_271,N_1);
nand U231 (N_231,N_131,In_393);
and U232 (N_232,In_182,In_264);
nand U233 (N_233,N_32,N_33);
nor U234 (N_234,In_231,N_102);
nor U235 (N_235,In_585,N_158);
nor U236 (N_236,In_230,N_56);
nand U237 (N_237,In_744,N_5);
nand U238 (N_238,In_548,In_309);
or U239 (N_239,In_246,N_55);
nand U240 (N_240,In_320,N_148);
or U241 (N_241,In_71,In_577);
nor U242 (N_242,In_329,In_345);
and U243 (N_243,In_568,In_172);
nor U244 (N_244,N_156,In_503);
nand U245 (N_245,In_580,In_241);
nor U246 (N_246,N_15,In_527);
xor U247 (N_247,In_183,N_62);
and U248 (N_248,In_652,In_470);
or U249 (N_249,In_289,N_150);
and U250 (N_250,In_123,N_70);
nor U251 (N_251,In_94,N_152);
nand U252 (N_252,N_121,In_681);
nor U253 (N_253,In_683,N_80);
and U254 (N_254,N_138,In_692);
nor U255 (N_255,In_279,N_17);
or U256 (N_256,In_447,N_135);
or U257 (N_257,N_7,In_19);
nor U258 (N_258,In_390,In_440);
xnor U259 (N_259,In_623,N_194);
and U260 (N_260,N_94,In_370);
and U261 (N_261,In_486,In_8);
or U262 (N_262,N_126,N_127);
or U263 (N_263,N_144,In_645);
nor U264 (N_264,In_456,N_13);
or U265 (N_265,In_175,N_8);
nand U266 (N_266,N_191,In_262);
nor U267 (N_267,In_364,In_38);
nand U268 (N_268,In_249,In_48);
or U269 (N_269,In_494,N_36);
and U270 (N_270,In_433,In_515);
and U271 (N_271,In_145,In_534);
or U272 (N_272,In_732,N_143);
or U273 (N_273,In_6,In_708);
nor U274 (N_274,In_489,In_285);
or U275 (N_275,In_214,N_19);
or U276 (N_276,In_510,N_162);
nand U277 (N_277,In_487,N_71);
or U278 (N_278,N_9,In_237);
and U279 (N_279,In_205,In_415);
nand U280 (N_280,In_324,In_259);
and U281 (N_281,In_586,N_173);
nand U282 (N_282,N_14,In_501);
and U283 (N_283,In_111,In_157);
or U284 (N_284,In_201,N_175);
nor U285 (N_285,In_649,In_646);
nand U286 (N_286,In_286,N_60);
nor U287 (N_287,N_111,N_154);
nor U288 (N_288,In_239,In_62);
and U289 (N_289,In_647,In_385);
or U290 (N_290,In_464,In_13);
nand U291 (N_291,In_465,In_332);
nor U292 (N_292,In_547,N_22);
nand U293 (N_293,In_454,In_610);
and U294 (N_294,In_165,In_311);
nand U295 (N_295,In_446,In_66);
or U296 (N_296,In_745,N_176);
or U297 (N_297,N_24,In_293);
nand U298 (N_298,In_482,N_170);
and U299 (N_299,In_697,In_99);
nand U300 (N_300,N_181,In_561);
nor U301 (N_301,In_480,N_42);
nor U302 (N_302,N_140,In_17);
nor U303 (N_303,In_662,In_443);
or U304 (N_304,In_195,In_461);
nand U305 (N_305,In_669,In_134);
nor U306 (N_306,N_96,In_224);
nand U307 (N_307,In_709,In_101);
nor U308 (N_308,In_68,In_169);
nand U309 (N_309,In_722,In_661);
and U310 (N_310,In_555,N_99);
nor U311 (N_311,In_100,N_66);
and U312 (N_312,In_187,In_739);
or U313 (N_313,In_459,In_426);
or U314 (N_314,In_206,In_78);
and U315 (N_315,In_44,N_146);
and U316 (N_316,In_326,N_87);
nand U317 (N_317,In_51,In_431);
or U318 (N_318,In_717,In_740);
or U319 (N_319,In_263,N_54);
nor U320 (N_320,N_184,In_255);
and U321 (N_321,In_581,N_88);
nand U322 (N_322,N_105,In_104);
and U323 (N_323,N_95,N_171);
or U324 (N_324,In_127,In_724);
nand U325 (N_325,In_408,In_583);
nand U326 (N_326,In_620,In_278);
nor U327 (N_327,In_79,N_89);
nand U328 (N_328,N_104,In_595);
nor U329 (N_329,N_86,In_619);
nand U330 (N_330,N_116,N_52);
nand U331 (N_331,N_147,In_70);
and U332 (N_332,In_711,N_2);
nand U333 (N_333,N_37,N_174);
nand U334 (N_334,N_97,In_10);
and U335 (N_335,N_157,In_342);
or U336 (N_336,In_593,N_93);
nand U337 (N_337,N_26,In_76);
or U338 (N_338,In_220,In_287);
nand U339 (N_339,N_92,N_20);
and U340 (N_340,N_68,In_609);
nor U341 (N_341,In_143,In_667);
nor U342 (N_342,In_222,N_166);
nor U343 (N_343,In_713,In_193);
and U344 (N_344,In_305,N_145);
nor U345 (N_345,N_25,In_641);
and U346 (N_346,In_627,In_253);
nor U347 (N_347,In_347,In_720);
and U348 (N_348,N_192,In_392);
nor U349 (N_349,In_383,In_397);
nor U350 (N_350,In_635,In_260);
nor U351 (N_351,In_541,In_582);
nand U352 (N_352,In_166,In_55);
nand U353 (N_353,In_746,N_155);
nor U354 (N_354,N_109,In_199);
and U355 (N_355,In_118,In_299);
or U356 (N_356,In_151,In_457);
nand U357 (N_357,N_169,In_306);
nor U358 (N_358,In_88,In_594);
and U359 (N_359,N_29,In_291);
or U360 (N_360,In_558,In_572);
and U361 (N_361,In_574,N_40);
nand U362 (N_362,In_727,In_471);
or U363 (N_363,N_47,N_183);
or U364 (N_364,In_671,N_177);
nor U365 (N_365,In_689,In_356);
nand U366 (N_366,In_618,N_11);
and U367 (N_367,N_78,In_675);
and U368 (N_368,In_73,In_550);
nor U369 (N_369,In_92,In_96);
nor U370 (N_370,In_304,In_41);
and U371 (N_371,In_379,In_43);
nor U372 (N_372,In_63,In_504);
or U373 (N_373,N_100,In_565);
and U374 (N_374,In_210,N_129);
or U375 (N_375,N_31,N_165);
or U376 (N_376,In_327,N_113);
and U377 (N_377,N_132,N_4);
nand U378 (N_378,N_58,In_130);
and U379 (N_379,In_450,In_69);
nand U380 (N_380,N_38,N_163);
nor U381 (N_381,N_115,In_269);
nand U382 (N_382,In_156,N_122);
nand U383 (N_383,N_136,In_116);
and U384 (N_384,In_82,In_90);
and U385 (N_385,N_114,In_91);
nand U386 (N_386,In_60,N_167);
or U387 (N_387,In_476,N_28);
and U388 (N_388,N_188,In_656);
or U389 (N_389,In_188,N_76);
and U390 (N_390,In_369,In_544);
nand U391 (N_391,In_307,In_625);
nand U392 (N_392,In_710,N_189);
nand U393 (N_393,N_139,In_124);
or U394 (N_394,In_557,N_197);
and U395 (N_395,N_3,N_65);
nor U396 (N_396,N_27,In_444);
nor U397 (N_397,In_539,N_16);
and U398 (N_398,In_367,N_108);
and U399 (N_399,In_417,N_43);
nand U400 (N_400,N_161,N_223);
nor U401 (N_401,N_281,N_265);
or U402 (N_402,In_575,In_344);
or U403 (N_403,N_241,N_119);
nor U404 (N_404,N_249,N_75);
or U405 (N_405,N_352,In_335);
nand U406 (N_406,N_353,In_358);
nor U407 (N_407,In_442,In_295);
nand U408 (N_408,N_124,N_260);
nand U409 (N_409,N_386,N_326);
nand U410 (N_410,In_336,N_378);
nand U411 (N_411,N_219,N_250);
and U412 (N_412,N_85,In_602);
and U413 (N_413,N_313,In_325);
and U414 (N_414,N_289,N_247);
and U415 (N_415,N_51,N_21);
and U416 (N_416,In_366,N_237);
nor U417 (N_417,N_271,N_330);
or U418 (N_418,In_164,In_563);
or U419 (N_419,N_235,N_370);
or U420 (N_420,N_252,In_316);
or U421 (N_421,N_282,In_463);
and U422 (N_422,N_344,N_354);
and U423 (N_423,In_562,N_210);
nand U424 (N_424,N_351,N_345);
nand U425 (N_425,N_216,N_153);
nor U426 (N_426,N_324,N_302);
or U427 (N_427,N_212,N_397);
nor U428 (N_428,In_120,N_375);
and U429 (N_429,N_376,N_343);
nand U430 (N_430,N_205,N_225);
or U431 (N_431,N_303,N_243);
nor U432 (N_432,N_264,In_559);
nor U433 (N_433,N_385,N_310);
nor U434 (N_434,N_23,In_227);
or U435 (N_435,In_294,In_407);
nor U436 (N_436,In_128,In_411);
and U437 (N_437,N_128,N_342);
and U438 (N_438,N_196,N_263);
or U439 (N_439,In_163,In_680);
or U440 (N_440,N_276,N_279);
nor U441 (N_441,N_59,N_256);
nand U442 (N_442,In_535,N_67);
nand U443 (N_443,N_283,N_73);
or U444 (N_444,N_199,In_676);
and U445 (N_445,N_50,N_329);
nor U446 (N_446,N_214,N_284);
nor U447 (N_447,N_295,In_530);
nor U448 (N_448,N_399,N_83);
nand U449 (N_449,N_358,N_338);
nand U450 (N_450,N_206,N_317);
and U451 (N_451,N_379,In_492);
or U452 (N_452,N_164,N_236);
nor U453 (N_453,N_288,N_74);
nand U454 (N_454,N_290,N_201);
nand U455 (N_455,N_287,N_239);
and U456 (N_456,N_323,N_103);
nor U457 (N_457,N_259,N_244);
nor U458 (N_458,In_176,In_274);
nor U459 (N_459,N_200,N_312);
nor U460 (N_460,N_380,N_190);
or U461 (N_461,N_286,N_91);
or U462 (N_462,N_322,N_364);
or U463 (N_463,N_298,N_72);
or U464 (N_464,N_203,N_266);
nor U465 (N_465,In_373,In_452);
or U466 (N_466,In_288,N_275);
and U467 (N_467,N_346,N_278);
and U468 (N_468,N_34,In_81);
nor U469 (N_469,N_44,N_49);
and U470 (N_470,In_178,N_328);
nor U471 (N_471,N_381,In_83);
and U472 (N_472,N_395,N_251);
nor U473 (N_473,N_334,N_384);
or U474 (N_474,N_142,N_293);
nor U475 (N_475,In_589,In_655);
xor U476 (N_476,N_333,N_308);
and U477 (N_477,N_337,N_234);
or U478 (N_478,N_211,In_95);
nand U479 (N_479,N_226,N_359);
nand U480 (N_480,N_269,In_677);
nor U481 (N_481,N_368,In_67);
nor U482 (N_482,In_52,N_382);
nor U483 (N_483,N_82,In_517);
nand U484 (N_484,N_141,In_42);
or U485 (N_485,In_578,N_377);
or U486 (N_486,N_274,N_365);
nand U487 (N_487,N_117,N_292);
or U488 (N_488,N_195,N_217);
or U489 (N_489,N_41,N_149);
nor U490 (N_490,N_187,N_253);
or U491 (N_491,N_215,In_428);
nand U492 (N_492,N_178,In_372);
and U493 (N_493,In_518,In_493);
and U494 (N_494,N_391,N_305);
and U495 (N_495,In_242,N_349);
and U496 (N_496,N_48,N_314);
or U497 (N_497,N_306,N_296);
or U498 (N_498,N_258,N_357);
nor U499 (N_499,In_477,N_304);
and U500 (N_500,In_97,In_632);
or U501 (N_501,N_262,In_430);
and U502 (N_502,N_112,N_207);
nand U503 (N_503,N_394,N_396);
or U504 (N_504,N_309,N_61);
or U505 (N_505,N_350,N_81);
nand U506 (N_506,In_1,N_90);
or U507 (N_507,N_388,In_668);
or U508 (N_508,N_46,N_130);
and U509 (N_509,N_213,N_222);
nor U510 (N_510,In_247,N_340);
and U511 (N_511,N_327,N_341);
or U512 (N_512,N_231,N_392);
and U513 (N_513,N_245,In_628);
nand U514 (N_514,N_387,N_230);
and U515 (N_515,N_356,N_373);
nor U516 (N_516,N_371,N_220);
nand U517 (N_517,N_307,N_285);
nor U518 (N_518,N_248,In_341);
and U519 (N_519,N_228,N_254);
or U520 (N_520,N_272,In_738);
nor U521 (N_521,In_154,In_401);
nand U522 (N_522,N_257,N_347);
nor U523 (N_523,N_355,In_102);
nor U524 (N_524,N_348,N_311);
nand U525 (N_525,N_332,N_360);
and U526 (N_526,N_390,N_268);
nor U527 (N_527,N_369,N_77);
or U528 (N_528,In_49,N_45);
nor U529 (N_529,N_242,N_372);
nor U530 (N_530,In_159,N_106);
nor U531 (N_531,In_705,N_221);
xor U532 (N_532,In_303,In_601);
or U533 (N_533,N_227,In_270);
or U534 (N_534,In_716,N_204);
nand U535 (N_535,N_393,N_374);
nor U536 (N_536,N_363,N_240);
and U537 (N_537,N_180,N_398);
nor U538 (N_538,N_335,In_211);
and U539 (N_539,N_316,N_18);
or U540 (N_540,N_120,N_366);
nor U541 (N_541,In_624,In_406);
nor U542 (N_542,N_218,N_198);
or U543 (N_543,In_39,N_331);
nand U544 (N_544,In_741,N_336);
nand U545 (N_545,N_361,N_321);
or U546 (N_546,N_224,N_383);
nor U547 (N_547,N_209,N_179);
nand U548 (N_548,N_57,N_137);
nand U549 (N_549,In_598,N_246);
or U550 (N_550,In_89,N_39);
nand U551 (N_551,In_191,In_564);
nor U552 (N_552,N_53,N_63);
nand U553 (N_553,N_301,N_367);
and U554 (N_554,N_389,N_291);
nand U555 (N_555,N_233,In_532);
nand U556 (N_556,N_229,N_299);
nor U557 (N_557,N_255,In_229);
nor U558 (N_558,N_273,N_270);
nand U559 (N_559,In_107,In_142);
or U560 (N_560,N_320,N_297);
or U561 (N_561,N_261,N_339);
and U562 (N_562,N_315,In_221);
nor U563 (N_563,N_319,In_566);
or U564 (N_564,N_123,In_719);
or U565 (N_565,In_108,N_325);
nor U566 (N_566,N_208,In_712);
nor U567 (N_567,N_267,In_160);
nand U568 (N_568,N_300,N_134);
nand U569 (N_569,N_238,In_59);
nor U570 (N_570,N_280,N_362);
nor U571 (N_571,N_277,N_318);
nor U572 (N_572,N_232,N_294);
or U573 (N_573,N_202,In_155);
or U574 (N_574,In_382,In_228);
nor U575 (N_575,In_341,In_142);
nor U576 (N_576,N_216,N_354);
or U577 (N_577,N_57,N_204);
and U578 (N_578,N_235,N_134);
nor U579 (N_579,In_530,N_211);
or U580 (N_580,N_361,N_241);
nand U581 (N_581,N_216,N_314);
or U582 (N_582,N_336,N_233);
and U583 (N_583,N_281,N_266);
nor U584 (N_584,N_239,N_332);
and U585 (N_585,N_306,N_263);
and U586 (N_586,N_236,N_372);
and U587 (N_587,N_235,N_336);
and U588 (N_588,N_216,N_90);
nor U589 (N_589,N_221,N_212);
and U590 (N_590,N_264,N_232);
nor U591 (N_591,N_85,N_308);
and U592 (N_592,N_297,N_387);
or U593 (N_593,N_240,N_376);
nand U594 (N_594,N_304,In_566);
and U595 (N_595,N_202,N_63);
or U596 (N_596,N_391,N_296);
xor U597 (N_597,In_176,N_330);
and U598 (N_598,N_281,N_344);
and U599 (N_599,In_242,In_716);
and U600 (N_600,N_557,N_429);
and U601 (N_601,N_546,N_520);
or U602 (N_602,N_423,N_535);
nor U603 (N_603,N_474,N_444);
or U604 (N_604,N_565,N_538);
or U605 (N_605,N_587,N_445);
nand U606 (N_606,N_481,N_564);
or U607 (N_607,N_487,N_446);
nor U608 (N_608,N_456,N_488);
nor U609 (N_609,N_454,N_575);
xor U610 (N_610,N_586,N_553);
nor U611 (N_611,N_509,N_483);
nand U612 (N_612,N_568,N_437);
and U613 (N_613,N_584,N_518);
nand U614 (N_614,N_415,N_545);
or U615 (N_615,N_405,N_489);
or U616 (N_616,N_526,N_473);
nor U617 (N_617,N_468,N_599);
or U618 (N_618,N_537,N_562);
nor U619 (N_619,N_581,N_469);
nand U620 (N_620,N_560,N_515);
or U621 (N_621,N_530,N_470);
or U622 (N_622,N_531,N_578);
nor U623 (N_623,N_449,N_567);
and U624 (N_624,N_506,N_577);
nand U625 (N_625,N_508,N_579);
nor U626 (N_626,N_410,N_421);
and U627 (N_627,N_582,N_401);
and U628 (N_628,N_559,N_527);
or U629 (N_629,N_458,N_498);
and U630 (N_630,N_556,N_490);
nand U631 (N_631,N_521,N_590);
nor U632 (N_632,N_541,N_433);
and U633 (N_633,N_514,N_532);
or U634 (N_634,N_496,N_406);
nand U635 (N_635,N_419,N_432);
nor U636 (N_636,N_443,N_576);
nand U637 (N_637,N_480,N_510);
nand U638 (N_638,N_476,N_484);
nand U639 (N_639,N_422,N_402);
nand U640 (N_640,N_430,N_563);
nor U641 (N_641,N_462,N_504);
or U642 (N_642,N_549,N_441);
or U643 (N_643,N_598,N_517);
and U644 (N_644,N_452,N_569);
and U645 (N_645,N_589,N_417);
or U646 (N_646,N_511,N_548);
or U647 (N_647,N_595,N_447);
nor U648 (N_648,N_594,N_501);
or U649 (N_649,N_466,N_551);
and U650 (N_650,N_412,N_425);
nand U651 (N_651,N_555,N_588);
xor U652 (N_652,N_475,N_513);
nor U653 (N_653,N_516,N_591);
or U654 (N_654,N_547,N_438);
and U655 (N_655,N_550,N_479);
nand U656 (N_656,N_492,N_558);
nor U657 (N_657,N_583,N_554);
nand U658 (N_658,N_497,N_457);
and U659 (N_659,N_442,N_570);
nor U660 (N_660,N_525,N_596);
nor U661 (N_661,N_536,N_428);
or U662 (N_662,N_539,N_420);
or U663 (N_663,N_523,N_505);
nand U664 (N_664,N_404,N_580);
or U665 (N_665,N_407,N_574);
or U666 (N_666,N_403,N_413);
or U667 (N_667,N_435,N_471);
and U668 (N_668,N_512,N_571);
nor U669 (N_669,N_540,N_459);
nand U670 (N_670,N_464,N_500);
nor U671 (N_671,N_585,N_409);
and U672 (N_672,N_593,N_478);
nand U673 (N_673,N_440,N_528);
nor U674 (N_674,N_450,N_461);
nor U675 (N_675,N_529,N_534);
and U676 (N_676,N_542,N_424);
nand U677 (N_677,N_485,N_411);
nand U678 (N_678,N_426,N_453);
nand U679 (N_679,N_482,N_436);
xnor U680 (N_680,N_431,N_499);
or U681 (N_681,N_455,N_486);
nand U682 (N_682,N_472,N_427);
nand U683 (N_683,N_463,N_522);
and U684 (N_684,N_503,N_494);
and U685 (N_685,N_448,N_414);
nand U686 (N_686,N_566,N_434);
nand U687 (N_687,N_495,N_533);
xnor U688 (N_688,N_418,N_460);
or U689 (N_689,N_543,N_544);
nand U690 (N_690,N_451,N_592);
nor U691 (N_691,N_524,N_416);
or U692 (N_692,N_467,N_493);
nor U693 (N_693,N_561,N_502);
nand U694 (N_694,N_597,N_552);
or U695 (N_695,N_572,N_477);
or U696 (N_696,N_465,N_519);
nor U697 (N_697,N_439,N_408);
nand U698 (N_698,N_573,N_507);
nand U699 (N_699,N_491,N_400);
nor U700 (N_700,N_576,N_410);
nor U701 (N_701,N_509,N_468);
or U702 (N_702,N_432,N_595);
nor U703 (N_703,N_590,N_430);
or U704 (N_704,N_484,N_506);
or U705 (N_705,N_561,N_483);
nor U706 (N_706,N_462,N_485);
and U707 (N_707,N_471,N_478);
nand U708 (N_708,N_453,N_436);
or U709 (N_709,N_538,N_552);
and U710 (N_710,N_481,N_577);
nor U711 (N_711,N_404,N_513);
nor U712 (N_712,N_586,N_427);
and U713 (N_713,N_526,N_530);
and U714 (N_714,N_433,N_571);
nor U715 (N_715,N_403,N_478);
nand U716 (N_716,N_555,N_519);
or U717 (N_717,N_571,N_526);
or U718 (N_718,N_498,N_471);
nand U719 (N_719,N_422,N_417);
nand U720 (N_720,N_490,N_510);
nor U721 (N_721,N_532,N_441);
nor U722 (N_722,N_515,N_412);
nand U723 (N_723,N_447,N_543);
or U724 (N_724,N_471,N_567);
or U725 (N_725,N_517,N_512);
nor U726 (N_726,N_596,N_401);
and U727 (N_727,N_453,N_423);
nor U728 (N_728,N_519,N_565);
nor U729 (N_729,N_462,N_598);
and U730 (N_730,N_582,N_596);
nand U731 (N_731,N_466,N_573);
nand U732 (N_732,N_451,N_552);
nor U733 (N_733,N_476,N_491);
or U734 (N_734,N_568,N_483);
or U735 (N_735,N_569,N_553);
nor U736 (N_736,N_478,N_416);
nor U737 (N_737,N_459,N_448);
and U738 (N_738,N_563,N_471);
or U739 (N_739,N_563,N_476);
nor U740 (N_740,N_427,N_492);
or U741 (N_741,N_575,N_405);
nand U742 (N_742,N_422,N_497);
and U743 (N_743,N_486,N_442);
and U744 (N_744,N_438,N_543);
nor U745 (N_745,N_545,N_522);
nor U746 (N_746,N_489,N_521);
and U747 (N_747,N_431,N_412);
and U748 (N_748,N_493,N_411);
and U749 (N_749,N_407,N_451);
or U750 (N_750,N_549,N_463);
nand U751 (N_751,N_432,N_492);
nand U752 (N_752,N_590,N_536);
and U753 (N_753,N_539,N_498);
nor U754 (N_754,N_574,N_417);
and U755 (N_755,N_518,N_476);
or U756 (N_756,N_448,N_468);
and U757 (N_757,N_512,N_521);
and U758 (N_758,N_530,N_438);
nand U759 (N_759,N_506,N_575);
and U760 (N_760,N_558,N_556);
or U761 (N_761,N_518,N_578);
nor U762 (N_762,N_595,N_505);
and U763 (N_763,N_539,N_508);
or U764 (N_764,N_501,N_542);
nand U765 (N_765,N_580,N_429);
nor U766 (N_766,N_535,N_451);
or U767 (N_767,N_561,N_542);
nand U768 (N_768,N_488,N_524);
and U769 (N_769,N_407,N_505);
nand U770 (N_770,N_593,N_568);
nor U771 (N_771,N_435,N_502);
nor U772 (N_772,N_507,N_588);
or U773 (N_773,N_408,N_426);
nand U774 (N_774,N_404,N_542);
nor U775 (N_775,N_540,N_550);
nand U776 (N_776,N_512,N_481);
or U777 (N_777,N_515,N_462);
or U778 (N_778,N_405,N_492);
nand U779 (N_779,N_429,N_536);
nor U780 (N_780,N_495,N_565);
and U781 (N_781,N_571,N_572);
nand U782 (N_782,N_579,N_553);
or U783 (N_783,N_568,N_534);
and U784 (N_784,N_572,N_565);
nand U785 (N_785,N_488,N_490);
or U786 (N_786,N_505,N_442);
nand U787 (N_787,N_573,N_481);
or U788 (N_788,N_574,N_522);
or U789 (N_789,N_596,N_543);
nor U790 (N_790,N_411,N_566);
nand U791 (N_791,N_596,N_455);
nand U792 (N_792,N_400,N_447);
nor U793 (N_793,N_506,N_457);
and U794 (N_794,N_411,N_539);
nand U795 (N_795,N_537,N_478);
nor U796 (N_796,N_428,N_513);
nor U797 (N_797,N_598,N_590);
and U798 (N_798,N_446,N_424);
or U799 (N_799,N_462,N_572);
nand U800 (N_800,N_727,N_606);
and U801 (N_801,N_797,N_607);
or U802 (N_802,N_616,N_765);
nand U803 (N_803,N_745,N_671);
nand U804 (N_804,N_736,N_624);
nand U805 (N_805,N_785,N_655);
and U806 (N_806,N_631,N_724);
nand U807 (N_807,N_691,N_653);
and U808 (N_808,N_641,N_642);
and U809 (N_809,N_608,N_696);
nand U810 (N_810,N_714,N_749);
nor U811 (N_811,N_798,N_794);
nand U812 (N_812,N_661,N_725);
nand U813 (N_813,N_738,N_726);
or U814 (N_814,N_698,N_778);
nand U815 (N_815,N_796,N_731);
nor U816 (N_816,N_650,N_699);
or U817 (N_817,N_654,N_790);
nand U818 (N_818,N_741,N_649);
nor U819 (N_819,N_625,N_768);
nand U820 (N_820,N_611,N_733);
and U821 (N_821,N_629,N_759);
nand U822 (N_822,N_767,N_603);
and U823 (N_823,N_667,N_651);
nor U824 (N_824,N_619,N_735);
or U825 (N_825,N_648,N_670);
xor U826 (N_826,N_688,N_678);
nand U827 (N_827,N_638,N_780);
and U828 (N_828,N_690,N_763);
nor U829 (N_829,N_739,N_746);
nor U830 (N_830,N_769,N_743);
and U831 (N_831,N_633,N_766);
and U832 (N_832,N_721,N_637);
nor U833 (N_833,N_612,N_636);
and U834 (N_834,N_600,N_709);
nor U835 (N_835,N_789,N_757);
or U836 (N_836,N_728,N_750);
and U837 (N_837,N_604,N_740);
nor U838 (N_838,N_621,N_617);
nor U839 (N_839,N_700,N_626);
nor U840 (N_840,N_723,N_664);
nor U841 (N_841,N_729,N_646);
or U842 (N_842,N_630,N_618);
nor U843 (N_843,N_610,N_602);
and U844 (N_844,N_656,N_627);
nor U845 (N_845,N_640,N_705);
or U846 (N_846,N_628,N_615);
nand U847 (N_847,N_711,N_719);
nand U848 (N_848,N_776,N_752);
nor U849 (N_849,N_793,N_657);
nand U850 (N_850,N_716,N_717);
or U851 (N_851,N_751,N_660);
and U852 (N_852,N_701,N_676);
nand U853 (N_853,N_707,N_737);
and U854 (N_854,N_692,N_792);
nand U855 (N_855,N_687,N_703);
and U856 (N_856,N_704,N_754);
nor U857 (N_857,N_781,N_684);
and U858 (N_858,N_710,N_718);
and U859 (N_859,N_791,N_668);
and U860 (N_860,N_786,N_753);
and U861 (N_861,N_613,N_755);
nand U862 (N_862,N_799,N_635);
and U863 (N_863,N_734,N_695);
and U864 (N_864,N_783,N_715);
nand U865 (N_865,N_669,N_756);
nand U866 (N_866,N_747,N_644);
nor U867 (N_867,N_762,N_777);
xor U868 (N_868,N_720,N_774);
nor U869 (N_869,N_742,N_779);
nor U870 (N_870,N_693,N_744);
nor U871 (N_871,N_677,N_713);
or U872 (N_872,N_680,N_675);
and U873 (N_873,N_748,N_634);
or U874 (N_874,N_758,N_771);
nor U875 (N_875,N_772,N_685);
or U876 (N_876,N_645,N_659);
nor U877 (N_877,N_673,N_694);
xnor U878 (N_878,N_722,N_708);
nand U879 (N_879,N_666,N_601);
nand U880 (N_880,N_620,N_681);
xnor U881 (N_881,N_761,N_605);
nand U882 (N_882,N_672,N_697);
nand U883 (N_883,N_665,N_775);
and U884 (N_884,N_662,N_623);
and U885 (N_885,N_609,N_682);
nand U886 (N_886,N_674,N_622);
or U887 (N_887,N_663,N_760);
or U888 (N_888,N_795,N_706);
nand U889 (N_889,N_712,N_764);
nor U890 (N_890,N_784,N_686);
and U891 (N_891,N_773,N_782);
or U892 (N_892,N_647,N_652);
nor U893 (N_893,N_702,N_632);
or U894 (N_894,N_732,N_643);
and U895 (N_895,N_639,N_683);
nand U896 (N_896,N_788,N_614);
nor U897 (N_897,N_658,N_689);
nor U898 (N_898,N_787,N_730);
nand U899 (N_899,N_679,N_770);
or U900 (N_900,N_747,N_773);
xnor U901 (N_901,N_663,N_688);
nor U902 (N_902,N_779,N_780);
and U903 (N_903,N_788,N_607);
and U904 (N_904,N_775,N_781);
and U905 (N_905,N_648,N_780);
nor U906 (N_906,N_781,N_645);
and U907 (N_907,N_729,N_734);
or U908 (N_908,N_612,N_619);
or U909 (N_909,N_715,N_759);
and U910 (N_910,N_669,N_769);
and U911 (N_911,N_644,N_660);
nor U912 (N_912,N_636,N_754);
nand U913 (N_913,N_637,N_687);
or U914 (N_914,N_789,N_659);
or U915 (N_915,N_713,N_722);
nor U916 (N_916,N_787,N_714);
and U917 (N_917,N_720,N_662);
nor U918 (N_918,N_619,N_626);
or U919 (N_919,N_770,N_601);
nand U920 (N_920,N_639,N_791);
nor U921 (N_921,N_609,N_757);
nand U922 (N_922,N_630,N_743);
nand U923 (N_923,N_799,N_662);
and U924 (N_924,N_656,N_778);
nand U925 (N_925,N_728,N_770);
and U926 (N_926,N_699,N_682);
nand U927 (N_927,N_617,N_663);
or U928 (N_928,N_636,N_708);
nand U929 (N_929,N_681,N_754);
or U930 (N_930,N_620,N_605);
or U931 (N_931,N_760,N_649);
nor U932 (N_932,N_616,N_606);
and U933 (N_933,N_679,N_601);
or U934 (N_934,N_674,N_794);
nand U935 (N_935,N_693,N_758);
or U936 (N_936,N_646,N_668);
nor U937 (N_937,N_719,N_794);
nor U938 (N_938,N_699,N_622);
nand U939 (N_939,N_765,N_737);
nand U940 (N_940,N_759,N_678);
nand U941 (N_941,N_612,N_650);
nand U942 (N_942,N_640,N_758);
and U943 (N_943,N_755,N_703);
or U944 (N_944,N_755,N_692);
or U945 (N_945,N_705,N_651);
nor U946 (N_946,N_725,N_711);
nand U947 (N_947,N_672,N_704);
nor U948 (N_948,N_721,N_624);
or U949 (N_949,N_643,N_742);
nor U950 (N_950,N_682,N_780);
or U951 (N_951,N_727,N_710);
and U952 (N_952,N_796,N_682);
or U953 (N_953,N_770,N_611);
or U954 (N_954,N_680,N_789);
nand U955 (N_955,N_736,N_797);
or U956 (N_956,N_711,N_772);
or U957 (N_957,N_706,N_691);
nor U958 (N_958,N_603,N_739);
nand U959 (N_959,N_750,N_621);
nand U960 (N_960,N_654,N_700);
and U961 (N_961,N_714,N_741);
and U962 (N_962,N_706,N_647);
nor U963 (N_963,N_726,N_635);
or U964 (N_964,N_758,N_700);
or U965 (N_965,N_760,N_720);
nor U966 (N_966,N_620,N_656);
or U967 (N_967,N_769,N_760);
or U968 (N_968,N_730,N_783);
nand U969 (N_969,N_723,N_719);
and U970 (N_970,N_705,N_639);
nor U971 (N_971,N_695,N_662);
or U972 (N_972,N_776,N_714);
or U973 (N_973,N_678,N_764);
nor U974 (N_974,N_722,N_717);
or U975 (N_975,N_776,N_675);
xor U976 (N_976,N_739,N_658);
nand U977 (N_977,N_728,N_793);
xnor U978 (N_978,N_694,N_691);
or U979 (N_979,N_757,N_667);
and U980 (N_980,N_660,N_637);
nor U981 (N_981,N_639,N_770);
nand U982 (N_982,N_654,N_707);
xor U983 (N_983,N_720,N_787);
or U984 (N_984,N_670,N_642);
nor U985 (N_985,N_711,N_710);
or U986 (N_986,N_716,N_605);
and U987 (N_987,N_690,N_721);
xnor U988 (N_988,N_673,N_787);
and U989 (N_989,N_638,N_742);
and U990 (N_990,N_743,N_627);
nand U991 (N_991,N_632,N_726);
and U992 (N_992,N_632,N_756);
and U993 (N_993,N_738,N_768);
nor U994 (N_994,N_634,N_635);
or U995 (N_995,N_661,N_726);
or U996 (N_996,N_653,N_721);
nand U997 (N_997,N_784,N_616);
and U998 (N_998,N_731,N_793);
or U999 (N_999,N_617,N_772);
nor U1000 (N_1000,N_917,N_827);
nand U1001 (N_1001,N_857,N_872);
nand U1002 (N_1002,N_817,N_828);
nand U1003 (N_1003,N_987,N_970);
nand U1004 (N_1004,N_913,N_908);
or U1005 (N_1005,N_883,N_851);
nor U1006 (N_1006,N_999,N_898);
nand U1007 (N_1007,N_818,N_996);
or U1008 (N_1008,N_888,N_859);
nor U1009 (N_1009,N_990,N_920);
and U1010 (N_1010,N_985,N_862);
or U1011 (N_1011,N_816,N_833);
nand U1012 (N_1012,N_809,N_983);
and U1013 (N_1013,N_967,N_834);
or U1014 (N_1014,N_890,N_948);
or U1015 (N_1015,N_936,N_820);
nand U1016 (N_1016,N_986,N_847);
xor U1017 (N_1017,N_854,N_950);
nand U1018 (N_1018,N_853,N_937);
or U1019 (N_1019,N_848,N_994);
and U1020 (N_1020,N_943,N_957);
nand U1021 (N_1021,N_867,N_823);
and U1022 (N_1022,N_988,N_959);
nor U1023 (N_1023,N_866,N_933);
nor U1024 (N_1024,N_964,N_830);
nor U1025 (N_1025,N_947,N_929);
nand U1026 (N_1026,N_870,N_800);
or U1027 (N_1027,N_839,N_856);
nor U1028 (N_1028,N_922,N_811);
and U1029 (N_1029,N_951,N_916);
xnor U1030 (N_1030,N_840,N_865);
nand U1031 (N_1031,N_882,N_829);
nor U1032 (N_1032,N_801,N_984);
nor U1033 (N_1033,N_860,N_930);
or U1034 (N_1034,N_807,N_914);
nand U1035 (N_1035,N_963,N_842);
and U1036 (N_1036,N_978,N_918);
or U1037 (N_1037,N_938,N_819);
and U1038 (N_1038,N_899,N_954);
and U1039 (N_1039,N_923,N_934);
and U1040 (N_1040,N_993,N_926);
or U1041 (N_1041,N_982,N_886);
nor U1042 (N_1042,N_885,N_892);
nor U1043 (N_1043,N_861,N_989);
or U1044 (N_1044,N_941,N_919);
and U1045 (N_1045,N_997,N_911);
and U1046 (N_1046,N_846,N_826);
and U1047 (N_1047,N_924,N_969);
nor U1048 (N_1048,N_932,N_991);
or U1049 (N_1049,N_871,N_884);
and U1050 (N_1050,N_921,N_901);
or U1051 (N_1051,N_852,N_831);
nor U1052 (N_1052,N_965,N_971);
nor U1053 (N_1053,N_975,N_900);
or U1054 (N_1054,N_881,N_887);
and U1055 (N_1055,N_925,N_945);
or U1056 (N_1056,N_972,N_909);
nand U1057 (N_1057,N_906,N_973);
or U1058 (N_1058,N_824,N_927);
and U1059 (N_1059,N_873,N_949);
or U1060 (N_1060,N_974,N_891);
or U1061 (N_1061,N_907,N_814);
or U1062 (N_1062,N_902,N_832);
nand U1063 (N_1063,N_998,N_939);
and U1064 (N_1064,N_981,N_895);
and U1065 (N_1065,N_812,N_992);
or U1066 (N_1066,N_995,N_855);
and U1067 (N_1067,N_944,N_889);
nand U1068 (N_1068,N_880,N_962);
nand U1069 (N_1069,N_835,N_815);
and U1070 (N_1070,N_912,N_928);
and U1071 (N_1071,N_876,N_869);
and U1072 (N_1072,N_813,N_850);
and U1073 (N_1073,N_810,N_875);
or U1074 (N_1074,N_803,N_903);
and U1075 (N_1075,N_879,N_976);
or U1076 (N_1076,N_897,N_877);
nand U1077 (N_1077,N_953,N_825);
and U1078 (N_1078,N_893,N_864);
or U1079 (N_1079,N_806,N_931);
nand U1080 (N_1080,N_837,N_843);
or U1081 (N_1081,N_838,N_946);
or U1082 (N_1082,N_977,N_858);
and U1083 (N_1083,N_878,N_961);
nand U1084 (N_1084,N_956,N_805);
or U1085 (N_1085,N_910,N_966);
or U1086 (N_1086,N_802,N_845);
nand U1087 (N_1087,N_905,N_980);
and U1088 (N_1088,N_942,N_844);
nor U1089 (N_1089,N_822,N_868);
and U1090 (N_1090,N_904,N_863);
nor U1091 (N_1091,N_952,N_960);
and U1092 (N_1092,N_836,N_874);
nand U1093 (N_1093,N_955,N_808);
or U1094 (N_1094,N_935,N_915);
nand U1095 (N_1095,N_958,N_979);
or U1096 (N_1096,N_841,N_896);
or U1097 (N_1097,N_968,N_894);
nor U1098 (N_1098,N_804,N_849);
nand U1099 (N_1099,N_821,N_940);
and U1100 (N_1100,N_925,N_939);
nor U1101 (N_1101,N_923,N_974);
and U1102 (N_1102,N_974,N_961);
and U1103 (N_1103,N_990,N_841);
or U1104 (N_1104,N_962,N_882);
or U1105 (N_1105,N_866,N_905);
xor U1106 (N_1106,N_814,N_980);
and U1107 (N_1107,N_950,N_867);
nor U1108 (N_1108,N_880,N_854);
or U1109 (N_1109,N_881,N_954);
or U1110 (N_1110,N_948,N_961);
and U1111 (N_1111,N_823,N_947);
and U1112 (N_1112,N_950,N_883);
or U1113 (N_1113,N_943,N_885);
nor U1114 (N_1114,N_942,N_947);
and U1115 (N_1115,N_984,N_930);
nor U1116 (N_1116,N_954,N_982);
nor U1117 (N_1117,N_887,N_880);
nand U1118 (N_1118,N_853,N_897);
nor U1119 (N_1119,N_850,N_879);
or U1120 (N_1120,N_999,N_877);
and U1121 (N_1121,N_887,N_828);
nor U1122 (N_1122,N_819,N_884);
or U1123 (N_1123,N_817,N_802);
nand U1124 (N_1124,N_896,N_960);
nor U1125 (N_1125,N_912,N_959);
nor U1126 (N_1126,N_909,N_835);
and U1127 (N_1127,N_918,N_921);
nand U1128 (N_1128,N_813,N_880);
nor U1129 (N_1129,N_939,N_901);
nand U1130 (N_1130,N_915,N_848);
or U1131 (N_1131,N_971,N_827);
nor U1132 (N_1132,N_909,N_943);
or U1133 (N_1133,N_832,N_903);
and U1134 (N_1134,N_984,N_939);
or U1135 (N_1135,N_937,N_941);
nand U1136 (N_1136,N_990,N_994);
and U1137 (N_1137,N_994,N_864);
and U1138 (N_1138,N_901,N_991);
nor U1139 (N_1139,N_894,N_979);
or U1140 (N_1140,N_958,N_954);
nand U1141 (N_1141,N_824,N_880);
and U1142 (N_1142,N_869,N_896);
nor U1143 (N_1143,N_983,N_901);
and U1144 (N_1144,N_924,N_951);
or U1145 (N_1145,N_959,N_800);
nand U1146 (N_1146,N_866,N_895);
and U1147 (N_1147,N_832,N_853);
nand U1148 (N_1148,N_924,N_995);
or U1149 (N_1149,N_929,N_916);
or U1150 (N_1150,N_914,N_886);
or U1151 (N_1151,N_863,N_888);
nor U1152 (N_1152,N_897,N_872);
nand U1153 (N_1153,N_939,N_948);
or U1154 (N_1154,N_917,N_922);
nor U1155 (N_1155,N_866,N_903);
or U1156 (N_1156,N_869,N_847);
xnor U1157 (N_1157,N_956,N_890);
and U1158 (N_1158,N_945,N_938);
and U1159 (N_1159,N_957,N_841);
nor U1160 (N_1160,N_838,N_930);
nor U1161 (N_1161,N_865,N_875);
nor U1162 (N_1162,N_937,N_988);
nand U1163 (N_1163,N_998,N_977);
or U1164 (N_1164,N_905,N_846);
and U1165 (N_1165,N_976,N_980);
and U1166 (N_1166,N_801,N_854);
and U1167 (N_1167,N_902,N_814);
nor U1168 (N_1168,N_981,N_967);
nor U1169 (N_1169,N_972,N_869);
nor U1170 (N_1170,N_874,N_824);
and U1171 (N_1171,N_979,N_880);
nand U1172 (N_1172,N_884,N_904);
and U1173 (N_1173,N_806,N_825);
or U1174 (N_1174,N_912,N_933);
nand U1175 (N_1175,N_826,N_930);
or U1176 (N_1176,N_839,N_925);
nand U1177 (N_1177,N_884,N_988);
or U1178 (N_1178,N_923,N_870);
nand U1179 (N_1179,N_897,N_986);
nor U1180 (N_1180,N_876,N_872);
xnor U1181 (N_1181,N_987,N_920);
or U1182 (N_1182,N_859,N_849);
nor U1183 (N_1183,N_802,N_941);
and U1184 (N_1184,N_883,N_985);
nand U1185 (N_1185,N_891,N_915);
and U1186 (N_1186,N_991,N_813);
or U1187 (N_1187,N_959,N_998);
nand U1188 (N_1188,N_885,N_877);
and U1189 (N_1189,N_904,N_912);
or U1190 (N_1190,N_911,N_919);
nor U1191 (N_1191,N_931,N_964);
and U1192 (N_1192,N_924,N_946);
and U1193 (N_1193,N_854,N_860);
nand U1194 (N_1194,N_923,N_869);
nor U1195 (N_1195,N_828,N_848);
and U1196 (N_1196,N_965,N_907);
and U1197 (N_1197,N_887,N_813);
or U1198 (N_1198,N_948,N_985);
nor U1199 (N_1199,N_828,N_917);
and U1200 (N_1200,N_1158,N_1173);
nand U1201 (N_1201,N_1065,N_1167);
and U1202 (N_1202,N_1141,N_1043);
nand U1203 (N_1203,N_1102,N_1082);
nor U1204 (N_1204,N_1150,N_1094);
nor U1205 (N_1205,N_1067,N_1007);
nand U1206 (N_1206,N_1099,N_1055);
and U1207 (N_1207,N_1077,N_1138);
nor U1208 (N_1208,N_1097,N_1186);
nor U1209 (N_1209,N_1156,N_1103);
nor U1210 (N_1210,N_1198,N_1061);
nor U1211 (N_1211,N_1171,N_1121);
or U1212 (N_1212,N_1075,N_1093);
and U1213 (N_1213,N_1002,N_1071);
and U1214 (N_1214,N_1177,N_1159);
or U1215 (N_1215,N_1100,N_1073);
and U1216 (N_1216,N_1176,N_1136);
and U1217 (N_1217,N_1026,N_1046);
and U1218 (N_1218,N_1196,N_1106);
or U1219 (N_1219,N_1111,N_1142);
nor U1220 (N_1220,N_1057,N_1036);
nor U1221 (N_1221,N_1045,N_1029);
nand U1222 (N_1222,N_1048,N_1020);
and U1223 (N_1223,N_1070,N_1021);
nor U1224 (N_1224,N_1014,N_1072);
nand U1225 (N_1225,N_1139,N_1025);
nor U1226 (N_1226,N_1076,N_1179);
or U1227 (N_1227,N_1080,N_1117);
nor U1228 (N_1228,N_1134,N_1155);
or U1229 (N_1229,N_1010,N_1009);
nor U1230 (N_1230,N_1133,N_1145);
and U1231 (N_1231,N_1088,N_1000);
or U1232 (N_1232,N_1068,N_1022);
nand U1233 (N_1233,N_1189,N_1104);
nand U1234 (N_1234,N_1039,N_1028);
nand U1235 (N_1235,N_1063,N_1113);
or U1236 (N_1236,N_1084,N_1165);
xnor U1237 (N_1237,N_1183,N_1125);
nand U1238 (N_1238,N_1164,N_1116);
or U1239 (N_1239,N_1115,N_1033);
nor U1240 (N_1240,N_1192,N_1149);
nand U1241 (N_1241,N_1105,N_1052);
or U1242 (N_1242,N_1041,N_1053);
or U1243 (N_1243,N_1058,N_1078);
or U1244 (N_1244,N_1144,N_1051);
nor U1245 (N_1245,N_1147,N_1016);
nor U1246 (N_1246,N_1187,N_1098);
or U1247 (N_1247,N_1180,N_1037);
nand U1248 (N_1248,N_1008,N_1013);
or U1249 (N_1249,N_1087,N_1185);
and U1250 (N_1250,N_1095,N_1130);
or U1251 (N_1251,N_1152,N_1003);
nand U1252 (N_1252,N_1027,N_1166);
and U1253 (N_1253,N_1091,N_1127);
nand U1254 (N_1254,N_1066,N_1194);
nand U1255 (N_1255,N_1175,N_1184);
nand U1256 (N_1256,N_1197,N_1131);
nand U1257 (N_1257,N_1132,N_1018);
nor U1258 (N_1258,N_1140,N_1040);
nand U1259 (N_1259,N_1129,N_1015);
and U1260 (N_1260,N_1006,N_1042);
and U1261 (N_1261,N_1109,N_1188);
nand U1262 (N_1262,N_1024,N_1178);
nor U1263 (N_1263,N_1181,N_1162);
nor U1264 (N_1264,N_1054,N_1034);
or U1265 (N_1265,N_1108,N_1135);
and U1266 (N_1266,N_1035,N_1060);
nand U1267 (N_1267,N_1118,N_1182);
and U1268 (N_1268,N_1161,N_1050);
and U1269 (N_1269,N_1112,N_1011);
and U1270 (N_1270,N_1101,N_1032);
and U1271 (N_1271,N_1031,N_1092);
nand U1272 (N_1272,N_1047,N_1086);
and U1273 (N_1273,N_1079,N_1170);
and U1274 (N_1274,N_1089,N_1085);
and U1275 (N_1275,N_1096,N_1004);
nand U1276 (N_1276,N_1012,N_1168);
nor U1277 (N_1277,N_1137,N_1157);
or U1278 (N_1278,N_1191,N_1120);
nand U1279 (N_1279,N_1123,N_1190);
or U1280 (N_1280,N_1146,N_1001);
and U1281 (N_1281,N_1160,N_1172);
nor U1282 (N_1282,N_1154,N_1017);
nand U1283 (N_1283,N_1195,N_1056);
nor U1284 (N_1284,N_1019,N_1038);
and U1285 (N_1285,N_1069,N_1081);
nand U1286 (N_1286,N_1030,N_1174);
nor U1287 (N_1287,N_1044,N_1023);
nor U1288 (N_1288,N_1199,N_1128);
nor U1289 (N_1289,N_1122,N_1062);
nor U1290 (N_1290,N_1153,N_1169);
nor U1291 (N_1291,N_1083,N_1119);
nand U1292 (N_1292,N_1107,N_1059);
and U1293 (N_1293,N_1124,N_1163);
nor U1294 (N_1294,N_1143,N_1005);
nor U1295 (N_1295,N_1064,N_1110);
or U1296 (N_1296,N_1126,N_1090);
and U1297 (N_1297,N_1074,N_1114);
or U1298 (N_1298,N_1193,N_1148);
xnor U1299 (N_1299,N_1049,N_1151);
or U1300 (N_1300,N_1143,N_1090);
and U1301 (N_1301,N_1079,N_1077);
and U1302 (N_1302,N_1183,N_1016);
or U1303 (N_1303,N_1085,N_1040);
nor U1304 (N_1304,N_1092,N_1046);
nand U1305 (N_1305,N_1108,N_1173);
nand U1306 (N_1306,N_1023,N_1188);
xor U1307 (N_1307,N_1116,N_1156);
or U1308 (N_1308,N_1027,N_1065);
nand U1309 (N_1309,N_1055,N_1114);
and U1310 (N_1310,N_1179,N_1137);
and U1311 (N_1311,N_1064,N_1132);
and U1312 (N_1312,N_1055,N_1107);
nand U1313 (N_1313,N_1020,N_1053);
nand U1314 (N_1314,N_1030,N_1143);
and U1315 (N_1315,N_1139,N_1102);
and U1316 (N_1316,N_1103,N_1195);
or U1317 (N_1317,N_1172,N_1009);
nor U1318 (N_1318,N_1138,N_1098);
nor U1319 (N_1319,N_1136,N_1088);
nand U1320 (N_1320,N_1049,N_1051);
nand U1321 (N_1321,N_1110,N_1109);
nand U1322 (N_1322,N_1010,N_1038);
xor U1323 (N_1323,N_1115,N_1062);
nand U1324 (N_1324,N_1101,N_1017);
nand U1325 (N_1325,N_1024,N_1027);
nor U1326 (N_1326,N_1093,N_1034);
and U1327 (N_1327,N_1190,N_1079);
nand U1328 (N_1328,N_1022,N_1188);
nor U1329 (N_1329,N_1187,N_1190);
nand U1330 (N_1330,N_1144,N_1181);
nor U1331 (N_1331,N_1079,N_1013);
nand U1332 (N_1332,N_1138,N_1129);
nor U1333 (N_1333,N_1033,N_1110);
nor U1334 (N_1334,N_1079,N_1148);
nand U1335 (N_1335,N_1141,N_1163);
or U1336 (N_1336,N_1166,N_1045);
and U1337 (N_1337,N_1122,N_1176);
nand U1338 (N_1338,N_1156,N_1081);
and U1339 (N_1339,N_1161,N_1168);
or U1340 (N_1340,N_1130,N_1149);
and U1341 (N_1341,N_1183,N_1126);
nand U1342 (N_1342,N_1168,N_1164);
nand U1343 (N_1343,N_1109,N_1163);
nor U1344 (N_1344,N_1145,N_1070);
or U1345 (N_1345,N_1179,N_1167);
or U1346 (N_1346,N_1156,N_1157);
or U1347 (N_1347,N_1084,N_1020);
nand U1348 (N_1348,N_1087,N_1018);
nor U1349 (N_1349,N_1120,N_1007);
nand U1350 (N_1350,N_1005,N_1054);
nand U1351 (N_1351,N_1075,N_1179);
or U1352 (N_1352,N_1112,N_1195);
nand U1353 (N_1353,N_1080,N_1065);
nand U1354 (N_1354,N_1008,N_1191);
nand U1355 (N_1355,N_1005,N_1077);
or U1356 (N_1356,N_1079,N_1023);
or U1357 (N_1357,N_1057,N_1034);
nand U1358 (N_1358,N_1190,N_1054);
and U1359 (N_1359,N_1065,N_1003);
or U1360 (N_1360,N_1058,N_1174);
nand U1361 (N_1361,N_1007,N_1115);
nand U1362 (N_1362,N_1049,N_1096);
nand U1363 (N_1363,N_1049,N_1025);
nor U1364 (N_1364,N_1120,N_1091);
and U1365 (N_1365,N_1093,N_1066);
and U1366 (N_1366,N_1148,N_1184);
nand U1367 (N_1367,N_1110,N_1138);
and U1368 (N_1368,N_1133,N_1151);
and U1369 (N_1369,N_1031,N_1103);
or U1370 (N_1370,N_1194,N_1010);
nand U1371 (N_1371,N_1020,N_1182);
and U1372 (N_1372,N_1106,N_1011);
nand U1373 (N_1373,N_1186,N_1114);
or U1374 (N_1374,N_1158,N_1097);
or U1375 (N_1375,N_1094,N_1032);
nand U1376 (N_1376,N_1158,N_1014);
nor U1377 (N_1377,N_1147,N_1138);
nand U1378 (N_1378,N_1024,N_1047);
nor U1379 (N_1379,N_1025,N_1140);
xnor U1380 (N_1380,N_1064,N_1094);
nand U1381 (N_1381,N_1026,N_1109);
or U1382 (N_1382,N_1198,N_1085);
nor U1383 (N_1383,N_1157,N_1019);
or U1384 (N_1384,N_1180,N_1029);
and U1385 (N_1385,N_1142,N_1151);
nor U1386 (N_1386,N_1083,N_1056);
nor U1387 (N_1387,N_1016,N_1018);
and U1388 (N_1388,N_1105,N_1098);
nand U1389 (N_1389,N_1189,N_1182);
or U1390 (N_1390,N_1122,N_1054);
xor U1391 (N_1391,N_1019,N_1076);
and U1392 (N_1392,N_1197,N_1148);
nand U1393 (N_1393,N_1184,N_1112);
nor U1394 (N_1394,N_1003,N_1198);
and U1395 (N_1395,N_1075,N_1146);
or U1396 (N_1396,N_1176,N_1027);
or U1397 (N_1397,N_1065,N_1047);
or U1398 (N_1398,N_1069,N_1115);
nor U1399 (N_1399,N_1067,N_1170);
xnor U1400 (N_1400,N_1310,N_1312);
nor U1401 (N_1401,N_1382,N_1252);
nor U1402 (N_1402,N_1320,N_1271);
or U1403 (N_1403,N_1203,N_1226);
nand U1404 (N_1404,N_1332,N_1327);
nand U1405 (N_1405,N_1379,N_1250);
and U1406 (N_1406,N_1251,N_1354);
or U1407 (N_1407,N_1297,N_1227);
nand U1408 (N_1408,N_1342,N_1334);
nand U1409 (N_1409,N_1344,N_1374);
and U1410 (N_1410,N_1290,N_1266);
or U1411 (N_1411,N_1211,N_1348);
or U1412 (N_1412,N_1204,N_1302);
or U1413 (N_1413,N_1336,N_1207);
nand U1414 (N_1414,N_1304,N_1277);
nor U1415 (N_1415,N_1247,N_1341);
nand U1416 (N_1416,N_1284,N_1347);
nand U1417 (N_1417,N_1373,N_1324);
nand U1418 (N_1418,N_1392,N_1202);
nand U1419 (N_1419,N_1280,N_1352);
nand U1420 (N_1420,N_1268,N_1291);
nand U1421 (N_1421,N_1386,N_1258);
nor U1422 (N_1422,N_1300,N_1314);
nor U1423 (N_1423,N_1267,N_1274);
nor U1424 (N_1424,N_1323,N_1316);
nand U1425 (N_1425,N_1393,N_1303);
or U1426 (N_1426,N_1225,N_1276);
nor U1427 (N_1427,N_1398,N_1216);
or U1428 (N_1428,N_1322,N_1235);
or U1429 (N_1429,N_1285,N_1208);
nand U1430 (N_1430,N_1261,N_1333);
or U1431 (N_1431,N_1306,N_1218);
and U1432 (N_1432,N_1358,N_1381);
nor U1433 (N_1433,N_1318,N_1237);
nor U1434 (N_1434,N_1248,N_1321);
and U1435 (N_1435,N_1395,N_1330);
and U1436 (N_1436,N_1307,N_1234);
nor U1437 (N_1437,N_1338,N_1372);
nor U1438 (N_1438,N_1396,N_1308);
nor U1439 (N_1439,N_1223,N_1366);
and U1440 (N_1440,N_1388,N_1328);
or U1441 (N_1441,N_1289,N_1368);
nor U1442 (N_1442,N_1313,N_1294);
and U1443 (N_1443,N_1287,N_1356);
or U1444 (N_1444,N_1353,N_1259);
or U1445 (N_1445,N_1305,N_1273);
and U1446 (N_1446,N_1229,N_1299);
nor U1447 (N_1447,N_1351,N_1309);
nor U1448 (N_1448,N_1377,N_1263);
nor U1449 (N_1449,N_1212,N_1293);
or U1450 (N_1450,N_1265,N_1275);
nor U1451 (N_1451,N_1205,N_1298);
nand U1452 (N_1452,N_1397,N_1239);
or U1453 (N_1453,N_1384,N_1385);
nand U1454 (N_1454,N_1375,N_1253);
nor U1455 (N_1455,N_1362,N_1325);
and U1456 (N_1456,N_1249,N_1264);
nor U1457 (N_1457,N_1399,N_1278);
and U1458 (N_1458,N_1210,N_1295);
and U1459 (N_1459,N_1340,N_1331);
and U1460 (N_1460,N_1260,N_1296);
nor U1461 (N_1461,N_1364,N_1245);
nand U1462 (N_1462,N_1389,N_1383);
nor U1463 (N_1463,N_1359,N_1254);
nor U1464 (N_1464,N_1288,N_1357);
nor U1465 (N_1465,N_1241,N_1209);
or U1466 (N_1466,N_1232,N_1215);
nor U1467 (N_1467,N_1228,N_1349);
or U1468 (N_1468,N_1346,N_1390);
nand U1469 (N_1469,N_1282,N_1391);
and U1470 (N_1470,N_1363,N_1339);
and U1471 (N_1471,N_1286,N_1329);
and U1472 (N_1472,N_1345,N_1236);
nand U1473 (N_1473,N_1230,N_1311);
nor U1474 (N_1474,N_1380,N_1335);
nor U1475 (N_1475,N_1240,N_1370);
nor U1476 (N_1476,N_1238,N_1256);
and U1477 (N_1477,N_1262,N_1326);
nor U1478 (N_1478,N_1292,N_1213);
nand U1479 (N_1479,N_1217,N_1233);
nor U1480 (N_1480,N_1371,N_1343);
or U1481 (N_1481,N_1337,N_1387);
nor U1482 (N_1482,N_1224,N_1361);
nor U1483 (N_1483,N_1317,N_1270);
nand U1484 (N_1484,N_1257,N_1201);
and U1485 (N_1485,N_1242,N_1367);
nor U1486 (N_1486,N_1219,N_1376);
nand U1487 (N_1487,N_1231,N_1315);
nand U1488 (N_1488,N_1360,N_1206);
or U1489 (N_1489,N_1246,N_1365);
or U1490 (N_1490,N_1244,N_1355);
or U1491 (N_1491,N_1222,N_1255);
nand U1492 (N_1492,N_1394,N_1281);
or U1493 (N_1493,N_1283,N_1279);
and U1494 (N_1494,N_1269,N_1221);
or U1495 (N_1495,N_1220,N_1243);
and U1496 (N_1496,N_1319,N_1378);
nand U1497 (N_1497,N_1301,N_1272);
nor U1498 (N_1498,N_1214,N_1200);
nor U1499 (N_1499,N_1369,N_1350);
or U1500 (N_1500,N_1225,N_1376);
and U1501 (N_1501,N_1399,N_1285);
nor U1502 (N_1502,N_1295,N_1270);
nand U1503 (N_1503,N_1348,N_1215);
or U1504 (N_1504,N_1208,N_1216);
and U1505 (N_1505,N_1229,N_1230);
and U1506 (N_1506,N_1391,N_1302);
nor U1507 (N_1507,N_1377,N_1321);
xor U1508 (N_1508,N_1358,N_1293);
and U1509 (N_1509,N_1368,N_1349);
nand U1510 (N_1510,N_1347,N_1239);
and U1511 (N_1511,N_1337,N_1350);
nand U1512 (N_1512,N_1300,N_1240);
nor U1513 (N_1513,N_1384,N_1312);
or U1514 (N_1514,N_1387,N_1278);
nor U1515 (N_1515,N_1385,N_1336);
nor U1516 (N_1516,N_1256,N_1385);
nor U1517 (N_1517,N_1271,N_1290);
and U1518 (N_1518,N_1286,N_1269);
nor U1519 (N_1519,N_1334,N_1350);
nor U1520 (N_1520,N_1214,N_1267);
nor U1521 (N_1521,N_1333,N_1215);
or U1522 (N_1522,N_1270,N_1287);
and U1523 (N_1523,N_1363,N_1331);
nand U1524 (N_1524,N_1202,N_1319);
or U1525 (N_1525,N_1312,N_1246);
nor U1526 (N_1526,N_1384,N_1329);
nor U1527 (N_1527,N_1307,N_1396);
and U1528 (N_1528,N_1324,N_1260);
nor U1529 (N_1529,N_1336,N_1396);
and U1530 (N_1530,N_1379,N_1238);
nand U1531 (N_1531,N_1334,N_1277);
or U1532 (N_1532,N_1258,N_1202);
or U1533 (N_1533,N_1256,N_1320);
or U1534 (N_1534,N_1353,N_1298);
nor U1535 (N_1535,N_1386,N_1330);
nand U1536 (N_1536,N_1365,N_1366);
and U1537 (N_1537,N_1342,N_1351);
or U1538 (N_1538,N_1255,N_1350);
nand U1539 (N_1539,N_1275,N_1358);
and U1540 (N_1540,N_1293,N_1310);
and U1541 (N_1541,N_1368,N_1231);
or U1542 (N_1542,N_1266,N_1297);
and U1543 (N_1543,N_1240,N_1267);
nand U1544 (N_1544,N_1388,N_1209);
nor U1545 (N_1545,N_1353,N_1380);
nor U1546 (N_1546,N_1287,N_1228);
nor U1547 (N_1547,N_1270,N_1251);
nor U1548 (N_1548,N_1301,N_1321);
nor U1549 (N_1549,N_1387,N_1297);
or U1550 (N_1550,N_1298,N_1237);
nor U1551 (N_1551,N_1220,N_1326);
nor U1552 (N_1552,N_1299,N_1218);
nor U1553 (N_1553,N_1234,N_1336);
or U1554 (N_1554,N_1209,N_1353);
nand U1555 (N_1555,N_1277,N_1273);
nor U1556 (N_1556,N_1344,N_1207);
and U1557 (N_1557,N_1355,N_1328);
and U1558 (N_1558,N_1278,N_1252);
nand U1559 (N_1559,N_1328,N_1255);
and U1560 (N_1560,N_1296,N_1321);
nor U1561 (N_1561,N_1202,N_1211);
and U1562 (N_1562,N_1280,N_1291);
and U1563 (N_1563,N_1304,N_1274);
and U1564 (N_1564,N_1237,N_1379);
and U1565 (N_1565,N_1202,N_1346);
or U1566 (N_1566,N_1211,N_1336);
nor U1567 (N_1567,N_1259,N_1267);
or U1568 (N_1568,N_1258,N_1382);
nor U1569 (N_1569,N_1393,N_1235);
xor U1570 (N_1570,N_1396,N_1248);
or U1571 (N_1571,N_1371,N_1312);
nor U1572 (N_1572,N_1370,N_1211);
and U1573 (N_1573,N_1235,N_1215);
nand U1574 (N_1574,N_1327,N_1270);
nand U1575 (N_1575,N_1256,N_1390);
nand U1576 (N_1576,N_1207,N_1282);
nand U1577 (N_1577,N_1290,N_1312);
and U1578 (N_1578,N_1358,N_1235);
nand U1579 (N_1579,N_1379,N_1281);
nor U1580 (N_1580,N_1267,N_1224);
and U1581 (N_1581,N_1224,N_1360);
nand U1582 (N_1582,N_1269,N_1285);
nand U1583 (N_1583,N_1297,N_1276);
or U1584 (N_1584,N_1382,N_1225);
nand U1585 (N_1585,N_1336,N_1283);
and U1586 (N_1586,N_1332,N_1248);
nand U1587 (N_1587,N_1305,N_1369);
nand U1588 (N_1588,N_1321,N_1365);
and U1589 (N_1589,N_1235,N_1356);
or U1590 (N_1590,N_1266,N_1216);
nor U1591 (N_1591,N_1315,N_1233);
nor U1592 (N_1592,N_1205,N_1387);
or U1593 (N_1593,N_1363,N_1216);
or U1594 (N_1594,N_1243,N_1278);
nor U1595 (N_1595,N_1345,N_1220);
or U1596 (N_1596,N_1234,N_1285);
and U1597 (N_1597,N_1335,N_1222);
xnor U1598 (N_1598,N_1298,N_1286);
or U1599 (N_1599,N_1355,N_1346);
xnor U1600 (N_1600,N_1595,N_1439);
nand U1601 (N_1601,N_1487,N_1545);
nand U1602 (N_1602,N_1430,N_1412);
and U1603 (N_1603,N_1565,N_1551);
nand U1604 (N_1604,N_1494,N_1592);
nor U1605 (N_1605,N_1593,N_1527);
and U1606 (N_1606,N_1578,N_1549);
and U1607 (N_1607,N_1400,N_1423);
nand U1608 (N_1608,N_1402,N_1510);
and U1609 (N_1609,N_1480,N_1552);
and U1610 (N_1610,N_1415,N_1457);
nor U1611 (N_1611,N_1484,N_1591);
and U1612 (N_1612,N_1512,N_1424);
nand U1613 (N_1613,N_1467,N_1564);
and U1614 (N_1614,N_1479,N_1517);
and U1615 (N_1615,N_1449,N_1535);
nand U1616 (N_1616,N_1472,N_1525);
nand U1617 (N_1617,N_1529,N_1590);
nand U1618 (N_1618,N_1505,N_1406);
nand U1619 (N_1619,N_1405,N_1440);
or U1620 (N_1620,N_1532,N_1417);
nand U1621 (N_1621,N_1500,N_1456);
or U1622 (N_1622,N_1498,N_1434);
nand U1623 (N_1623,N_1420,N_1550);
nand U1624 (N_1624,N_1488,N_1594);
or U1625 (N_1625,N_1534,N_1579);
and U1626 (N_1626,N_1432,N_1503);
nor U1627 (N_1627,N_1443,N_1451);
nor U1628 (N_1628,N_1530,N_1486);
or U1629 (N_1629,N_1458,N_1422);
and U1630 (N_1630,N_1459,N_1468);
and U1631 (N_1631,N_1514,N_1460);
or U1632 (N_1632,N_1522,N_1463);
nand U1633 (N_1633,N_1543,N_1576);
and U1634 (N_1634,N_1419,N_1533);
nor U1635 (N_1635,N_1448,N_1548);
and U1636 (N_1636,N_1560,N_1582);
nand U1637 (N_1637,N_1569,N_1556);
and U1638 (N_1638,N_1520,N_1597);
nand U1639 (N_1639,N_1499,N_1554);
nor U1640 (N_1640,N_1539,N_1567);
nand U1641 (N_1641,N_1476,N_1513);
nor U1642 (N_1642,N_1586,N_1544);
nand U1643 (N_1643,N_1573,N_1584);
or U1644 (N_1644,N_1446,N_1497);
xor U1645 (N_1645,N_1435,N_1566);
nor U1646 (N_1646,N_1453,N_1465);
nand U1647 (N_1647,N_1438,N_1414);
and U1648 (N_1648,N_1425,N_1466);
nor U1649 (N_1649,N_1496,N_1477);
or U1650 (N_1650,N_1429,N_1538);
and U1651 (N_1651,N_1507,N_1495);
and U1652 (N_1652,N_1416,N_1485);
or U1653 (N_1653,N_1492,N_1516);
nor U1654 (N_1654,N_1403,N_1431);
nor U1655 (N_1655,N_1561,N_1559);
or U1656 (N_1656,N_1427,N_1553);
or U1657 (N_1657,N_1445,N_1475);
and U1658 (N_1658,N_1518,N_1599);
or U1659 (N_1659,N_1464,N_1511);
nand U1660 (N_1660,N_1469,N_1574);
nor U1661 (N_1661,N_1509,N_1501);
or U1662 (N_1662,N_1404,N_1504);
nand U1663 (N_1663,N_1409,N_1461);
nand U1664 (N_1664,N_1428,N_1437);
nand U1665 (N_1665,N_1452,N_1542);
nor U1666 (N_1666,N_1555,N_1583);
and U1667 (N_1667,N_1455,N_1562);
and U1668 (N_1668,N_1490,N_1471);
or U1669 (N_1669,N_1568,N_1557);
and U1670 (N_1670,N_1478,N_1519);
nand U1671 (N_1671,N_1521,N_1589);
nand U1672 (N_1672,N_1407,N_1540);
nor U1673 (N_1673,N_1444,N_1441);
nand U1674 (N_1674,N_1536,N_1526);
nor U1675 (N_1675,N_1411,N_1483);
and U1676 (N_1676,N_1524,N_1418);
nand U1677 (N_1677,N_1587,N_1426);
and U1678 (N_1678,N_1546,N_1491);
nand U1679 (N_1679,N_1489,N_1572);
nand U1680 (N_1680,N_1577,N_1581);
nand U1681 (N_1681,N_1528,N_1481);
nand U1682 (N_1682,N_1588,N_1473);
or U1683 (N_1683,N_1433,N_1541);
nor U1684 (N_1684,N_1408,N_1570);
or U1685 (N_1685,N_1450,N_1563);
and U1686 (N_1686,N_1580,N_1474);
nor U1687 (N_1687,N_1531,N_1454);
and U1688 (N_1688,N_1502,N_1462);
nor U1689 (N_1689,N_1447,N_1571);
or U1690 (N_1690,N_1558,N_1413);
and U1691 (N_1691,N_1506,N_1547);
or U1692 (N_1692,N_1508,N_1598);
nor U1693 (N_1693,N_1410,N_1575);
and U1694 (N_1694,N_1482,N_1470);
nor U1695 (N_1695,N_1515,N_1585);
nand U1696 (N_1696,N_1523,N_1421);
nor U1697 (N_1697,N_1442,N_1596);
or U1698 (N_1698,N_1537,N_1401);
nor U1699 (N_1699,N_1493,N_1436);
and U1700 (N_1700,N_1408,N_1458);
and U1701 (N_1701,N_1582,N_1555);
or U1702 (N_1702,N_1528,N_1431);
or U1703 (N_1703,N_1434,N_1420);
and U1704 (N_1704,N_1502,N_1582);
nand U1705 (N_1705,N_1442,N_1563);
and U1706 (N_1706,N_1540,N_1487);
or U1707 (N_1707,N_1490,N_1548);
nand U1708 (N_1708,N_1596,N_1551);
or U1709 (N_1709,N_1547,N_1562);
nand U1710 (N_1710,N_1536,N_1489);
nor U1711 (N_1711,N_1557,N_1419);
and U1712 (N_1712,N_1403,N_1548);
or U1713 (N_1713,N_1591,N_1570);
nor U1714 (N_1714,N_1403,N_1450);
or U1715 (N_1715,N_1583,N_1438);
and U1716 (N_1716,N_1573,N_1582);
nor U1717 (N_1717,N_1597,N_1556);
nor U1718 (N_1718,N_1569,N_1543);
nor U1719 (N_1719,N_1425,N_1499);
and U1720 (N_1720,N_1596,N_1513);
or U1721 (N_1721,N_1488,N_1554);
and U1722 (N_1722,N_1515,N_1441);
or U1723 (N_1723,N_1474,N_1509);
nor U1724 (N_1724,N_1527,N_1569);
or U1725 (N_1725,N_1417,N_1436);
nor U1726 (N_1726,N_1567,N_1553);
and U1727 (N_1727,N_1420,N_1567);
or U1728 (N_1728,N_1458,N_1503);
or U1729 (N_1729,N_1425,N_1463);
nand U1730 (N_1730,N_1409,N_1468);
nand U1731 (N_1731,N_1503,N_1552);
or U1732 (N_1732,N_1532,N_1412);
or U1733 (N_1733,N_1556,N_1560);
or U1734 (N_1734,N_1580,N_1565);
and U1735 (N_1735,N_1436,N_1527);
or U1736 (N_1736,N_1515,N_1543);
nor U1737 (N_1737,N_1567,N_1467);
or U1738 (N_1738,N_1549,N_1431);
nand U1739 (N_1739,N_1542,N_1514);
and U1740 (N_1740,N_1490,N_1426);
nor U1741 (N_1741,N_1538,N_1482);
nor U1742 (N_1742,N_1543,N_1518);
nor U1743 (N_1743,N_1547,N_1453);
nand U1744 (N_1744,N_1466,N_1441);
and U1745 (N_1745,N_1599,N_1441);
nor U1746 (N_1746,N_1451,N_1516);
or U1747 (N_1747,N_1488,N_1528);
nor U1748 (N_1748,N_1566,N_1512);
nand U1749 (N_1749,N_1590,N_1478);
nor U1750 (N_1750,N_1564,N_1589);
nor U1751 (N_1751,N_1465,N_1595);
and U1752 (N_1752,N_1469,N_1549);
nand U1753 (N_1753,N_1563,N_1499);
nand U1754 (N_1754,N_1547,N_1479);
nand U1755 (N_1755,N_1430,N_1441);
nor U1756 (N_1756,N_1411,N_1482);
and U1757 (N_1757,N_1518,N_1481);
nand U1758 (N_1758,N_1589,N_1501);
or U1759 (N_1759,N_1474,N_1414);
or U1760 (N_1760,N_1576,N_1527);
nand U1761 (N_1761,N_1580,N_1502);
nor U1762 (N_1762,N_1463,N_1547);
nor U1763 (N_1763,N_1410,N_1586);
and U1764 (N_1764,N_1554,N_1489);
nand U1765 (N_1765,N_1436,N_1447);
and U1766 (N_1766,N_1594,N_1453);
nor U1767 (N_1767,N_1517,N_1551);
nor U1768 (N_1768,N_1402,N_1555);
and U1769 (N_1769,N_1580,N_1528);
and U1770 (N_1770,N_1447,N_1408);
nand U1771 (N_1771,N_1528,N_1524);
or U1772 (N_1772,N_1462,N_1534);
xnor U1773 (N_1773,N_1594,N_1483);
nand U1774 (N_1774,N_1567,N_1548);
or U1775 (N_1775,N_1457,N_1493);
or U1776 (N_1776,N_1434,N_1541);
and U1777 (N_1777,N_1549,N_1507);
or U1778 (N_1778,N_1507,N_1470);
nor U1779 (N_1779,N_1468,N_1423);
and U1780 (N_1780,N_1479,N_1485);
or U1781 (N_1781,N_1408,N_1479);
nand U1782 (N_1782,N_1539,N_1591);
nor U1783 (N_1783,N_1473,N_1464);
nor U1784 (N_1784,N_1467,N_1474);
nor U1785 (N_1785,N_1563,N_1545);
nand U1786 (N_1786,N_1521,N_1448);
and U1787 (N_1787,N_1473,N_1543);
nand U1788 (N_1788,N_1522,N_1598);
nor U1789 (N_1789,N_1543,N_1544);
and U1790 (N_1790,N_1546,N_1542);
nor U1791 (N_1791,N_1463,N_1493);
and U1792 (N_1792,N_1541,N_1461);
nor U1793 (N_1793,N_1461,N_1497);
or U1794 (N_1794,N_1514,N_1506);
nor U1795 (N_1795,N_1598,N_1529);
nand U1796 (N_1796,N_1452,N_1524);
nor U1797 (N_1797,N_1459,N_1567);
nor U1798 (N_1798,N_1458,N_1514);
nor U1799 (N_1799,N_1572,N_1528);
nand U1800 (N_1800,N_1710,N_1636);
nand U1801 (N_1801,N_1660,N_1784);
nand U1802 (N_1802,N_1733,N_1709);
or U1803 (N_1803,N_1721,N_1681);
nor U1804 (N_1804,N_1651,N_1705);
nand U1805 (N_1805,N_1747,N_1672);
and U1806 (N_1806,N_1758,N_1675);
and U1807 (N_1807,N_1745,N_1754);
and U1808 (N_1808,N_1700,N_1623);
or U1809 (N_1809,N_1771,N_1735);
and U1810 (N_1810,N_1634,N_1650);
or U1811 (N_1811,N_1673,N_1679);
nand U1812 (N_1812,N_1618,N_1755);
or U1813 (N_1813,N_1770,N_1738);
or U1814 (N_1814,N_1702,N_1730);
nand U1815 (N_1815,N_1637,N_1706);
nor U1816 (N_1816,N_1604,N_1778);
nor U1817 (N_1817,N_1787,N_1704);
nor U1818 (N_1818,N_1646,N_1612);
or U1819 (N_1819,N_1764,N_1707);
nor U1820 (N_1820,N_1668,N_1657);
or U1821 (N_1821,N_1677,N_1666);
or U1822 (N_1822,N_1688,N_1664);
and U1823 (N_1823,N_1712,N_1765);
nand U1824 (N_1824,N_1614,N_1797);
and U1825 (N_1825,N_1615,N_1678);
and U1826 (N_1826,N_1772,N_1686);
or U1827 (N_1827,N_1661,N_1719);
and U1828 (N_1828,N_1619,N_1725);
xnor U1829 (N_1829,N_1760,N_1785);
nor U1830 (N_1830,N_1741,N_1625);
nor U1831 (N_1831,N_1740,N_1622);
and U1832 (N_1832,N_1663,N_1626);
and U1833 (N_1833,N_1689,N_1790);
nand U1834 (N_1834,N_1602,N_1701);
or U1835 (N_1835,N_1699,N_1682);
nand U1836 (N_1836,N_1611,N_1749);
nand U1837 (N_1837,N_1684,N_1696);
and U1838 (N_1838,N_1671,N_1766);
nand U1839 (N_1839,N_1609,N_1676);
and U1840 (N_1840,N_1674,N_1685);
nor U1841 (N_1841,N_1703,N_1690);
or U1842 (N_1842,N_1748,N_1723);
nand U1843 (N_1843,N_1786,N_1670);
and U1844 (N_1844,N_1794,N_1714);
nor U1845 (N_1845,N_1742,N_1662);
or U1846 (N_1846,N_1621,N_1759);
or U1847 (N_1847,N_1796,N_1647);
nand U1848 (N_1848,N_1694,N_1736);
nand U1849 (N_1849,N_1642,N_1716);
and U1850 (N_1850,N_1708,N_1720);
and U1851 (N_1851,N_1627,N_1781);
or U1852 (N_1852,N_1680,N_1630);
nor U1853 (N_1853,N_1620,N_1613);
and U1854 (N_1854,N_1669,N_1629);
nor U1855 (N_1855,N_1783,N_1665);
nor U1856 (N_1856,N_1792,N_1722);
or U1857 (N_1857,N_1791,N_1632);
or U1858 (N_1858,N_1649,N_1610);
nor U1859 (N_1859,N_1658,N_1753);
nand U1860 (N_1860,N_1644,N_1628);
nor U1861 (N_1861,N_1732,N_1752);
or U1862 (N_1862,N_1667,N_1774);
nor U1863 (N_1863,N_1683,N_1737);
nor U1864 (N_1864,N_1743,N_1635);
or U1865 (N_1865,N_1640,N_1633);
and U1866 (N_1866,N_1711,N_1643);
xnor U1867 (N_1867,N_1779,N_1695);
or U1868 (N_1868,N_1645,N_1653);
or U1869 (N_1869,N_1655,N_1769);
nand U1870 (N_1870,N_1789,N_1698);
nand U1871 (N_1871,N_1601,N_1780);
and U1872 (N_1872,N_1729,N_1756);
nand U1873 (N_1873,N_1746,N_1693);
nor U1874 (N_1874,N_1691,N_1603);
or U1875 (N_1875,N_1798,N_1793);
nand U1876 (N_1876,N_1762,N_1788);
nor U1877 (N_1877,N_1731,N_1638);
and U1878 (N_1878,N_1795,N_1654);
or U1879 (N_1879,N_1751,N_1608);
nor U1880 (N_1880,N_1606,N_1777);
or U1881 (N_1881,N_1724,N_1631);
nand U1882 (N_1882,N_1734,N_1775);
and U1883 (N_1883,N_1768,N_1761);
and U1884 (N_1884,N_1744,N_1659);
or U1885 (N_1885,N_1728,N_1692);
nor U1886 (N_1886,N_1641,N_1648);
nand U1887 (N_1887,N_1750,N_1652);
nand U1888 (N_1888,N_1617,N_1718);
and U1889 (N_1889,N_1607,N_1799);
and U1890 (N_1890,N_1624,N_1605);
or U1891 (N_1891,N_1616,N_1782);
or U1892 (N_1892,N_1713,N_1656);
nor U1893 (N_1893,N_1739,N_1763);
or U1894 (N_1894,N_1727,N_1717);
and U1895 (N_1895,N_1776,N_1687);
or U1896 (N_1896,N_1767,N_1726);
nand U1897 (N_1897,N_1639,N_1757);
nor U1898 (N_1898,N_1773,N_1715);
nand U1899 (N_1899,N_1600,N_1697);
or U1900 (N_1900,N_1726,N_1755);
and U1901 (N_1901,N_1795,N_1613);
nor U1902 (N_1902,N_1614,N_1740);
nor U1903 (N_1903,N_1798,N_1656);
nor U1904 (N_1904,N_1730,N_1765);
nand U1905 (N_1905,N_1752,N_1790);
or U1906 (N_1906,N_1732,N_1670);
nand U1907 (N_1907,N_1744,N_1729);
and U1908 (N_1908,N_1692,N_1705);
nor U1909 (N_1909,N_1758,N_1678);
nor U1910 (N_1910,N_1797,N_1759);
nand U1911 (N_1911,N_1745,N_1744);
and U1912 (N_1912,N_1692,N_1612);
nand U1913 (N_1913,N_1685,N_1663);
or U1914 (N_1914,N_1692,N_1690);
nor U1915 (N_1915,N_1733,N_1797);
nand U1916 (N_1916,N_1762,N_1748);
or U1917 (N_1917,N_1617,N_1736);
nor U1918 (N_1918,N_1619,N_1674);
and U1919 (N_1919,N_1683,N_1779);
nand U1920 (N_1920,N_1610,N_1670);
or U1921 (N_1921,N_1769,N_1762);
or U1922 (N_1922,N_1757,N_1673);
or U1923 (N_1923,N_1757,N_1658);
or U1924 (N_1924,N_1740,N_1653);
nand U1925 (N_1925,N_1688,N_1756);
nor U1926 (N_1926,N_1731,N_1672);
nand U1927 (N_1927,N_1600,N_1741);
or U1928 (N_1928,N_1791,N_1794);
and U1929 (N_1929,N_1773,N_1726);
and U1930 (N_1930,N_1774,N_1704);
nand U1931 (N_1931,N_1777,N_1771);
nor U1932 (N_1932,N_1652,N_1636);
nand U1933 (N_1933,N_1771,N_1631);
and U1934 (N_1934,N_1759,N_1747);
nand U1935 (N_1935,N_1623,N_1629);
nor U1936 (N_1936,N_1729,N_1703);
nor U1937 (N_1937,N_1702,N_1716);
nand U1938 (N_1938,N_1611,N_1776);
nand U1939 (N_1939,N_1661,N_1646);
and U1940 (N_1940,N_1701,N_1601);
nand U1941 (N_1941,N_1735,N_1665);
nand U1942 (N_1942,N_1629,N_1634);
and U1943 (N_1943,N_1752,N_1741);
and U1944 (N_1944,N_1773,N_1643);
and U1945 (N_1945,N_1687,N_1725);
and U1946 (N_1946,N_1754,N_1664);
or U1947 (N_1947,N_1740,N_1746);
nor U1948 (N_1948,N_1664,N_1641);
nand U1949 (N_1949,N_1644,N_1780);
or U1950 (N_1950,N_1700,N_1770);
or U1951 (N_1951,N_1721,N_1770);
or U1952 (N_1952,N_1769,N_1657);
nor U1953 (N_1953,N_1644,N_1716);
or U1954 (N_1954,N_1746,N_1633);
xnor U1955 (N_1955,N_1677,N_1634);
nor U1956 (N_1956,N_1774,N_1770);
or U1957 (N_1957,N_1761,N_1783);
nand U1958 (N_1958,N_1766,N_1726);
nor U1959 (N_1959,N_1798,N_1695);
nand U1960 (N_1960,N_1647,N_1780);
or U1961 (N_1961,N_1722,N_1777);
and U1962 (N_1962,N_1652,N_1775);
and U1963 (N_1963,N_1707,N_1775);
nor U1964 (N_1964,N_1671,N_1651);
or U1965 (N_1965,N_1795,N_1614);
nand U1966 (N_1966,N_1602,N_1694);
and U1967 (N_1967,N_1616,N_1798);
nand U1968 (N_1968,N_1604,N_1637);
or U1969 (N_1969,N_1747,N_1727);
nand U1970 (N_1970,N_1621,N_1723);
and U1971 (N_1971,N_1645,N_1689);
nor U1972 (N_1972,N_1612,N_1606);
nor U1973 (N_1973,N_1717,N_1791);
xnor U1974 (N_1974,N_1750,N_1738);
nand U1975 (N_1975,N_1605,N_1636);
and U1976 (N_1976,N_1693,N_1642);
or U1977 (N_1977,N_1753,N_1709);
nand U1978 (N_1978,N_1747,N_1790);
or U1979 (N_1979,N_1756,N_1733);
nor U1980 (N_1980,N_1612,N_1697);
nor U1981 (N_1981,N_1792,N_1621);
or U1982 (N_1982,N_1657,N_1778);
or U1983 (N_1983,N_1732,N_1617);
nor U1984 (N_1984,N_1775,N_1638);
nand U1985 (N_1985,N_1764,N_1636);
nor U1986 (N_1986,N_1607,N_1684);
or U1987 (N_1987,N_1782,N_1792);
or U1988 (N_1988,N_1740,N_1780);
nand U1989 (N_1989,N_1764,N_1738);
and U1990 (N_1990,N_1702,N_1711);
or U1991 (N_1991,N_1617,N_1637);
and U1992 (N_1992,N_1789,N_1685);
nor U1993 (N_1993,N_1795,N_1737);
nor U1994 (N_1994,N_1649,N_1781);
nand U1995 (N_1995,N_1785,N_1618);
nor U1996 (N_1996,N_1647,N_1746);
and U1997 (N_1997,N_1707,N_1625);
nor U1998 (N_1998,N_1685,N_1600);
nor U1999 (N_1999,N_1649,N_1618);
or U2000 (N_2000,N_1970,N_1889);
and U2001 (N_2001,N_1823,N_1953);
and U2002 (N_2002,N_1902,N_1838);
nand U2003 (N_2003,N_1991,N_1843);
nor U2004 (N_2004,N_1972,N_1956);
or U2005 (N_2005,N_1811,N_1816);
nor U2006 (N_2006,N_1813,N_1982);
or U2007 (N_2007,N_1895,N_1867);
and U2008 (N_2008,N_1948,N_1877);
or U2009 (N_2009,N_1942,N_1806);
nor U2010 (N_2010,N_1907,N_1818);
nand U2011 (N_2011,N_1883,N_1820);
nand U2012 (N_2012,N_1801,N_1891);
xnor U2013 (N_2013,N_1910,N_1926);
nand U2014 (N_2014,N_1934,N_1861);
nor U2015 (N_2015,N_1921,N_1832);
nand U2016 (N_2016,N_1914,N_1929);
or U2017 (N_2017,N_1957,N_1947);
and U2018 (N_2018,N_1879,N_1866);
nor U2019 (N_2019,N_1880,N_1938);
nand U2020 (N_2020,N_1872,N_1846);
or U2021 (N_2021,N_1939,N_1984);
and U2022 (N_2022,N_1807,N_1884);
and U2023 (N_2023,N_1988,N_1821);
or U2024 (N_2024,N_1836,N_1903);
and U2025 (N_2025,N_1845,N_1997);
and U2026 (N_2026,N_1999,N_1887);
and U2027 (N_2027,N_1898,N_1847);
nor U2028 (N_2028,N_1949,N_1854);
or U2029 (N_2029,N_1943,N_1940);
or U2030 (N_2030,N_1951,N_1840);
nand U2031 (N_2031,N_1905,N_1875);
nand U2032 (N_2032,N_1876,N_1977);
or U2033 (N_2033,N_1804,N_1828);
and U2034 (N_2034,N_1841,N_1975);
nand U2035 (N_2035,N_1901,N_1928);
or U2036 (N_2036,N_1993,N_1826);
nor U2037 (N_2037,N_1944,N_1871);
xor U2038 (N_2038,N_1817,N_1918);
and U2039 (N_2039,N_1955,N_1892);
or U2040 (N_2040,N_1800,N_1878);
nand U2041 (N_2041,N_1978,N_1976);
or U2042 (N_2042,N_1965,N_1857);
nor U2043 (N_2043,N_1844,N_1853);
and U2044 (N_2044,N_1995,N_1859);
or U2045 (N_2045,N_1924,N_1873);
nand U2046 (N_2046,N_1908,N_1868);
nand U2047 (N_2047,N_1916,N_1930);
nand U2048 (N_2048,N_1860,N_1852);
and U2049 (N_2049,N_1858,N_1969);
nand U2050 (N_2050,N_1885,N_1945);
and U2051 (N_2051,N_1959,N_1909);
nor U2052 (N_2052,N_1912,N_1899);
nor U2053 (N_2053,N_1837,N_1835);
or U2054 (N_2054,N_1923,N_1961);
nor U2055 (N_2055,N_1960,N_1958);
nand U2056 (N_2056,N_1863,N_1981);
nand U2057 (N_2057,N_1937,N_1986);
nor U2058 (N_2058,N_1815,N_1897);
or U2059 (N_2059,N_1998,N_1882);
and U2060 (N_2060,N_1808,N_1812);
nor U2061 (N_2061,N_1946,N_1849);
or U2062 (N_2062,N_1810,N_1850);
and U2063 (N_2063,N_1855,N_1893);
xor U2064 (N_2064,N_1856,N_1966);
nand U2065 (N_2065,N_1874,N_1830);
nor U2066 (N_2066,N_1941,N_1839);
or U2067 (N_2067,N_1869,N_1831);
nor U2068 (N_2068,N_1829,N_1979);
nand U2069 (N_2069,N_1862,N_1805);
and U2070 (N_2070,N_1915,N_1996);
nor U2071 (N_2071,N_1967,N_1971);
xnor U2072 (N_2072,N_1824,N_1927);
or U2073 (N_2073,N_1950,N_1919);
nand U2074 (N_2074,N_1925,N_1913);
nor U2075 (N_2075,N_1989,N_1900);
or U2076 (N_2076,N_1890,N_1933);
and U2077 (N_2077,N_1848,N_1833);
or U2078 (N_2078,N_1894,N_1911);
and U2079 (N_2079,N_1822,N_1992);
or U2080 (N_2080,N_1888,N_1851);
nand U2081 (N_2081,N_1803,N_1819);
nor U2082 (N_2082,N_1932,N_1864);
or U2083 (N_2083,N_1865,N_1802);
or U2084 (N_2084,N_1987,N_1842);
or U2085 (N_2085,N_1870,N_1968);
nand U2086 (N_2086,N_1983,N_1922);
nand U2087 (N_2087,N_1904,N_1990);
or U2088 (N_2088,N_1962,N_1931);
and U2089 (N_2089,N_1920,N_1952);
or U2090 (N_2090,N_1834,N_1896);
or U2091 (N_2091,N_1963,N_1917);
nor U2092 (N_2092,N_1994,N_1964);
nor U2093 (N_2093,N_1809,N_1974);
xor U2094 (N_2094,N_1881,N_1980);
nand U2095 (N_2095,N_1985,N_1886);
or U2096 (N_2096,N_1954,N_1827);
or U2097 (N_2097,N_1936,N_1906);
nand U2098 (N_2098,N_1825,N_1973);
nand U2099 (N_2099,N_1935,N_1814);
and U2100 (N_2100,N_1850,N_1933);
and U2101 (N_2101,N_1849,N_1825);
and U2102 (N_2102,N_1951,N_1867);
nor U2103 (N_2103,N_1841,N_1863);
and U2104 (N_2104,N_1895,N_1816);
and U2105 (N_2105,N_1805,N_1831);
or U2106 (N_2106,N_1849,N_1837);
nand U2107 (N_2107,N_1900,N_1990);
or U2108 (N_2108,N_1858,N_1954);
or U2109 (N_2109,N_1974,N_1808);
or U2110 (N_2110,N_1851,N_1974);
and U2111 (N_2111,N_1839,N_1891);
and U2112 (N_2112,N_1853,N_1821);
nand U2113 (N_2113,N_1993,N_1806);
and U2114 (N_2114,N_1810,N_1802);
or U2115 (N_2115,N_1996,N_1816);
or U2116 (N_2116,N_1878,N_1815);
nor U2117 (N_2117,N_1817,N_1860);
nand U2118 (N_2118,N_1819,N_1946);
nor U2119 (N_2119,N_1980,N_1933);
nand U2120 (N_2120,N_1951,N_1895);
nor U2121 (N_2121,N_1991,N_1826);
nand U2122 (N_2122,N_1957,N_1807);
or U2123 (N_2123,N_1907,N_1967);
and U2124 (N_2124,N_1896,N_1930);
nand U2125 (N_2125,N_1846,N_1935);
nand U2126 (N_2126,N_1993,N_1998);
nand U2127 (N_2127,N_1875,N_1979);
nor U2128 (N_2128,N_1871,N_1973);
and U2129 (N_2129,N_1911,N_1877);
and U2130 (N_2130,N_1851,N_1939);
nand U2131 (N_2131,N_1810,N_1984);
nor U2132 (N_2132,N_1952,N_1968);
nand U2133 (N_2133,N_1893,N_1822);
or U2134 (N_2134,N_1833,N_1930);
and U2135 (N_2135,N_1925,N_1885);
nand U2136 (N_2136,N_1810,N_1970);
nand U2137 (N_2137,N_1939,N_1848);
and U2138 (N_2138,N_1822,N_1826);
nand U2139 (N_2139,N_1829,N_1936);
and U2140 (N_2140,N_1813,N_1869);
nor U2141 (N_2141,N_1874,N_1909);
nor U2142 (N_2142,N_1876,N_1818);
nor U2143 (N_2143,N_1956,N_1896);
nor U2144 (N_2144,N_1935,N_1816);
and U2145 (N_2145,N_1805,N_1965);
nor U2146 (N_2146,N_1895,N_1943);
and U2147 (N_2147,N_1873,N_1912);
or U2148 (N_2148,N_1858,N_1906);
nor U2149 (N_2149,N_1801,N_1888);
and U2150 (N_2150,N_1867,N_1825);
nand U2151 (N_2151,N_1807,N_1961);
nor U2152 (N_2152,N_1913,N_1995);
nor U2153 (N_2153,N_1834,N_1830);
or U2154 (N_2154,N_1955,N_1838);
nor U2155 (N_2155,N_1948,N_1978);
nand U2156 (N_2156,N_1957,N_1894);
nand U2157 (N_2157,N_1803,N_1937);
or U2158 (N_2158,N_1890,N_1800);
or U2159 (N_2159,N_1956,N_1977);
nand U2160 (N_2160,N_1852,N_1992);
or U2161 (N_2161,N_1898,N_1930);
and U2162 (N_2162,N_1977,N_1867);
and U2163 (N_2163,N_1801,N_1912);
or U2164 (N_2164,N_1966,N_1910);
or U2165 (N_2165,N_1986,N_1893);
or U2166 (N_2166,N_1992,N_1862);
nor U2167 (N_2167,N_1856,N_1883);
or U2168 (N_2168,N_1824,N_1961);
nand U2169 (N_2169,N_1990,N_1864);
or U2170 (N_2170,N_1904,N_1941);
and U2171 (N_2171,N_1839,N_1956);
and U2172 (N_2172,N_1813,N_1877);
nor U2173 (N_2173,N_1880,N_1937);
or U2174 (N_2174,N_1803,N_1907);
nor U2175 (N_2175,N_1837,N_1818);
nor U2176 (N_2176,N_1947,N_1833);
or U2177 (N_2177,N_1973,N_1942);
nor U2178 (N_2178,N_1827,N_1921);
nor U2179 (N_2179,N_1856,N_1982);
nor U2180 (N_2180,N_1956,N_1907);
nand U2181 (N_2181,N_1915,N_1989);
or U2182 (N_2182,N_1811,N_1952);
nand U2183 (N_2183,N_1926,N_1804);
and U2184 (N_2184,N_1967,N_1865);
nor U2185 (N_2185,N_1890,N_1809);
nand U2186 (N_2186,N_1959,N_1889);
and U2187 (N_2187,N_1816,N_1894);
nor U2188 (N_2188,N_1993,N_1914);
and U2189 (N_2189,N_1836,N_1908);
nand U2190 (N_2190,N_1907,N_1972);
nand U2191 (N_2191,N_1801,N_1842);
nand U2192 (N_2192,N_1885,N_1944);
and U2193 (N_2193,N_1939,N_1962);
or U2194 (N_2194,N_1818,N_1859);
and U2195 (N_2195,N_1874,N_1970);
nand U2196 (N_2196,N_1948,N_1981);
nor U2197 (N_2197,N_1997,N_1979);
nor U2198 (N_2198,N_1848,N_1868);
nand U2199 (N_2199,N_1885,N_1815);
and U2200 (N_2200,N_2082,N_2056);
nor U2201 (N_2201,N_2144,N_2073);
or U2202 (N_2202,N_2122,N_2064);
nand U2203 (N_2203,N_2126,N_2023);
or U2204 (N_2204,N_2098,N_2184);
nor U2205 (N_2205,N_2183,N_2119);
nand U2206 (N_2206,N_2032,N_2015);
nand U2207 (N_2207,N_2191,N_2132);
nor U2208 (N_2208,N_2103,N_2146);
nand U2209 (N_2209,N_2190,N_2020);
nand U2210 (N_2210,N_2050,N_2158);
nor U2211 (N_2211,N_2016,N_2070);
nand U2212 (N_2212,N_2072,N_2051);
nor U2213 (N_2213,N_2149,N_2186);
or U2214 (N_2214,N_2108,N_2067);
nor U2215 (N_2215,N_2076,N_2196);
nand U2216 (N_2216,N_2054,N_2038);
or U2217 (N_2217,N_2083,N_2057);
or U2218 (N_2218,N_2091,N_2141);
nor U2219 (N_2219,N_2000,N_2112);
and U2220 (N_2220,N_2048,N_2148);
and U2221 (N_2221,N_2100,N_2024);
nand U2222 (N_2222,N_2171,N_2173);
and U2223 (N_2223,N_2130,N_2081);
and U2224 (N_2224,N_2143,N_2089);
or U2225 (N_2225,N_2116,N_2153);
and U2226 (N_2226,N_2071,N_2147);
or U2227 (N_2227,N_2195,N_2140);
or U2228 (N_2228,N_2027,N_2181);
or U2229 (N_2229,N_2055,N_2011);
or U2230 (N_2230,N_2008,N_2097);
nor U2231 (N_2231,N_2075,N_2018);
nor U2232 (N_2232,N_2193,N_2155);
or U2233 (N_2233,N_2077,N_2017);
nand U2234 (N_2234,N_2175,N_2036);
or U2235 (N_2235,N_2078,N_2159);
nand U2236 (N_2236,N_2106,N_2022);
or U2237 (N_2237,N_2131,N_2165);
nand U2238 (N_2238,N_2188,N_2026);
or U2239 (N_2239,N_2066,N_2162);
nand U2240 (N_2240,N_2128,N_2139);
nor U2241 (N_2241,N_2010,N_2194);
nand U2242 (N_2242,N_2142,N_2198);
nor U2243 (N_2243,N_2102,N_2125);
nor U2244 (N_2244,N_2160,N_2154);
nor U2245 (N_2245,N_2185,N_2172);
or U2246 (N_2246,N_2180,N_2136);
nor U2247 (N_2247,N_2123,N_2189);
or U2248 (N_2248,N_2034,N_2033);
nor U2249 (N_2249,N_2019,N_2029);
nor U2250 (N_2250,N_2174,N_2065);
or U2251 (N_2251,N_2021,N_2151);
or U2252 (N_2252,N_2135,N_2093);
and U2253 (N_2253,N_2028,N_2035);
nand U2254 (N_2254,N_2170,N_2007);
nor U2255 (N_2255,N_2152,N_2012);
nor U2256 (N_2256,N_2031,N_2133);
and U2257 (N_2257,N_2005,N_2134);
or U2258 (N_2258,N_2177,N_2013);
nor U2259 (N_2259,N_2052,N_2163);
and U2260 (N_2260,N_2124,N_2061);
and U2261 (N_2261,N_2101,N_2182);
nor U2262 (N_2262,N_2009,N_2058);
and U2263 (N_2263,N_2085,N_2059);
or U2264 (N_2264,N_2129,N_2117);
and U2265 (N_2265,N_2063,N_2178);
nand U2266 (N_2266,N_2045,N_2192);
nand U2267 (N_2267,N_2169,N_2004);
xnor U2268 (N_2268,N_2105,N_2114);
nand U2269 (N_2269,N_2039,N_2113);
and U2270 (N_2270,N_2109,N_2006);
xor U2271 (N_2271,N_2069,N_2086);
nand U2272 (N_2272,N_2044,N_2167);
nand U2273 (N_2273,N_2176,N_2041);
or U2274 (N_2274,N_2120,N_2042);
nor U2275 (N_2275,N_2040,N_2092);
or U2276 (N_2276,N_2030,N_2079);
or U2277 (N_2277,N_2107,N_2001);
nand U2278 (N_2278,N_2037,N_2087);
nand U2279 (N_2279,N_2090,N_2121);
nand U2280 (N_2280,N_2145,N_2168);
or U2281 (N_2281,N_2047,N_2014);
nor U2282 (N_2282,N_2138,N_2049);
and U2283 (N_2283,N_2150,N_2197);
or U2284 (N_2284,N_2164,N_2157);
nand U2285 (N_2285,N_2003,N_2110);
nor U2286 (N_2286,N_2074,N_2095);
nand U2287 (N_2287,N_2096,N_2068);
and U2288 (N_2288,N_2025,N_2094);
or U2289 (N_2289,N_2053,N_2127);
or U2290 (N_2290,N_2161,N_2043);
and U2291 (N_2291,N_2156,N_2104);
nor U2292 (N_2292,N_2199,N_2002);
nor U2293 (N_2293,N_2084,N_2118);
nor U2294 (N_2294,N_2166,N_2099);
nand U2295 (N_2295,N_2062,N_2080);
and U2296 (N_2296,N_2088,N_2187);
and U2297 (N_2297,N_2179,N_2046);
or U2298 (N_2298,N_2111,N_2060);
nand U2299 (N_2299,N_2137,N_2115);
nand U2300 (N_2300,N_2190,N_2126);
nor U2301 (N_2301,N_2049,N_2173);
nor U2302 (N_2302,N_2164,N_2171);
nor U2303 (N_2303,N_2111,N_2108);
nand U2304 (N_2304,N_2120,N_2080);
or U2305 (N_2305,N_2062,N_2094);
or U2306 (N_2306,N_2111,N_2084);
nor U2307 (N_2307,N_2183,N_2016);
and U2308 (N_2308,N_2148,N_2179);
nor U2309 (N_2309,N_2199,N_2089);
nand U2310 (N_2310,N_2083,N_2196);
nor U2311 (N_2311,N_2089,N_2090);
nor U2312 (N_2312,N_2084,N_2099);
and U2313 (N_2313,N_2086,N_2147);
or U2314 (N_2314,N_2045,N_2109);
or U2315 (N_2315,N_2167,N_2050);
and U2316 (N_2316,N_2094,N_2127);
nand U2317 (N_2317,N_2046,N_2064);
nand U2318 (N_2318,N_2002,N_2095);
and U2319 (N_2319,N_2080,N_2162);
and U2320 (N_2320,N_2054,N_2128);
and U2321 (N_2321,N_2143,N_2054);
or U2322 (N_2322,N_2087,N_2162);
nand U2323 (N_2323,N_2114,N_2133);
nor U2324 (N_2324,N_2153,N_2171);
nand U2325 (N_2325,N_2159,N_2129);
or U2326 (N_2326,N_2033,N_2140);
nor U2327 (N_2327,N_2113,N_2178);
nand U2328 (N_2328,N_2011,N_2160);
nand U2329 (N_2329,N_2173,N_2168);
nor U2330 (N_2330,N_2097,N_2081);
and U2331 (N_2331,N_2043,N_2158);
and U2332 (N_2332,N_2047,N_2038);
nand U2333 (N_2333,N_2011,N_2162);
xor U2334 (N_2334,N_2187,N_2120);
nand U2335 (N_2335,N_2132,N_2058);
nor U2336 (N_2336,N_2155,N_2184);
nand U2337 (N_2337,N_2008,N_2125);
nand U2338 (N_2338,N_2138,N_2083);
and U2339 (N_2339,N_2051,N_2075);
and U2340 (N_2340,N_2154,N_2142);
nand U2341 (N_2341,N_2000,N_2132);
or U2342 (N_2342,N_2161,N_2097);
nor U2343 (N_2343,N_2110,N_2064);
nor U2344 (N_2344,N_2090,N_2192);
and U2345 (N_2345,N_2151,N_2014);
or U2346 (N_2346,N_2192,N_2098);
nor U2347 (N_2347,N_2029,N_2091);
and U2348 (N_2348,N_2160,N_2134);
nor U2349 (N_2349,N_2169,N_2081);
or U2350 (N_2350,N_2125,N_2018);
nor U2351 (N_2351,N_2150,N_2142);
nor U2352 (N_2352,N_2165,N_2105);
and U2353 (N_2353,N_2108,N_2138);
nor U2354 (N_2354,N_2156,N_2004);
nand U2355 (N_2355,N_2023,N_2173);
nor U2356 (N_2356,N_2098,N_2195);
or U2357 (N_2357,N_2014,N_2146);
and U2358 (N_2358,N_2072,N_2155);
nor U2359 (N_2359,N_2192,N_2017);
or U2360 (N_2360,N_2105,N_2123);
or U2361 (N_2361,N_2126,N_2032);
nand U2362 (N_2362,N_2149,N_2052);
or U2363 (N_2363,N_2126,N_2138);
nand U2364 (N_2364,N_2189,N_2007);
nand U2365 (N_2365,N_2018,N_2173);
and U2366 (N_2366,N_2109,N_2196);
or U2367 (N_2367,N_2154,N_2004);
and U2368 (N_2368,N_2048,N_2068);
nor U2369 (N_2369,N_2149,N_2085);
nand U2370 (N_2370,N_2033,N_2081);
nand U2371 (N_2371,N_2170,N_2084);
nand U2372 (N_2372,N_2101,N_2074);
nand U2373 (N_2373,N_2189,N_2014);
nand U2374 (N_2374,N_2088,N_2084);
nand U2375 (N_2375,N_2001,N_2104);
nor U2376 (N_2376,N_2189,N_2099);
and U2377 (N_2377,N_2164,N_2127);
or U2378 (N_2378,N_2114,N_2130);
nor U2379 (N_2379,N_2036,N_2109);
and U2380 (N_2380,N_2156,N_2035);
or U2381 (N_2381,N_2108,N_2129);
and U2382 (N_2382,N_2053,N_2082);
nand U2383 (N_2383,N_2070,N_2021);
and U2384 (N_2384,N_2086,N_2074);
nand U2385 (N_2385,N_2075,N_2191);
nand U2386 (N_2386,N_2151,N_2169);
nand U2387 (N_2387,N_2114,N_2163);
nor U2388 (N_2388,N_2078,N_2007);
or U2389 (N_2389,N_2198,N_2140);
and U2390 (N_2390,N_2166,N_2067);
nand U2391 (N_2391,N_2134,N_2099);
and U2392 (N_2392,N_2194,N_2104);
or U2393 (N_2393,N_2128,N_2084);
and U2394 (N_2394,N_2044,N_2164);
nand U2395 (N_2395,N_2084,N_2065);
nand U2396 (N_2396,N_2148,N_2156);
and U2397 (N_2397,N_2009,N_2137);
and U2398 (N_2398,N_2021,N_2044);
nor U2399 (N_2399,N_2114,N_2158);
and U2400 (N_2400,N_2229,N_2236);
and U2401 (N_2401,N_2367,N_2304);
or U2402 (N_2402,N_2230,N_2346);
nor U2403 (N_2403,N_2328,N_2355);
nand U2404 (N_2404,N_2205,N_2335);
and U2405 (N_2405,N_2246,N_2212);
nor U2406 (N_2406,N_2286,N_2253);
nand U2407 (N_2407,N_2359,N_2273);
and U2408 (N_2408,N_2203,N_2329);
nor U2409 (N_2409,N_2370,N_2323);
nand U2410 (N_2410,N_2245,N_2351);
or U2411 (N_2411,N_2298,N_2318);
and U2412 (N_2412,N_2218,N_2306);
or U2413 (N_2413,N_2310,N_2297);
nor U2414 (N_2414,N_2248,N_2373);
nor U2415 (N_2415,N_2295,N_2316);
nand U2416 (N_2416,N_2385,N_2281);
nand U2417 (N_2417,N_2381,N_2266);
and U2418 (N_2418,N_2380,N_2209);
or U2419 (N_2419,N_2233,N_2361);
nand U2420 (N_2420,N_2338,N_2302);
and U2421 (N_2421,N_2326,N_2276);
nor U2422 (N_2422,N_2348,N_2382);
and U2423 (N_2423,N_2208,N_2368);
nor U2424 (N_2424,N_2223,N_2264);
or U2425 (N_2425,N_2312,N_2268);
nor U2426 (N_2426,N_2299,N_2340);
nand U2427 (N_2427,N_2331,N_2337);
nor U2428 (N_2428,N_2239,N_2307);
nor U2429 (N_2429,N_2219,N_2360);
and U2430 (N_2430,N_2272,N_2242);
or U2431 (N_2431,N_2365,N_2345);
nand U2432 (N_2432,N_2263,N_2349);
or U2433 (N_2433,N_2293,N_2213);
nand U2434 (N_2434,N_2224,N_2366);
and U2435 (N_2435,N_2332,N_2291);
nor U2436 (N_2436,N_2265,N_2249);
nand U2437 (N_2437,N_2371,N_2280);
nand U2438 (N_2438,N_2217,N_2251);
nand U2439 (N_2439,N_2398,N_2358);
or U2440 (N_2440,N_2319,N_2261);
and U2441 (N_2441,N_2391,N_2247);
nand U2442 (N_2442,N_2379,N_2388);
nor U2443 (N_2443,N_2221,N_2389);
nand U2444 (N_2444,N_2336,N_2288);
or U2445 (N_2445,N_2339,N_2262);
nand U2446 (N_2446,N_2311,N_2383);
or U2447 (N_2447,N_2200,N_2308);
and U2448 (N_2448,N_2322,N_2238);
or U2449 (N_2449,N_2216,N_2395);
and U2450 (N_2450,N_2271,N_2354);
and U2451 (N_2451,N_2243,N_2227);
nand U2452 (N_2452,N_2282,N_2300);
and U2453 (N_2453,N_2237,N_2378);
nand U2454 (N_2454,N_2364,N_2325);
nor U2455 (N_2455,N_2285,N_2244);
and U2456 (N_2456,N_2397,N_2347);
and U2457 (N_2457,N_2270,N_2374);
or U2458 (N_2458,N_2204,N_2235);
and U2459 (N_2459,N_2240,N_2215);
and U2460 (N_2460,N_2343,N_2384);
or U2461 (N_2461,N_2254,N_2377);
and U2462 (N_2462,N_2225,N_2241);
and U2463 (N_2463,N_2301,N_2258);
nand U2464 (N_2464,N_2375,N_2320);
and U2465 (N_2465,N_2290,N_2260);
and U2466 (N_2466,N_2369,N_2287);
nor U2467 (N_2467,N_2390,N_2267);
or U2468 (N_2468,N_2330,N_2333);
nor U2469 (N_2469,N_2392,N_2283);
nor U2470 (N_2470,N_2334,N_2372);
and U2471 (N_2471,N_2314,N_2211);
nor U2472 (N_2472,N_2206,N_2393);
nor U2473 (N_2473,N_2363,N_2234);
nand U2474 (N_2474,N_2292,N_2269);
nand U2475 (N_2475,N_2294,N_2362);
nor U2476 (N_2476,N_2207,N_2231);
nand U2477 (N_2477,N_2387,N_2317);
nand U2478 (N_2478,N_2327,N_2394);
and U2479 (N_2479,N_2344,N_2202);
nand U2480 (N_2480,N_2352,N_2396);
or U2481 (N_2481,N_2210,N_2321);
nand U2482 (N_2482,N_2257,N_2350);
and U2483 (N_2483,N_2232,N_2305);
or U2484 (N_2484,N_2315,N_2222);
nor U2485 (N_2485,N_2303,N_2278);
nor U2486 (N_2486,N_2342,N_2275);
and U2487 (N_2487,N_2214,N_2353);
or U2488 (N_2488,N_2386,N_2277);
xnor U2489 (N_2489,N_2256,N_2279);
nor U2490 (N_2490,N_2220,N_2376);
nand U2491 (N_2491,N_2252,N_2356);
nor U2492 (N_2492,N_2313,N_2399);
nand U2493 (N_2493,N_2296,N_2324);
nor U2494 (N_2494,N_2201,N_2284);
and U2495 (N_2495,N_2309,N_2255);
and U2496 (N_2496,N_2341,N_2228);
nor U2497 (N_2497,N_2274,N_2289);
or U2498 (N_2498,N_2259,N_2250);
or U2499 (N_2499,N_2357,N_2226);
nor U2500 (N_2500,N_2212,N_2236);
nand U2501 (N_2501,N_2236,N_2280);
nand U2502 (N_2502,N_2327,N_2255);
or U2503 (N_2503,N_2387,N_2382);
nor U2504 (N_2504,N_2353,N_2209);
or U2505 (N_2505,N_2397,N_2337);
nand U2506 (N_2506,N_2244,N_2395);
nor U2507 (N_2507,N_2343,N_2264);
nor U2508 (N_2508,N_2359,N_2212);
xor U2509 (N_2509,N_2354,N_2336);
nor U2510 (N_2510,N_2368,N_2375);
or U2511 (N_2511,N_2358,N_2300);
and U2512 (N_2512,N_2261,N_2323);
nor U2513 (N_2513,N_2349,N_2361);
and U2514 (N_2514,N_2266,N_2238);
nand U2515 (N_2515,N_2305,N_2371);
and U2516 (N_2516,N_2358,N_2311);
nand U2517 (N_2517,N_2262,N_2313);
nor U2518 (N_2518,N_2398,N_2204);
or U2519 (N_2519,N_2324,N_2399);
nor U2520 (N_2520,N_2320,N_2361);
nor U2521 (N_2521,N_2308,N_2317);
nor U2522 (N_2522,N_2245,N_2260);
nor U2523 (N_2523,N_2358,N_2227);
nor U2524 (N_2524,N_2318,N_2296);
and U2525 (N_2525,N_2264,N_2390);
or U2526 (N_2526,N_2285,N_2215);
or U2527 (N_2527,N_2313,N_2212);
or U2528 (N_2528,N_2313,N_2210);
and U2529 (N_2529,N_2350,N_2363);
nand U2530 (N_2530,N_2344,N_2336);
or U2531 (N_2531,N_2239,N_2220);
nor U2532 (N_2532,N_2303,N_2287);
and U2533 (N_2533,N_2278,N_2220);
nand U2534 (N_2534,N_2276,N_2322);
or U2535 (N_2535,N_2293,N_2227);
nand U2536 (N_2536,N_2390,N_2230);
nand U2537 (N_2537,N_2354,N_2385);
nand U2538 (N_2538,N_2305,N_2238);
nand U2539 (N_2539,N_2248,N_2333);
or U2540 (N_2540,N_2291,N_2285);
and U2541 (N_2541,N_2323,N_2250);
and U2542 (N_2542,N_2235,N_2247);
nor U2543 (N_2543,N_2209,N_2255);
nand U2544 (N_2544,N_2388,N_2209);
nand U2545 (N_2545,N_2340,N_2335);
nor U2546 (N_2546,N_2329,N_2383);
nand U2547 (N_2547,N_2256,N_2324);
nand U2548 (N_2548,N_2391,N_2307);
and U2549 (N_2549,N_2298,N_2237);
nor U2550 (N_2550,N_2316,N_2233);
nand U2551 (N_2551,N_2255,N_2366);
nor U2552 (N_2552,N_2324,N_2249);
nor U2553 (N_2553,N_2213,N_2274);
xnor U2554 (N_2554,N_2277,N_2338);
nand U2555 (N_2555,N_2352,N_2322);
nand U2556 (N_2556,N_2329,N_2336);
and U2557 (N_2557,N_2208,N_2299);
xnor U2558 (N_2558,N_2247,N_2263);
and U2559 (N_2559,N_2295,N_2234);
or U2560 (N_2560,N_2205,N_2272);
nand U2561 (N_2561,N_2318,N_2378);
or U2562 (N_2562,N_2217,N_2366);
nand U2563 (N_2563,N_2362,N_2221);
nand U2564 (N_2564,N_2278,N_2262);
nor U2565 (N_2565,N_2213,N_2369);
nand U2566 (N_2566,N_2348,N_2255);
and U2567 (N_2567,N_2295,N_2349);
and U2568 (N_2568,N_2296,N_2373);
nor U2569 (N_2569,N_2275,N_2329);
nor U2570 (N_2570,N_2354,N_2335);
nor U2571 (N_2571,N_2249,N_2352);
or U2572 (N_2572,N_2342,N_2263);
nor U2573 (N_2573,N_2367,N_2238);
nor U2574 (N_2574,N_2241,N_2290);
or U2575 (N_2575,N_2392,N_2296);
nor U2576 (N_2576,N_2362,N_2332);
and U2577 (N_2577,N_2203,N_2389);
or U2578 (N_2578,N_2258,N_2253);
and U2579 (N_2579,N_2235,N_2350);
nand U2580 (N_2580,N_2347,N_2236);
nor U2581 (N_2581,N_2258,N_2316);
and U2582 (N_2582,N_2266,N_2285);
nor U2583 (N_2583,N_2216,N_2224);
nor U2584 (N_2584,N_2316,N_2376);
and U2585 (N_2585,N_2257,N_2277);
nand U2586 (N_2586,N_2306,N_2395);
or U2587 (N_2587,N_2377,N_2394);
nand U2588 (N_2588,N_2256,N_2215);
and U2589 (N_2589,N_2304,N_2362);
and U2590 (N_2590,N_2332,N_2264);
nand U2591 (N_2591,N_2277,N_2311);
nand U2592 (N_2592,N_2227,N_2366);
or U2593 (N_2593,N_2399,N_2292);
and U2594 (N_2594,N_2209,N_2250);
nand U2595 (N_2595,N_2220,N_2261);
nand U2596 (N_2596,N_2306,N_2237);
and U2597 (N_2597,N_2217,N_2383);
or U2598 (N_2598,N_2315,N_2269);
and U2599 (N_2599,N_2341,N_2291);
nor U2600 (N_2600,N_2469,N_2551);
and U2601 (N_2601,N_2510,N_2459);
nor U2602 (N_2602,N_2499,N_2512);
or U2603 (N_2603,N_2425,N_2516);
and U2604 (N_2604,N_2568,N_2585);
or U2605 (N_2605,N_2534,N_2525);
and U2606 (N_2606,N_2414,N_2485);
nand U2607 (N_2607,N_2579,N_2564);
nand U2608 (N_2608,N_2589,N_2448);
nand U2609 (N_2609,N_2515,N_2432);
and U2610 (N_2610,N_2419,N_2488);
or U2611 (N_2611,N_2490,N_2595);
and U2612 (N_2612,N_2555,N_2536);
or U2613 (N_2613,N_2550,N_2545);
and U2614 (N_2614,N_2497,N_2524);
nor U2615 (N_2615,N_2539,N_2484);
and U2616 (N_2616,N_2558,N_2500);
nor U2617 (N_2617,N_2434,N_2476);
or U2618 (N_2618,N_2491,N_2503);
nor U2619 (N_2619,N_2466,N_2535);
nor U2620 (N_2620,N_2482,N_2412);
nor U2621 (N_2621,N_2592,N_2546);
nand U2622 (N_2622,N_2454,N_2439);
or U2623 (N_2623,N_2410,N_2544);
or U2624 (N_2624,N_2526,N_2517);
nor U2625 (N_2625,N_2438,N_2580);
or U2626 (N_2626,N_2446,N_2547);
nand U2627 (N_2627,N_2511,N_2505);
or U2628 (N_2628,N_2553,N_2540);
nand U2629 (N_2629,N_2417,N_2496);
nor U2630 (N_2630,N_2538,N_2554);
nand U2631 (N_2631,N_2479,N_2567);
and U2632 (N_2632,N_2571,N_2495);
nor U2633 (N_2633,N_2584,N_2501);
nand U2634 (N_2634,N_2472,N_2478);
nor U2635 (N_2635,N_2442,N_2561);
and U2636 (N_2636,N_2541,N_2480);
or U2637 (N_2637,N_2444,N_2427);
or U2638 (N_2638,N_2455,N_2556);
xnor U2639 (N_2639,N_2424,N_2532);
nand U2640 (N_2640,N_2401,N_2477);
or U2641 (N_2641,N_2441,N_2514);
and U2642 (N_2642,N_2586,N_2519);
or U2643 (N_2643,N_2489,N_2423);
and U2644 (N_2644,N_2506,N_2529);
or U2645 (N_2645,N_2440,N_2431);
nand U2646 (N_2646,N_2436,N_2576);
or U2647 (N_2647,N_2404,N_2471);
nor U2648 (N_2648,N_2418,N_2578);
nor U2649 (N_2649,N_2437,N_2569);
or U2650 (N_2650,N_2572,N_2493);
nor U2651 (N_2651,N_2527,N_2559);
nor U2652 (N_2652,N_2597,N_2457);
or U2653 (N_2653,N_2599,N_2582);
or U2654 (N_2654,N_2447,N_2530);
and U2655 (N_2655,N_2591,N_2461);
nor U2656 (N_2656,N_2420,N_2502);
and U2657 (N_2657,N_2468,N_2449);
or U2658 (N_2658,N_2407,N_2481);
or U2659 (N_2659,N_2533,N_2543);
and U2660 (N_2660,N_2473,N_2464);
or U2661 (N_2661,N_2422,N_2537);
and U2662 (N_2662,N_2542,N_2594);
and U2663 (N_2663,N_2426,N_2460);
and U2664 (N_2664,N_2549,N_2400);
nor U2665 (N_2665,N_2596,N_2415);
nand U2666 (N_2666,N_2433,N_2557);
nand U2667 (N_2667,N_2452,N_2451);
nand U2668 (N_2668,N_2590,N_2416);
nand U2669 (N_2669,N_2507,N_2494);
nor U2670 (N_2670,N_2483,N_2453);
and U2671 (N_2671,N_2456,N_2518);
nand U2672 (N_2672,N_2562,N_2560);
or U2673 (N_2673,N_2552,N_2548);
nand U2674 (N_2674,N_2563,N_2587);
and U2675 (N_2675,N_2509,N_2570);
and U2676 (N_2676,N_2575,N_2450);
and U2677 (N_2677,N_2435,N_2598);
nor U2678 (N_2678,N_2593,N_2465);
nand U2679 (N_2679,N_2405,N_2467);
nor U2680 (N_2680,N_2430,N_2486);
and U2681 (N_2681,N_2521,N_2492);
nand U2682 (N_2682,N_2522,N_2411);
or U2683 (N_2683,N_2445,N_2531);
nand U2684 (N_2684,N_2470,N_2528);
and U2685 (N_2685,N_2463,N_2574);
or U2686 (N_2686,N_2428,N_2588);
nor U2687 (N_2687,N_2583,N_2487);
nor U2688 (N_2688,N_2513,N_2508);
and U2689 (N_2689,N_2581,N_2577);
or U2690 (N_2690,N_2406,N_2566);
nand U2691 (N_2691,N_2474,N_2573);
nor U2692 (N_2692,N_2408,N_2409);
and U2693 (N_2693,N_2523,N_2504);
nand U2694 (N_2694,N_2413,N_2443);
and U2695 (N_2695,N_2462,N_2429);
nor U2696 (N_2696,N_2475,N_2498);
nand U2697 (N_2697,N_2421,N_2402);
nand U2698 (N_2698,N_2458,N_2520);
and U2699 (N_2699,N_2403,N_2565);
nor U2700 (N_2700,N_2408,N_2519);
nor U2701 (N_2701,N_2552,N_2479);
or U2702 (N_2702,N_2431,N_2439);
and U2703 (N_2703,N_2532,N_2591);
nor U2704 (N_2704,N_2489,N_2523);
nand U2705 (N_2705,N_2482,N_2483);
or U2706 (N_2706,N_2431,N_2455);
and U2707 (N_2707,N_2517,N_2428);
nor U2708 (N_2708,N_2494,N_2529);
nand U2709 (N_2709,N_2537,N_2435);
nor U2710 (N_2710,N_2590,N_2519);
nand U2711 (N_2711,N_2486,N_2539);
or U2712 (N_2712,N_2572,N_2571);
or U2713 (N_2713,N_2555,N_2453);
nand U2714 (N_2714,N_2525,N_2477);
or U2715 (N_2715,N_2533,N_2507);
nor U2716 (N_2716,N_2499,N_2506);
or U2717 (N_2717,N_2452,N_2417);
or U2718 (N_2718,N_2552,N_2476);
or U2719 (N_2719,N_2443,N_2521);
or U2720 (N_2720,N_2594,N_2491);
or U2721 (N_2721,N_2428,N_2509);
or U2722 (N_2722,N_2589,N_2402);
and U2723 (N_2723,N_2496,N_2510);
nor U2724 (N_2724,N_2498,N_2566);
nor U2725 (N_2725,N_2494,N_2599);
nor U2726 (N_2726,N_2543,N_2498);
or U2727 (N_2727,N_2434,N_2556);
nand U2728 (N_2728,N_2407,N_2593);
and U2729 (N_2729,N_2549,N_2485);
or U2730 (N_2730,N_2522,N_2541);
nand U2731 (N_2731,N_2506,N_2433);
nand U2732 (N_2732,N_2567,N_2499);
nor U2733 (N_2733,N_2565,N_2400);
or U2734 (N_2734,N_2420,N_2493);
nand U2735 (N_2735,N_2425,N_2413);
nor U2736 (N_2736,N_2471,N_2405);
and U2737 (N_2737,N_2556,N_2514);
nor U2738 (N_2738,N_2510,N_2439);
nand U2739 (N_2739,N_2405,N_2475);
and U2740 (N_2740,N_2483,N_2559);
or U2741 (N_2741,N_2511,N_2566);
nor U2742 (N_2742,N_2432,N_2499);
nor U2743 (N_2743,N_2515,N_2441);
xor U2744 (N_2744,N_2452,N_2569);
nor U2745 (N_2745,N_2441,N_2588);
xnor U2746 (N_2746,N_2464,N_2576);
and U2747 (N_2747,N_2572,N_2494);
nand U2748 (N_2748,N_2445,N_2570);
and U2749 (N_2749,N_2553,N_2470);
or U2750 (N_2750,N_2514,N_2561);
or U2751 (N_2751,N_2526,N_2425);
nor U2752 (N_2752,N_2435,N_2494);
or U2753 (N_2753,N_2532,N_2416);
nor U2754 (N_2754,N_2538,N_2509);
nor U2755 (N_2755,N_2407,N_2514);
nor U2756 (N_2756,N_2472,N_2471);
and U2757 (N_2757,N_2550,N_2448);
nand U2758 (N_2758,N_2462,N_2582);
or U2759 (N_2759,N_2524,N_2560);
nor U2760 (N_2760,N_2570,N_2462);
or U2761 (N_2761,N_2570,N_2553);
nand U2762 (N_2762,N_2584,N_2425);
or U2763 (N_2763,N_2546,N_2473);
and U2764 (N_2764,N_2511,N_2466);
nor U2765 (N_2765,N_2478,N_2447);
or U2766 (N_2766,N_2422,N_2532);
nor U2767 (N_2767,N_2519,N_2559);
nand U2768 (N_2768,N_2413,N_2532);
and U2769 (N_2769,N_2522,N_2449);
or U2770 (N_2770,N_2514,N_2446);
or U2771 (N_2771,N_2472,N_2588);
nand U2772 (N_2772,N_2493,N_2579);
nor U2773 (N_2773,N_2526,N_2459);
or U2774 (N_2774,N_2496,N_2457);
or U2775 (N_2775,N_2468,N_2438);
and U2776 (N_2776,N_2462,N_2492);
nor U2777 (N_2777,N_2453,N_2470);
nor U2778 (N_2778,N_2575,N_2531);
or U2779 (N_2779,N_2582,N_2579);
and U2780 (N_2780,N_2515,N_2526);
or U2781 (N_2781,N_2450,N_2424);
or U2782 (N_2782,N_2517,N_2496);
xor U2783 (N_2783,N_2576,N_2405);
nand U2784 (N_2784,N_2584,N_2526);
nor U2785 (N_2785,N_2587,N_2500);
or U2786 (N_2786,N_2571,N_2452);
and U2787 (N_2787,N_2500,N_2514);
and U2788 (N_2788,N_2457,N_2487);
nor U2789 (N_2789,N_2464,N_2501);
and U2790 (N_2790,N_2419,N_2553);
nor U2791 (N_2791,N_2576,N_2561);
nand U2792 (N_2792,N_2455,N_2428);
or U2793 (N_2793,N_2567,N_2571);
nor U2794 (N_2794,N_2487,N_2566);
and U2795 (N_2795,N_2445,N_2447);
nor U2796 (N_2796,N_2470,N_2412);
or U2797 (N_2797,N_2563,N_2570);
nand U2798 (N_2798,N_2588,N_2407);
and U2799 (N_2799,N_2561,N_2590);
or U2800 (N_2800,N_2749,N_2724);
or U2801 (N_2801,N_2706,N_2619);
or U2802 (N_2802,N_2602,N_2697);
and U2803 (N_2803,N_2636,N_2726);
nor U2804 (N_2804,N_2674,N_2649);
nor U2805 (N_2805,N_2797,N_2677);
nor U2806 (N_2806,N_2623,N_2730);
and U2807 (N_2807,N_2746,N_2750);
nor U2808 (N_2808,N_2688,N_2661);
and U2809 (N_2809,N_2668,N_2625);
and U2810 (N_2810,N_2616,N_2716);
nand U2811 (N_2811,N_2765,N_2679);
nand U2812 (N_2812,N_2759,N_2747);
nand U2813 (N_2813,N_2685,N_2709);
or U2814 (N_2814,N_2736,N_2645);
nor U2815 (N_2815,N_2711,N_2784);
and U2816 (N_2816,N_2775,N_2631);
nand U2817 (N_2817,N_2703,N_2639);
nor U2818 (N_2818,N_2614,N_2753);
and U2819 (N_2819,N_2792,N_2712);
nand U2820 (N_2820,N_2624,N_2774);
nor U2821 (N_2821,N_2657,N_2764);
and U2822 (N_2822,N_2637,N_2666);
nor U2823 (N_2823,N_2717,N_2606);
or U2824 (N_2824,N_2683,N_2618);
nand U2825 (N_2825,N_2720,N_2741);
or U2826 (N_2826,N_2723,N_2684);
and U2827 (N_2827,N_2795,N_2762);
nor U2828 (N_2828,N_2693,N_2605);
and U2829 (N_2829,N_2781,N_2700);
nor U2830 (N_2830,N_2787,N_2669);
nor U2831 (N_2831,N_2760,N_2651);
or U2832 (N_2832,N_2673,N_2650);
or U2833 (N_2833,N_2632,N_2773);
nor U2834 (N_2834,N_2601,N_2788);
or U2835 (N_2835,N_2662,N_2740);
and U2836 (N_2836,N_2748,N_2702);
and U2837 (N_2837,N_2718,N_2676);
and U2838 (N_2838,N_2745,N_2769);
and U2839 (N_2839,N_2627,N_2611);
nand U2840 (N_2840,N_2600,N_2660);
and U2841 (N_2841,N_2667,N_2794);
and U2842 (N_2842,N_2691,N_2656);
nand U2843 (N_2843,N_2768,N_2786);
and U2844 (N_2844,N_2729,N_2613);
nand U2845 (N_2845,N_2728,N_2744);
or U2846 (N_2846,N_2752,N_2675);
or U2847 (N_2847,N_2789,N_2755);
or U2848 (N_2848,N_2622,N_2798);
nand U2849 (N_2849,N_2687,N_2761);
nand U2850 (N_2850,N_2756,N_2643);
and U2851 (N_2851,N_2626,N_2680);
nor U2852 (N_2852,N_2767,N_2612);
or U2853 (N_2853,N_2790,N_2725);
nand U2854 (N_2854,N_2791,N_2771);
nor U2855 (N_2855,N_2715,N_2694);
or U2856 (N_2856,N_2690,N_2772);
nor U2857 (N_2857,N_2727,N_2739);
and U2858 (N_2858,N_2705,N_2743);
and U2859 (N_2859,N_2799,N_2692);
or U2860 (N_2860,N_2737,N_2701);
and U2861 (N_2861,N_2665,N_2608);
nand U2862 (N_2862,N_2681,N_2628);
nor U2863 (N_2863,N_2695,N_2793);
nor U2864 (N_2864,N_2763,N_2610);
or U2865 (N_2865,N_2713,N_2607);
nor U2866 (N_2866,N_2640,N_2732);
and U2867 (N_2867,N_2766,N_2617);
and U2868 (N_2868,N_2641,N_2609);
nor U2869 (N_2869,N_2630,N_2664);
nand U2870 (N_2870,N_2777,N_2646);
nor U2871 (N_2871,N_2604,N_2655);
and U2872 (N_2872,N_2722,N_2686);
nor U2873 (N_2873,N_2654,N_2704);
nor U2874 (N_2874,N_2696,N_2714);
nor U2875 (N_2875,N_2778,N_2735);
and U2876 (N_2876,N_2707,N_2731);
nand U2877 (N_2877,N_2708,N_2621);
or U2878 (N_2878,N_2629,N_2672);
or U2879 (N_2879,N_2734,N_2783);
nor U2880 (N_2880,N_2671,N_2682);
nand U2881 (N_2881,N_2758,N_2742);
nor U2882 (N_2882,N_2782,N_2751);
or U2883 (N_2883,N_2603,N_2754);
or U2884 (N_2884,N_2642,N_2678);
nor U2885 (N_2885,N_2738,N_2653);
or U2886 (N_2886,N_2615,N_2652);
and U2887 (N_2887,N_2659,N_2620);
or U2888 (N_2888,N_2663,N_2780);
or U2889 (N_2889,N_2796,N_2647);
nand U2890 (N_2890,N_2644,N_2670);
or U2891 (N_2891,N_2634,N_2699);
nand U2892 (N_2892,N_2698,N_2785);
and U2893 (N_2893,N_2689,N_2770);
and U2894 (N_2894,N_2635,N_2757);
and U2895 (N_2895,N_2658,N_2733);
nand U2896 (N_2896,N_2721,N_2776);
nand U2897 (N_2897,N_2648,N_2633);
nand U2898 (N_2898,N_2710,N_2779);
or U2899 (N_2899,N_2719,N_2638);
or U2900 (N_2900,N_2770,N_2752);
nor U2901 (N_2901,N_2671,N_2755);
and U2902 (N_2902,N_2790,N_2695);
nor U2903 (N_2903,N_2661,N_2604);
nor U2904 (N_2904,N_2786,N_2745);
nand U2905 (N_2905,N_2638,N_2637);
nand U2906 (N_2906,N_2648,N_2730);
nand U2907 (N_2907,N_2729,N_2714);
nor U2908 (N_2908,N_2709,N_2744);
nand U2909 (N_2909,N_2660,N_2664);
nand U2910 (N_2910,N_2773,N_2643);
nand U2911 (N_2911,N_2646,N_2766);
nand U2912 (N_2912,N_2728,N_2672);
or U2913 (N_2913,N_2799,N_2774);
or U2914 (N_2914,N_2747,N_2651);
nand U2915 (N_2915,N_2622,N_2632);
or U2916 (N_2916,N_2654,N_2773);
or U2917 (N_2917,N_2603,N_2671);
or U2918 (N_2918,N_2636,N_2655);
and U2919 (N_2919,N_2764,N_2790);
or U2920 (N_2920,N_2673,N_2714);
and U2921 (N_2921,N_2656,N_2711);
and U2922 (N_2922,N_2683,N_2646);
nor U2923 (N_2923,N_2736,N_2752);
nor U2924 (N_2924,N_2748,N_2759);
nand U2925 (N_2925,N_2794,N_2783);
nor U2926 (N_2926,N_2673,N_2718);
nand U2927 (N_2927,N_2627,N_2677);
or U2928 (N_2928,N_2796,N_2753);
nand U2929 (N_2929,N_2725,N_2743);
and U2930 (N_2930,N_2710,N_2714);
or U2931 (N_2931,N_2751,N_2613);
nand U2932 (N_2932,N_2764,N_2693);
nand U2933 (N_2933,N_2745,N_2691);
or U2934 (N_2934,N_2791,N_2676);
or U2935 (N_2935,N_2690,N_2615);
or U2936 (N_2936,N_2725,N_2721);
nor U2937 (N_2937,N_2782,N_2633);
nor U2938 (N_2938,N_2645,N_2782);
or U2939 (N_2939,N_2601,N_2774);
and U2940 (N_2940,N_2739,N_2654);
nor U2941 (N_2941,N_2719,N_2697);
nor U2942 (N_2942,N_2770,N_2701);
nor U2943 (N_2943,N_2672,N_2663);
nand U2944 (N_2944,N_2770,N_2749);
or U2945 (N_2945,N_2666,N_2716);
nor U2946 (N_2946,N_2681,N_2748);
nor U2947 (N_2947,N_2676,N_2741);
or U2948 (N_2948,N_2759,N_2674);
nor U2949 (N_2949,N_2605,N_2682);
and U2950 (N_2950,N_2608,N_2617);
nor U2951 (N_2951,N_2672,N_2799);
or U2952 (N_2952,N_2600,N_2738);
nand U2953 (N_2953,N_2649,N_2699);
nand U2954 (N_2954,N_2717,N_2709);
or U2955 (N_2955,N_2656,N_2737);
nor U2956 (N_2956,N_2787,N_2672);
nand U2957 (N_2957,N_2643,N_2749);
nand U2958 (N_2958,N_2766,N_2799);
nor U2959 (N_2959,N_2682,N_2610);
nor U2960 (N_2960,N_2675,N_2630);
or U2961 (N_2961,N_2789,N_2758);
and U2962 (N_2962,N_2791,N_2749);
nand U2963 (N_2963,N_2711,N_2776);
or U2964 (N_2964,N_2657,N_2752);
and U2965 (N_2965,N_2697,N_2670);
or U2966 (N_2966,N_2782,N_2677);
or U2967 (N_2967,N_2692,N_2748);
nand U2968 (N_2968,N_2669,N_2658);
xnor U2969 (N_2969,N_2726,N_2667);
and U2970 (N_2970,N_2760,N_2655);
nand U2971 (N_2971,N_2781,N_2738);
nand U2972 (N_2972,N_2722,N_2643);
and U2973 (N_2973,N_2620,N_2746);
or U2974 (N_2974,N_2713,N_2690);
and U2975 (N_2975,N_2648,N_2665);
nor U2976 (N_2976,N_2620,N_2608);
or U2977 (N_2977,N_2611,N_2678);
and U2978 (N_2978,N_2715,N_2731);
nor U2979 (N_2979,N_2692,N_2643);
nand U2980 (N_2980,N_2694,N_2740);
nand U2981 (N_2981,N_2657,N_2616);
and U2982 (N_2982,N_2715,N_2644);
and U2983 (N_2983,N_2661,N_2680);
and U2984 (N_2984,N_2620,N_2634);
nor U2985 (N_2985,N_2647,N_2714);
nand U2986 (N_2986,N_2799,N_2613);
nand U2987 (N_2987,N_2753,N_2663);
nand U2988 (N_2988,N_2760,N_2648);
and U2989 (N_2989,N_2633,N_2693);
nand U2990 (N_2990,N_2638,N_2681);
or U2991 (N_2991,N_2645,N_2794);
and U2992 (N_2992,N_2788,N_2744);
nand U2993 (N_2993,N_2613,N_2774);
nand U2994 (N_2994,N_2703,N_2689);
nand U2995 (N_2995,N_2629,N_2740);
nor U2996 (N_2996,N_2736,N_2669);
nor U2997 (N_2997,N_2757,N_2783);
nor U2998 (N_2998,N_2689,N_2660);
and U2999 (N_2999,N_2694,N_2755);
or U3000 (N_3000,N_2847,N_2917);
or U3001 (N_3001,N_2832,N_2849);
or U3002 (N_3002,N_2900,N_2853);
or U3003 (N_3003,N_2930,N_2944);
and U3004 (N_3004,N_2845,N_2989);
nor U3005 (N_3005,N_2863,N_2966);
or U3006 (N_3006,N_2843,N_2830);
nand U3007 (N_3007,N_2954,N_2820);
and U3008 (N_3008,N_2866,N_2840);
and U3009 (N_3009,N_2943,N_2864);
nor U3010 (N_3010,N_2920,N_2877);
nand U3011 (N_3011,N_2945,N_2922);
nor U3012 (N_3012,N_2803,N_2899);
or U3013 (N_3013,N_2878,N_2862);
nor U3014 (N_3014,N_2857,N_2859);
and U3015 (N_3015,N_2875,N_2910);
nor U3016 (N_3016,N_2809,N_2971);
or U3017 (N_3017,N_2938,N_2984);
nor U3018 (N_3018,N_2992,N_2886);
or U3019 (N_3019,N_2928,N_2981);
nor U3020 (N_3020,N_2897,N_2978);
xnor U3021 (N_3021,N_2986,N_2942);
nor U3022 (N_3022,N_2879,N_2894);
nor U3023 (N_3023,N_2860,N_2896);
and U3024 (N_3024,N_2939,N_2818);
nor U3025 (N_3025,N_2888,N_2881);
nor U3026 (N_3026,N_2850,N_2958);
and U3027 (N_3027,N_2977,N_2976);
nand U3028 (N_3028,N_2858,N_2957);
nand U3029 (N_3029,N_2951,N_2831);
nor U3030 (N_3030,N_2835,N_2825);
or U3031 (N_3031,N_2880,N_2924);
nand U3032 (N_3032,N_2839,N_2911);
or U3033 (N_3033,N_2868,N_2991);
and U3034 (N_3034,N_2932,N_2996);
nand U3035 (N_3035,N_2994,N_2901);
nand U3036 (N_3036,N_2974,N_2908);
nor U3037 (N_3037,N_2870,N_2969);
nor U3038 (N_3038,N_2885,N_2801);
nor U3039 (N_3039,N_2874,N_2952);
nor U3040 (N_3040,N_2844,N_2872);
nor U3041 (N_3041,N_2972,N_2947);
and U3042 (N_3042,N_2893,N_2964);
xnor U3043 (N_3043,N_2834,N_2995);
nor U3044 (N_3044,N_2842,N_2923);
and U3045 (N_3045,N_2833,N_2817);
nand U3046 (N_3046,N_2869,N_2876);
nand U3047 (N_3047,N_2882,N_2927);
and U3048 (N_3048,N_2925,N_2946);
or U3049 (N_3049,N_2823,N_2916);
nand U3050 (N_3050,N_2967,N_2889);
nor U3051 (N_3051,N_2987,N_2913);
and U3052 (N_3052,N_2884,N_2919);
or U3053 (N_3053,N_2887,N_2931);
or U3054 (N_3054,N_2811,N_2812);
and U3055 (N_3055,N_2970,N_2993);
and U3056 (N_3056,N_2813,N_2965);
and U3057 (N_3057,N_2960,N_2814);
nor U3058 (N_3058,N_2982,N_2963);
or U3059 (N_3059,N_2904,N_2822);
nor U3060 (N_3060,N_2937,N_2940);
nor U3061 (N_3061,N_2968,N_2936);
nor U3062 (N_3062,N_2929,N_2975);
nand U3063 (N_3063,N_2935,N_2979);
nand U3064 (N_3064,N_2829,N_2997);
and U3065 (N_3065,N_2819,N_2949);
nand U3066 (N_3066,N_2912,N_2837);
nor U3067 (N_3067,N_2873,N_2890);
or U3068 (N_3068,N_2804,N_2800);
or U3069 (N_3069,N_2883,N_2961);
nand U3070 (N_3070,N_2852,N_2851);
or U3071 (N_3071,N_2906,N_2836);
and U3072 (N_3072,N_2815,N_2918);
and U3073 (N_3073,N_2806,N_2821);
or U3074 (N_3074,N_2816,N_2861);
nor U3075 (N_3075,N_2865,N_2921);
nand U3076 (N_3076,N_2828,N_2948);
or U3077 (N_3077,N_2915,N_2962);
nand U3078 (N_3078,N_2956,N_2955);
or U3079 (N_3079,N_2807,N_2838);
or U3080 (N_3080,N_2808,N_2934);
nor U3081 (N_3081,N_2914,N_2854);
nand U3082 (N_3082,N_2891,N_2990);
nor U3083 (N_3083,N_2999,N_2902);
nor U3084 (N_3084,N_2907,N_2826);
nor U3085 (N_3085,N_2824,N_2841);
or U3086 (N_3086,N_2980,N_2855);
and U3087 (N_3087,N_2867,N_2985);
or U3088 (N_3088,N_2933,N_2892);
nand U3089 (N_3089,N_2959,N_2810);
and U3090 (N_3090,N_2905,N_2941);
or U3091 (N_3091,N_2895,N_2848);
nand U3092 (N_3092,N_2983,N_2988);
nor U3093 (N_3093,N_2871,N_2846);
nor U3094 (N_3094,N_2805,N_2953);
nor U3095 (N_3095,N_2903,N_2827);
nand U3096 (N_3096,N_2909,N_2998);
and U3097 (N_3097,N_2856,N_2950);
and U3098 (N_3098,N_2926,N_2898);
nand U3099 (N_3099,N_2973,N_2802);
and U3100 (N_3100,N_2930,N_2974);
and U3101 (N_3101,N_2999,N_2822);
and U3102 (N_3102,N_2950,N_2998);
and U3103 (N_3103,N_2830,N_2859);
and U3104 (N_3104,N_2934,N_2896);
xor U3105 (N_3105,N_2978,N_2803);
nand U3106 (N_3106,N_2961,N_2948);
or U3107 (N_3107,N_2835,N_2947);
nor U3108 (N_3108,N_2808,N_2954);
nand U3109 (N_3109,N_2856,N_2978);
nor U3110 (N_3110,N_2966,N_2850);
and U3111 (N_3111,N_2840,N_2868);
or U3112 (N_3112,N_2992,N_2845);
nand U3113 (N_3113,N_2902,N_2992);
or U3114 (N_3114,N_2861,N_2879);
or U3115 (N_3115,N_2825,N_2877);
xnor U3116 (N_3116,N_2869,N_2920);
nand U3117 (N_3117,N_2964,N_2902);
nand U3118 (N_3118,N_2850,N_2979);
nand U3119 (N_3119,N_2964,N_2859);
and U3120 (N_3120,N_2888,N_2869);
or U3121 (N_3121,N_2851,N_2822);
nor U3122 (N_3122,N_2984,N_2876);
nor U3123 (N_3123,N_2810,N_2981);
nand U3124 (N_3124,N_2881,N_2972);
nand U3125 (N_3125,N_2926,N_2999);
or U3126 (N_3126,N_2922,N_2873);
and U3127 (N_3127,N_2954,N_2899);
and U3128 (N_3128,N_2882,N_2995);
nand U3129 (N_3129,N_2807,N_2884);
or U3130 (N_3130,N_2820,N_2885);
nor U3131 (N_3131,N_2852,N_2992);
nor U3132 (N_3132,N_2958,N_2881);
nor U3133 (N_3133,N_2949,N_2897);
or U3134 (N_3134,N_2968,N_2978);
and U3135 (N_3135,N_2895,N_2990);
nor U3136 (N_3136,N_2889,N_2911);
nor U3137 (N_3137,N_2919,N_2951);
nor U3138 (N_3138,N_2823,N_2894);
nor U3139 (N_3139,N_2885,N_2981);
nor U3140 (N_3140,N_2980,N_2880);
and U3141 (N_3141,N_2900,N_2891);
nor U3142 (N_3142,N_2901,N_2938);
nor U3143 (N_3143,N_2818,N_2931);
nand U3144 (N_3144,N_2849,N_2916);
xor U3145 (N_3145,N_2932,N_2902);
nor U3146 (N_3146,N_2932,N_2900);
and U3147 (N_3147,N_2866,N_2963);
nand U3148 (N_3148,N_2945,N_2863);
nor U3149 (N_3149,N_2986,N_2990);
or U3150 (N_3150,N_2823,N_2879);
and U3151 (N_3151,N_2929,N_2802);
or U3152 (N_3152,N_2825,N_2981);
or U3153 (N_3153,N_2805,N_2800);
or U3154 (N_3154,N_2855,N_2898);
and U3155 (N_3155,N_2988,N_2845);
nand U3156 (N_3156,N_2813,N_2881);
nand U3157 (N_3157,N_2972,N_2840);
or U3158 (N_3158,N_2856,N_2893);
nor U3159 (N_3159,N_2964,N_2868);
nor U3160 (N_3160,N_2954,N_2889);
or U3161 (N_3161,N_2802,N_2874);
or U3162 (N_3162,N_2881,N_2932);
and U3163 (N_3163,N_2914,N_2807);
and U3164 (N_3164,N_2823,N_2931);
or U3165 (N_3165,N_2971,N_2804);
nor U3166 (N_3166,N_2953,N_2973);
nand U3167 (N_3167,N_2906,N_2844);
nor U3168 (N_3168,N_2971,N_2845);
and U3169 (N_3169,N_2971,N_2974);
nand U3170 (N_3170,N_2866,N_2919);
nand U3171 (N_3171,N_2804,N_2895);
nand U3172 (N_3172,N_2971,N_2967);
nor U3173 (N_3173,N_2839,N_2804);
nand U3174 (N_3174,N_2846,N_2994);
or U3175 (N_3175,N_2902,N_2986);
nand U3176 (N_3176,N_2869,N_2985);
or U3177 (N_3177,N_2867,N_2997);
or U3178 (N_3178,N_2937,N_2870);
and U3179 (N_3179,N_2987,N_2995);
or U3180 (N_3180,N_2916,N_2911);
nor U3181 (N_3181,N_2831,N_2983);
or U3182 (N_3182,N_2975,N_2847);
and U3183 (N_3183,N_2912,N_2967);
and U3184 (N_3184,N_2827,N_2802);
and U3185 (N_3185,N_2950,N_2844);
nor U3186 (N_3186,N_2968,N_2851);
nor U3187 (N_3187,N_2840,N_2879);
or U3188 (N_3188,N_2919,N_2897);
and U3189 (N_3189,N_2862,N_2912);
or U3190 (N_3190,N_2897,N_2987);
and U3191 (N_3191,N_2812,N_2901);
nand U3192 (N_3192,N_2833,N_2964);
and U3193 (N_3193,N_2823,N_2968);
or U3194 (N_3194,N_2966,N_2881);
or U3195 (N_3195,N_2923,N_2888);
nand U3196 (N_3196,N_2829,N_2956);
nand U3197 (N_3197,N_2828,N_2830);
nor U3198 (N_3198,N_2882,N_2936);
or U3199 (N_3199,N_2811,N_2826);
nand U3200 (N_3200,N_3179,N_3110);
nor U3201 (N_3201,N_3007,N_3128);
nor U3202 (N_3202,N_3061,N_3038);
nor U3203 (N_3203,N_3191,N_3084);
nor U3204 (N_3204,N_3127,N_3171);
nor U3205 (N_3205,N_3169,N_3013);
or U3206 (N_3206,N_3103,N_3176);
and U3207 (N_3207,N_3075,N_3139);
nand U3208 (N_3208,N_3014,N_3121);
or U3209 (N_3209,N_3035,N_3122);
and U3210 (N_3210,N_3158,N_3147);
nor U3211 (N_3211,N_3159,N_3184);
and U3212 (N_3212,N_3046,N_3093);
and U3213 (N_3213,N_3145,N_3140);
or U3214 (N_3214,N_3117,N_3064);
or U3215 (N_3215,N_3006,N_3153);
nand U3216 (N_3216,N_3107,N_3030);
or U3217 (N_3217,N_3050,N_3009);
or U3218 (N_3218,N_3119,N_3194);
and U3219 (N_3219,N_3090,N_3073);
nand U3220 (N_3220,N_3005,N_3161);
nor U3221 (N_3221,N_3181,N_3144);
and U3222 (N_3222,N_3018,N_3183);
nand U3223 (N_3223,N_3077,N_3146);
and U3224 (N_3224,N_3136,N_3026);
nand U3225 (N_3225,N_3059,N_3199);
or U3226 (N_3226,N_3097,N_3137);
and U3227 (N_3227,N_3094,N_3164);
or U3228 (N_3228,N_3126,N_3174);
and U3229 (N_3229,N_3133,N_3045);
or U3230 (N_3230,N_3081,N_3180);
nand U3231 (N_3231,N_3079,N_3108);
and U3232 (N_3232,N_3098,N_3125);
or U3233 (N_3233,N_3172,N_3095);
or U3234 (N_3234,N_3010,N_3091);
nand U3235 (N_3235,N_3196,N_3019);
and U3236 (N_3236,N_3056,N_3032);
and U3237 (N_3237,N_3142,N_3027);
nand U3238 (N_3238,N_3085,N_3012);
or U3239 (N_3239,N_3175,N_3148);
or U3240 (N_3240,N_3155,N_3023);
and U3241 (N_3241,N_3082,N_3021);
nor U3242 (N_3242,N_3020,N_3182);
nor U3243 (N_3243,N_3000,N_3074);
and U3244 (N_3244,N_3157,N_3165);
or U3245 (N_3245,N_3063,N_3105);
and U3246 (N_3246,N_3055,N_3186);
nand U3247 (N_3247,N_3067,N_3120);
nand U3248 (N_3248,N_3188,N_3129);
or U3249 (N_3249,N_3192,N_3187);
and U3250 (N_3250,N_3034,N_3111);
nor U3251 (N_3251,N_3170,N_3015);
and U3252 (N_3252,N_3162,N_3124);
nand U3253 (N_3253,N_3160,N_3022);
or U3254 (N_3254,N_3195,N_3143);
and U3255 (N_3255,N_3053,N_3069);
and U3256 (N_3256,N_3189,N_3011);
nor U3257 (N_3257,N_3047,N_3101);
or U3258 (N_3258,N_3154,N_3112);
or U3259 (N_3259,N_3193,N_3100);
nor U3260 (N_3260,N_3113,N_3151);
or U3261 (N_3261,N_3123,N_3138);
nand U3262 (N_3262,N_3198,N_3062);
and U3263 (N_3263,N_3092,N_3163);
nor U3264 (N_3264,N_3068,N_3166);
nand U3265 (N_3265,N_3025,N_3118);
nand U3266 (N_3266,N_3043,N_3116);
nor U3267 (N_3267,N_3049,N_3044);
and U3268 (N_3268,N_3099,N_3054);
and U3269 (N_3269,N_3048,N_3152);
nand U3270 (N_3270,N_3060,N_3173);
or U3271 (N_3271,N_3185,N_3040);
nand U3272 (N_3272,N_3150,N_3130);
and U3273 (N_3273,N_3168,N_3135);
nand U3274 (N_3274,N_3037,N_3096);
nor U3275 (N_3275,N_3033,N_3070);
nor U3276 (N_3276,N_3076,N_3104);
and U3277 (N_3277,N_3149,N_3102);
nor U3278 (N_3278,N_3106,N_3134);
nand U3279 (N_3279,N_3083,N_3008);
or U3280 (N_3280,N_3024,N_3028);
or U3281 (N_3281,N_3039,N_3190);
and U3282 (N_3282,N_3078,N_3058);
and U3283 (N_3283,N_3042,N_3080);
and U3284 (N_3284,N_3052,N_3001);
and U3285 (N_3285,N_3002,N_3072);
or U3286 (N_3286,N_3004,N_3088);
or U3287 (N_3287,N_3041,N_3086);
or U3288 (N_3288,N_3089,N_3036);
or U3289 (N_3289,N_3114,N_3017);
or U3290 (N_3290,N_3197,N_3131);
nand U3291 (N_3291,N_3178,N_3167);
and U3292 (N_3292,N_3029,N_3016);
nand U3293 (N_3293,N_3057,N_3132);
and U3294 (N_3294,N_3109,N_3141);
or U3295 (N_3295,N_3115,N_3003);
nor U3296 (N_3296,N_3065,N_3156);
and U3297 (N_3297,N_3177,N_3031);
and U3298 (N_3298,N_3087,N_3066);
nor U3299 (N_3299,N_3051,N_3071);
or U3300 (N_3300,N_3158,N_3122);
or U3301 (N_3301,N_3178,N_3044);
nand U3302 (N_3302,N_3142,N_3028);
nand U3303 (N_3303,N_3097,N_3065);
nand U3304 (N_3304,N_3156,N_3068);
nor U3305 (N_3305,N_3010,N_3041);
nand U3306 (N_3306,N_3048,N_3192);
nand U3307 (N_3307,N_3155,N_3001);
and U3308 (N_3308,N_3156,N_3015);
nand U3309 (N_3309,N_3085,N_3017);
and U3310 (N_3310,N_3048,N_3063);
or U3311 (N_3311,N_3153,N_3146);
nor U3312 (N_3312,N_3034,N_3050);
nand U3313 (N_3313,N_3174,N_3032);
nand U3314 (N_3314,N_3004,N_3197);
or U3315 (N_3315,N_3122,N_3172);
nor U3316 (N_3316,N_3090,N_3078);
and U3317 (N_3317,N_3132,N_3156);
nand U3318 (N_3318,N_3028,N_3053);
or U3319 (N_3319,N_3195,N_3012);
nand U3320 (N_3320,N_3014,N_3132);
nor U3321 (N_3321,N_3009,N_3099);
nor U3322 (N_3322,N_3084,N_3073);
nor U3323 (N_3323,N_3153,N_3111);
nand U3324 (N_3324,N_3153,N_3079);
nor U3325 (N_3325,N_3196,N_3047);
nand U3326 (N_3326,N_3083,N_3134);
nor U3327 (N_3327,N_3183,N_3058);
or U3328 (N_3328,N_3094,N_3112);
and U3329 (N_3329,N_3177,N_3062);
and U3330 (N_3330,N_3190,N_3138);
and U3331 (N_3331,N_3139,N_3199);
or U3332 (N_3332,N_3009,N_3057);
nor U3333 (N_3333,N_3145,N_3177);
nand U3334 (N_3334,N_3164,N_3079);
and U3335 (N_3335,N_3022,N_3111);
nand U3336 (N_3336,N_3164,N_3168);
nand U3337 (N_3337,N_3049,N_3021);
and U3338 (N_3338,N_3132,N_3127);
nand U3339 (N_3339,N_3190,N_3045);
and U3340 (N_3340,N_3134,N_3088);
or U3341 (N_3341,N_3142,N_3183);
xnor U3342 (N_3342,N_3119,N_3000);
xnor U3343 (N_3343,N_3196,N_3005);
nor U3344 (N_3344,N_3131,N_3090);
nand U3345 (N_3345,N_3098,N_3075);
and U3346 (N_3346,N_3113,N_3072);
or U3347 (N_3347,N_3192,N_3160);
or U3348 (N_3348,N_3123,N_3172);
and U3349 (N_3349,N_3155,N_3018);
or U3350 (N_3350,N_3037,N_3030);
nand U3351 (N_3351,N_3121,N_3027);
nor U3352 (N_3352,N_3131,N_3024);
nor U3353 (N_3353,N_3002,N_3188);
nor U3354 (N_3354,N_3025,N_3099);
or U3355 (N_3355,N_3198,N_3166);
nor U3356 (N_3356,N_3120,N_3146);
or U3357 (N_3357,N_3185,N_3028);
or U3358 (N_3358,N_3084,N_3087);
or U3359 (N_3359,N_3165,N_3004);
nand U3360 (N_3360,N_3178,N_3091);
nand U3361 (N_3361,N_3034,N_3174);
nand U3362 (N_3362,N_3168,N_3009);
nor U3363 (N_3363,N_3081,N_3055);
nand U3364 (N_3364,N_3083,N_3165);
nand U3365 (N_3365,N_3168,N_3084);
or U3366 (N_3366,N_3161,N_3165);
nand U3367 (N_3367,N_3193,N_3051);
nand U3368 (N_3368,N_3059,N_3052);
nand U3369 (N_3369,N_3031,N_3139);
nand U3370 (N_3370,N_3099,N_3036);
or U3371 (N_3371,N_3122,N_3197);
or U3372 (N_3372,N_3088,N_3075);
nor U3373 (N_3373,N_3041,N_3196);
or U3374 (N_3374,N_3194,N_3059);
or U3375 (N_3375,N_3122,N_3097);
and U3376 (N_3376,N_3162,N_3138);
nand U3377 (N_3377,N_3152,N_3181);
or U3378 (N_3378,N_3103,N_3158);
and U3379 (N_3379,N_3060,N_3093);
or U3380 (N_3380,N_3039,N_3154);
and U3381 (N_3381,N_3066,N_3070);
nand U3382 (N_3382,N_3076,N_3152);
nor U3383 (N_3383,N_3137,N_3068);
nor U3384 (N_3384,N_3006,N_3111);
nor U3385 (N_3385,N_3169,N_3177);
nor U3386 (N_3386,N_3115,N_3067);
or U3387 (N_3387,N_3059,N_3007);
nand U3388 (N_3388,N_3009,N_3162);
nand U3389 (N_3389,N_3106,N_3005);
and U3390 (N_3390,N_3081,N_3157);
and U3391 (N_3391,N_3026,N_3020);
and U3392 (N_3392,N_3149,N_3052);
or U3393 (N_3393,N_3137,N_3169);
or U3394 (N_3394,N_3155,N_3060);
nand U3395 (N_3395,N_3129,N_3039);
nand U3396 (N_3396,N_3072,N_3064);
nand U3397 (N_3397,N_3043,N_3047);
and U3398 (N_3398,N_3035,N_3051);
and U3399 (N_3399,N_3137,N_3129);
or U3400 (N_3400,N_3247,N_3233);
nor U3401 (N_3401,N_3265,N_3367);
or U3402 (N_3402,N_3364,N_3237);
and U3403 (N_3403,N_3375,N_3399);
nor U3404 (N_3404,N_3266,N_3281);
nor U3405 (N_3405,N_3303,N_3395);
nor U3406 (N_3406,N_3398,N_3294);
or U3407 (N_3407,N_3396,N_3338);
nor U3408 (N_3408,N_3336,N_3278);
nor U3409 (N_3409,N_3334,N_3390);
nand U3410 (N_3410,N_3355,N_3275);
or U3411 (N_3411,N_3296,N_3304);
nand U3412 (N_3412,N_3345,N_3330);
nand U3413 (N_3413,N_3246,N_3222);
or U3414 (N_3414,N_3309,N_3202);
xor U3415 (N_3415,N_3212,N_3220);
and U3416 (N_3416,N_3308,N_3332);
nand U3417 (N_3417,N_3259,N_3239);
or U3418 (N_3418,N_3290,N_3201);
and U3419 (N_3419,N_3317,N_3384);
and U3420 (N_3420,N_3350,N_3370);
or U3421 (N_3421,N_3279,N_3238);
and U3422 (N_3422,N_3274,N_3319);
nor U3423 (N_3423,N_3357,N_3366);
nand U3424 (N_3424,N_3219,N_3272);
or U3425 (N_3425,N_3335,N_3223);
and U3426 (N_3426,N_3292,N_3311);
and U3427 (N_3427,N_3245,N_3268);
nand U3428 (N_3428,N_3287,N_3363);
or U3429 (N_3429,N_3249,N_3273);
nand U3430 (N_3430,N_3374,N_3283);
and U3431 (N_3431,N_3313,N_3295);
nand U3432 (N_3432,N_3230,N_3228);
or U3433 (N_3433,N_3288,N_3326);
nand U3434 (N_3434,N_3381,N_3299);
or U3435 (N_3435,N_3214,N_3280);
nand U3436 (N_3436,N_3235,N_3277);
nand U3437 (N_3437,N_3234,N_3379);
nor U3438 (N_3438,N_3221,N_3389);
nor U3439 (N_3439,N_3354,N_3373);
nor U3440 (N_3440,N_3253,N_3276);
nor U3441 (N_3441,N_3205,N_3376);
or U3442 (N_3442,N_3300,N_3206);
and U3443 (N_3443,N_3263,N_3397);
nand U3444 (N_3444,N_3252,N_3359);
and U3445 (N_3445,N_3227,N_3209);
or U3446 (N_3446,N_3318,N_3360);
nor U3447 (N_3447,N_3341,N_3371);
xor U3448 (N_3448,N_3226,N_3346);
nand U3449 (N_3449,N_3358,N_3255);
and U3450 (N_3450,N_3314,N_3307);
nor U3451 (N_3451,N_3322,N_3385);
nand U3452 (N_3452,N_3215,N_3306);
or U3453 (N_3453,N_3264,N_3333);
or U3454 (N_3454,N_3380,N_3285);
nand U3455 (N_3455,N_3327,N_3337);
or U3456 (N_3456,N_3340,N_3394);
nor U3457 (N_3457,N_3291,N_3297);
nand U3458 (N_3458,N_3231,N_3353);
and U3459 (N_3459,N_3267,N_3232);
and U3460 (N_3460,N_3260,N_3254);
nor U3461 (N_3461,N_3388,N_3325);
or U3462 (N_3462,N_3352,N_3282);
or U3463 (N_3463,N_3286,N_3207);
nor U3464 (N_3464,N_3269,N_3216);
nor U3465 (N_3465,N_3236,N_3356);
and U3466 (N_3466,N_3344,N_3377);
nand U3467 (N_3467,N_3250,N_3368);
and U3468 (N_3468,N_3293,N_3200);
or U3469 (N_3469,N_3323,N_3315);
or U3470 (N_3470,N_3392,N_3244);
nor U3471 (N_3471,N_3347,N_3270);
nor U3472 (N_3472,N_3316,N_3203);
nor U3473 (N_3473,N_3218,N_3372);
or U3474 (N_3474,N_3258,N_3331);
and U3475 (N_3475,N_3284,N_3298);
and U3476 (N_3476,N_3210,N_3256);
and U3477 (N_3477,N_3208,N_3378);
and U3478 (N_3478,N_3301,N_3217);
nor U3479 (N_3479,N_3349,N_3362);
nand U3480 (N_3480,N_3324,N_3391);
nand U3481 (N_3481,N_3312,N_3224);
or U3482 (N_3482,N_3302,N_3289);
and U3483 (N_3483,N_3211,N_3251);
nor U3484 (N_3484,N_3339,N_3242);
and U3485 (N_3485,N_3310,N_3342);
nor U3486 (N_3486,N_3348,N_3393);
nor U3487 (N_3487,N_3361,N_3321);
and U3488 (N_3488,N_3261,N_3365);
nor U3489 (N_3489,N_3241,N_3240);
and U3490 (N_3490,N_3225,N_3213);
nor U3491 (N_3491,N_3271,N_3387);
or U3492 (N_3492,N_3382,N_3328);
or U3493 (N_3493,N_3369,N_3229);
and U3494 (N_3494,N_3243,N_3386);
or U3495 (N_3495,N_3329,N_3305);
nand U3496 (N_3496,N_3257,N_3248);
and U3497 (N_3497,N_3383,N_3204);
nor U3498 (N_3498,N_3262,N_3343);
nand U3499 (N_3499,N_3351,N_3320);
and U3500 (N_3500,N_3278,N_3327);
and U3501 (N_3501,N_3320,N_3302);
nor U3502 (N_3502,N_3355,N_3362);
nand U3503 (N_3503,N_3331,N_3312);
nand U3504 (N_3504,N_3229,N_3342);
or U3505 (N_3505,N_3316,N_3347);
nor U3506 (N_3506,N_3307,N_3228);
and U3507 (N_3507,N_3259,N_3327);
nor U3508 (N_3508,N_3275,N_3253);
or U3509 (N_3509,N_3298,N_3387);
and U3510 (N_3510,N_3319,N_3383);
nand U3511 (N_3511,N_3267,N_3272);
and U3512 (N_3512,N_3399,N_3265);
nor U3513 (N_3513,N_3293,N_3319);
and U3514 (N_3514,N_3334,N_3233);
nand U3515 (N_3515,N_3347,N_3215);
nor U3516 (N_3516,N_3334,N_3345);
nor U3517 (N_3517,N_3208,N_3333);
and U3518 (N_3518,N_3310,N_3258);
or U3519 (N_3519,N_3267,N_3315);
nor U3520 (N_3520,N_3369,N_3213);
nor U3521 (N_3521,N_3274,N_3324);
nor U3522 (N_3522,N_3340,N_3290);
nor U3523 (N_3523,N_3301,N_3269);
nand U3524 (N_3524,N_3250,N_3202);
nor U3525 (N_3525,N_3249,N_3359);
nor U3526 (N_3526,N_3394,N_3207);
or U3527 (N_3527,N_3224,N_3215);
nor U3528 (N_3528,N_3334,N_3270);
nand U3529 (N_3529,N_3395,N_3218);
and U3530 (N_3530,N_3226,N_3265);
or U3531 (N_3531,N_3289,N_3311);
or U3532 (N_3532,N_3219,N_3236);
and U3533 (N_3533,N_3274,N_3286);
or U3534 (N_3534,N_3207,N_3247);
and U3535 (N_3535,N_3390,N_3257);
nand U3536 (N_3536,N_3256,N_3387);
or U3537 (N_3537,N_3321,N_3373);
and U3538 (N_3538,N_3200,N_3284);
nand U3539 (N_3539,N_3285,N_3210);
nor U3540 (N_3540,N_3322,N_3346);
nor U3541 (N_3541,N_3316,N_3253);
and U3542 (N_3542,N_3333,N_3275);
nand U3543 (N_3543,N_3288,N_3369);
nor U3544 (N_3544,N_3269,N_3297);
or U3545 (N_3545,N_3341,N_3377);
and U3546 (N_3546,N_3312,N_3359);
and U3547 (N_3547,N_3360,N_3366);
nand U3548 (N_3548,N_3371,N_3306);
or U3549 (N_3549,N_3202,N_3383);
nor U3550 (N_3550,N_3302,N_3379);
nor U3551 (N_3551,N_3239,N_3305);
nor U3552 (N_3552,N_3386,N_3367);
nor U3553 (N_3553,N_3299,N_3207);
and U3554 (N_3554,N_3370,N_3333);
nor U3555 (N_3555,N_3304,N_3316);
nor U3556 (N_3556,N_3260,N_3392);
and U3557 (N_3557,N_3229,N_3328);
nand U3558 (N_3558,N_3314,N_3299);
nor U3559 (N_3559,N_3336,N_3382);
or U3560 (N_3560,N_3347,N_3268);
or U3561 (N_3561,N_3355,N_3219);
and U3562 (N_3562,N_3364,N_3390);
and U3563 (N_3563,N_3299,N_3268);
or U3564 (N_3564,N_3225,N_3387);
or U3565 (N_3565,N_3235,N_3320);
and U3566 (N_3566,N_3329,N_3269);
and U3567 (N_3567,N_3205,N_3273);
or U3568 (N_3568,N_3225,N_3293);
or U3569 (N_3569,N_3236,N_3229);
nor U3570 (N_3570,N_3289,N_3201);
and U3571 (N_3571,N_3299,N_3352);
nand U3572 (N_3572,N_3360,N_3343);
and U3573 (N_3573,N_3386,N_3332);
or U3574 (N_3574,N_3208,N_3216);
and U3575 (N_3575,N_3286,N_3394);
or U3576 (N_3576,N_3295,N_3294);
xnor U3577 (N_3577,N_3343,N_3304);
and U3578 (N_3578,N_3350,N_3358);
nor U3579 (N_3579,N_3350,N_3300);
or U3580 (N_3580,N_3389,N_3373);
or U3581 (N_3581,N_3348,N_3225);
nand U3582 (N_3582,N_3308,N_3276);
nand U3583 (N_3583,N_3204,N_3309);
and U3584 (N_3584,N_3349,N_3345);
or U3585 (N_3585,N_3233,N_3326);
and U3586 (N_3586,N_3287,N_3397);
and U3587 (N_3587,N_3211,N_3210);
or U3588 (N_3588,N_3284,N_3249);
xor U3589 (N_3589,N_3394,N_3338);
and U3590 (N_3590,N_3308,N_3382);
or U3591 (N_3591,N_3252,N_3315);
nand U3592 (N_3592,N_3303,N_3226);
nand U3593 (N_3593,N_3379,N_3259);
and U3594 (N_3594,N_3227,N_3331);
or U3595 (N_3595,N_3333,N_3330);
nor U3596 (N_3596,N_3236,N_3383);
and U3597 (N_3597,N_3220,N_3255);
and U3598 (N_3598,N_3216,N_3354);
nor U3599 (N_3599,N_3374,N_3291);
or U3600 (N_3600,N_3558,N_3456);
or U3601 (N_3601,N_3448,N_3519);
and U3602 (N_3602,N_3518,N_3470);
nand U3603 (N_3603,N_3534,N_3503);
and U3604 (N_3604,N_3597,N_3572);
nand U3605 (N_3605,N_3552,N_3439);
nor U3606 (N_3606,N_3464,N_3514);
or U3607 (N_3607,N_3405,N_3563);
and U3608 (N_3608,N_3560,N_3400);
nand U3609 (N_3609,N_3447,N_3596);
and U3610 (N_3610,N_3494,N_3530);
nand U3611 (N_3611,N_3551,N_3504);
xnor U3612 (N_3612,N_3463,N_3495);
nand U3613 (N_3613,N_3580,N_3480);
nor U3614 (N_3614,N_3564,N_3491);
or U3615 (N_3615,N_3487,N_3543);
nand U3616 (N_3616,N_3542,N_3509);
nand U3617 (N_3617,N_3516,N_3481);
nor U3618 (N_3618,N_3550,N_3525);
and U3619 (N_3619,N_3513,N_3581);
or U3620 (N_3620,N_3546,N_3541);
nand U3621 (N_3621,N_3523,N_3576);
and U3622 (N_3622,N_3425,N_3469);
or U3623 (N_3623,N_3445,N_3512);
or U3624 (N_3624,N_3515,N_3562);
nand U3625 (N_3625,N_3402,N_3436);
nand U3626 (N_3626,N_3467,N_3593);
nand U3627 (N_3627,N_3529,N_3462);
and U3628 (N_3628,N_3461,N_3561);
nand U3629 (N_3629,N_3521,N_3422);
nand U3630 (N_3630,N_3549,N_3404);
nor U3631 (N_3631,N_3417,N_3585);
nor U3632 (N_3632,N_3424,N_3465);
or U3633 (N_3633,N_3511,N_3468);
and U3634 (N_3634,N_3486,N_3489);
or U3635 (N_3635,N_3432,N_3505);
or U3636 (N_3636,N_3472,N_3547);
and U3637 (N_3637,N_3440,N_3420);
nor U3638 (N_3638,N_3437,N_3450);
nand U3639 (N_3639,N_3459,N_3570);
or U3640 (N_3640,N_3508,N_3526);
or U3641 (N_3641,N_3449,N_3442);
nor U3642 (N_3642,N_3453,N_3497);
nand U3643 (N_3643,N_3455,N_3435);
nand U3644 (N_3644,N_3429,N_3446);
and U3645 (N_3645,N_3476,N_3531);
nor U3646 (N_3646,N_3433,N_3428);
or U3647 (N_3647,N_3595,N_3579);
and U3648 (N_3648,N_3507,N_3587);
nor U3649 (N_3649,N_3554,N_3522);
or U3650 (N_3650,N_3538,N_3427);
or U3651 (N_3651,N_3466,N_3548);
nand U3652 (N_3652,N_3568,N_3419);
nor U3653 (N_3653,N_3478,N_3520);
or U3654 (N_3654,N_3458,N_3413);
nand U3655 (N_3655,N_3575,N_3484);
or U3656 (N_3656,N_3599,N_3501);
nor U3657 (N_3657,N_3498,N_3475);
and U3658 (N_3658,N_3409,N_3567);
nor U3659 (N_3659,N_3532,N_3490);
nand U3660 (N_3660,N_3416,N_3407);
and U3661 (N_3661,N_3569,N_3408);
nor U3662 (N_3662,N_3479,N_3415);
nand U3663 (N_3663,N_3488,N_3438);
or U3664 (N_3664,N_3577,N_3499);
or U3665 (N_3665,N_3527,N_3582);
or U3666 (N_3666,N_3571,N_3540);
nor U3667 (N_3667,N_3443,N_3598);
or U3668 (N_3668,N_3403,N_3544);
nand U3669 (N_3669,N_3460,N_3477);
nand U3670 (N_3670,N_3586,N_3557);
and U3671 (N_3671,N_3457,N_3500);
nor U3672 (N_3672,N_3493,N_3583);
xnor U3673 (N_3673,N_3412,N_3553);
nand U3674 (N_3674,N_3533,N_3441);
nor U3675 (N_3675,N_3588,N_3545);
nor U3676 (N_3676,N_3535,N_3430);
and U3677 (N_3677,N_3485,N_3426);
or U3678 (N_3678,N_3506,N_3592);
or U3679 (N_3679,N_3474,N_3584);
or U3680 (N_3680,N_3517,N_3573);
or U3681 (N_3681,N_3473,N_3492);
or U3682 (N_3682,N_3483,N_3410);
or U3683 (N_3683,N_3471,N_3496);
nor U3684 (N_3684,N_3565,N_3556);
and U3685 (N_3685,N_3401,N_3418);
or U3686 (N_3686,N_3537,N_3539);
nor U3687 (N_3687,N_3559,N_3423);
nor U3688 (N_3688,N_3590,N_3536);
or U3689 (N_3689,N_3524,N_3482);
or U3690 (N_3690,N_3411,N_3566);
or U3691 (N_3691,N_3502,N_3444);
or U3692 (N_3692,N_3555,N_3578);
and U3693 (N_3693,N_3451,N_3454);
nand U3694 (N_3694,N_3594,N_3434);
nor U3695 (N_3695,N_3406,N_3589);
or U3696 (N_3696,N_3528,N_3452);
nand U3697 (N_3697,N_3421,N_3591);
nand U3698 (N_3698,N_3431,N_3510);
or U3699 (N_3699,N_3574,N_3414);
and U3700 (N_3700,N_3454,N_3435);
nor U3701 (N_3701,N_3559,N_3400);
nor U3702 (N_3702,N_3571,N_3535);
nand U3703 (N_3703,N_3597,N_3508);
nor U3704 (N_3704,N_3495,N_3404);
nor U3705 (N_3705,N_3452,N_3488);
or U3706 (N_3706,N_3413,N_3521);
nand U3707 (N_3707,N_3593,N_3473);
nor U3708 (N_3708,N_3401,N_3588);
and U3709 (N_3709,N_3528,N_3443);
nor U3710 (N_3710,N_3473,N_3509);
nand U3711 (N_3711,N_3405,N_3582);
or U3712 (N_3712,N_3575,N_3592);
or U3713 (N_3713,N_3443,N_3563);
nor U3714 (N_3714,N_3491,N_3524);
nor U3715 (N_3715,N_3464,N_3581);
nand U3716 (N_3716,N_3407,N_3589);
nand U3717 (N_3717,N_3532,N_3548);
or U3718 (N_3718,N_3515,N_3510);
or U3719 (N_3719,N_3496,N_3572);
nor U3720 (N_3720,N_3536,N_3453);
or U3721 (N_3721,N_3562,N_3510);
nand U3722 (N_3722,N_3497,N_3411);
and U3723 (N_3723,N_3521,N_3462);
nand U3724 (N_3724,N_3482,N_3588);
and U3725 (N_3725,N_3529,N_3404);
nand U3726 (N_3726,N_3584,N_3571);
nor U3727 (N_3727,N_3569,N_3570);
nor U3728 (N_3728,N_3544,N_3417);
or U3729 (N_3729,N_3548,N_3556);
nor U3730 (N_3730,N_3409,N_3543);
nand U3731 (N_3731,N_3571,N_3463);
or U3732 (N_3732,N_3514,N_3570);
nor U3733 (N_3733,N_3513,N_3436);
and U3734 (N_3734,N_3496,N_3487);
nor U3735 (N_3735,N_3405,N_3407);
and U3736 (N_3736,N_3598,N_3582);
and U3737 (N_3737,N_3500,N_3592);
or U3738 (N_3738,N_3564,N_3434);
and U3739 (N_3739,N_3444,N_3540);
or U3740 (N_3740,N_3431,N_3567);
or U3741 (N_3741,N_3438,N_3407);
xnor U3742 (N_3742,N_3537,N_3463);
or U3743 (N_3743,N_3503,N_3572);
or U3744 (N_3744,N_3426,N_3512);
nor U3745 (N_3745,N_3449,N_3493);
or U3746 (N_3746,N_3505,N_3458);
and U3747 (N_3747,N_3558,N_3479);
or U3748 (N_3748,N_3413,N_3533);
or U3749 (N_3749,N_3436,N_3568);
and U3750 (N_3750,N_3412,N_3406);
and U3751 (N_3751,N_3555,N_3410);
and U3752 (N_3752,N_3428,N_3578);
and U3753 (N_3753,N_3400,N_3404);
nor U3754 (N_3754,N_3550,N_3508);
nor U3755 (N_3755,N_3403,N_3591);
or U3756 (N_3756,N_3556,N_3540);
nand U3757 (N_3757,N_3531,N_3447);
nor U3758 (N_3758,N_3515,N_3434);
or U3759 (N_3759,N_3409,N_3538);
nand U3760 (N_3760,N_3501,N_3424);
nand U3761 (N_3761,N_3550,N_3457);
or U3762 (N_3762,N_3460,N_3465);
nor U3763 (N_3763,N_3593,N_3419);
and U3764 (N_3764,N_3593,N_3414);
and U3765 (N_3765,N_3424,N_3481);
or U3766 (N_3766,N_3598,N_3581);
nand U3767 (N_3767,N_3408,N_3418);
nand U3768 (N_3768,N_3521,N_3476);
or U3769 (N_3769,N_3470,N_3503);
or U3770 (N_3770,N_3590,N_3417);
nor U3771 (N_3771,N_3490,N_3488);
nand U3772 (N_3772,N_3485,N_3401);
or U3773 (N_3773,N_3599,N_3568);
nor U3774 (N_3774,N_3476,N_3427);
or U3775 (N_3775,N_3478,N_3418);
nor U3776 (N_3776,N_3597,N_3521);
or U3777 (N_3777,N_3431,N_3494);
nor U3778 (N_3778,N_3584,N_3555);
nand U3779 (N_3779,N_3521,N_3418);
nor U3780 (N_3780,N_3551,N_3427);
and U3781 (N_3781,N_3538,N_3578);
nand U3782 (N_3782,N_3504,N_3515);
nand U3783 (N_3783,N_3500,N_3488);
and U3784 (N_3784,N_3484,N_3565);
nand U3785 (N_3785,N_3545,N_3469);
and U3786 (N_3786,N_3499,N_3404);
and U3787 (N_3787,N_3446,N_3567);
nand U3788 (N_3788,N_3498,N_3471);
and U3789 (N_3789,N_3559,N_3461);
and U3790 (N_3790,N_3431,N_3558);
nand U3791 (N_3791,N_3523,N_3573);
and U3792 (N_3792,N_3584,N_3563);
nor U3793 (N_3793,N_3599,N_3571);
nand U3794 (N_3794,N_3425,N_3535);
and U3795 (N_3795,N_3458,N_3437);
or U3796 (N_3796,N_3582,N_3571);
or U3797 (N_3797,N_3598,N_3473);
or U3798 (N_3798,N_3557,N_3414);
and U3799 (N_3799,N_3536,N_3478);
nand U3800 (N_3800,N_3608,N_3727);
nand U3801 (N_3801,N_3784,N_3712);
and U3802 (N_3802,N_3769,N_3796);
nor U3803 (N_3803,N_3667,N_3650);
nor U3804 (N_3804,N_3674,N_3724);
and U3805 (N_3805,N_3654,N_3626);
or U3806 (N_3806,N_3640,N_3788);
nor U3807 (N_3807,N_3781,N_3718);
or U3808 (N_3808,N_3621,N_3719);
nor U3809 (N_3809,N_3678,N_3658);
and U3810 (N_3810,N_3692,N_3791);
nand U3811 (N_3811,N_3601,N_3761);
nor U3812 (N_3812,N_3703,N_3700);
and U3813 (N_3813,N_3680,N_3664);
and U3814 (N_3814,N_3662,N_3749);
or U3815 (N_3815,N_3641,N_3697);
or U3816 (N_3816,N_3715,N_3652);
nand U3817 (N_3817,N_3636,N_3647);
nor U3818 (N_3818,N_3631,N_3795);
nor U3819 (N_3819,N_3763,N_3698);
and U3820 (N_3820,N_3684,N_3695);
or U3821 (N_3821,N_3747,N_3670);
nand U3822 (N_3822,N_3794,N_3611);
or U3823 (N_3823,N_3775,N_3633);
and U3824 (N_3824,N_3661,N_3754);
or U3825 (N_3825,N_3606,N_3797);
nor U3826 (N_3826,N_3683,N_3771);
nand U3827 (N_3827,N_3786,N_3744);
and U3828 (N_3828,N_3701,N_3702);
nand U3829 (N_3829,N_3738,N_3714);
or U3830 (N_3830,N_3639,N_3688);
nor U3831 (N_3831,N_3753,N_3630);
and U3832 (N_3832,N_3665,N_3735);
nand U3833 (N_3833,N_3629,N_3799);
or U3834 (N_3834,N_3721,N_3765);
nor U3835 (N_3835,N_3634,N_3711);
nor U3836 (N_3836,N_3745,N_3774);
and U3837 (N_3837,N_3691,N_3779);
and U3838 (N_3838,N_3609,N_3699);
and U3839 (N_3839,N_3750,N_3676);
and U3840 (N_3840,N_3704,N_3655);
or U3841 (N_3841,N_3644,N_3717);
or U3842 (N_3842,N_3677,N_3748);
or U3843 (N_3843,N_3663,N_3635);
nand U3844 (N_3844,N_3778,N_3681);
nor U3845 (N_3845,N_3660,N_3758);
or U3846 (N_3846,N_3659,N_3798);
or U3847 (N_3847,N_3657,N_3739);
or U3848 (N_3848,N_3666,N_3615);
nand U3849 (N_3849,N_3736,N_3734);
nor U3850 (N_3850,N_3776,N_3642);
and U3851 (N_3851,N_3746,N_3730);
or U3852 (N_3852,N_3731,N_3725);
nor U3853 (N_3853,N_3637,N_3716);
or U3854 (N_3854,N_3645,N_3612);
nand U3855 (N_3855,N_3643,N_3679);
and U3856 (N_3856,N_3671,N_3624);
nor U3857 (N_3857,N_3696,N_3766);
nor U3858 (N_3858,N_3760,N_3751);
nand U3859 (N_3859,N_3782,N_3772);
or U3860 (N_3860,N_3607,N_3675);
nor U3861 (N_3861,N_3741,N_3618);
and U3862 (N_3862,N_3619,N_3785);
or U3863 (N_3863,N_3617,N_3705);
and U3864 (N_3864,N_3768,N_3669);
and U3865 (N_3865,N_3722,N_3729);
nor U3866 (N_3866,N_3602,N_3743);
and U3867 (N_3867,N_3689,N_3726);
nor U3868 (N_3868,N_3777,N_3780);
or U3869 (N_3869,N_3600,N_3756);
nand U3870 (N_3870,N_3686,N_3614);
or U3871 (N_3871,N_3653,N_3685);
or U3872 (N_3872,N_3604,N_3710);
nand U3873 (N_3873,N_3690,N_3787);
nor U3874 (N_3874,N_3628,N_3622);
and U3875 (N_3875,N_3733,N_3790);
and U3876 (N_3876,N_3732,N_3673);
nand U3877 (N_3877,N_3672,N_3737);
nand U3878 (N_3878,N_3759,N_3762);
nand U3879 (N_3879,N_3740,N_3755);
and U3880 (N_3880,N_3638,N_3783);
nor U3881 (N_3881,N_3651,N_3720);
nand U3882 (N_3882,N_3649,N_3728);
nor U3883 (N_3883,N_3632,N_3613);
or U3884 (N_3884,N_3767,N_3793);
nor U3885 (N_3885,N_3625,N_3707);
nand U3886 (N_3886,N_3656,N_3694);
and U3887 (N_3887,N_3742,N_3764);
or U3888 (N_3888,N_3693,N_3708);
nor U3889 (N_3889,N_3603,N_3616);
and U3890 (N_3890,N_3620,N_3623);
or U3891 (N_3891,N_3757,N_3709);
or U3892 (N_3892,N_3770,N_3792);
or U3893 (N_3893,N_3605,N_3773);
and U3894 (N_3894,N_3610,N_3706);
or U3895 (N_3895,N_3713,N_3682);
nand U3896 (N_3896,N_3646,N_3789);
nand U3897 (N_3897,N_3627,N_3752);
or U3898 (N_3898,N_3648,N_3723);
nand U3899 (N_3899,N_3687,N_3668);
or U3900 (N_3900,N_3752,N_3603);
nand U3901 (N_3901,N_3708,N_3614);
nand U3902 (N_3902,N_3682,N_3702);
nand U3903 (N_3903,N_3736,N_3781);
nand U3904 (N_3904,N_3601,N_3688);
and U3905 (N_3905,N_3620,N_3722);
or U3906 (N_3906,N_3682,N_3777);
nand U3907 (N_3907,N_3776,N_3797);
or U3908 (N_3908,N_3704,N_3625);
xnor U3909 (N_3909,N_3679,N_3692);
nor U3910 (N_3910,N_3664,N_3682);
or U3911 (N_3911,N_3622,N_3646);
and U3912 (N_3912,N_3778,N_3689);
and U3913 (N_3913,N_3647,N_3603);
nand U3914 (N_3914,N_3741,N_3743);
nand U3915 (N_3915,N_3777,N_3738);
nand U3916 (N_3916,N_3621,N_3645);
and U3917 (N_3917,N_3792,N_3674);
and U3918 (N_3918,N_3731,N_3601);
or U3919 (N_3919,N_3680,N_3616);
and U3920 (N_3920,N_3712,N_3700);
nor U3921 (N_3921,N_3737,N_3613);
or U3922 (N_3922,N_3608,N_3774);
and U3923 (N_3923,N_3721,N_3747);
nand U3924 (N_3924,N_3660,N_3653);
nor U3925 (N_3925,N_3710,N_3766);
or U3926 (N_3926,N_3634,N_3714);
nand U3927 (N_3927,N_3678,N_3691);
nor U3928 (N_3928,N_3696,N_3730);
and U3929 (N_3929,N_3625,N_3795);
or U3930 (N_3930,N_3730,N_3718);
or U3931 (N_3931,N_3713,N_3749);
or U3932 (N_3932,N_3765,N_3729);
or U3933 (N_3933,N_3647,N_3655);
and U3934 (N_3934,N_3736,N_3674);
and U3935 (N_3935,N_3796,N_3704);
nor U3936 (N_3936,N_3753,N_3710);
nand U3937 (N_3937,N_3617,N_3725);
and U3938 (N_3938,N_3735,N_3709);
or U3939 (N_3939,N_3741,N_3760);
and U3940 (N_3940,N_3613,N_3603);
and U3941 (N_3941,N_3713,N_3672);
and U3942 (N_3942,N_3648,N_3685);
or U3943 (N_3943,N_3642,N_3738);
or U3944 (N_3944,N_3798,N_3643);
nand U3945 (N_3945,N_3671,N_3678);
and U3946 (N_3946,N_3655,N_3703);
nand U3947 (N_3947,N_3653,N_3707);
or U3948 (N_3948,N_3759,N_3698);
and U3949 (N_3949,N_3642,N_3619);
nor U3950 (N_3950,N_3700,N_3739);
and U3951 (N_3951,N_3745,N_3686);
or U3952 (N_3952,N_3745,N_3645);
and U3953 (N_3953,N_3719,N_3625);
or U3954 (N_3954,N_3643,N_3783);
or U3955 (N_3955,N_3689,N_3743);
or U3956 (N_3956,N_3795,N_3655);
nand U3957 (N_3957,N_3607,N_3667);
nor U3958 (N_3958,N_3792,N_3799);
or U3959 (N_3959,N_3657,N_3682);
nor U3960 (N_3960,N_3728,N_3673);
nand U3961 (N_3961,N_3774,N_3712);
nand U3962 (N_3962,N_3736,N_3761);
or U3963 (N_3963,N_3688,N_3649);
or U3964 (N_3964,N_3777,N_3664);
nor U3965 (N_3965,N_3671,N_3737);
and U3966 (N_3966,N_3697,N_3606);
nor U3967 (N_3967,N_3700,N_3644);
and U3968 (N_3968,N_3729,N_3723);
nor U3969 (N_3969,N_3635,N_3657);
nand U3970 (N_3970,N_3714,N_3719);
and U3971 (N_3971,N_3783,N_3633);
and U3972 (N_3972,N_3684,N_3631);
nand U3973 (N_3973,N_3760,N_3792);
nor U3974 (N_3974,N_3784,N_3676);
nand U3975 (N_3975,N_3662,N_3796);
nor U3976 (N_3976,N_3741,N_3647);
and U3977 (N_3977,N_3705,N_3760);
nor U3978 (N_3978,N_3783,N_3722);
or U3979 (N_3979,N_3618,N_3795);
nand U3980 (N_3980,N_3794,N_3646);
nand U3981 (N_3981,N_3647,N_3607);
and U3982 (N_3982,N_3628,N_3777);
nor U3983 (N_3983,N_3705,N_3771);
nor U3984 (N_3984,N_3747,N_3644);
nand U3985 (N_3985,N_3625,N_3695);
or U3986 (N_3986,N_3610,N_3643);
and U3987 (N_3987,N_3601,N_3641);
nand U3988 (N_3988,N_3738,N_3711);
nor U3989 (N_3989,N_3749,N_3654);
and U3990 (N_3990,N_3792,N_3791);
or U3991 (N_3991,N_3682,N_3753);
nor U3992 (N_3992,N_3692,N_3788);
nor U3993 (N_3993,N_3641,N_3667);
or U3994 (N_3994,N_3722,N_3792);
nand U3995 (N_3995,N_3681,N_3679);
or U3996 (N_3996,N_3654,N_3774);
nand U3997 (N_3997,N_3782,N_3640);
and U3998 (N_3998,N_3651,N_3795);
or U3999 (N_3999,N_3795,N_3780);
and U4000 (N_4000,N_3986,N_3882);
nand U4001 (N_4001,N_3958,N_3800);
or U4002 (N_4002,N_3931,N_3850);
or U4003 (N_4003,N_3943,N_3859);
and U4004 (N_4004,N_3916,N_3938);
nand U4005 (N_4005,N_3904,N_3894);
nor U4006 (N_4006,N_3851,N_3948);
or U4007 (N_4007,N_3923,N_3997);
nor U4008 (N_4008,N_3906,N_3818);
and U4009 (N_4009,N_3987,N_3806);
and U4010 (N_4010,N_3813,N_3905);
and U4011 (N_4011,N_3954,N_3885);
and U4012 (N_4012,N_3982,N_3804);
nor U4013 (N_4013,N_3828,N_3893);
or U4014 (N_4014,N_3830,N_3929);
nand U4015 (N_4015,N_3815,N_3845);
nor U4016 (N_4016,N_3844,N_3953);
or U4017 (N_4017,N_3877,N_3913);
nand U4018 (N_4018,N_3952,N_3874);
or U4019 (N_4019,N_3937,N_3903);
nand U4020 (N_4020,N_3942,N_3846);
and U4021 (N_4021,N_3848,N_3915);
nand U4022 (N_4022,N_3865,N_3867);
nand U4023 (N_4023,N_3925,N_3901);
and U4024 (N_4024,N_3963,N_3852);
and U4025 (N_4025,N_3896,N_3898);
or U4026 (N_4026,N_3983,N_3989);
or U4027 (N_4027,N_3979,N_3817);
and U4028 (N_4028,N_3823,N_3808);
nor U4029 (N_4029,N_3847,N_3810);
xor U4030 (N_4030,N_3886,N_3928);
or U4031 (N_4031,N_3863,N_3957);
nor U4032 (N_4032,N_3837,N_3866);
nor U4033 (N_4033,N_3856,N_3889);
nand U4034 (N_4034,N_3926,N_3879);
nand U4035 (N_4035,N_3939,N_3861);
or U4036 (N_4036,N_3914,N_3843);
nor U4037 (N_4037,N_3908,N_3839);
nand U4038 (N_4038,N_3968,N_3860);
and U4039 (N_4039,N_3827,N_3940);
or U4040 (N_4040,N_3890,N_3842);
nand U4041 (N_4041,N_3835,N_3883);
or U4042 (N_4042,N_3973,N_3972);
nand U4043 (N_4043,N_3870,N_3961);
nor U4044 (N_4044,N_3871,N_3829);
and U4045 (N_4045,N_3966,N_3918);
and U4046 (N_4046,N_3819,N_3814);
or U4047 (N_4047,N_3977,N_3909);
or U4048 (N_4048,N_3930,N_3911);
or U4049 (N_4049,N_3801,N_3994);
nor U4050 (N_4050,N_3951,N_3821);
or U4051 (N_4051,N_3981,N_3920);
nor U4052 (N_4052,N_3872,N_3947);
and U4053 (N_4053,N_3964,N_3864);
and U4054 (N_4054,N_3807,N_3878);
nor U4055 (N_4055,N_3965,N_3812);
nor U4056 (N_4056,N_3857,N_3811);
and U4057 (N_4057,N_3962,N_3836);
and U4058 (N_4058,N_3975,N_3825);
and U4059 (N_4059,N_3891,N_3881);
and U4060 (N_4060,N_3824,N_3853);
or U4061 (N_4061,N_3955,N_3924);
nand U4062 (N_4062,N_3946,N_3945);
and U4063 (N_4063,N_3999,N_3831);
or U4064 (N_4064,N_3809,N_3996);
and U4065 (N_4065,N_3834,N_3970);
nor U4066 (N_4066,N_3956,N_3820);
or U4067 (N_4067,N_3949,N_3849);
and U4068 (N_4068,N_3900,N_3907);
and U4069 (N_4069,N_3935,N_3988);
or U4070 (N_4070,N_3910,N_3880);
and U4071 (N_4071,N_3895,N_3933);
nor U4072 (N_4072,N_3927,N_3822);
nand U4073 (N_4073,N_3934,N_3833);
or U4074 (N_4074,N_3993,N_3941);
and U4075 (N_4075,N_3816,N_3917);
and U4076 (N_4076,N_3932,N_3950);
or U4077 (N_4077,N_3984,N_3869);
nor U4078 (N_4078,N_3912,N_3803);
nor U4079 (N_4079,N_3921,N_3868);
and U4080 (N_4080,N_3974,N_3919);
and U4081 (N_4081,N_3832,N_3876);
nor U4082 (N_4082,N_3992,N_3838);
nor U4083 (N_4083,N_3855,N_3969);
nor U4084 (N_4084,N_3854,N_3902);
nor U4085 (N_4085,N_3805,N_3959);
or U4086 (N_4086,N_3960,N_3990);
nand U4087 (N_4087,N_3884,N_3840);
or U4088 (N_4088,N_3841,N_3995);
nor U4089 (N_4089,N_3887,N_3922);
nand U4090 (N_4090,N_3971,N_3998);
nor U4091 (N_4091,N_3978,N_3862);
nor U4092 (N_4092,N_3985,N_3826);
or U4093 (N_4093,N_3888,N_3991);
nand U4094 (N_4094,N_3899,N_3802);
or U4095 (N_4095,N_3892,N_3980);
nand U4096 (N_4096,N_3936,N_3873);
or U4097 (N_4097,N_3875,N_3897);
and U4098 (N_4098,N_3976,N_3858);
or U4099 (N_4099,N_3967,N_3944);
or U4100 (N_4100,N_3865,N_3827);
and U4101 (N_4101,N_3874,N_3839);
nor U4102 (N_4102,N_3938,N_3939);
and U4103 (N_4103,N_3851,N_3915);
and U4104 (N_4104,N_3973,N_3832);
and U4105 (N_4105,N_3842,N_3964);
or U4106 (N_4106,N_3886,N_3936);
and U4107 (N_4107,N_3899,N_3957);
or U4108 (N_4108,N_3940,N_3953);
or U4109 (N_4109,N_3918,N_3866);
or U4110 (N_4110,N_3937,N_3958);
nand U4111 (N_4111,N_3974,N_3936);
nand U4112 (N_4112,N_3981,N_3935);
nor U4113 (N_4113,N_3833,N_3987);
and U4114 (N_4114,N_3931,N_3972);
nand U4115 (N_4115,N_3884,N_3817);
nand U4116 (N_4116,N_3842,N_3936);
and U4117 (N_4117,N_3802,N_3848);
or U4118 (N_4118,N_3890,N_3987);
nand U4119 (N_4119,N_3803,N_3903);
nand U4120 (N_4120,N_3859,N_3954);
or U4121 (N_4121,N_3927,N_3903);
or U4122 (N_4122,N_3937,N_3851);
or U4123 (N_4123,N_3819,N_3988);
or U4124 (N_4124,N_3942,N_3879);
nand U4125 (N_4125,N_3832,N_3830);
and U4126 (N_4126,N_3826,N_3994);
nor U4127 (N_4127,N_3804,N_3857);
or U4128 (N_4128,N_3935,N_3857);
nor U4129 (N_4129,N_3842,N_3978);
nor U4130 (N_4130,N_3957,N_3810);
nand U4131 (N_4131,N_3963,N_3874);
or U4132 (N_4132,N_3985,N_3928);
and U4133 (N_4133,N_3897,N_3879);
xnor U4134 (N_4134,N_3838,N_3964);
nand U4135 (N_4135,N_3862,N_3801);
or U4136 (N_4136,N_3960,N_3998);
or U4137 (N_4137,N_3877,N_3982);
nor U4138 (N_4138,N_3869,N_3809);
nor U4139 (N_4139,N_3845,N_3862);
nand U4140 (N_4140,N_3803,N_3854);
and U4141 (N_4141,N_3802,N_3930);
and U4142 (N_4142,N_3971,N_3878);
and U4143 (N_4143,N_3839,N_3932);
nor U4144 (N_4144,N_3874,N_3943);
nor U4145 (N_4145,N_3942,N_3941);
and U4146 (N_4146,N_3809,N_3998);
nor U4147 (N_4147,N_3901,N_3959);
or U4148 (N_4148,N_3991,N_3919);
and U4149 (N_4149,N_3869,N_3944);
nand U4150 (N_4150,N_3937,N_3890);
or U4151 (N_4151,N_3874,N_3808);
and U4152 (N_4152,N_3932,N_3903);
nand U4153 (N_4153,N_3943,N_3837);
or U4154 (N_4154,N_3857,N_3945);
and U4155 (N_4155,N_3841,N_3844);
nand U4156 (N_4156,N_3812,N_3912);
nand U4157 (N_4157,N_3942,N_3865);
and U4158 (N_4158,N_3851,N_3959);
nor U4159 (N_4159,N_3878,N_3969);
nor U4160 (N_4160,N_3921,N_3860);
or U4161 (N_4161,N_3815,N_3802);
nor U4162 (N_4162,N_3862,N_3958);
and U4163 (N_4163,N_3950,N_3997);
and U4164 (N_4164,N_3849,N_3986);
nand U4165 (N_4165,N_3912,N_3996);
nor U4166 (N_4166,N_3887,N_3849);
nor U4167 (N_4167,N_3939,N_3964);
or U4168 (N_4168,N_3831,N_3982);
nor U4169 (N_4169,N_3860,N_3812);
nor U4170 (N_4170,N_3869,N_3980);
nor U4171 (N_4171,N_3958,N_3871);
nand U4172 (N_4172,N_3893,N_3960);
nor U4173 (N_4173,N_3915,N_3824);
or U4174 (N_4174,N_3987,N_3939);
nor U4175 (N_4175,N_3947,N_3815);
or U4176 (N_4176,N_3891,N_3929);
or U4177 (N_4177,N_3932,N_3870);
or U4178 (N_4178,N_3908,N_3837);
nand U4179 (N_4179,N_3919,N_3868);
or U4180 (N_4180,N_3808,N_3973);
or U4181 (N_4181,N_3827,N_3981);
nor U4182 (N_4182,N_3807,N_3963);
and U4183 (N_4183,N_3886,N_3841);
or U4184 (N_4184,N_3895,N_3943);
or U4185 (N_4185,N_3879,N_3881);
or U4186 (N_4186,N_3861,N_3904);
nor U4187 (N_4187,N_3989,N_3837);
nand U4188 (N_4188,N_3966,N_3993);
nand U4189 (N_4189,N_3847,N_3970);
and U4190 (N_4190,N_3993,N_3884);
or U4191 (N_4191,N_3835,N_3852);
nor U4192 (N_4192,N_3821,N_3830);
and U4193 (N_4193,N_3969,N_3909);
and U4194 (N_4194,N_3983,N_3893);
nor U4195 (N_4195,N_3991,N_3849);
and U4196 (N_4196,N_3910,N_3899);
nor U4197 (N_4197,N_3870,N_3931);
or U4198 (N_4198,N_3958,N_3910);
nand U4199 (N_4199,N_3864,N_3971);
nor U4200 (N_4200,N_4026,N_4099);
and U4201 (N_4201,N_4182,N_4161);
or U4202 (N_4202,N_4007,N_4109);
nand U4203 (N_4203,N_4148,N_4064);
or U4204 (N_4204,N_4005,N_4142);
or U4205 (N_4205,N_4153,N_4195);
or U4206 (N_4206,N_4016,N_4119);
nor U4207 (N_4207,N_4128,N_4145);
nand U4208 (N_4208,N_4107,N_4038);
xor U4209 (N_4209,N_4024,N_4097);
nand U4210 (N_4210,N_4150,N_4100);
nand U4211 (N_4211,N_4076,N_4091);
or U4212 (N_4212,N_4046,N_4037);
or U4213 (N_4213,N_4051,N_4065);
and U4214 (N_4214,N_4177,N_4066);
nand U4215 (N_4215,N_4055,N_4168);
nor U4216 (N_4216,N_4163,N_4179);
or U4217 (N_4217,N_4041,N_4090);
and U4218 (N_4218,N_4120,N_4196);
or U4219 (N_4219,N_4127,N_4030);
nor U4220 (N_4220,N_4158,N_4042);
nor U4221 (N_4221,N_4108,N_4075);
or U4222 (N_4222,N_4093,N_4040);
nor U4223 (N_4223,N_4193,N_4011);
nor U4224 (N_4224,N_4073,N_4146);
nand U4225 (N_4225,N_4085,N_4001);
and U4226 (N_4226,N_4126,N_4162);
nand U4227 (N_4227,N_4077,N_4124);
nand U4228 (N_4228,N_4106,N_4058);
or U4229 (N_4229,N_4169,N_4003);
and U4230 (N_4230,N_4172,N_4114);
or U4231 (N_4231,N_4014,N_4031);
nand U4232 (N_4232,N_4167,N_4134);
nor U4233 (N_4233,N_4000,N_4171);
and U4234 (N_4234,N_4082,N_4015);
nand U4235 (N_4235,N_4139,N_4012);
or U4236 (N_4236,N_4187,N_4068);
nand U4237 (N_4237,N_4101,N_4054);
or U4238 (N_4238,N_4079,N_4095);
nor U4239 (N_4239,N_4188,N_4165);
nor U4240 (N_4240,N_4141,N_4059);
nand U4241 (N_4241,N_4170,N_4063);
nor U4242 (N_4242,N_4049,N_4029);
or U4243 (N_4243,N_4071,N_4131);
nand U4244 (N_4244,N_4140,N_4133);
and U4245 (N_4245,N_4089,N_4019);
and U4246 (N_4246,N_4192,N_4098);
or U4247 (N_4247,N_4136,N_4034);
or U4248 (N_4248,N_4018,N_4023);
nand U4249 (N_4249,N_4080,N_4022);
nand U4250 (N_4250,N_4086,N_4118);
nor U4251 (N_4251,N_4190,N_4039);
nor U4252 (N_4252,N_4020,N_4044);
and U4253 (N_4253,N_4081,N_4074);
or U4254 (N_4254,N_4173,N_4102);
nor U4255 (N_4255,N_4137,N_4062);
nor U4256 (N_4256,N_4008,N_4027);
or U4257 (N_4257,N_4006,N_4194);
or U4258 (N_4258,N_4123,N_4184);
or U4259 (N_4259,N_4147,N_4160);
or U4260 (N_4260,N_4197,N_4151);
and U4261 (N_4261,N_4010,N_4047);
nand U4262 (N_4262,N_4186,N_4180);
or U4263 (N_4263,N_4094,N_4103);
nor U4264 (N_4264,N_4174,N_4116);
nor U4265 (N_4265,N_4189,N_4060);
nand U4266 (N_4266,N_4070,N_4112);
and U4267 (N_4267,N_4175,N_4154);
or U4268 (N_4268,N_4056,N_4152);
nand U4269 (N_4269,N_4155,N_4083);
or U4270 (N_4270,N_4105,N_4028);
or U4271 (N_4271,N_4032,N_4025);
and U4272 (N_4272,N_4166,N_4092);
or U4273 (N_4273,N_4087,N_4104);
nor U4274 (N_4274,N_4088,N_4185);
nand U4275 (N_4275,N_4069,N_4129);
nand U4276 (N_4276,N_4096,N_4143);
nor U4277 (N_4277,N_4004,N_4110);
or U4278 (N_4278,N_4009,N_4176);
and U4279 (N_4279,N_4157,N_4121);
and U4280 (N_4280,N_4117,N_4138);
nand U4281 (N_4281,N_4135,N_4199);
and U4282 (N_4282,N_4053,N_4130);
nor U4283 (N_4283,N_4159,N_4013);
or U4284 (N_4284,N_4078,N_4057);
or U4285 (N_4285,N_4191,N_4072);
nor U4286 (N_4286,N_4132,N_4061);
nand U4287 (N_4287,N_4178,N_4149);
nand U4288 (N_4288,N_4002,N_4045);
or U4289 (N_4289,N_4017,N_4052);
or U4290 (N_4290,N_4156,N_4084);
and U4291 (N_4291,N_4198,N_4144);
nand U4292 (N_4292,N_4181,N_4067);
nand U4293 (N_4293,N_4122,N_4033);
and U4294 (N_4294,N_4164,N_4021);
and U4295 (N_4295,N_4035,N_4048);
and U4296 (N_4296,N_4043,N_4050);
and U4297 (N_4297,N_4036,N_4111);
xnor U4298 (N_4298,N_4125,N_4115);
and U4299 (N_4299,N_4183,N_4113);
or U4300 (N_4300,N_4087,N_4189);
nand U4301 (N_4301,N_4084,N_4172);
or U4302 (N_4302,N_4017,N_4143);
or U4303 (N_4303,N_4115,N_4001);
xnor U4304 (N_4304,N_4040,N_4068);
and U4305 (N_4305,N_4161,N_4132);
and U4306 (N_4306,N_4176,N_4137);
or U4307 (N_4307,N_4178,N_4139);
nor U4308 (N_4308,N_4089,N_4107);
or U4309 (N_4309,N_4066,N_4193);
nor U4310 (N_4310,N_4124,N_4007);
and U4311 (N_4311,N_4051,N_4199);
nand U4312 (N_4312,N_4122,N_4119);
nand U4313 (N_4313,N_4168,N_4074);
nor U4314 (N_4314,N_4197,N_4110);
nor U4315 (N_4315,N_4149,N_4106);
and U4316 (N_4316,N_4021,N_4148);
and U4317 (N_4317,N_4195,N_4109);
nand U4318 (N_4318,N_4198,N_4061);
or U4319 (N_4319,N_4080,N_4144);
nand U4320 (N_4320,N_4134,N_4029);
nor U4321 (N_4321,N_4124,N_4010);
nand U4322 (N_4322,N_4083,N_4100);
nand U4323 (N_4323,N_4055,N_4005);
and U4324 (N_4324,N_4013,N_4118);
nand U4325 (N_4325,N_4057,N_4062);
or U4326 (N_4326,N_4009,N_4046);
nand U4327 (N_4327,N_4147,N_4170);
nor U4328 (N_4328,N_4182,N_4100);
or U4329 (N_4329,N_4082,N_4153);
nor U4330 (N_4330,N_4009,N_4179);
nor U4331 (N_4331,N_4088,N_4112);
nor U4332 (N_4332,N_4172,N_4170);
nand U4333 (N_4333,N_4176,N_4149);
nor U4334 (N_4334,N_4140,N_4012);
nand U4335 (N_4335,N_4022,N_4032);
and U4336 (N_4336,N_4091,N_4058);
nand U4337 (N_4337,N_4103,N_4184);
and U4338 (N_4338,N_4191,N_4046);
nand U4339 (N_4339,N_4136,N_4026);
nand U4340 (N_4340,N_4175,N_4177);
nand U4341 (N_4341,N_4195,N_4093);
nor U4342 (N_4342,N_4198,N_4173);
or U4343 (N_4343,N_4119,N_4041);
and U4344 (N_4344,N_4121,N_4008);
or U4345 (N_4345,N_4123,N_4135);
and U4346 (N_4346,N_4099,N_4157);
nor U4347 (N_4347,N_4160,N_4154);
or U4348 (N_4348,N_4014,N_4106);
nand U4349 (N_4349,N_4114,N_4188);
nand U4350 (N_4350,N_4013,N_4015);
nand U4351 (N_4351,N_4152,N_4141);
nor U4352 (N_4352,N_4012,N_4066);
and U4353 (N_4353,N_4119,N_4015);
nand U4354 (N_4354,N_4130,N_4043);
and U4355 (N_4355,N_4116,N_4070);
nand U4356 (N_4356,N_4025,N_4024);
nor U4357 (N_4357,N_4017,N_4098);
nor U4358 (N_4358,N_4020,N_4178);
and U4359 (N_4359,N_4002,N_4185);
and U4360 (N_4360,N_4093,N_4106);
nor U4361 (N_4361,N_4118,N_4089);
and U4362 (N_4362,N_4046,N_4126);
and U4363 (N_4363,N_4026,N_4015);
nor U4364 (N_4364,N_4035,N_4159);
or U4365 (N_4365,N_4127,N_4106);
nor U4366 (N_4366,N_4119,N_4077);
or U4367 (N_4367,N_4158,N_4057);
nand U4368 (N_4368,N_4033,N_4044);
or U4369 (N_4369,N_4016,N_4034);
nor U4370 (N_4370,N_4028,N_4123);
or U4371 (N_4371,N_4145,N_4180);
nand U4372 (N_4372,N_4164,N_4105);
and U4373 (N_4373,N_4037,N_4001);
or U4374 (N_4374,N_4085,N_4191);
nand U4375 (N_4375,N_4082,N_4062);
nor U4376 (N_4376,N_4168,N_4141);
nand U4377 (N_4377,N_4043,N_4196);
or U4378 (N_4378,N_4181,N_4008);
or U4379 (N_4379,N_4039,N_4156);
and U4380 (N_4380,N_4033,N_4109);
nor U4381 (N_4381,N_4098,N_4126);
nor U4382 (N_4382,N_4169,N_4149);
and U4383 (N_4383,N_4179,N_4055);
and U4384 (N_4384,N_4052,N_4055);
or U4385 (N_4385,N_4073,N_4074);
nor U4386 (N_4386,N_4098,N_4107);
nand U4387 (N_4387,N_4194,N_4009);
or U4388 (N_4388,N_4181,N_4195);
or U4389 (N_4389,N_4180,N_4160);
nor U4390 (N_4390,N_4067,N_4057);
nor U4391 (N_4391,N_4141,N_4058);
and U4392 (N_4392,N_4194,N_4162);
nor U4393 (N_4393,N_4093,N_4109);
or U4394 (N_4394,N_4188,N_4036);
and U4395 (N_4395,N_4152,N_4095);
nor U4396 (N_4396,N_4185,N_4100);
nor U4397 (N_4397,N_4068,N_4132);
nor U4398 (N_4398,N_4081,N_4103);
nand U4399 (N_4399,N_4164,N_4046);
nand U4400 (N_4400,N_4317,N_4326);
nand U4401 (N_4401,N_4340,N_4359);
nor U4402 (N_4402,N_4209,N_4235);
or U4403 (N_4403,N_4256,N_4299);
and U4404 (N_4404,N_4388,N_4384);
and U4405 (N_4405,N_4308,N_4271);
nand U4406 (N_4406,N_4239,N_4363);
nor U4407 (N_4407,N_4258,N_4306);
nand U4408 (N_4408,N_4369,N_4365);
and U4409 (N_4409,N_4204,N_4313);
nand U4410 (N_4410,N_4353,N_4349);
or U4411 (N_4411,N_4288,N_4249);
and U4412 (N_4412,N_4309,N_4356);
nor U4413 (N_4413,N_4337,N_4207);
or U4414 (N_4414,N_4240,N_4331);
or U4415 (N_4415,N_4364,N_4358);
and U4416 (N_4416,N_4279,N_4312);
and U4417 (N_4417,N_4243,N_4229);
nor U4418 (N_4418,N_4254,N_4233);
and U4419 (N_4419,N_4389,N_4341);
and U4420 (N_4420,N_4293,N_4302);
nor U4421 (N_4421,N_4371,N_4310);
and U4422 (N_4422,N_4325,N_4395);
nand U4423 (N_4423,N_4230,N_4355);
nand U4424 (N_4424,N_4231,N_4269);
nand U4425 (N_4425,N_4361,N_4321);
nor U4426 (N_4426,N_4390,N_4398);
nor U4427 (N_4427,N_4339,N_4290);
nand U4428 (N_4428,N_4200,N_4387);
or U4429 (N_4429,N_4266,N_4316);
nor U4430 (N_4430,N_4373,N_4304);
nor U4431 (N_4431,N_4203,N_4227);
or U4432 (N_4432,N_4228,N_4328);
or U4433 (N_4433,N_4296,N_4367);
and U4434 (N_4434,N_4292,N_4297);
and U4435 (N_4435,N_4260,N_4305);
and U4436 (N_4436,N_4255,N_4338);
nor U4437 (N_4437,N_4330,N_4345);
nor U4438 (N_4438,N_4307,N_4267);
nor U4439 (N_4439,N_4377,N_4357);
nand U4440 (N_4440,N_4242,N_4346);
or U4441 (N_4441,N_4270,N_4211);
xor U4442 (N_4442,N_4300,N_4327);
nor U4443 (N_4443,N_4393,N_4276);
and U4444 (N_4444,N_4343,N_4352);
and U4445 (N_4445,N_4298,N_4379);
nor U4446 (N_4446,N_4382,N_4237);
and U4447 (N_4447,N_4360,N_4392);
or U4448 (N_4448,N_4215,N_4381);
nor U4449 (N_4449,N_4324,N_4259);
nor U4450 (N_4450,N_4277,N_4265);
nor U4451 (N_4451,N_4287,N_4350);
nand U4452 (N_4452,N_4248,N_4375);
nand U4453 (N_4453,N_4333,N_4273);
nand U4454 (N_4454,N_4247,N_4354);
nor U4455 (N_4455,N_4391,N_4251);
and U4456 (N_4456,N_4222,N_4336);
and U4457 (N_4457,N_4286,N_4329);
nor U4458 (N_4458,N_4214,N_4234);
nand U4459 (N_4459,N_4383,N_4268);
nor U4460 (N_4460,N_4323,N_4362);
and U4461 (N_4461,N_4232,N_4280);
nor U4462 (N_4462,N_4201,N_4241);
and U4463 (N_4463,N_4319,N_4342);
and U4464 (N_4464,N_4244,N_4322);
and U4465 (N_4465,N_4295,N_4217);
nand U4466 (N_4466,N_4394,N_4399);
or U4467 (N_4467,N_4213,N_4219);
and U4468 (N_4468,N_4252,N_4368);
or U4469 (N_4469,N_4202,N_4210);
or U4470 (N_4470,N_4224,N_4278);
nor U4471 (N_4471,N_4283,N_4261);
or U4472 (N_4472,N_4397,N_4225);
nor U4473 (N_4473,N_4311,N_4263);
nor U4474 (N_4474,N_4386,N_4374);
and U4475 (N_4475,N_4246,N_4291);
nor U4476 (N_4476,N_4294,N_4245);
nor U4477 (N_4477,N_4218,N_4220);
nand U4478 (N_4478,N_4262,N_4285);
and U4479 (N_4479,N_4385,N_4275);
or U4480 (N_4480,N_4378,N_4257);
nand U4481 (N_4481,N_4335,N_4205);
nand U4482 (N_4482,N_4396,N_4303);
or U4483 (N_4483,N_4380,N_4250);
and U4484 (N_4484,N_4226,N_4376);
nand U4485 (N_4485,N_4264,N_4281);
and U4486 (N_4486,N_4348,N_4366);
nor U4487 (N_4487,N_4282,N_4253);
xnor U4488 (N_4488,N_4212,N_4216);
or U4489 (N_4489,N_4208,N_4274);
nand U4490 (N_4490,N_4272,N_4351);
nand U4491 (N_4491,N_4289,N_4370);
and U4492 (N_4492,N_4236,N_4372);
nor U4493 (N_4493,N_4301,N_4284);
nor U4494 (N_4494,N_4347,N_4315);
or U4495 (N_4495,N_4332,N_4344);
nor U4496 (N_4496,N_4320,N_4314);
nor U4497 (N_4497,N_4221,N_4206);
nor U4498 (N_4498,N_4334,N_4223);
xnor U4499 (N_4499,N_4318,N_4238);
nand U4500 (N_4500,N_4320,N_4275);
or U4501 (N_4501,N_4357,N_4248);
nand U4502 (N_4502,N_4293,N_4334);
nor U4503 (N_4503,N_4320,N_4356);
and U4504 (N_4504,N_4214,N_4352);
and U4505 (N_4505,N_4344,N_4312);
nand U4506 (N_4506,N_4262,N_4274);
or U4507 (N_4507,N_4379,N_4361);
xor U4508 (N_4508,N_4238,N_4234);
nand U4509 (N_4509,N_4234,N_4362);
and U4510 (N_4510,N_4279,N_4280);
and U4511 (N_4511,N_4337,N_4363);
nand U4512 (N_4512,N_4381,N_4318);
nand U4513 (N_4513,N_4367,N_4307);
nor U4514 (N_4514,N_4371,N_4220);
nand U4515 (N_4515,N_4385,N_4329);
or U4516 (N_4516,N_4392,N_4387);
and U4517 (N_4517,N_4242,N_4343);
nor U4518 (N_4518,N_4390,N_4203);
nand U4519 (N_4519,N_4213,N_4284);
nand U4520 (N_4520,N_4258,N_4234);
or U4521 (N_4521,N_4339,N_4243);
and U4522 (N_4522,N_4367,N_4274);
and U4523 (N_4523,N_4368,N_4212);
nor U4524 (N_4524,N_4267,N_4308);
nor U4525 (N_4525,N_4330,N_4395);
and U4526 (N_4526,N_4394,N_4343);
nand U4527 (N_4527,N_4351,N_4247);
nor U4528 (N_4528,N_4284,N_4274);
or U4529 (N_4529,N_4234,N_4206);
and U4530 (N_4530,N_4235,N_4230);
nand U4531 (N_4531,N_4301,N_4267);
nor U4532 (N_4532,N_4257,N_4277);
nor U4533 (N_4533,N_4332,N_4363);
or U4534 (N_4534,N_4344,N_4364);
nor U4535 (N_4535,N_4260,N_4295);
nand U4536 (N_4536,N_4386,N_4314);
or U4537 (N_4537,N_4268,N_4367);
nand U4538 (N_4538,N_4298,N_4246);
nor U4539 (N_4539,N_4257,N_4363);
and U4540 (N_4540,N_4292,N_4240);
and U4541 (N_4541,N_4347,N_4358);
and U4542 (N_4542,N_4386,N_4296);
or U4543 (N_4543,N_4255,N_4233);
and U4544 (N_4544,N_4252,N_4288);
nand U4545 (N_4545,N_4262,N_4303);
or U4546 (N_4546,N_4312,N_4320);
nand U4547 (N_4547,N_4289,N_4315);
or U4548 (N_4548,N_4221,N_4365);
nand U4549 (N_4549,N_4367,N_4238);
or U4550 (N_4550,N_4314,N_4214);
and U4551 (N_4551,N_4334,N_4355);
nand U4552 (N_4552,N_4391,N_4353);
nand U4553 (N_4553,N_4226,N_4375);
or U4554 (N_4554,N_4217,N_4274);
nor U4555 (N_4555,N_4296,N_4304);
or U4556 (N_4556,N_4202,N_4329);
or U4557 (N_4557,N_4345,N_4225);
and U4558 (N_4558,N_4222,N_4231);
and U4559 (N_4559,N_4229,N_4352);
or U4560 (N_4560,N_4388,N_4294);
nor U4561 (N_4561,N_4221,N_4237);
nor U4562 (N_4562,N_4265,N_4323);
or U4563 (N_4563,N_4258,N_4298);
nand U4564 (N_4564,N_4339,N_4395);
and U4565 (N_4565,N_4291,N_4275);
nor U4566 (N_4566,N_4375,N_4353);
and U4567 (N_4567,N_4377,N_4356);
nor U4568 (N_4568,N_4263,N_4366);
nand U4569 (N_4569,N_4360,N_4362);
nor U4570 (N_4570,N_4277,N_4319);
and U4571 (N_4571,N_4262,N_4221);
or U4572 (N_4572,N_4222,N_4351);
nand U4573 (N_4573,N_4201,N_4288);
and U4574 (N_4574,N_4370,N_4271);
and U4575 (N_4575,N_4311,N_4274);
and U4576 (N_4576,N_4285,N_4259);
or U4577 (N_4577,N_4275,N_4373);
or U4578 (N_4578,N_4250,N_4255);
or U4579 (N_4579,N_4340,N_4387);
xnor U4580 (N_4580,N_4332,N_4261);
and U4581 (N_4581,N_4219,N_4330);
nand U4582 (N_4582,N_4247,N_4212);
and U4583 (N_4583,N_4228,N_4249);
and U4584 (N_4584,N_4354,N_4217);
or U4585 (N_4585,N_4238,N_4288);
nand U4586 (N_4586,N_4388,N_4366);
nand U4587 (N_4587,N_4262,N_4337);
and U4588 (N_4588,N_4380,N_4211);
nor U4589 (N_4589,N_4284,N_4201);
or U4590 (N_4590,N_4333,N_4397);
nand U4591 (N_4591,N_4286,N_4379);
nor U4592 (N_4592,N_4316,N_4201);
or U4593 (N_4593,N_4367,N_4298);
nor U4594 (N_4594,N_4247,N_4265);
nor U4595 (N_4595,N_4239,N_4221);
nor U4596 (N_4596,N_4332,N_4209);
and U4597 (N_4597,N_4220,N_4299);
or U4598 (N_4598,N_4375,N_4292);
or U4599 (N_4599,N_4304,N_4397);
nand U4600 (N_4600,N_4571,N_4470);
nand U4601 (N_4601,N_4443,N_4459);
nor U4602 (N_4602,N_4475,N_4409);
nand U4603 (N_4603,N_4404,N_4442);
and U4604 (N_4604,N_4546,N_4584);
xor U4605 (N_4605,N_4501,N_4446);
and U4606 (N_4606,N_4563,N_4541);
nor U4607 (N_4607,N_4462,N_4424);
nor U4608 (N_4608,N_4453,N_4410);
nor U4609 (N_4609,N_4498,N_4489);
nor U4610 (N_4610,N_4492,N_4429);
nor U4611 (N_4611,N_4539,N_4529);
nand U4612 (N_4612,N_4469,N_4414);
or U4613 (N_4613,N_4569,N_4561);
nand U4614 (N_4614,N_4532,N_4454);
and U4615 (N_4615,N_4494,N_4436);
or U4616 (N_4616,N_4595,N_4576);
nor U4617 (N_4617,N_4435,N_4497);
or U4618 (N_4618,N_4438,N_4551);
nand U4619 (N_4619,N_4412,N_4553);
nand U4620 (N_4620,N_4420,N_4549);
nor U4621 (N_4621,N_4586,N_4554);
nor U4622 (N_4622,N_4568,N_4559);
or U4623 (N_4623,N_4510,N_4535);
nor U4624 (N_4624,N_4522,N_4540);
and U4625 (N_4625,N_4426,N_4480);
nor U4626 (N_4626,N_4573,N_4543);
nand U4627 (N_4627,N_4574,N_4450);
nand U4628 (N_4628,N_4428,N_4468);
or U4629 (N_4629,N_4548,N_4422);
nand U4630 (N_4630,N_4457,N_4523);
nor U4631 (N_4631,N_4467,N_4562);
and U4632 (N_4632,N_4486,N_4527);
or U4633 (N_4633,N_4403,N_4531);
or U4634 (N_4634,N_4484,N_4407);
nor U4635 (N_4635,N_4550,N_4525);
and U4636 (N_4636,N_4558,N_4476);
or U4637 (N_4637,N_4502,N_4417);
or U4638 (N_4638,N_4589,N_4472);
or U4639 (N_4639,N_4533,N_4594);
nor U4640 (N_4640,N_4405,N_4514);
and U4641 (N_4641,N_4499,N_4490);
or U4642 (N_4642,N_4534,N_4432);
or U4643 (N_4643,N_4597,N_4425);
nand U4644 (N_4644,N_4463,N_4590);
nand U4645 (N_4645,N_4505,N_4521);
nor U4646 (N_4646,N_4481,N_4465);
or U4647 (N_4647,N_4482,N_4439);
or U4648 (N_4648,N_4448,N_4579);
or U4649 (N_4649,N_4528,N_4455);
or U4650 (N_4650,N_4418,N_4560);
and U4651 (N_4651,N_4440,N_4449);
nor U4652 (N_4652,N_4513,N_4402);
nor U4653 (N_4653,N_4536,N_4466);
nand U4654 (N_4654,N_4542,N_4580);
nor U4655 (N_4655,N_4503,N_4473);
nand U4656 (N_4656,N_4508,N_4415);
or U4657 (N_4657,N_4427,N_4461);
nor U4658 (N_4658,N_4570,N_4413);
nand U4659 (N_4659,N_4488,N_4447);
nand U4660 (N_4660,N_4556,N_4566);
or U4661 (N_4661,N_4477,N_4416);
and U4662 (N_4662,N_4408,N_4441);
and U4663 (N_4663,N_4591,N_4419);
and U4664 (N_4664,N_4524,N_4575);
nand U4665 (N_4665,N_4504,N_4509);
or U4666 (N_4666,N_4452,N_4496);
and U4667 (N_4667,N_4592,N_4507);
or U4668 (N_4668,N_4406,N_4437);
nor U4669 (N_4669,N_4460,N_4458);
nand U4670 (N_4670,N_4585,N_4511);
nand U4671 (N_4671,N_4565,N_4493);
nor U4672 (N_4672,N_4564,N_4519);
nand U4673 (N_4673,N_4500,N_4487);
and U4674 (N_4674,N_4555,N_4485);
nor U4675 (N_4675,N_4433,N_4483);
or U4676 (N_4676,N_4430,N_4479);
and U4677 (N_4677,N_4423,N_4530);
and U4678 (N_4678,N_4567,N_4552);
and U4679 (N_4679,N_4581,N_4444);
or U4680 (N_4680,N_4587,N_4471);
or U4681 (N_4681,N_4451,N_4515);
or U4682 (N_4682,N_4596,N_4478);
or U4683 (N_4683,N_4518,N_4578);
nand U4684 (N_4684,N_4464,N_4538);
nand U4685 (N_4685,N_4474,N_4491);
xnor U4686 (N_4686,N_4495,N_4434);
and U4687 (N_4687,N_4456,N_4411);
nand U4688 (N_4688,N_4506,N_4599);
and U4689 (N_4689,N_4512,N_4431);
or U4690 (N_4690,N_4593,N_4544);
and U4691 (N_4691,N_4583,N_4526);
and U4692 (N_4692,N_4572,N_4557);
and U4693 (N_4693,N_4537,N_4517);
and U4694 (N_4694,N_4588,N_4401);
nor U4695 (N_4695,N_4520,N_4421);
nand U4696 (N_4696,N_4545,N_4400);
and U4697 (N_4697,N_4516,N_4598);
or U4698 (N_4698,N_4577,N_4547);
nand U4699 (N_4699,N_4445,N_4582);
nor U4700 (N_4700,N_4535,N_4444);
nor U4701 (N_4701,N_4592,N_4543);
nand U4702 (N_4702,N_4534,N_4415);
and U4703 (N_4703,N_4559,N_4439);
nand U4704 (N_4704,N_4507,N_4450);
nand U4705 (N_4705,N_4484,N_4533);
or U4706 (N_4706,N_4585,N_4566);
or U4707 (N_4707,N_4547,N_4535);
or U4708 (N_4708,N_4517,N_4573);
and U4709 (N_4709,N_4495,N_4488);
or U4710 (N_4710,N_4445,N_4580);
nor U4711 (N_4711,N_4443,N_4417);
and U4712 (N_4712,N_4420,N_4562);
and U4713 (N_4713,N_4446,N_4484);
nor U4714 (N_4714,N_4563,N_4503);
or U4715 (N_4715,N_4568,N_4457);
or U4716 (N_4716,N_4461,N_4432);
and U4717 (N_4717,N_4506,N_4573);
or U4718 (N_4718,N_4447,N_4444);
nand U4719 (N_4719,N_4488,N_4492);
and U4720 (N_4720,N_4590,N_4431);
or U4721 (N_4721,N_4400,N_4530);
nor U4722 (N_4722,N_4557,N_4562);
and U4723 (N_4723,N_4480,N_4436);
nor U4724 (N_4724,N_4538,N_4479);
nor U4725 (N_4725,N_4528,N_4474);
or U4726 (N_4726,N_4404,N_4468);
or U4727 (N_4727,N_4476,N_4541);
nand U4728 (N_4728,N_4485,N_4498);
nand U4729 (N_4729,N_4454,N_4404);
and U4730 (N_4730,N_4562,N_4487);
and U4731 (N_4731,N_4547,N_4537);
or U4732 (N_4732,N_4555,N_4421);
nand U4733 (N_4733,N_4488,N_4599);
nor U4734 (N_4734,N_4598,N_4465);
nor U4735 (N_4735,N_4418,N_4471);
nand U4736 (N_4736,N_4464,N_4510);
nor U4737 (N_4737,N_4585,N_4534);
or U4738 (N_4738,N_4558,N_4522);
and U4739 (N_4739,N_4521,N_4532);
and U4740 (N_4740,N_4445,N_4594);
and U4741 (N_4741,N_4490,N_4502);
and U4742 (N_4742,N_4509,N_4517);
or U4743 (N_4743,N_4498,N_4528);
nor U4744 (N_4744,N_4432,N_4565);
nand U4745 (N_4745,N_4575,N_4537);
and U4746 (N_4746,N_4515,N_4576);
nor U4747 (N_4747,N_4412,N_4540);
nor U4748 (N_4748,N_4493,N_4443);
nor U4749 (N_4749,N_4538,N_4550);
nor U4750 (N_4750,N_4599,N_4510);
nor U4751 (N_4751,N_4501,N_4530);
nor U4752 (N_4752,N_4407,N_4453);
and U4753 (N_4753,N_4557,N_4463);
nand U4754 (N_4754,N_4569,N_4538);
nor U4755 (N_4755,N_4588,N_4441);
and U4756 (N_4756,N_4426,N_4437);
nor U4757 (N_4757,N_4455,N_4494);
nor U4758 (N_4758,N_4589,N_4549);
nor U4759 (N_4759,N_4400,N_4481);
nand U4760 (N_4760,N_4463,N_4542);
nand U4761 (N_4761,N_4486,N_4550);
nand U4762 (N_4762,N_4574,N_4539);
or U4763 (N_4763,N_4591,N_4577);
and U4764 (N_4764,N_4466,N_4531);
nor U4765 (N_4765,N_4536,N_4469);
and U4766 (N_4766,N_4587,N_4407);
or U4767 (N_4767,N_4593,N_4564);
nand U4768 (N_4768,N_4596,N_4540);
nor U4769 (N_4769,N_4522,N_4419);
nand U4770 (N_4770,N_4459,N_4514);
or U4771 (N_4771,N_4583,N_4439);
nor U4772 (N_4772,N_4459,N_4582);
nor U4773 (N_4773,N_4590,N_4518);
nor U4774 (N_4774,N_4437,N_4444);
or U4775 (N_4775,N_4513,N_4511);
or U4776 (N_4776,N_4474,N_4561);
or U4777 (N_4777,N_4554,N_4411);
and U4778 (N_4778,N_4580,N_4435);
and U4779 (N_4779,N_4584,N_4470);
and U4780 (N_4780,N_4445,N_4456);
or U4781 (N_4781,N_4428,N_4413);
nand U4782 (N_4782,N_4586,N_4400);
and U4783 (N_4783,N_4463,N_4464);
and U4784 (N_4784,N_4446,N_4430);
nand U4785 (N_4785,N_4406,N_4475);
or U4786 (N_4786,N_4463,N_4473);
nand U4787 (N_4787,N_4517,N_4439);
or U4788 (N_4788,N_4597,N_4587);
and U4789 (N_4789,N_4552,N_4579);
and U4790 (N_4790,N_4410,N_4482);
nand U4791 (N_4791,N_4541,N_4490);
or U4792 (N_4792,N_4482,N_4495);
nand U4793 (N_4793,N_4571,N_4401);
nand U4794 (N_4794,N_4405,N_4501);
and U4795 (N_4795,N_4406,N_4487);
nand U4796 (N_4796,N_4488,N_4593);
nor U4797 (N_4797,N_4453,N_4582);
nor U4798 (N_4798,N_4584,N_4532);
nor U4799 (N_4799,N_4575,N_4525);
nand U4800 (N_4800,N_4626,N_4724);
nor U4801 (N_4801,N_4652,N_4671);
nand U4802 (N_4802,N_4682,N_4794);
or U4803 (N_4803,N_4709,N_4642);
and U4804 (N_4804,N_4744,N_4788);
nor U4805 (N_4805,N_4753,N_4714);
or U4806 (N_4806,N_4631,N_4646);
nor U4807 (N_4807,N_4607,N_4613);
or U4808 (N_4808,N_4658,N_4758);
nor U4809 (N_4809,N_4657,N_4731);
and U4810 (N_4810,N_4689,N_4601);
and U4811 (N_4811,N_4690,N_4693);
or U4812 (N_4812,N_4697,N_4787);
or U4813 (N_4813,N_4659,N_4694);
and U4814 (N_4814,N_4701,N_4737);
and U4815 (N_4815,N_4750,N_4654);
nand U4816 (N_4816,N_4799,N_4624);
or U4817 (N_4817,N_4727,N_4645);
nand U4818 (N_4818,N_4778,N_4691);
and U4819 (N_4819,N_4795,N_4656);
and U4820 (N_4820,N_4749,N_4718);
nand U4821 (N_4821,N_4666,N_4776);
nor U4822 (N_4822,N_4755,N_4619);
and U4823 (N_4823,N_4710,N_4650);
or U4824 (N_4824,N_4633,N_4777);
nand U4825 (N_4825,N_4635,N_4751);
and U4826 (N_4826,N_4669,N_4707);
and U4827 (N_4827,N_4637,N_4617);
nor U4828 (N_4828,N_4747,N_4785);
or U4829 (N_4829,N_4764,N_4786);
and U4830 (N_4830,N_4640,N_4621);
and U4831 (N_4831,N_4668,N_4632);
nor U4832 (N_4832,N_4674,N_4615);
or U4833 (N_4833,N_4702,N_4670);
or U4834 (N_4834,N_4684,N_4660);
or U4835 (N_4835,N_4729,N_4752);
nor U4836 (N_4836,N_4771,N_4603);
or U4837 (N_4837,N_4622,N_4790);
and U4838 (N_4838,N_4616,N_4728);
nor U4839 (N_4839,N_4716,N_4732);
and U4840 (N_4840,N_4757,N_4653);
nor U4841 (N_4841,N_4667,N_4704);
nor U4842 (N_4842,N_4779,N_4734);
or U4843 (N_4843,N_4706,N_4677);
and U4844 (N_4844,N_4698,N_4717);
and U4845 (N_4845,N_4708,N_4756);
nor U4846 (N_4846,N_4781,N_4748);
nor U4847 (N_4847,N_4796,N_4726);
nand U4848 (N_4848,N_4611,N_4792);
nor U4849 (N_4849,N_4797,N_4720);
or U4850 (N_4850,N_4745,N_4606);
nor U4851 (N_4851,N_4688,N_4696);
nor U4852 (N_4852,N_4614,N_4649);
nand U4853 (N_4853,N_4761,N_4648);
and U4854 (N_4854,N_4742,N_4695);
nor U4855 (N_4855,N_4686,N_4672);
nand U4856 (N_4856,N_4620,N_4628);
or U4857 (N_4857,N_4740,N_4673);
and U4858 (N_4858,N_4765,N_4791);
or U4859 (N_4859,N_4636,N_4627);
or U4860 (N_4860,N_4641,N_4738);
nand U4861 (N_4861,N_4722,N_4700);
nor U4862 (N_4862,N_4625,N_4676);
or U4863 (N_4863,N_4772,N_4664);
or U4864 (N_4864,N_4634,N_4651);
nor U4865 (N_4865,N_4767,N_4612);
nand U4866 (N_4866,N_4623,N_4768);
or U4867 (N_4867,N_4766,N_4730);
nor U4868 (N_4868,N_4638,N_4712);
and U4869 (N_4869,N_4680,N_4675);
nand U4870 (N_4870,N_4743,N_4643);
nand U4871 (N_4871,N_4608,N_4647);
or U4872 (N_4872,N_4774,N_4679);
and U4873 (N_4873,N_4735,N_4741);
and U4874 (N_4874,N_4665,N_4687);
nor U4875 (N_4875,N_4602,N_4605);
nand U4876 (N_4876,N_4759,N_4692);
nor U4877 (N_4877,N_4629,N_4610);
nor U4878 (N_4878,N_4798,N_4683);
and U4879 (N_4879,N_4733,N_4639);
and U4880 (N_4880,N_4644,N_4661);
or U4881 (N_4881,N_4782,N_4773);
or U4882 (N_4882,N_4703,N_4678);
nor U4883 (N_4883,N_4739,N_4719);
and U4884 (N_4884,N_4780,N_4769);
nand U4885 (N_4885,N_4763,N_4630);
or U4886 (N_4886,N_4783,N_4762);
or U4887 (N_4887,N_4663,N_4760);
xor U4888 (N_4888,N_4715,N_4789);
nand U4889 (N_4889,N_4600,N_4604);
or U4890 (N_4890,N_4723,N_4754);
and U4891 (N_4891,N_4746,N_4775);
nand U4892 (N_4892,N_4784,N_4662);
and U4893 (N_4893,N_4725,N_4655);
and U4894 (N_4894,N_4736,N_4681);
or U4895 (N_4895,N_4793,N_4711);
or U4896 (N_4896,N_4609,N_4770);
nand U4897 (N_4897,N_4713,N_4685);
nor U4898 (N_4898,N_4721,N_4699);
nor U4899 (N_4899,N_4705,N_4618);
and U4900 (N_4900,N_4797,N_4768);
and U4901 (N_4901,N_4647,N_4793);
or U4902 (N_4902,N_4727,N_4736);
and U4903 (N_4903,N_4628,N_4666);
and U4904 (N_4904,N_4783,N_4758);
and U4905 (N_4905,N_4678,N_4719);
or U4906 (N_4906,N_4625,N_4684);
nor U4907 (N_4907,N_4622,N_4719);
or U4908 (N_4908,N_4779,N_4633);
nor U4909 (N_4909,N_4796,N_4753);
nand U4910 (N_4910,N_4628,N_4721);
nor U4911 (N_4911,N_4727,N_4791);
and U4912 (N_4912,N_4621,N_4753);
and U4913 (N_4913,N_4669,N_4794);
nor U4914 (N_4914,N_4651,N_4641);
nand U4915 (N_4915,N_4628,N_4645);
or U4916 (N_4916,N_4661,N_4777);
or U4917 (N_4917,N_4693,N_4606);
or U4918 (N_4918,N_4721,N_4609);
or U4919 (N_4919,N_4655,N_4680);
nand U4920 (N_4920,N_4713,N_4735);
and U4921 (N_4921,N_4753,N_4762);
and U4922 (N_4922,N_4741,N_4655);
nor U4923 (N_4923,N_4770,N_4709);
and U4924 (N_4924,N_4673,N_4779);
or U4925 (N_4925,N_4695,N_4744);
nand U4926 (N_4926,N_4688,N_4739);
or U4927 (N_4927,N_4732,N_4743);
nor U4928 (N_4928,N_4644,N_4676);
nor U4929 (N_4929,N_4765,N_4747);
or U4930 (N_4930,N_4710,N_4769);
or U4931 (N_4931,N_4780,N_4610);
nand U4932 (N_4932,N_4631,N_4690);
nor U4933 (N_4933,N_4652,N_4713);
or U4934 (N_4934,N_4705,N_4614);
nor U4935 (N_4935,N_4680,N_4747);
nand U4936 (N_4936,N_4615,N_4679);
and U4937 (N_4937,N_4603,N_4680);
nand U4938 (N_4938,N_4646,N_4641);
nand U4939 (N_4939,N_4626,N_4711);
and U4940 (N_4940,N_4717,N_4710);
nor U4941 (N_4941,N_4734,N_4619);
and U4942 (N_4942,N_4623,N_4699);
and U4943 (N_4943,N_4742,N_4635);
or U4944 (N_4944,N_4649,N_4694);
or U4945 (N_4945,N_4605,N_4796);
nor U4946 (N_4946,N_4751,N_4625);
nand U4947 (N_4947,N_4648,N_4654);
or U4948 (N_4948,N_4764,N_4737);
or U4949 (N_4949,N_4615,N_4631);
and U4950 (N_4950,N_4632,N_4705);
or U4951 (N_4951,N_4603,N_4684);
or U4952 (N_4952,N_4754,N_4720);
and U4953 (N_4953,N_4701,N_4765);
nor U4954 (N_4954,N_4625,N_4674);
nand U4955 (N_4955,N_4758,N_4662);
and U4956 (N_4956,N_4614,N_4748);
nor U4957 (N_4957,N_4734,N_4642);
and U4958 (N_4958,N_4746,N_4686);
nand U4959 (N_4959,N_4645,N_4693);
nor U4960 (N_4960,N_4746,N_4711);
and U4961 (N_4961,N_4777,N_4718);
and U4962 (N_4962,N_4621,N_4641);
or U4963 (N_4963,N_4716,N_4625);
or U4964 (N_4964,N_4719,N_4687);
nand U4965 (N_4965,N_4725,N_4701);
and U4966 (N_4966,N_4782,N_4621);
and U4967 (N_4967,N_4623,N_4654);
or U4968 (N_4968,N_4690,N_4751);
and U4969 (N_4969,N_4736,N_4712);
or U4970 (N_4970,N_4731,N_4722);
and U4971 (N_4971,N_4645,N_4752);
nand U4972 (N_4972,N_4727,N_4641);
nor U4973 (N_4973,N_4724,N_4746);
nor U4974 (N_4974,N_4756,N_4723);
and U4975 (N_4975,N_4671,N_4752);
and U4976 (N_4976,N_4740,N_4679);
nand U4977 (N_4977,N_4759,N_4630);
and U4978 (N_4978,N_4789,N_4624);
nand U4979 (N_4979,N_4774,N_4719);
or U4980 (N_4980,N_4726,N_4779);
nand U4981 (N_4981,N_4666,N_4730);
nor U4982 (N_4982,N_4792,N_4748);
nand U4983 (N_4983,N_4683,N_4784);
or U4984 (N_4984,N_4620,N_4771);
nor U4985 (N_4985,N_4693,N_4642);
and U4986 (N_4986,N_4657,N_4617);
or U4987 (N_4987,N_4707,N_4715);
or U4988 (N_4988,N_4710,N_4724);
nand U4989 (N_4989,N_4792,N_4702);
and U4990 (N_4990,N_4659,N_4741);
nand U4991 (N_4991,N_4766,N_4676);
nor U4992 (N_4992,N_4678,N_4662);
nor U4993 (N_4993,N_4610,N_4678);
or U4994 (N_4994,N_4601,N_4626);
or U4995 (N_4995,N_4777,N_4606);
nor U4996 (N_4996,N_4750,N_4797);
and U4997 (N_4997,N_4730,N_4717);
or U4998 (N_4998,N_4647,N_4764);
nand U4999 (N_4999,N_4653,N_4797);
and UO_0 (O_0,N_4910,N_4854);
or UO_1 (O_1,N_4875,N_4889);
nand UO_2 (O_2,N_4815,N_4995);
or UO_3 (O_3,N_4879,N_4918);
nor UO_4 (O_4,N_4803,N_4829);
nand UO_5 (O_5,N_4836,N_4984);
nor UO_6 (O_6,N_4823,N_4979);
or UO_7 (O_7,N_4804,N_4852);
nor UO_8 (O_8,N_4837,N_4980);
nand UO_9 (O_9,N_4880,N_4973);
nand UO_10 (O_10,N_4814,N_4811);
and UO_11 (O_11,N_4808,N_4849);
or UO_12 (O_12,N_4869,N_4857);
or UO_13 (O_13,N_4926,N_4839);
nor UO_14 (O_14,N_4820,N_4967);
nor UO_15 (O_15,N_4920,N_4903);
nor UO_16 (O_16,N_4913,N_4818);
nand UO_17 (O_17,N_4847,N_4873);
nor UO_18 (O_18,N_4883,N_4897);
and UO_19 (O_19,N_4871,N_4891);
nor UO_20 (O_20,N_4835,N_4916);
and UO_21 (O_21,N_4959,N_4862);
and UO_22 (O_22,N_4987,N_4939);
nor UO_23 (O_23,N_4986,N_4905);
nand UO_24 (O_24,N_4914,N_4930);
and UO_25 (O_25,N_4821,N_4977);
or UO_26 (O_26,N_4828,N_4867);
nand UO_27 (O_27,N_4813,N_4841);
nand UO_28 (O_28,N_4825,N_4990);
and UO_29 (O_29,N_4864,N_4812);
nand UO_30 (O_30,N_4944,N_4800);
or UO_31 (O_31,N_4966,N_4898);
nand UO_32 (O_32,N_4831,N_4983);
and UO_33 (O_33,N_4893,N_4943);
nor UO_34 (O_34,N_4950,N_4861);
nand UO_35 (O_35,N_4992,N_4947);
nor UO_36 (O_36,N_4985,N_4958);
nand UO_37 (O_37,N_4809,N_4838);
nor UO_38 (O_38,N_4817,N_4832);
nor UO_39 (O_39,N_4952,N_4919);
xor UO_40 (O_40,N_4969,N_4885);
or UO_41 (O_41,N_4901,N_4940);
nand UO_42 (O_42,N_4801,N_4922);
nor UO_43 (O_43,N_4846,N_4964);
nand UO_44 (O_44,N_4865,N_4834);
nand UO_45 (O_45,N_4863,N_4842);
or UO_46 (O_46,N_4954,N_4927);
nand UO_47 (O_47,N_4965,N_4909);
nor UO_48 (O_48,N_4884,N_4868);
nor UO_49 (O_49,N_4877,N_4997);
and UO_50 (O_50,N_4970,N_4911);
or UO_51 (O_51,N_4906,N_4826);
nand UO_52 (O_52,N_4945,N_4996);
nand UO_53 (O_53,N_4933,N_4802);
or UO_54 (O_54,N_4936,N_4824);
and UO_55 (O_55,N_4816,N_4982);
nand UO_56 (O_56,N_4928,N_4935);
nor UO_57 (O_57,N_4899,N_4878);
or UO_58 (O_58,N_4872,N_4874);
or UO_59 (O_59,N_4998,N_4830);
and UO_60 (O_60,N_4851,N_4953);
and UO_61 (O_61,N_4886,N_4917);
nor UO_62 (O_62,N_4855,N_4866);
or UO_63 (O_63,N_4931,N_4843);
or UO_64 (O_64,N_4887,N_4925);
or UO_65 (O_65,N_4921,N_4963);
nor UO_66 (O_66,N_4907,N_4948);
nor UO_67 (O_67,N_4856,N_4946);
nor UO_68 (O_68,N_4908,N_4938);
or UO_69 (O_69,N_4962,N_4853);
nor UO_70 (O_70,N_4819,N_4974);
and UO_71 (O_71,N_4902,N_4924);
and UO_72 (O_72,N_4858,N_4961);
nand UO_73 (O_73,N_4932,N_4929);
or UO_74 (O_74,N_4942,N_4993);
or UO_75 (O_75,N_4972,N_4895);
and UO_76 (O_76,N_4999,N_4960);
nand UO_77 (O_77,N_4827,N_4989);
nor UO_78 (O_78,N_4955,N_4949);
or UO_79 (O_79,N_4975,N_4805);
nand UO_80 (O_80,N_4848,N_4988);
nor UO_81 (O_81,N_4976,N_4941);
nor UO_82 (O_82,N_4822,N_4904);
nor UO_83 (O_83,N_4971,N_4860);
nand UO_84 (O_84,N_4956,N_4934);
nor UO_85 (O_85,N_4915,N_4859);
nand UO_86 (O_86,N_4888,N_4912);
nand UO_87 (O_87,N_4870,N_4850);
or UO_88 (O_88,N_4882,N_4994);
or UO_89 (O_89,N_4981,N_4968);
nor UO_90 (O_90,N_4894,N_4978);
nor UO_91 (O_91,N_4876,N_4896);
or UO_92 (O_92,N_4806,N_4991);
and UO_93 (O_93,N_4844,N_4810);
and UO_94 (O_94,N_4890,N_4833);
or UO_95 (O_95,N_4923,N_4881);
xnor UO_96 (O_96,N_4845,N_4807);
nand UO_97 (O_97,N_4840,N_4892);
and UO_98 (O_98,N_4900,N_4957);
or UO_99 (O_99,N_4951,N_4937);
nand UO_100 (O_100,N_4963,N_4837);
nand UO_101 (O_101,N_4916,N_4959);
and UO_102 (O_102,N_4815,N_4800);
nand UO_103 (O_103,N_4928,N_4803);
nand UO_104 (O_104,N_4999,N_4936);
nand UO_105 (O_105,N_4881,N_4908);
nor UO_106 (O_106,N_4980,N_4849);
nand UO_107 (O_107,N_4892,N_4823);
nand UO_108 (O_108,N_4994,N_4811);
or UO_109 (O_109,N_4939,N_4808);
nor UO_110 (O_110,N_4973,N_4976);
or UO_111 (O_111,N_4975,N_4808);
nor UO_112 (O_112,N_4875,N_4964);
nor UO_113 (O_113,N_4910,N_4881);
and UO_114 (O_114,N_4949,N_4870);
or UO_115 (O_115,N_4834,N_4937);
or UO_116 (O_116,N_4983,N_4805);
or UO_117 (O_117,N_4996,N_4833);
nor UO_118 (O_118,N_4811,N_4937);
nor UO_119 (O_119,N_4860,N_4811);
nand UO_120 (O_120,N_4947,N_4901);
nand UO_121 (O_121,N_4975,N_4883);
nand UO_122 (O_122,N_4895,N_4829);
nor UO_123 (O_123,N_4870,N_4966);
or UO_124 (O_124,N_4870,N_4874);
nor UO_125 (O_125,N_4894,N_4807);
or UO_126 (O_126,N_4908,N_4854);
nor UO_127 (O_127,N_4998,N_4977);
or UO_128 (O_128,N_4846,N_4836);
nand UO_129 (O_129,N_4872,N_4950);
nor UO_130 (O_130,N_4853,N_4835);
nor UO_131 (O_131,N_4854,N_4994);
and UO_132 (O_132,N_4851,N_4804);
nand UO_133 (O_133,N_4824,N_4964);
nor UO_134 (O_134,N_4975,N_4978);
and UO_135 (O_135,N_4801,N_4837);
and UO_136 (O_136,N_4907,N_4874);
and UO_137 (O_137,N_4882,N_4969);
nand UO_138 (O_138,N_4959,N_4867);
nand UO_139 (O_139,N_4882,N_4854);
nor UO_140 (O_140,N_4956,N_4826);
nand UO_141 (O_141,N_4960,N_4913);
and UO_142 (O_142,N_4946,N_4828);
nor UO_143 (O_143,N_4914,N_4895);
nor UO_144 (O_144,N_4881,N_4882);
nor UO_145 (O_145,N_4967,N_4955);
or UO_146 (O_146,N_4857,N_4803);
or UO_147 (O_147,N_4804,N_4978);
and UO_148 (O_148,N_4842,N_4911);
nor UO_149 (O_149,N_4919,N_4917);
and UO_150 (O_150,N_4979,N_4966);
nand UO_151 (O_151,N_4987,N_4915);
nor UO_152 (O_152,N_4920,N_4877);
nand UO_153 (O_153,N_4870,N_4866);
nand UO_154 (O_154,N_4936,N_4816);
nand UO_155 (O_155,N_4941,N_4985);
and UO_156 (O_156,N_4953,N_4946);
and UO_157 (O_157,N_4980,N_4864);
nand UO_158 (O_158,N_4950,N_4866);
nand UO_159 (O_159,N_4866,N_4960);
nor UO_160 (O_160,N_4996,N_4977);
or UO_161 (O_161,N_4960,N_4949);
nand UO_162 (O_162,N_4929,N_4890);
or UO_163 (O_163,N_4917,N_4888);
and UO_164 (O_164,N_4809,N_4837);
or UO_165 (O_165,N_4837,N_4954);
nand UO_166 (O_166,N_4971,N_4992);
or UO_167 (O_167,N_4846,N_4860);
or UO_168 (O_168,N_4873,N_4805);
or UO_169 (O_169,N_4977,N_4921);
and UO_170 (O_170,N_4832,N_4990);
nor UO_171 (O_171,N_4855,N_4846);
or UO_172 (O_172,N_4827,N_4810);
and UO_173 (O_173,N_4811,N_4962);
or UO_174 (O_174,N_4856,N_4912);
or UO_175 (O_175,N_4910,N_4927);
nor UO_176 (O_176,N_4980,N_4846);
nand UO_177 (O_177,N_4975,N_4814);
or UO_178 (O_178,N_4848,N_4820);
and UO_179 (O_179,N_4939,N_4897);
nand UO_180 (O_180,N_4895,N_4897);
nor UO_181 (O_181,N_4942,N_4845);
nand UO_182 (O_182,N_4999,N_4813);
nor UO_183 (O_183,N_4985,N_4827);
or UO_184 (O_184,N_4811,N_4895);
and UO_185 (O_185,N_4968,N_4823);
or UO_186 (O_186,N_4870,N_4881);
or UO_187 (O_187,N_4823,N_4910);
nor UO_188 (O_188,N_4826,N_4835);
or UO_189 (O_189,N_4818,N_4838);
nor UO_190 (O_190,N_4946,N_4852);
nor UO_191 (O_191,N_4862,N_4902);
nor UO_192 (O_192,N_4808,N_4998);
or UO_193 (O_193,N_4886,N_4950);
nand UO_194 (O_194,N_4870,N_4884);
and UO_195 (O_195,N_4881,N_4883);
and UO_196 (O_196,N_4888,N_4937);
or UO_197 (O_197,N_4888,N_4859);
and UO_198 (O_198,N_4964,N_4871);
or UO_199 (O_199,N_4872,N_4913);
or UO_200 (O_200,N_4851,N_4833);
nand UO_201 (O_201,N_4850,N_4966);
and UO_202 (O_202,N_4874,N_4961);
nor UO_203 (O_203,N_4801,N_4800);
or UO_204 (O_204,N_4915,N_4908);
nor UO_205 (O_205,N_4897,N_4906);
or UO_206 (O_206,N_4861,N_4850);
nor UO_207 (O_207,N_4958,N_4965);
or UO_208 (O_208,N_4956,N_4807);
or UO_209 (O_209,N_4850,N_4842);
nor UO_210 (O_210,N_4866,N_4905);
or UO_211 (O_211,N_4841,N_4920);
or UO_212 (O_212,N_4980,N_4918);
nand UO_213 (O_213,N_4964,N_4985);
or UO_214 (O_214,N_4865,N_4830);
and UO_215 (O_215,N_4992,N_4886);
xor UO_216 (O_216,N_4952,N_4893);
or UO_217 (O_217,N_4835,N_4818);
nand UO_218 (O_218,N_4955,N_4911);
or UO_219 (O_219,N_4811,N_4883);
nand UO_220 (O_220,N_4979,N_4868);
and UO_221 (O_221,N_4867,N_4868);
or UO_222 (O_222,N_4952,N_4942);
and UO_223 (O_223,N_4801,N_4821);
xnor UO_224 (O_224,N_4908,N_4808);
nand UO_225 (O_225,N_4805,N_4898);
nor UO_226 (O_226,N_4937,N_4886);
nand UO_227 (O_227,N_4962,N_4998);
and UO_228 (O_228,N_4884,N_4933);
and UO_229 (O_229,N_4903,N_4958);
nand UO_230 (O_230,N_4980,N_4824);
or UO_231 (O_231,N_4939,N_4904);
or UO_232 (O_232,N_4914,N_4849);
or UO_233 (O_233,N_4842,N_4815);
nand UO_234 (O_234,N_4942,N_4977);
or UO_235 (O_235,N_4946,N_4811);
nor UO_236 (O_236,N_4951,N_4967);
nand UO_237 (O_237,N_4912,N_4839);
or UO_238 (O_238,N_4930,N_4873);
nand UO_239 (O_239,N_4803,N_4935);
and UO_240 (O_240,N_4947,N_4971);
nand UO_241 (O_241,N_4871,N_4873);
nand UO_242 (O_242,N_4917,N_4959);
or UO_243 (O_243,N_4852,N_4938);
nand UO_244 (O_244,N_4815,N_4984);
or UO_245 (O_245,N_4999,N_4966);
nor UO_246 (O_246,N_4875,N_4810);
or UO_247 (O_247,N_4983,N_4854);
nand UO_248 (O_248,N_4949,N_4948);
and UO_249 (O_249,N_4860,N_4869);
or UO_250 (O_250,N_4936,N_4896);
or UO_251 (O_251,N_4988,N_4863);
nor UO_252 (O_252,N_4927,N_4996);
and UO_253 (O_253,N_4878,N_4868);
or UO_254 (O_254,N_4874,N_4922);
or UO_255 (O_255,N_4945,N_4869);
or UO_256 (O_256,N_4917,N_4871);
nand UO_257 (O_257,N_4817,N_4855);
nor UO_258 (O_258,N_4828,N_4821);
or UO_259 (O_259,N_4901,N_4999);
or UO_260 (O_260,N_4927,N_4802);
nand UO_261 (O_261,N_4922,N_4833);
and UO_262 (O_262,N_4928,N_4946);
nor UO_263 (O_263,N_4991,N_4916);
or UO_264 (O_264,N_4807,N_4949);
or UO_265 (O_265,N_4955,N_4857);
nand UO_266 (O_266,N_4963,N_4942);
or UO_267 (O_267,N_4864,N_4840);
and UO_268 (O_268,N_4951,N_4932);
and UO_269 (O_269,N_4845,N_4856);
and UO_270 (O_270,N_4810,N_4996);
nand UO_271 (O_271,N_4968,N_4977);
nand UO_272 (O_272,N_4981,N_4909);
nor UO_273 (O_273,N_4836,N_4868);
nand UO_274 (O_274,N_4961,N_4811);
or UO_275 (O_275,N_4980,N_4851);
or UO_276 (O_276,N_4985,N_4907);
and UO_277 (O_277,N_4989,N_4916);
nand UO_278 (O_278,N_4888,N_4887);
nor UO_279 (O_279,N_4813,N_4842);
nand UO_280 (O_280,N_4946,N_4817);
nor UO_281 (O_281,N_4989,N_4889);
nand UO_282 (O_282,N_4837,N_4956);
and UO_283 (O_283,N_4867,N_4991);
nand UO_284 (O_284,N_4819,N_4858);
nand UO_285 (O_285,N_4997,N_4955);
nor UO_286 (O_286,N_4988,N_4978);
or UO_287 (O_287,N_4927,N_4892);
and UO_288 (O_288,N_4976,N_4864);
or UO_289 (O_289,N_4812,N_4819);
nand UO_290 (O_290,N_4802,N_4985);
and UO_291 (O_291,N_4801,N_4916);
and UO_292 (O_292,N_4837,N_4836);
or UO_293 (O_293,N_4908,N_4832);
and UO_294 (O_294,N_4946,N_4840);
or UO_295 (O_295,N_4944,N_4949);
and UO_296 (O_296,N_4971,N_4891);
nand UO_297 (O_297,N_4893,N_4906);
and UO_298 (O_298,N_4892,N_4817);
or UO_299 (O_299,N_4840,N_4815);
nor UO_300 (O_300,N_4821,N_4931);
nor UO_301 (O_301,N_4816,N_4871);
or UO_302 (O_302,N_4973,N_4988);
nand UO_303 (O_303,N_4973,N_4838);
nand UO_304 (O_304,N_4895,N_4863);
nand UO_305 (O_305,N_4896,N_4990);
nand UO_306 (O_306,N_4978,N_4821);
or UO_307 (O_307,N_4893,N_4841);
and UO_308 (O_308,N_4925,N_4935);
nand UO_309 (O_309,N_4869,N_4867);
nor UO_310 (O_310,N_4857,N_4817);
nor UO_311 (O_311,N_4858,N_4883);
nor UO_312 (O_312,N_4820,N_4943);
nand UO_313 (O_313,N_4990,N_4956);
nand UO_314 (O_314,N_4964,N_4864);
or UO_315 (O_315,N_4989,N_4848);
or UO_316 (O_316,N_4852,N_4928);
and UO_317 (O_317,N_4999,N_4899);
and UO_318 (O_318,N_4826,N_4893);
nor UO_319 (O_319,N_4901,N_4875);
nand UO_320 (O_320,N_4879,N_4937);
nor UO_321 (O_321,N_4823,N_4803);
or UO_322 (O_322,N_4900,N_4985);
nor UO_323 (O_323,N_4925,N_4848);
nor UO_324 (O_324,N_4919,N_4957);
nor UO_325 (O_325,N_4856,N_4848);
or UO_326 (O_326,N_4923,N_4972);
or UO_327 (O_327,N_4815,N_4986);
nor UO_328 (O_328,N_4857,N_4988);
nand UO_329 (O_329,N_4955,N_4953);
nand UO_330 (O_330,N_4923,N_4815);
or UO_331 (O_331,N_4930,N_4956);
or UO_332 (O_332,N_4869,N_4849);
and UO_333 (O_333,N_4863,N_4983);
and UO_334 (O_334,N_4878,N_4931);
or UO_335 (O_335,N_4914,N_4981);
nor UO_336 (O_336,N_4818,N_4968);
nor UO_337 (O_337,N_4874,N_4826);
nor UO_338 (O_338,N_4876,N_4998);
nand UO_339 (O_339,N_4970,N_4902);
and UO_340 (O_340,N_4927,N_4988);
or UO_341 (O_341,N_4858,N_4812);
nor UO_342 (O_342,N_4994,N_4858);
nor UO_343 (O_343,N_4965,N_4841);
nand UO_344 (O_344,N_4835,N_4977);
nand UO_345 (O_345,N_4941,N_4920);
and UO_346 (O_346,N_4932,N_4944);
and UO_347 (O_347,N_4866,N_4837);
or UO_348 (O_348,N_4955,N_4922);
and UO_349 (O_349,N_4939,N_4804);
nor UO_350 (O_350,N_4984,N_4863);
nand UO_351 (O_351,N_4814,N_4838);
nor UO_352 (O_352,N_4858,N_4837);
nor UO_353 (O_353,N_4925,N_4810);
or UO_354 (O_354,N_4870,N_4936);
and UO_355 (O_355,N_4966,N_4911);
or UO_356 (O_356,N_4949,N_4956);
and UO_357 (O_357,N_4903,N_4967);
and UO_358 (O_358,N_4846,N_4823);
nand UO_359 (O_359,N_4891,N_4895);
and UO_360 (O_360,N_4833,N_4933);
and UO_361 (O_361,N_4928,N_4867);
nor UO_362 (O_362,N_4877,N_4821);
or UO_363 (O_363,N_4859,N_4860);
xor UO_364 (O_364,N_4816,N_4806);
or UO_365 (O_365,N_4968,N_4850);
or UO_366 (O_366,N_4934,N_4907);
and UO_367 (O_367,N_4995,N_4824);
and UO_368 (O_368,N_4964,N_4826);
nand UO_369 (O_369,N_4937,N_4858);
or UO_370 (O_370,N_4904,N_4886);
nor UO_371 (O_371,N_4931,N_4849);
nand UO_372 (O_372,N_4929,N_4860);
nor UO_373 (O_373,N_4911,N_4845);
and UO_374 (O_374,N_4976,N_4970);
nand UO_375 (O_375,N_4958,N_4802);
nor UO_376 (O_376,N_4824,N_4814);
nor UO_377 (O_377,N_4992,N_4818);
nor UO_378 (O_378,N_4889,N_4854);
nand UO_379 (O_379,N_4970,N_4866);
nand UO_380 (O_380,N_4869,N_4991);
nor UO_381 (O_381,N_4976,N_4816);
or UO_382 (O_382,N_4999,N_4806);
nor UO_383 (O_383,N_4930,N_4936);
or UO_384 (O_384,N_4894,N_4874);
nor UO_385 (O_385,N_4817,N_4887);
nand UO_386 (O_386,N_4939,N_4902);
nand UO_387 (O_387,N_4948,N_4929);
and UO_388 (O_388,N_4843,N_4990);
xnor UO_389 (O_389,N_4956,N_4957);
and UO_390 (O_390,N_4807,N_4833);
nand UO_391 (O_391,N_4938,N_4987);
nand UO_392 (O_392,N_4847,N_4990);
or UO_393 (O_393,N_4973,N_4917);
and UO_394 (O_394,N_4967,N_4881);
nor UO_395 (O_395,N_4817,N_4807);
nor UO_396 (O_396,N_4898,N_4809);
or UO_397 (O_397,N_4831,N_4808);
and UO_398 (O_398,N_4989,N_4955);
nor UO_399 (O_399,N_4988,N_4969);
and UO_400 (O_400,N_4829,N_4884);
or UO_401 (O_401,N_4830,N_4928);
or UO_402 (O_402,N_4953,N_4850);
or UO_403 (O_403,N_4993,N_4935);
or UO_404 (O_404,N_4863,N_4954);
or UO_405 (O_405,N_4961,N_4980);
and UO_406 (O_406,N_4908,N_4928);
or UO_407 (O_407,N_4870,N_4983);
nor UO_408 (O_408,N_4943,N_4814);
nand UO_409 (O_409,N_4818,N_4990);
nand UO_410 (O_410,N_4997,N_4805);
xnor UO_411 (O_411,N_4940,N_4928);
and UO_412 (O_412,N_4907,N_4823);
or UO_413 (O_413,N_4931,N_4831);
nor UO_414 (O_414,N_4995,N_4937);
and UO_415 (O_415,N_4936,N_4859);
or UO_416 (O_416,N_4915,N_4821);
and UO_417 (O_417,N_4826,N_4944);
and UO_418 (O_418,N_4908,N_4886);
nand UO_419 (O_419,N_4909,N_4875);
and UO_420 (O_420,N_4906,N_4974);
nor UO_421 (O_421,N_4907,N_4940);
and UO_422 (O_422,N_4987,N_4964);
and UO_423 (O_423,N_4868,N_4891);
and UO_424 (O_424,N_4824,N_4928);
and UO_425 (O_425,N_4970,N_4977);
nor UO_426 (O_426,N_4970,N_4932);
and UO_427 (O_427,N_4845,N_4979);
nand UO_428 (O_428,N_4954,N_4908);
nand UO_429 (O_429,N_4916,N_4974);
nand UO_430 (O_430,N_4933,N_4943);
nor UO_431 (O_431,N_4919,N_4974);
or UO_432 (O_432,N_4802,N_4838);
nor UO_433 (O_433,N_4858,N_4891);
nor UO_434 (O_434,N_4995,N_4952);
and UO_435 (O_435,N_4864,N_4996);
nand UO_436 (O_436,N_4843,N_4940);
and UO_437 (O_437,N_4815,N_4839);
or UO_438 (O_438,N_4866,N_4948);
nand UO_439 (O_439,N_4971,N_4975);
nor UO_440 (O_440,N_4894,N_4959);
nand UO_441 (O_441,N_4913,N_4967);
nor UO_442 (O_442,N_4964,N_4902);
nor UO_443 (O_443,N_4814,N_4845);
nor UO_444 (O_444,N_4816,N_4863);
and UO_445 (O_445,N_4877,N_4827);
or UO_446 (O_446,N_4882,N_4842);
or UO_447 (O_447,N_4801,N_4893);
or UO_448 (O_448,N_4922,N_4846);
or UO_449 (O_449,N_4882,N_4926);
nand UO_450 (O_450,N_4877,N_4927);
nand UO_451 (O_451,N_4900,N_4871);
or UO_452 (O_452,N_4878,N_4934);
and UO_453 (O_453,N_4935,N_4980);
nand UO_454 (O_454,N_4869,N_4907);
nor UO_455 (O_455,N_4840,N_4965);
and UO_456 (O_456,N_4855,N_4843);
and UO_457 (O_457,N_4865,N_4920);
nor UO_458 (O_458,N_4864,N_4852);
and UO_459 (O_459,N_4837,N_4815);
or UO_460 (O_460,N_4898,N_4820);
nor UO_461 (O_461,N_4973,N_4989);
or UO_462 (O_462,N_4995,N_4901);
and UO_463 (O_463,N_4998,N_4980);
nand UO_464 (O_464,N_4888,N_4940);
nor UO_465 (O_465,N_4805,N_4826);
and UO_466 (O_466,N_4810,N_4977);
xor UO_467 (O_467,N_4945,N_4899);
nand UO_468 (O_468,N_4960,N_4962);
or UO_469 (O_469,N_4815,N_4854);
nor UO_470 (O_470,N_4802,N_4918);
nor UO_471 (O_471,N_4969,N_4820);
nor UO_472 (O_472,N_4878,N_4986);
nand UO_473 (O_473,N_4916,N_4802);
nor UO_474 (O_474,N_4939,N_4964);
nor UO_475 (O_475,N_4924,N_4982);
nand UO_476 (O_476,N_4952,N_4854);
or UO_477 (O_477,N_4919,N_4970);
or UO_478 (O_478,N_4903,N_4950);
nand UO_479 (O_479,N_4937,N_4941);
nor UO_480 (O_480,N_4870,N_4818);
nand UO_481 (O_481,N_4899,N_4926);
and UO_482 (O_482,N_4839,N_4952);
nor UO_483 (O_483,N_4944,N_4809);
or UO_484 (O_484,N_4805,N_4837);
nor UO_485 (O_485,N_4846,N_4850);
and UO_486 (O_486,N_4844,N_4980);
or UO_487 (O_487,N_4979,N_4878);
or UO_488 (O_488,N_4911,N_4914);
and UO_489 (O_489,N_4887,N_4870);
and UO_490 (O_490,N_4901,N_4921);
or UO_491 (O_491,N_4817,N_4891);
or UO_492 (O_492,N_4974,N_4932);
or UO_493 (O_493,N_4897,N_4839);
and UO_494 (O_494,N_4819,N_4888);
nor UO_495 (O_495,N_4900,N_4936);
nand UO_496 (O_496,N_4856,N_4943);
nor UO_497 (O_497,N_4910,N_4837);
or UO_498 (O_498,N_4989,N_4971);
and UO_499 (O_499,N_4913,N_4831);
nand UO_500 (O_500,N_4865,N_4890);
and UO_501 (O_501,N_4925,N_4937);
or UO_502 (O_502,N_4972,N_4838);
nor UO_503 (O_503,N_4887,N_4915);
nand UO_504 (O_504,N_4856,N_4901);
nand UO_505 (O_505,N_4918,N_4853);
nand UO_506 (O_506,N_4975,N_4995);
nand UO_507 (O_507,N_4955,N_4964);
and UO_508 (O_508,N_4910,N_4981);
and UO_509 (O_509,N_4827,N_4934);
nor UO_510 (O_510,N_4916,N_4958);
nand UO_511 (O_511,N_4949,N_4886);
nand UO_512 (O_512,N_4860,N_4853);
nor UO_513 (O_513,N_4891,N_4957);
nand UO_514 (O_514,N_4910,N_4967);
or UO_515 (O_515,N_4943,N_4865);
nor UO_516 (O_516,N_4970,N_4926);
or UO_517 (O_517,N_4887,N_4946);
nand UO_518 (O_518,N_4926,N_4813);
nor UO_519 (O_519,N_4909,N_4995);
nor UO_520 (O_520,N_4950,N_4996);
and UO_521 (O_521,N_4967,N_4854);
nor UO_522 (O_522,N_4855,N_4877);
and UO_523 (O_523,N_4924,N_4957);
and UO_524 (O_524,N_4966,N_4960);
nand UO_525 (O_525,N_4955,N_4988);
or UO_526 (O_526,N_4903,N_4946);
nor UO_527 (O_527,N_4806,N_4949);
or UO_528 (O_528,N_4983,N_4998);
nand UO_529 (O_529,N_4815,N_4918);
nor UO_530 (O_530,N_4908,N_4956);
or UO_531 (O_531,N_4823,N_4822);
xnor UO_532 (O_532,N_4923,N_4929);
and UO_533 (O_533,N_4850,N_4892);
nor UO_534 (O_534,N_4893,N_4975);
nor UO_535 (O_535,N_4936,N_4880);
or UO_536 (O_536,N_4874,N_4927);
nor UO_537 (O_537,N_4884,N_4843);
and UO_538 (O_538,N_4930,N_4910);
nand UO_539 (O_539,N_4857,N_4826);
or UO_540 (O_540,N_4824,N_4893);
nand UO_541 (O_541,N_4923,N_4975);
or UO_542 (O_542,N_4828,N_4885);
nor UO_543 (O_543,N_4944,N_4837);
and UO_544 (O_544,N_4998,N_4863);
nor UO_545 (O_545,N_4808,N_4983);
nand UO_546 (O_546,N_4947,N_4879);
and UO_547 (O_547,N_4821,N_4809);
nor UO_548 (O_548,N_4842,N_4996);
and UO_549 (O_549,N_4832,N_4812);
or UO_550 (O_550,N_4922,N_4881);
or UO_551 (O_551,N_4916,N_4876);
or UO_552 (O_552,N_4848,N_4990);
nor UO_553 (O_553,N_4982,N_4903);
or UO_554 (O_554,N_4801,N_4953);
or UO_555 (O_555,N_4847,N_4879);
or UO_556 (O_556,N_4866,N_4802);
xor UO_557 (O_557,N_4990,N_4826);
nor UO_558 (O_558,N_4812,N_4863);
and UO_559 (O_559,N_4870,N_4817);
or UO_560 (O_560,N_4858,N_4977);
and UO_561 (O_561,N_4908,N_4974);
xnor UO_562 (O_562,N_4931,N_4964);
nor UO_563 (O_563,N_4924,N_4876);
or UO_564 (O_564,N_4924,N_4807);
nor UO_565 (O_565,N_4883,N_4859);
nor UO_566 (O_566,N_4996,N_4902);
nor UO_567 (O_567,N_4831,N_4887);
nand UO_568 (O_568,N_4940,N_4966);
nand UO_569 (O_569,N_4970,N_4813);
or UO_570 (O_570,N_4874,N_4918);
and UO_571 (O_571,N_4880,N_4878);
nand UO_572 (O_572,N_4908,N_4979);
and UO_573 (O_573,N_4832,N_4975);
nand UO_574 (O_574,N_4993,N_4876);
or UO_575 (O_575,N_4803,N_4902);
nand UO_576 (O_576,N_4882,N_4816);
nor UO_577 (O_577,N_4971,N_4916);
nor UO_578 (O_578,N_4978,N_4950);
or UO_579 (O_579,N_4903,N_4854);
and UO_580 (O_580,N_4951,N_4836);
nand UO_581 (O_581,N_4869,N_4895);
or UO_582 (O_582,N_4833,N_4888);
or UO_583 (O_583,N_4987,N_4821);
or UO_584 (O_584,N_4978,N_4995);
nand UO_585 (O_585,N_4821,N_4951);
nor UO_586 (O_586,N_4967,N_4858);
and UO_587 (O_587,N_4872,N_4987);
or UO_588 (O_588,N_4888,N_4981);
and UO_589 (O_589,N_4881,N_4838);
and UO_590 (O_590,N_4832,N_4935);
and UO_591 (O_591,N_4974,N_4943);
and UO_592 (O_592,N_4843,N_4804);
nand UO_593 (O_593,N_4950,N_4809);
nor UO_594 (O_594,N_4935,N_4952);
or UO_595 (O_595,N_4857,N_4958);
nand UO_596 (O_596,N_4807,N_4959);
nor UO_597 (O_597,N_4985,N_4949);
nor UO_598 (O_598,N_4915,N_4953);
nor UO_599 (O_599,N_4870,N_4880);
nor UO_600 (O_600,N_4911,N_4833);
and UO_601 (O_601,N_4864,N_4969);
nor UO_602 (O_602,N_4886,N_4934);
or UO_603 (O_603,N_4840,N_4985);
and UO_604 (O_604,N_4922,N_4828);
nand UO_605 (O_605,N_4920,N_4942);
and UO_606 (O_606,N_4855,N_4961);
nor UO_607 (O_607,N_4839,N_4923);
nor UO_608 (O_608,N_4817,N_4907);
or UO_609 (O_609,N_4828,N_4993);
or UO_610 (O_610,N_4921,N_4806);
or UO_611 (O_611,N_4923,N_4880);
or UO_612 (O_612,N_4998,N_4858);
nand UO_613 (O_613,N_4987,N_4937);
and UO_614 (O_614,N_4802,N_4903);
and UO_615 (O_615,N_4943,N_4982);
or UO_616 (O_616,N_4808,N_4996);
or UO_617 (O_617,N_4958,N_4865);
and UO_618 (O_618,N_4992,N_4817);
or UO_619 (O_619,N_4862,N_4897);
or UO_620 (O_620,N_4948,N_4881);
nor UO_621 (O_621,N_4804,N_4872);
nor UO_622 (O_622,N_4913,N_4813);
or UO_623 (O_623,N_4955,N_4926);
or UO_624 (O_624,N_4833,N_4934);
and UO_625 (O_625,N_4922,N_4938);
or UO_626 (O_626,N_4805,N_4957);
nor UO_627 (O_627,N_4951,N_4949);
or UO_628 (O_628,N_4818,N_4806);
and UO_629 (O_629,N_4834,N_4800);
or UO_630 (O_630,N_4847,N_4973);
and UO_631 (O_631,N_4974,N_4877);
nor UO_632 (O_632,N_4893,N_4806);
nand UO_633 (O_633,N_4909,N_4857);
nor UO_634 (O_634,N_4891,N_4916);
nor UO_635 (O_635,N_4874,N_4944);
or UO_636 (O_636,N_4954,N_4826);
nor UO_637 (O_637,N_4956,N_4895);
nor UO_638 (O_638,N_4871,N_4985);
and UO_639 (O_639,N_4966,N_4925);
nand UO_640 (O_640,N_4812,N_4946);
nor UO_641 (O_641,N_4932,N_4910);
and UO_642 (O_642,N_4838,N_4834);
nand UO_643 (O_643,N_4924,N_4997);
nand UO_644 (O_644,N_4910,N_4812);
and UO_645 (O_645,N_4829,N_4956);
nor UO_646 (O_646,N_4871,N_4911);
nand UO_647 (O_647,N_4952,N_4914);
nor UO_648 (O_648,N_4881,N_4956);
and UO_649 (O_649,N_4807,N_4947);
nand UO_650 (O_650,N_4936,N_4942);
and UO_651 (O_651,N_4818,N_4875);
or UO_652 (O_652,N_4882,N_4971);
nand UO_653 (O_653,N_4840,N_4802);
nand UO_654 (O_654,N_4922,N_4985);
and UO_655 (O_655,N_4914,N_4946);
and UO_656 (O_656,N_4859,N_4998);
nor UO_657 (O_657,N_4995,N_4972);
and UO_658 (O_658,N_4982,N_4880);
nand UO_659 (O_659,N_4827,N_4825);
and UO_660 (O_660,N_4986,N_4949);
and UO_661 (O_661,N_4978,N_4944);
and UO_662 (O_662,N_4929,N_4812);
or UO_663 (O_663,N_4907,N_4856);
nand UO_664 (O_664,N_4905,N_4973);
nand UO_665 (O_665,N_4964,N_4807);
nand UO_666 (O_666,N_4807,N_4946);
xor UO_667 (O_667,N_4968,N_4923);
nor UO_668 (O_668,N_4803,N_4909);
nand UO_669 (O_669,N_4852,N_4914);
or UO_670 (O_670,N_4847,N_4951);
and UO_671 (O_671,N_4927,N_4936);
or UO_672 (O_672,N_4973,N_4911);
or UO_673 (O_673,N_4950,N_4930);
and UO_674 (O_674,N_4882,N_4905);
or UO_675 (O_675,N_4849,N_4801);
or UO_676 (O_676,N_4965,N_4847);
and UO_677 (O_677,N_4800,N_4876);
or UO_678 (O_678,N_4823,N_4830);
or UO_679 (O_679,N_4961,N_4824);
and UO_680 (O_680,N_4814,N_4986);
nor UO_681 (O_681,N_4952,N_4975);
and UO_682 (O_682,N_4856,N_4859);
or UO_683 (O_683,N_4976,N_4884);
nand UO_684 (O_684,N_4918,N_4861);
and UO_685 (O_685,N_4896,N_4940);
and UO_686 (O_686,N_4862,N_4900);
nor UO_687 (O_687,N_4993,N_4913);
nor UO_688 (O_688,N_4940,N_4969);
and UO_689 (O_689,N_4849,N_4897);
nand UO_690 (O_690,N_4858,N_4814);
or UO_691 (O_691,N_4972,N_4951);
and UO_692 (O_692,N_4818,N_4914);
nor UO_693 (O_693,N_4986,N_4999);
or UO_694 (O_694,N_4976,N_4877);
or UO_695 (O_695,N_4835,N_4965);
and UO_696 (O_696,N_4832,N_4836);
and UO_697 (O_697,N_4864,N_4884);
and UO_698 (O_698,N_4871,N_4861);
nor UO_699 (O_699,N_4922,N_4870);
nand UO_700 (O_700,N_4832,N_4883);
and UO_701 (O_701,N_4867,N_4983);
and UO_702 (O_702,N_4861,N_4940);
nand UO_703 (O_703,N_4851,N_4829);
or UO_704 (O_704,N_4846,N_4915);
and UO_705 (O_705,N_4959,N_4981);
or UO_706 (O_706,N_4955,N_4904);
nand UO_707 (O_707,N_4816,N_4934);
or UO_708 (O_708,N_4955,N_4993);
and UO_709 (O_709,N_4964,N_4802);
and UO_710 (O_710,N_4944,N_4919);
or UO_711 (O_711,N_4813,N_4978);
nand UO_712 (O_712,N_4902,N_4896);
nand UO_713 (O_713,N_4997,N_4966);
nand UO_714 (O_714,N_4926,N_4903);
or UO_715 (O_715,N_4922,N_4848);
nand UO_716 (O_716,N_4809,N_4878);
nor UO_717 (O_717,N_4982,N_4963);
nor UO_718 (O_718,N_4983,N_4803);
nor UO_719 (O_719,N_4935,N_4813);
nand UO_720 (O_720,N_4909,N_4808);
nand UO_721 (O_721,N_4886,N_4885);
and UO_722 (O_722,N_4896,N_4803);
and UO_723 (O_723,N_4905,N_4833);
nand UO_724 (O_724,N_4943,N_4838);
or UO_725 (O_725,N_4841,N_4850);
or UO_726 (O_726,N_4867,N_4961);
nand UO_727 (O_727,N_4809,N_4924);
or UO_728 (O_728,N_4876,N_4827);
nand UO_729 (O_729,N_4964,N_4936);
or UO_730 (O_730,N_4885,N_4872);
nor UO_731 (O_731,N_4841,N_4845);
and UO_732 (O_732,N_4959,N_4804);
or UO_733 (O_733,N_4804,N_4955);
nand UO_734 (O_734,N_4931,N_4984);
and UO_735 (O_735,N_4960,N_4839);
and UO_736 (O_736,N_4942,N_4864);
nand UO_737 (O_737,N_4941,N_4832);
nor UO_738 (O_738,N_4842,N_4967);
or UO_739 (O_739,N_4806,N_4946);
and UO_740 (O_740,N_4888,N_4943);
nand UO_741 (O_741,N_4831,N_4943);
nand UO_742 (O_742,N_4995,N_4856);
nor UO_743 (O_743,N_4869,N_4856);
nor UO_744 (O_744,N_4826,N_4971);
nor UO_745 (O_745,N_4974,N_4923);
or UO_746 (O_746,N_4916,N_4804);
or UO_747 (O_747,N_4848,N_4832);
and UO_748 (O_748,N_4987,N_4980);
nor UO_749 (O_749,N_4950,N_4804);
nor UO_750 (O_750,N_4874,N_4839);
and UO_751 (O_751,N_4968,N_4913);
nand UO_752 (O_752,N_4896,N_4955);
nand UO_753 (O_753,N_4939,N_4914);
or UO_754 (O_754,N_4840,N_4974);
nor UO_755 (O_755,N_4937,N_4840);
and UO_756 (O_756,N_4906,N_4932);
or UO_757 (O_757,N_4970,N_4849);
and UO_758 (O_758,N_4826,N_4947);
nor UO_759 (O_759,N_4978,N_4882);
and UO_760 (O_760,N_4839,N_4988);
nand UO_761 (O_761,N_4904,N_4876);
or UO_762 (O_762,N_4964,N_4981);
nor UO_763 (O_763,N_4826,N_4852);
nand UO_764 (O_764,N_4874,N_4830);
and UO_765 (O_765,N_4886,N_4845);
and UO_766 (O_766,N_4886,N_4953);
and UO_767 (O_767,N_4954,N_4817);
nor UO_768 (O_768,N_4974,N_4960);
or UO_769 (O_769,N_4950,N_4973);
nor UO_770 (O_770,N_4987,N_4899);
nor UO_771 (O_771,N_4885,N_4968);
or UO_772 (O_772,N_4824,N_4895);
nor UO_773 (O_773,N_4995,N_4907);
nor UO_774 (O_774,N_4838,N_4879);
nor UO_775 (O_775,N_4982,N_4810);
or UO_776 (O_776,N_4924,N_4838);
and UO_777 (O_777,N_4828,N_4965);
nand UO_778 (O_778,N_4878,N_4992);
and UO_779 (O_779,N_4950,N_4884);
or UO_780 (O_780,N_4834,N_4891);
and UO_781 (O_781,N_4924,N_4979);
or UO_782 (O_782,N_4844,N_4899);
or UO_783 (O_783,N_4966,N_4826);
nand UO_784 (O_784,N_4812,N_4870);
or UO_785 (O_785,N_4840,N_4860);
or UO_786 (O_786,N_4820,N_4872);
nor UO_787 (O_787,N_4820,N_4948);
and UO_788 (O_788,N_4841,N_4871);
or UO_789 (O_789,N_4931,N_4871);
and UO_790 (O_790,N_4817,N_4900);
nand UO_791 (O_791,N_4915,N_4982);
nor UO_792 (O_792,N_4950,N_4993);
or UO_793 (O_793,N_4911,N_4865);
and UO_794 (O_794,N_4919,N_4922);
nor UO_795 (O_795,N_4842,N_4805);
nand UO_796 (O_796,N_4871,N_4986);
nand UO_797 (O_797,N_4924,N_4806);
or UO_798 (O_798,N_4862,N_4818);
or UO_799 (O_799,N_4964,N_4922);
or UO_800 (O_800,N_4979,N_4863);
and UO_801 (O_801,N_4963,N_4876);
nor UO_802 (O_802,N_4832,N_4813);
nand UO_803 (O_803,N_4802,N_4898);
and UO_804 (O_804,N_4910,N_4993);
nand UO_805 (O_805,N_4967,N_4975);
or UO_806 (O_806,N_4851,N_4914);
nor UO_807 (O_807,N_4909,N_4830);
nor UO_808 (O_808,N_4885,N_4913);
or UO_809 (O_809,N_4888,N_4988);
nor UO_810 (O_810,N_4908,N_4804);
or UO_811 (O_811,N_4915,N_4838);
nand UO_812 (O_812,N_4887,N_4960);
nand UO_813 (O_813,N_4858,N_4931);
nand UO_814 (O_814,N_4944,N_4991);
nand UO_815 (O_815,N_4896,N_4948);
nor UO_816 (O_816,N_4857,N_4819);
nor UO_817 (O_817,N_4870,N_4821);
nor UO_818 (O_818,N_4838,N_4846);
nor UO_819 (O_819,N_4829,N_4835);
nor UO_820 (O_820,N_4875,N_4886);
and UO_821 (O_821,N_4862,N_4836);
and UO_822 (O_822,N_4982,N_4821);
nor UO_823 (O_823,N_4936,N_4954);
and UO_824 (O_824,N_4856,N_4866);
xor UO_825 (O_825,N_4918,N_4910);
and UO_826 (O_826,N_4852,N_4806);
or UO_827 (O_827,N_4875,N_4997);
and UO_828 (O_828,N_4853,N_4992);
xor UO_829 (O_829,N_4800,N_4816);
nand UO_830 (O_830,N_4868,N_4993);
nor UO_831 (O_831,N_4947,N_4917);
nand UO_832 (O_832,N_4957,N_4937);
and UO_833 (O_833,N_4905,N_4949);
or UO_834 (O_834,N_4977,N_4964);
and UO_835 (O_835,N_4824,N_4963);
nand UO_836 (O_836,N_4897,N_4997);
xor UO_837 (O_837,N_4911,N_4940);
nor UO_838 (O_838,N_4967,N_4800);
and UO_839 (O_839,N_4891,N_4919);
and UO_840 (O_840,N_4834,N_4977);
nand UO_841 (O_841,N_4987,N_4918);
and UO_842 (O_842,N_4997,N_4916);
nand UO_843 (O_843,N_4955,N_4801);
and UO_844 (O_844,N_4956,N_4810);
nand UO_845 (O_845,N_4932,N_4876);
or UO_846 (O_846,N_4862,N_4884);
and UO_847 (O_847,N_4822,N_4911);
or UO_848 (O_848,N_4990,N_4977);
and UO_849 (O_849,N_4817,N_4806);
or UO_850 (O_850,N_4999,N_4839);
nand UO_851 (O_851,N_4918,N_4840);
or UO_852 (O_852,N_4910,N_4836);
nand UO_853 (O_853,N_4838,N_4905);
nand UO_854 (O_854,N_4865,N_4908);
or UO_855 (O_855,N_4924,N_4976);
or UO_856 (O_856,N_4989,N_4870);
nand UO_857 (O_857,N_4820,N_4913);
and UO_858 (O_858,N_4861,N_4998);
or UO_859 (O_859,N_4984,N_4872);
nand UO_860 (O_860,N_4808,N_4994);
nand UO_861 (O_861,N_4935,N_4818);
nor UO_862 (O_862,N_4982,N_4908);
and UO_863 (O_863,N_4938,N_4814);
nand UO_864 (O_864,N_4953,N_4969);
and UO_865 (O_865,N_4822,N_4956);
or UO_866 (O_866,N_4885,N_4843);
and UO_867 (O_867,N_4949,N_4802);
nand UO_868 (O_868,N_4892,N_4919);
and UO_869 (O_869,N_4874,N_4803);
nor UO_870 (O_870,N_4995,N_4827);
nor UO_871 (O_871,N_4959,N_4918);
and UO_872 (O_872,N_4968,N_4960);
nor UO_873 (O_873,N_4962,N_4987);
and UO_874 (O_874,N_4985,N_4886);
nand UO_875 (O_875,N_4919,N_4936);
or UO_876 (O_876,N_4858,N_4992);
or UO_877 (O_877,N_4832,N_4825);
nor UO_878 (O_878,N_4962,N_4829);
nor UO_879 (O_879,N_4895,N_4943);
and UO_880 (O_880,N_4819,N_4837);
and UO_881 (O_881,N_4901,N_4853);
or UO_882 (O_882,N_4907,N_4873);
nand UO_883 (O_883,N_4918,N_4968);
or UO_884 (O_884,N_4897,N_4918);
and UO_885 (O_885,N_4903,N_4879);
nor UO_886 (O_886,N_4854,N_4831);
nand UO_887 (O_887,N_4978,N_4857);
nor UO_888 (O_888,N_4847,N_4999);
nand UO_889 (O_889,N_4945,N_4946);
nor UO_890 (O_890,N_4906,N_4919);
nand UO_891 (O_891,N_4821,N_4941);
or UO_892 (O_892,N_4810,N_4830);
nand UO_893 (O_893,N_4813,N_4878);
or UO_894 (O_894,N_4945,N_4917);
or UO_895 (O_895,N_4919,N_4837);
nor UO_896 (O_896,N_4922,N_4913);
or UO_897 (O_897,N_4883,N_4899);
nor UO_898 (O_898,N_4904,N_4933);
or UO_899 (O_899,N_4961,N_4810);
and UO_900 (O_900,N_4863,N_4901);
and UO_901 (O_901,N_4881,N_4965);
nor UO_902 (O_902,N_4852,N_4998);
nand UO_903 (O_903,N_4813,N_4993);
nand UO_904 (O_904,N_4896,N_4808);
and UO_905 (O_905,N_4831,N_4895);
and UO_906 (O_906,N_4815,N_4838);
nor UO_907 (O_907,N_4955,N_4973);
and UO_908 (O_908,N_4818,N_4973);
and UO_909 (O_909,N_4833,N_4965);
and UO_910 (O_910,N_4956,N_4882);
and UO_911 (O_911,N_4855,N_4947);
nand UO_912 (O_912,N_4878,N_4921);
nor UO_913 (O_913,N_4953,N_4963);
nor UO_914 (O_914,N_4944,N_4983);
nor UO_915 (O_915,N_4830,N_4960);
nor UO_916 (O_916,N_4820,N_4876);
or UO_917 (O_917,N_4962,N_4976);
nand UO_918 (O_918,N_4870,N_4895);
nor UO_919 (O_919,N_4940,N_4835);
nand UO_920 (O_920,N_4976,N_4947);
nor UO_921 (O_921,N_4893,N_4836);
and UO_922 (O_922,N_4984,N_4812);
or UO_923 (O_923,N_4998,N_4891);
xnor UO_924 (O_924,N_4915,N_4856);
or UO_925 (O_925,N_4890,N_4811);
nor UO_926 (O_926,N_4944,N_4807);
nand UO_927 (O_927,N_4818,N_4848);
or UO_928 (O_928,N_4825,N_4879);
nor UO_929 (O_929,N_4964,N_4887);
and UO_930 (O_930,N_4885,N_4997);
nor UO_931 (O_931,N_4933,N_4938);
nand UO_932 (O_932,N_4908,N_4910);
nand UO_933 (O_933,N_4940,N_4815);
nor UO_934 (O_934,N_4904,N_4844);
nor UO_935 (O_935,N_4821,N_4967);
or UO_936 (O_936,N_4986,N_4888);
or UO_937 (O_937,N_4977,N_4895);
nor UO_938 (O_938,N_4864,N_4907);
nor UO_939 (O_939,N_4896,N_4860);
or UO_940 (O_940,N_4887,N_4832);
or UO_941 (O_941,N_4969,N_4920);
and UO_942 (O_942,N_4890,N_4856);
nand UO_943 (O_943,N_4931,N_4950);
or UO_944 (O_944,N_4858,N_4875);
and UO_945 (O_945,N_4813,N_4843);
nand UO_946 (O_946,N_4822,N_4837);
and UO_947 (O_947,N_4835,N_4896);
nand UO_948 (O_948,N_4808,N_4912);
or UO_949 (O_949,N_4954,N_4929);
nand UO_950 (O_950,N_4952,N_4812);
nand UO_951 (O_951,N_4869,N_4890);
and UO_952 (O_952,N_4864,N_4971);
nand UO_953 (O_953,N_4868,N_4952);
nand UO_954 (O_954,N_4810,N_4842);
or UO_955 (O_955,N_4880,N_4907);
and UO_956 (O_956,N_4908,N_4983);
nor UO_957 (O_957,N_4895,N_4842);
and UO_958 (O_958,N_4835,N_4820);
and UO_959 (O_959,N_4845,N_4874);
and UO_960 (O_960,N_4979,N_4833);
and UO_961 (O_961,N_4955,N_4974);
nor UO_962 (O_962,N_4993,N_4917);
nand UO_963 (O_963,N_4825,N_4941);
nor UO_964 (O_964,N_4900,N_4960);
nand UO_965 (O_965,N_4936,N_4823);
and UO_966 (O_966,N_4926,N_4868);
nand UO_967 (O_967,N_4909,N_4960);
nand UO_968 (O_968,N_4826,N_4918);
nand UO_969 (O_969,N_4895,N_4885);
nor UO_970 (O_970,N_4821,N_4868);
and UO_971 (O_971,N_4899,N_4904);
or UO_972 (O_972,N_4848,N_4966);
nand UO_973 (O_973,N_4939,N_4852);
nor UO_974 (O_974,N_4941,N_4930);
nor UO_975 (O_975,N_4923,N_4897);
nand UO_976 (O_976,N_4944,N_4868);
or UO_977 (O_977,N_4839,N_4876);
nand UO_978 (O_978,N_4853,N_4899);
or UO_979 (O_979,N_4858,N_4887);
nor UO_980 (O_980,N_4870,N_4852);
and UO_981 (O_981,N_4906,N_4903);
nor UO_982 (O_982,N_4906,N_4927);
or UO_983 (O_983,N_4930,N_4949);
nand UO_984 (O_984,N_4976,N_4826);
or UO_985 (O_985,N_4909,N_4951);
or UO_986 (O_986,N_4801,N_4914);
or UO_987 (O_987,N_4909,N_4913);
and UO_988 (O_988,N_4951,N_4852);
nand UO_989 (O_989,N_4856,N_4904);
nand UO_990 (O_990,N_4956,N_4835);
and UO_991 (O_991,N_4910,N_4941);
nor UO_992 (O_992,N_4986,N_4861);
nor UO_993 (O_993,N_4991,N_4823);
nand UO_994 (O_994,N_4911,N_4840);
or UO_995 (O_995,N_4811,N_4834);
and UO_996 (O_996,N_4902,N_4906);
or UO_997 (O_997,N_4969,N_4897);
or UO_998 (O_998,N_4908,N_4905);
nor UO_999 (O_999,N_4932,N_4980);
endmodule