module basic_500_3000_500_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_52,In_404);
or U1 (N_1,In_376,In_296);
xnor U2 (N_2,In_108,In_110);
nand U3 (N_3,In_143,In_364);
and U4 (N_4,In_193,In_304);
and U5 (N_5,In_178,In_334);
nor U6 (N_6,In_139,In_244);
or U7 (N_7,In_17,In_74);
xor U8 (N_8,In_4,In_175);
nand U9 (N_9,In_303,In_202);
or U10 (N_10,In_323,In_236);
and U11 (N_11,In_148,In_430);
nand U12 (N_12,In_242,In_200);
nor U13 (N_13,In_109,In_125);
nand U14 (N_14,In_26,In_185);
xor U15 (N_15,In_259,In_232);
or U16 (N_16,In_499,In_219);
or U17 (N_17,In_497,In_260);
xnor U18 (N_18,In_402,In_336);
and U19 (N_19,In_186,In_136);
and U20 (N_20,In_373,In_162);
and U21 (N_21,In_37,In_25);
nand U22 (N_22,In_179,In_133);
xor U23 (N_23,In_152,In_89);
or U24 (N_24,In_115,In_121);
nand U25 (N_25,In_150,In_187);
nor U26 (N_26,In_378,In_463);
nand U27 (N_27,In_341,In_226);
xnor U28 (N_28,In_312,In_167);
xor U29 (N_29,In_331,In_380);
nor U30 (N_30,In_149,In_411);
nand U31 (N_31,In_194,In_469);
and U32 (N_32,In_72,In_158);
or U33 (N_33,In_263,In_9);
or U34 (N_34,In_225,In_145);
xor U35 (N_35,In_118,In_488);
xnor U36 (N_36,In_64,In_366);
nor U37 (N_37,In_416,In_16);
or U38 (N_38,In_486,In_410);
and U39 (N_39,In_38,In_473);
and U40 (N_40,In_314,In_7);
or U41 (N_41,In_395,In_298);
xor U42 (N_42,In_338,In_199);
nand U43 (N_43,In_113,In_262);
nor U44 (N_44,In_285,In_195);
nor U45 (N_45,In_326,In_28);
xor U46 (N_46,In_0,In_377);
nand U47 (N_47,In_83,In_127);
or U48 (N_48,In_292,In_392);
xor U49 (N_49,In_135,In_138);
nand U50 (N_50,In_434,In_413);
xnor U51 (N_51,In_224,In_360);
nand U52 (N_52,In_264,In_478);
and U53 (N_53,In_196,In_169);
nand U54 (N_54,In_154,In_254);
and U55 (N_55,In_151,In_69);
nor U56 (N_56,In_293,In_95);
and U57 (N_57,In_126,In_464);
xor U58 (N_58,In_405,In_182);
nand U59 (N_59,In_307,In_198);
or U60 (N_60,In_12,In_370);
nor U61 (N_61,In_471,N_20);
or U62 (N_62,In_197,In_278);
or U63 (N_63,In_99,In_493);
xnor U64 (N_64,In_369,In_129);
nand U65 (N_65,In_163,N_9);
nand U66 (N_66,N_13,In_213);
xor U67 (N_67,In_368,In_1);
nor U68 (N_68,In_418,In_170);
xor U69 (N_69,In_494,In_306);
or U70 (N_70,In_454,In_86);
and U71 (N_71,In_300,In_447);
xnor U72 (N_72,N_1,In_273);
and U73 (N_73,In_290,In_205);
or U74 (N_74,In_257,N_29);
nor U75 (N_75,N_57,In_192);
xor U76 (N_76,In_371,N_34);
nor U77 (N_77,In_267,N_0);
xnor U78 (N_78,In_428,In_209);
nor U79 (N_79,N_12,In_45);
and U80 (N_80,In_6,In_282);
and U81 (N_81,In_382,In_82);
nand U82 (N_82,In_350,In_498);
nor U83 (N_83,In_496,In_311);
nand U84 (N_84,In_355,In_98);
nor U85 (N_85,In_365,In_270);
xor U86 (N_86,In_91,In_190);
nand U87 (N_87,In_33,In_207);
or U88 (N_88,In_452,In_183);
nor U89 (N_89,In_36,In_397);
and U90 (N_90,In_217,In_39);
or U91 (N_91,In_495,In_246);
xnor U92 (N_92,In_344,N_39);
or U93 (N_93,In_31,In_385);
or U94 (N_94,N_17,In_329);
or U95 (N_95,In_315,In_295);
and U96 (N_96,In_432,In_346);
and U97 (N_97,In_318,In_436);
xor U98 (N_98,In_310,In_445);
and U99 (N_99,In_431,N_40);
and U100 (N_100,In_42,In_208);
nor U101 (N_101,In_339,In_168);
and U102 (N_102,In_173,In_287);
or U103 (N_103,In_362,In_122);
nand U104 (N_104,N_48,N_47);
and U105 (N_105,In_32,In_441);
or U106 (N_106,In_288,In_24);
xor U107 (N_107,In_390,N_45);
nor U108 (N_108,In_316,In_337);
nor U109 (N_109,In_424,In_41);
xnor U110 (N_110,In_490,In_132);
and U111 (N_111,N_2,In_375);
nor U112 (N_112,In_457,In_119);
or U113 (N_113,In_22,In_415);
nor U114 (N_114,In_321,In_313);
xor U115 (N_115,In_130,In_363);
nand U116 (N_116,In_446,In_101);
nor U117 (N_117,N_53,In_105);
or U118 (N_118,In_420,N_42);
nor U119 (N_119,In_201,In_5);
or U120 (N_120,In_348,In_358);
xnor U121 (N_121,In_8,In_230);
xor U122 (N_122,N_86,N_5);
and U123 (N_123,In_51,N_51);
or U124 (N_124,In_189,In_367);
or U125 (N_125,N_24,N_31);
and U126 (N_126,In_250,In_79);
or U127 (N_127,N_30,N_11);
xor U128 (N_128,N_65,N_98);
nand U129 (N_129,In_171,In_409);
or U130 (N_130,In_332,N_90);
and U131 (N_131,In_164,In_184);
xnor U132 (N_132,In_393,In_492);
nor U133 (N_133,In_309,In_455);
nor U134 (N_134,In_399,In_210);
nor U135 (N_135,In_212,N_7);
nand U136 (N_136,In_123,In_137);
nor U137 (N_137,N_62,In_439);
xor U138 (N_138,In_88,N_89);
and U139 (N_139,N_107,In_353);
xnor U140 (N_140,N_43,In_342);
or U141 (N_141,In_271,N_21);
nand U142 (N_142,In_426,In_90);
and U143 (N_143,In_396,In_94);
and U144 (N_144,N_16,In_87);
xor U145 (N_145,In_57,In_403);
and U146 (N_146,In_67,In_423);
xnor U147 (N_147,N_63,In_448);
nor U148 (N_148,In_477,N_116);
nand U149 (N_149,In_361,In_357);
or U150 (N_150,In_10,In_65);
nor U151 (N_151,In_317,In_13);
xnor U152 (N_152,In_21,In_484);
xnor U153 (N_153,In_256,In_84);
nand U154 (N_154,N_83,In_44);
and U155 (N_155,In_35,In_475);
or U156 (N_156,In_466,In_245);
and U157 (N_157,In_291,In_379);
and U158 (N_158,In_425,In_120);
nor U159 (N_159,In_359,In_29);
nor U160 (N_160,In_252,N_108);
and U161 (N_161,N_71,In_241);
nor U162 (N_162,In_374,In_289);
or U163 (N_163,In_414,N_87);
and U164 (N_164,N_102,In_156);
nor U165 (N_165,In_134,In_220);
nand U166 (N_166,In_474,In_104);
nor U167 (N_167,In_258,In_117);
nor U168 (N_168,N_95,In_147);
nor U169 (N_169,In_294,In_100);
xor U170 (N_170,In_215,In_20);
nor U171 (N_171,In_166,In_461);
xnor U172 (N_172,N_113,In_297);
and U173 (N_173,In_153,In_319);
xor U174 (N_174,In_48,In_372);
or U175 (N_175,In_333,In_284);
and U176 (N_176,In_49,N_93);
or U177 (N_177,In_235,In_479);
nor U178 (N_178,N_32,N_35);
xor U179 (N_179,N_111,N_73);
and U180 (N_180,In_324,In_2);
or U181 (N_181,In_470,In_406);
and U182 (N_182,In_255,N_50);
nand U183 (N_183,N_55,In_349);
and U184 (N_184,N_161,N_69);
or U185 (N_185,In_216,In_203);
xnor U186 (N_186,In_155,In_141);
or U187 (N_187,In_459,In_177);
and U188 (N_188,N_68,In_320);
xnor U189 (N_189,In_352,N_27);
or U190 (N_190,In_60,N_125);
nand U191 (N_191,N_18,N_146);
nand U192 (N_192,N_159,N_64);
and U193 (N_193,In_174,In_161);
and U194 (N_194,In_146,In_407);
or U195 (N_195,In_47,In_62);
nand U196 (N_196,N_56,In_421);
nor U197 (N_197,N_52,N_143);
or U198 (N_198,N_166,N_96);
nand U199 (N_199,In_322,N_74);
or U200 (N_200,In_237,N_115);
and U201 (N_201,N_114,In_160);
nand U202 (N_202,In_266,In_66);
nor U203 (N_203,In_46,N_91);
or U204 (N_204,In_61,In_325);
or U205 (N_205,N_38,N_132);
and U206 (N_206,N_80,In_299);
or U207 (N_207,In_176,In_180);
nor U208 (N_208,N_58,N_106);
or U209 (N_209,In_480,N_127);
and U210 (N_210,In_54,N_19);
or U211 (N_211,N_41,N_104);
or U212 (N_212,In_472,N_141);
or U213 (N_213,N_110,In_383);
and U214 (N_214,In_222,In_18);
nand U215 (N_215,In_56,N_4);
xnor U216 (N_216,In_356,In_78);
xnor U217 (N_217,In_240,In_327);
nand U218 (N_218,N_28,N_179);
xor U219 (N_219,N_148,In_116);
nand U220 (N_220,N_67,N_178);
xnor U221 (N_221,In_112,N_167);
or U222 (N_222,N_8,N_3);
and U223 (N_223,In_451,N_151);
xor U224 (N_224,In_223,In_412);
or U225 (N_225,In_305,N_36);
nor U226 (N_226,In_443,In_131);
or U227 (N_227,N_155,In_302);
and U228 (N_228,In_481,In_63);
xor U229 (N_229,In_280,In_238);
or U230 (N_230,In_485,In_283);
and U231 (N_231,In_106,In_308);
and U232 (N_232,In_144,In_191);
nand U233 (N_233,N_79,In_30);
and U234 (N_234,In_111,N_153);
or U235 (N_235,In_233,In_400);
and U236 (N_236,In_347,In_261);
nor U237 (N_237,N_145,In_231);
xnor U238 (N_238,In_59,In_437);
and U239 (N_239,In_75,N_162);
xnor U240 (N_240,N_165,In_85);
and U241 (N_241,N_235,In_343);
nor U242 (N_242,In_398,In_427);
or U243 (N_243,In_387,In_142);
nand U244 (N_244,N_81,N_149);
nor U245 (N_245,N_233,N_219);
xnor U246 (N_246,N_97,N_238);
or U247 (N_247,N_228,N_208);
or U248 (N_248,In_204,In_71);
nor U249 (N_249,In_58,N_195);
or U250 (N_250,In_476,In_442);
nor U251 (N_251,In_124,In_269);
xnor U252 (N_252,In_456,In_19);
or U253 (N_253,N_88,In_279);
xor U254 (N_254,In_458,N_198);
or U255 (N_255,N_72,In_43);
xnor U256 (N_256,N_15,In_340);
or U257 (N_257,In_408,In_330);
nand U258 (N_258,In_468,In_11);
and U259 (N_259,N_25,N_211);
and U260 (N_260,In_328,In_429);
and U261 (N_261,N_144,N_139);
nand U262 (N_262,N_123,N_122);
xor U263 (N_263,In_14,In_301);
xor U264 (N_264,N_78,N_158);
or U265 (N_265,N_221,N_168);
or U266 (N_266,N_152,In_249);
or U267 (N_267,N_6,In_247);
and U268 (N_268,In_114,N_225);
or U269 (N_269,N_186,In_53);
nor U270 (N_270,N_231,N_202);
or U271 (N_271,In_419,N_207);
or U272 (N_272,N_142,In_73);
and U273 (N_273,N_212,N_109);
nor U274 (N_274,In_276,N_164);
nand U275 (N_275,N_147,In_417);
xor U276 (N_276,N_171,In_234);
and U277 (N_277,In_391,N_176);
and U278 (N_278,In_70,N_130);
xor U279 (N_279,In_335,N_224);
or U280 (N_280,In_40,N_183);
or U281 (N_281,N_120,N_157);
and U282 (N_282,In_34,In_450);
or U283 (N_283,N_234,N_10);
nor U284 (N_284,In_218,N_121);
nor U285 (N_285,In_97,N_70);
nand U286 (N_286,In_55,N_205);
xnor U287 (N_287,N_173,In_384);
or U288 (N_288,N_134,N_99);
or U289 (N_289,N_94,N_100);
and U290 (N_290,N_75,In_462);
xnor U291 (N_291,In_286,In_487);
and U292 (N_292,In_76,N_226);
or U293 (N_293,N_22,N_37);
nor U294 (N_294,N_215,N_49);
or U295 (N_295,N_101,In_277);
nand U296 (N_296,N_223,N_118);
nor U297 (N_297,In_228,In_433);
nor U298 (N_298,In_438,In_206);
xor U299 (N_299,In_211,In_435);
xnor U300 (N_300,N_210,In_248);
or U301 (N_301,In_23,N_266);
and U302 (N_302,N_252,N_281);
and U303 (N_303,N_26,In_27);
xor U304 (N_304,In_465,In_351);
or U305 (N_305,In_268,N_61);
nand U306 (N_306,In_401,In_394);
and U307 (N_307,N_203,N_277);
and U308 (N_308,In_93,N_77);
xnor U309 (N_309,N_59,In_265);
and U310 (N_310,N_256,N_267);
nor U311 (N_311,N_206,N_60);
or U312 (N_312,N_175,N_135);
nor U313 (N_313,N_84,N_290);
or U314 (N_314,N_216,In_15);
and U315 (N_315,N_82,In_68);
xor U316 (N_316,N_163,N_112);
and U317 (N_317,N_258,N_156);
nor U318 (N_318,N_263,N_292);
and U319 (N_319,N_214,In_103);
nor U320 (N_320,N_275,N_180);
xor U321 (N_321,In_157,N_220);
and U322 (N_322,In_422,In_128);
and U323 (N_323,N_222,N_237);
or U324 (N_324,N_131,N_295);
or U325 (N_325,N_247,In_251);
and U326 (N_326,N_193,In_389);
nor U327 (N_327,In_491,N_23);
xor U328 (N_328,N_272,N_188);
nand U329 (N_329,N_76,N_260);
nand U330 (N_330,N_288,N_299);
and U331 (N_331,N_264,N_248);
or U332 (N_332,In_281,In_77);
xor U333 (N_333,N_199,In_275);
xor U334 (N_334,N_181,N_269);
or U335 (N_335,In_140,N_191);
or U336 (N_336,N_279,In_221);
and U337 (N_337,N_133,N_66);
and U338 (N_338,In_274,N_204);
nor U339 (N_339,In_102,N_189);
or U340 (N_340,In_460,N_259);
or U341 (N_341,N_297,N_246);
and U342 (N_342,N_194,In_482);
nand U343 (N_343,N_296,N_271);
nand U344 (N_344,N_250,N_241);
or U345 (N_345,N_150,N_140);
nor U346 (N_346,N_154,N_255);
and U347 (N_347,N_124,N_282);
nand U348 (N_348,N_137,In_386);
xnor U349 (N_349,N_117,N_197);
or U350 (N_350,N_44,N_240);
or U351 (N_351,N_92,N_265);
or U352 (N_352,N_242,N_177);
nand U353 (N_353,N_229,N_249);
nor U354 (N_354,In_229,In_381);
or U355 (N_355,N_239,In_81);
xnor U356 (N_356,N_105,N_291);
nand U357 (N_357,In_467,N_293);
and U358 (N_358,N_126,N_244);
and U359 (N_359,In_253,N_268);
nor U360 (N_360,N_236,N_253);
nand U361 (N_361,N_322,N_230);
and U362 (N_362,In_483,N_276);
nor U363 (N_363,N_317,N_232);
nor U364 (N_364,N_320,N_289);
and U365 (N_365,In_440,N_345);
and U366 (N_366,N_326,N_333);
or U367 (N_367,In_188,N_329);
and U368 (N_368,In_181,N_184);
nor U369 (N_369,N_262,N_358);
and U370 (N_370,N_160,N_330);
or U371 (N_371,N_261,N_287);
and U372 (N_372,N_301,N_351);
nor U373 (N_373,N_316,N_332);
nand U374 (N_374,N_33,N_217);
xor U375 (N_375,N_339,N_85);
and U376 (N_376,N_14,In_227);
nor U377 (N_377,N_218,N_182);
nor U378 (N_378,N_304,N_346);
nand U379 (N_379,N_319,N_314);
xnor U380 (N_380,N_170,In_354);
xnor U381 (N_381,N_318,N_300);
and U382 (N_382,N_348,In_3);
nand U383 (N_383,In_243,N_283);
xor U384 (N_384,N_336,N_356);
nor U385 (N_385,N_270,N_103);
nand U386 (N_386,N_285,N_328);
nor U387 (N_387,N_303,N_306);
nand U388 (N_388,N_187,In_172);
xnor U389 (N_389,In_80,In_239);
nor U390 (N_390,N_196,In_453);
xor U391 (N_391,N_343,N_129);
and U392 (N_392,In_96,N_185);
nand U393 (N_393,N_46,N_298);
or U394 (N_394,N_355,In_489);
nor U395 (N_395,N_350,In_449);
xor U396 (N_396,N_338,N_136);
and U397 (N_397,In_159,N_313);
or U398 (N_398,N_257,N_344);
nor U399 (N_399,N_327,N_335);
nor U400 (N_400,N_315,N_352);
nor U401 (N_401,N_245,N_128);
nor U402 (N_402,N_353,N_357);
nand U403 (N_403,N_349,N_169);
xnor U404 (N_404,In_214,N_280);
nand U405 (N_405,N_324,N_331);
xor U406 (N_406,N_359,N_174);
or U407 (N_407,N_172,N_200);
and U408 (N_408,N_337,In_165);
and U409 (N_409,In_107,N_323);
nor U410 (N_410,N_119,N_321);
xnor U411 (N_411,N_278,N_308);
nor U412 (N_412,N_284,N_138);
or U413 (N_413,N_310,N_274);
nand U414 (N_414,N_54,N_286);
nor U415 (N_415,N_311,N_273);
nand U416 (N_416,N_347,N_243);
nand U417 (N_417,N_227,N_254);
and U418 (N_418,N_190,In_272);
and U419 (N_419,N_302,In_92);
xor U420 (N_420,N_366,N_385);
nand U421 (N_421,N_201,N_402);
xnor U422 (N_422,N_391,N_341);
and U423 (N_423,N_370,N_192);
and U424 (N_424,N_384,N_379);
and U425 (N_425,N_367,N_375);
or U426 (N_426,N_363,N_389);
xnor U427 (N_427,N_213,In_388);
nand U428 (N_428,N_403,N_312);
nand U429 (N_429,In_444,N_354);
or U430 (N_430,N_209,N_373);
nor U431 (N_431,N_342,N_399);
nand U432 (N_432,N_396,N_418);
xnor U433 (N_433,N_368,N_380);
nor U434 (N_434,N_390,In_50);
xnor U435 (N_435,N_360,N_393);
xnor U436 (N_436,N_410,N_309);
or U437 (N_437,N_294,N_400);
or U438 (N_438,N_305,N_334);
nor U439 (N_439,N_411,N_415);
and U440 (N_440,N_417,N_419);
and U441 (N_441,N_374,N_407);
nand U442 (N_442,N_372,N_377);
nand U443 (N_443,N_408,N_371);
nor U444 (N_444,N_387,N_381);
nor U445 (N_445,N_369,N_414);
nand U446 (N_446,N_386,N_406);
nand U447 (N_447,N_405,N_325);
or U448 (N_448,N_397,N_392);
or U449 (N_449,N_382,N_412);
nor U450 (N_450,N_376,N_365);
and U451 (N_451,N_383,N_395);
nor U452 (N_452,N_362,N_251);
and U453 (N_453,N_409,In_345);
nor U454 (N_454,N_388,N_413);
xnor U455 (N_455,N_307,N_340);
xor U456 (N_456,N_398,N_364);
xor U457 (N_457,N_378,N_401);
nor U458 (N_458,N_394,N_361);
and U459 (N_459,N_416,N_404);
or U460 (N_460,N_393,N_377);
xor U461 (N_461,N_341,N_395);
or U462 (N_462,N_418,N_392);
nand U463 (N_463,N_380,N_307);
and U464 (N_464,N_401,N_368);
or U465 (N_465,N_192,N_383);
nor U466 (N_466,N_399,N_389);
nand U467 (N_467,N_395,N_385);
nand U468 (N_468,N_309,N_400);
nor U469 (N_469,N_374,N_411);
xor U470 (N_470,N_367,N_383);
nor U471 (N_471,N_367,N_392);
and U472 (N_472,N_412,N_390);
xor U473 (N_473,N_405,N_192);
and U474 (N_474,N_395,In_444);
and U475 (N_475,N_385,N_362);
nor U476 (N_476,N_395,N_379);
nor U477 (N_477,N_418,N_379);
xnor U478 (N_478,N_378,N_366);
xnor U479 (N_479,N_363,N_401);
nand U480 (N_480,N_452,N_466);
xnor U481 (N_481,N_448,N_430);
xnor U482 (N_482,N_425,N_443);
nor U483 (N_483,N_463,N_453);
nor U484 (N_484,N_437,N_461);
nand U485 (N_485,N_473,N_460);
and U486 (N_486,N_465,N_462);
nand U487 (N_487,N_434,N_428);
or U488 (N_488,N_464,N_474);
or U489 (N_489,N_420,N_468);
xor U490 (N_490,N_433,N_471);
or U491 (N_491,N_477,N_458);
nand U492 (N_492,N_442,N_459);
and U493 (N_493,N_472,N_470);
and U494 (N_494,N_436,N_421);
nor U495 (N_495,N_467,N_440);
nand U496 (N_496,N_479,N_432);
or U497 (N_497,N_445,N_438);
and U498 (N_498,N_457,N_431);
and U499 (N_499,N_429,N_478);
xor U500 (N_500,N_426,N_456);
nand U501 (N_501,N_427,N_449);
or U502 (N_502,N_435,N_455);
and U503 (N_503,N_454,N_446);
nor U504 (N_504,N_450,N_424);
nor U505 (N_505,N_444,N_451);
and U506 (N_506,N_475,N_476);
nand U507 (N_507,N_441,N_422);
and U508 (N_508,N_447,N_423);
nand U509 (N_509,N_469,N_439);
nor U510 (N_510,N_429,N_449);
nor U511 (N_511,N_424,N_436);
nand U512 (N_512,N_428,N_457);
and U513 (N_513,N_427,N_452);
xnor U514 (N_514,N_459,N_477);
and U515 (N_515,N_421,N_458);
and U516 (N_516,N_424,N_472);
or U517 (N_517,N_472,N_469);
xnor U518 (N_518,N_444,N_426);
or U519 (N_519,N_452,N_425);
or U520 (N_520,N_466,N_437);
or U521 (N_521,N_440,N_436);
and U522 (N_522,N_457,N_455);
nand U523 (N_523,N_424,N_439);
nor U524 (N_524,N_435,N_424);
xor U525 (N_525,N_465,N_421);
nor U526 (N_526,N_445,N_461);
or U527 (N_527,N_463,N_456);
and U528 (N_528,N_428,N_460);
and U529 (N_529,N_441,N_465);
or U530 (N_530,N_426,N_440);
xor U531 (N_531,N_464,N_459);
xor U532 (N_532,N_464,N_436);
or U533 (N_533,N_471,N_447);
nor U534 (N_534,N_464,N_468);
and U535 (N_535,N_436,N_479);
xnor U536 (N_536,N_433,N_472);
or U537 (N_537,N_445,N_451);
nand U538 (N_538,N_453,N_433);
xnor U539 (N_539,N_426,N_476);
and U540 (N_540,N_493,N_501);
nor U541 (N_541,N_515,N_496);
nand U542 (N_542,N_536,N_534);
and U543 (N_543,N_488,N_500);
or U544 (N_544,N_513,N_516);
nor U545 (N_545,N_504,N_522);
and U546 (N_546,N_507,N_505);
nand U547 (N_547,N_517,N_518);
nand U548 (N_548,N_485,N_537);
nor U549 (N_549,N_482,N_486);
and U550 (N_550,N_512,N_526);
nand U551 (N_551,N_494,N_511);
xnor U552 (N_552,N_495,N_519);
or U553 (N_553,N_527,N_524);
and U554 (N_554,N_484,N_509);
and U555 (N_555,N_490,N_531);
and U556 (N_556,N_525,N_508);
nor U557 (N_557,N_491,N_492);
and U558 (N_558,N_497,N_481);
nor U559 (N_559,N_523,N_529);
and U560 (N_560,N_480,N_532);
and U561 (N_561,N_483,N_535);
nand U562 (N_562,N_528,N_521);
xor U563 (N_563,N_538,N_539);
xor U564 (N_564,N_502,N_487);
nand U565 (N_565,N_520,N_503);
nor U566 (N_566,N_506,N_530);
or U567 (N_567,N_489,N_499);
or U568 (N_568,N_498,N_510);
or U569 (N_569,N_533,N_514);
or U570 (N_570,N_493,N_504);
xnor U571 (N_571,N_518,N_490);
xor U572 (N_572,N_528,N_501);
xnor U573 (N_573,N_512,N_536);
xor U574 (N_574,N_526,N_506);
and U575 (N_575,N_518,N_537);
xnor U576 (N_576,N_524,N_512);
xnor U577 (N_577,N_526,N_532);
xor U578 (N_578,N_509,N_518);
nor U579 (N_579,N_495,N_530);
or U580 (N_580,N_518,N_531);
or U581 (N_581,N_500,N_519);
nand U582 (N_582,N_510,N_493);
xnor U583 (N_583,N_517,N_503);
nand U584 (N_584,N_507,N_491);
and U585 (N_585,N_510,N_505);
or U586 (N_586,N_519,N_506);
xnor U587 (N_587,N_502,N_482);
or U588 (N_588,N_517,N_530);
nor U589 (N_589,N_503,N_488);
nand U590 (N_590,N_510,N_516);
and U591 (N_591,N_501,N_532);
xor U592 (N_592,N_505,N_529);
nor U593 (N_593,N_537,N_514);
nand U594 (N_594,N_518,N_529);
and U595 (N_595,N_492,N_533);
nor U596 (N_596,N_527,N_501);
xor U597 (N_597,N_535,N_515);
nor U598 (N_598,N_493,N_483);
or U599 (N_599,N_495,N_517);
and U600 (N_600,N_598,N_570);
nand U601 (N_601,N_589,N_549);
nand U602 (N_602,N_546,N_561);
nor U603 (N_603,N_556,N_550);
nand U604 (N_604,N_588,N_566);
nor U605 (N_605,N_596,N_585);
or U606 (N_606,N_583,N_593);
nand U607 (N_607,N_599,N_548);
nand U608 (N_608,N_562,N_554);
xor U609 (N_609,N_595,N_592);
nand U610 (N_610,N_547,N_577);
and U611 (N_611,N_568,N_563);
and U612 (N_612,N_564,N_591);
xor U613 (N_613,N_571,N_572);
nor U614 (N_614,N_544,N_575);
nand U615 (N_615,N_545,N_555);
or U616 (N_616,N_594,N_579);
nor U617 (N_617,N_576,N_582);
nor U618 (N_618,N_541,N_569);
nor U619 (N_619,N_578,N_590);
nand U620 (N_620,N_586,N_597);
nor U621 (N_621,N_580,N_543);
or U622 (N_622,N_551,N_584);
and U623 (N_623,N_565,N_558);
xor U624 (N_624,N_553,N_552);
and U625 (N_625,N_574,N_557);
nor U626 (N_626,N_573,N_542);
xor U627 (N_627,N_587,N_560);
and U628 (N_628,N_540,N_567);
xnor U629 (N_629,N_559,N_581);
nor U630 (N_630,N_580,N_569);
nor U631 (N_631,N_582,N_578);
nand U632 (N_632,N_592,N_575);
xor U633 (N_633,N_552,N_559);
nand U634 (N_634,N_555,N_582);
nor U635 (N_635,N_585,N_599);
xor U636 (N_636,N_543,N_578);
and U637 (N_637,N_540,N_549);
nor U638 (N_638,N_540,N_562);
or U639 (N_639,N_577,N_572);
nor U640 (N_640,N_551,N_567);
nand U641 (N_641,N_551,N_548);
nor U642 (N_642,N_594,N_546);
or U643 (N_643,N_545,N_556);
xnor U644 (N_644,N_550,N_588);
and U645 (N_645,N_569,N_592);
and U646 (N_646,N_599,N_595);
nor U647 (N_647,N_597,N_579);
nand U648 (N_648,N_576,N_570);
or U649 (N_649,N_545,N_562);
and U650 (N_650,N_569,N_586);
nor U651 (N_651,N_592,N_544);
and U652 (N_652,N_591,N_577);
xor U653 (N_653,N_569,N_574);
nor U654 (N_654,N_581,N_552);
and U655 (N_655,N_589,N_551);
xor U656 (N_656,N_560,N_568);
nand U657 (N_657,N_553,N_591);
and U658 (N_658,N_554,N_598);
and U659 (N_659,N_558,N_563);
and U660 (N_660,N_615,N_651);
and U661 (N_661,N_637,N_652);
xnor U662 (N_662,N_648,N_626);
xor U663 (N_663,N_603,N_630);
nand U664 (N_664,N_625,N_613);
and U665 (N_665,N_617,N_607);
nor U666 (N_666,N_653,N_632);
and U667 (N_667,N_643,N_611);
xor U668 (N_668,N_606,N_658);
or U669 (N_669,N_620,N_650);
nand U670 (N_670,N_608,N_654);
or U671 (N_671,N_639,N_619);
or U672 (N_672,N_647,N_640);
nand U673 (N_673,N_610,N_621);
and U674 (N_674,N_656,N_635);
and U675 (N_675,N_601,N_636);
and U676 (N_676,N_605,N_641);
nor U677 (N_677,N_629,N_602);
and U678 (N_678,N_657,N_659);
nor U679 (N_679,N_638,N_609);
nand U680 (N_680,N_618,N_614);
nand U681 (N_681,N_600,N_622);
and U682 (N_682,N_649,N_604);
or U683 (N_683,N_631,N_633);
and U684 (N_684,N_616,N_646);
nor U685 (N_685,N_624,N_645);
nor U686 (N_686,N_627,N_623);
nand U687 (N_687,N_628,N_642);
nor U688 (N_688,N_644,N_634);
xnor U689 (N_689,N_612,N_655);
or U690 (N_690,N_609,N_607);
or U691 (N_691,N_626,N_653);
or U692 (N_692,N_632,N_617);
nor U693 (N_693,N_613,N_626);
nand U694 (N_694,N_650,N_603);
nor U695 (N_695,N_631,N_607);
nand U696 (N_696,N_606,N_624);
or U697 (N_697,N_641,N_658);
nor U698 (N_698,N_625,N_640);
and U699 (N_699,N_656,N_602);
and U700 (N_700,N_618,N_608);
or U701 (N_701,N_634,N_623);
xnor U702 (N_702,N_625,N_647);
or U703 (N_703,N_638,N_619);
or U704 (N_704,N_646,N_621);
xnor U705 (N_705,N_635,N_639);
nor U706 (N_706,N_637,N_655);
nand U707 (N_707,N_635,N_624);
nor U708 (N_708,N_623,N_630);
xor U709 (N_709,N_602,N_658);
nor U710 (N_710,N_641,N_602);
xor U711 (N_711,N_625,N_624);
xnor U712 (N_712,N_638,N_604);
xor U713 (N_713,N_614,N_606);
nand U714 (N_714,N_618,N_640);
nand U715 (N_715,N_611,N_623);
xnor U716 (N_716,N_630,N_628);
or U717 (N_717,N_612,N_645);
and U718 (N_718,N_647,N_604);
nand U719 (N_719,N_617,N_608);
nor U720 (N_720,N_669,N_701);
or U721 (N_721,N_688,N_706);
or U722 (N_722,N_686,N_711);
nor U723 (N_723,N_698,N_677);
nand U724 (N_724,N_687,N_708);
nand U725 (N_725,N_667,N_666);
and U726 (N_726,N_704,N_676);
nand U727 (N_727,N_702,N_714);
or U728 (N_728,N_699,N_705);
xor U729 (N_729,N_709,N_695);
nand U730 (N_730,N_678,N_681);
nor U731 (N_731,N_717,N_719);
and U732 (N_732,N_715,N_692);
and U733 (N_733,N_684,N_703);
nand U734 (N_734,N_697,N_690);
nand U735 (N_735,N_668,N_683);
nand U736 (N_736,N_700,N_679);
nand U737 (N_737,N_663,N_660);
nand U738 (N_738,N_689,N_691);
xor U739 (N_739,N_670,N_696);
or U740 (N_740,N_682,N_713);
nor U741 (N_741,N_685,N_680);
xnor U742 (N_742,N_662,N_675);
nor U743 (N_743,N_671,N_694);
xnor U744 (N_744,N_665,N_672);
nand U745 (N_745,N_710,N_674);
and U746 (N_746,N_716,N_693);
xnor U747 (N_747,N_664,N_712);
xnor U748 (N_748,N_718,N_661);
or U749 (N_749,N_673,N_707);
and U750 (N_750,N_672,N_674);
nand U751 (N_751,N_714,N_701);
nor U752 (N_752,N_687,N_669);
or U753 (N_753,N_682,N_688);
xnor U754 (N_754,N_705,N_663);
nand U755 (N_755,N_681,N_684);
xor U756 (N_756,N_719,N_707);
xor U757 (N_757,N_675,N_716);
xnor U758 (N_758,N_675,N_706);
nor U759 (N_759,N_715,N_712);
or U760 (N_760,N_692,N_709);
or U761 (N_761,N_661,N_667);
nor U762 (N_762,N_662,N_682);
nor U763 (N_763,N_702,N_704);
xor U764 (N_764,N_717,N_709);
nor U765 (N_765,N_664,N_706);
or U766 (N_766,N_685,N_673);
nand U767 (N_767,N_706,N_702);
xor U768 (N_768,N_717,N_688);
and U769 (N_769,N_682,N_719);
nand U770 (N_770,N_666,N_660);
or U771 (N_771,N_705,N_671);
xnor U772 (N_772,N_702,N_665);
and U773 (N_773,N_686,N_688);
and U774 (N_774,N_665,N_699);
nor U775 (N_775,N_695,N_700);
nor U776 (N_776,N_715,N_667);
and U777 (N_777,N_705,N_674);
and U778 (N_778,N_661,N_673);
or U779 (N_779,N_708,N_661);
nand U780 (N_780,N_740,N_777);
nor U781 (N_781,N_747,N_760);
xor U782 (N_782,N_776,N_752);
nand U783 (N_783,N_720,N_744);
xnor U784 (N_784,N_755,N_764);
nand U785 (N_785,N_735,N_742);
and U786 (N_786,N_775,N_751);
xor U787 (N_787,N_753,N_766);
xor U788 (N_788,N_728,N_724);
xor U789 (N_789,N_739,N_761);
nor U790 (N_790,N_779,N_772);
nand U791 (N_791,N_727,N_730);
xor U792 (N_792,N_768,N_758);
nand U793 (N_793,N_757,N_771);
xor U794 (N_794,N_738,N_725);
nand U795 (N_795,N_745,N_746);
xnor U796 (N_796,N_726,N_754);
nand U797 (N_797,N_767,N_773);
or U798 (N_798,N_774,N_731);
nand U799 (N_799,N_741,N_737);
xnor U800 (N_800,N_729,N_736);
xnor U801 (N_801,N_733,N_750);
nor U802 (N_802,N_762,N_749);
and U803 (N_803,N_763,N_770);
or U804 (N_804,N_748,N_732);
nand U805 (N_805,N_756,N_765);
nor U806 (N_806,N_723,N_743);
nand U807 (N_807,N_734,N_722);
xnor U808 (N_808,N_778,N_759);
xnor U809 (N_809,N_769,N_721);
or U810 (N_810,N_731,N_746);
nand U811 (N_811,N_760,N_777);
or U812 (N_812,N_752,N_748);
and U813 (N_813,N_761,N_779);
nand U814 (N_814,N_732,N_774);
or U815 (N_815,N_772,N_741);
and U816 (N_816,N_770,N_722);
nand U817 (N_817,N_761,N_742);
and U818 (N_818,N_740,N_752);
and U819 (N_819,N_772,N_728);
or U820 (N_820,N_736,N_731);
nand U821 (N_821,N_729,N_750);
xor U822 (N_822,N_742,N_779);
or U823 (N_823,N_765,N_763);
nor U824 (N_824,N_746,N_772);
and U825 (N_825,N_762,N_751);
xor U826 (N_826,N_758,N_746);
nor U827 (N_827,N_765,N_731);
or U828 (N_828,N_762,N_758);
nand U829 (N_829,N_758,N_748);
nand U830 (N_830,N_749,N_747);
nor U831 (N_831,N_766,N_756);
or U832 (N_832,N_776,N_722);
xnor U833 (N_833,N_773,N_768);
nand U834 (N_834,N_721,N_743);
nand U835 (N_835,N_750,N_744);
or U836 (N_836,N_755,N_741);
xnor U837 (N_837,N_741,N_740);
nor U838 (N_838,N_746,N_742);
xor U839 (N_839,N_762,N_742);
and U840 (N_840,N_793,N_831);
or U841 (N_841,N_784,N_819);
nand U842 (N_842,N_782,N_781);
nor U843 (N_843,N_813,N_802);
xnor U844 (N_844,N_808,N_834);
nor U845 (N_845,N_791,N_823);
and U846 (N_846,N_797,N_804);
or U847 (N_847,N_825,N_795);
nand U848 (N_848,N_837,N_833);
xnor U849 (N_849,N_780,N_805);
or U850 (N_850,N_807,N_828);
xnor U851 (N_851,N_814,N_800);
xor U852 (N_852,N_798,N_822);
and U853 (N_853,N_821,N_815);
nand U854 (N_854,N_803,N_809);
or U855 (N_855,N_792,N_829);
nand U856 (N_856,N_818,N_806);
xnor U857 (N_857,N_801,N_788);
nand U858 (N_858,N_838,N_827);
xnor U859 (N_859,N_816,N_783);
xnor U860 (N_860,N_799,N_812);
or U861 (N_861,N_839,N_832);
or U862 (N_862,N_811,N_810);
nand U863 (N_863,N_817,N_796);
or U864 (N_864,N_785,N_835);
nand U865 (N_865,N_787,N_786);
xor U866 (N_866,N_830,N_794);
or U867 (N_867,N_790,N_824);
nand U868 (N_868,N_820,N_836);
nand U869 (N_869,N_789,N_826);
nand U870 (N_870,N_828,N_832);
and U871 (N_871,N_827,N_823);
nand U872 (N_872,N_814,N_837);
and U873 (N_873,N_814,N_810);
xor U874 (N_874,N_799,N_795);
nor U875 (N_875,N_833,N_813);
nor U876 (N_876,N_795,N_830);
nor U877 (N_877,N_807,N_811);
or U878 (N_878,N_833,N_787);
xor U879 (N_879,N_782,N_828);
or U880 (N_880,N_790,N_787);
nand U881 (N_881,N_789,N_792);
or U882 (N_882,N_834,N_803);
or U883 (N_883,N_824,N_782);
nor U884 (N_884,N_804,N_833);
xnor U885 (N_885,N_781,N_795);
nand U886 (N_886,N_787,N_825);
or U887 (N_887,N_838,N_818);
nor U888 (N_888,N_793,N_785);
or U889 (N_889,N_780,N_785);
xnor U890 (N_890,N_827,N_831);
nor U891 (N_891,N_810,N_787);
nand U892 (N_892,N_796,N_781);
nand U893 (N_893,N_824,N_804);
nand U894 (N_894,N_787,N_824);
or U895 (N_895,N_802,N_800);
xnor U896 (N_896,N_823,N_828);
nand U897 (N_897,N_794,N_787);
or U898 (N_898,N_826,N_806);
nor U899 (N_899,N_808,N_821);
xor U900 (N_900,N_872,N_881);
nand U901 (N_901,N_845,N_882);
and U902 (N_902,N_884,N_847);
nand U903 (N_903,N_871,N_874);
or U904 (N_904,N_875,N_892);
xor U905 (N_905,N_864,N_848);
xor U906 (N_906,N_862,N_898);
nand U907 (N_907,N_860,N_857);
xnor U908 (N_908,N_897,N_895);
and U909 (N_909,N_859,N_855);
and U910 (N_910,N_865,N_889);
xor U911 (N_911,N_850,N_891);
nand U912 (N_912,N_899,N_849);
nor U913 (N_913,N_842,N_844);
nand U914 (N_914,N_885,N_879);
or U915 (N_915,N_878,N_861);
and U916 (N_916,N_873,N_883);
nor U917 (N_917,N_863,N_868);
nor U918 (N_918,N_866,N_856);
nor U919 (N_919,N_869,N_853);
nor U920 (N_920,N_888,N_896);
xnor U921 (N_921,N_852,N_893);
nand U922 (N_922,N_894,N_840);
nor U923 (N_923,N_851,N_887);
or U924 (N_924,N_876,N_890);
and U925 (N_925,N_854,N_841);
xor U926 (N_926,N_886,N_870);
or U927 (N_927,N_846,N_880);
nor U928 (N_928,N_858,N_867);
and U929 (N_929,N_877,N_843);
nand U930 (N_930,N_891,N_892);
or U931 (N_931,N_859,N_865);
or U932 (N_932,N_873,N_874);
xor U933 (N_933,N_857,N_852);
or U934 (N_934,N_865,N_848);
xor U935 (N_935,N_842,N_877);
nand U936 (N_936,N_854,N_843);
and U937 (N_937,N_895,N_899);
nand U938 (N_938,N_872,N_866);
and U939 (N_939,N_872,N_846);
or U940 (N_940,N_898,N_847);
nor U941 (N_941,N_874,N_898);
nor U942 (N_942,N_885,N_878);
or U943 (N_943,N_848,N_887);
nand U944 (N_944,N_846,N_851);
or U945 (N_945,N_849,N_864);
nand U946 (N_946,N_850,N_869);
xnor U947 (N_947,N_886,N_846);
and U948 (N_948,N_876,N_894);
xnor U949 (N_949,N_850,N_848);
nor U950 (N_950,N_888,N_877);
nand U951 (N_951,N_840,N_850);
xnor U952 (N_952,N_856,N_881);
xnor U953 (N_953,N_861,N_849);
xnor U954 (N_954,N_869,N_860);
nor U955 (N_955,N_890,N_887);
or U956 (N_956,N_863,N_865);
and U957 (N_957,N_869,N_846);
and U958 (N_958,N_886,N_877);
nand U959 (N_959,N_857,N_883);
xnor U960 (N_960,N_942,N_957);
nand U961 (N_961,N_955,N_907);
and U962 (N_962,N_925,N_951);
or U963 (N_963,N_934,N_927);
xor U964 (N_964,N_938,N_919);
or U965 (N_965,N_921,N_902);
nand U966 (N_966,N_914,N_912);
xor U967 (N_967,N_901,N_909);
and U968 (N_968,N_924,N_915);
nand U969 (N_969,N_933,N_908);
or U970 (N_970,N_937,N_956);
or U971 (N_971,N_918,N_946);
and U972 (N_972,N_929,N_910);
nor U973 (N_973,N_950,N_906);
xor U974 (N_974,N_948,N_923);
and U975 (N_975,N_935,N_958);
and U976 (N_976,N_911,N_920);
and U977 (N_977,N_913,N_952);
nor U978 (N_978,N_905,N_928);
xnor U979 (N_979,N_943,N_944);
and U980 (N_980,N_947,N_954);
or U981 (N_981,N_939,N_904);
or U982 (N_982,N_916,N_945);
or U983 (N_983,N_959,N_940);
xor U984 (N_984,N_936,N_931);
xnor U985 (N_985,N_930,N_941);
xor U986 (N_986,N_903,N_949);
xnor U987 (N_987,N_953,N_926);
and U988 (N_988,N_900,N_922);
nor U989 (N_989,N_932,N_917);
or U990 (N_990,N_954,N_928);
nand U991 (N_991,N_953,N_915);
xor U992 (N_992,N_919,N_949);
nand U993 (N_993,N_928,N_935);
and U994 (N_994,N_904,N_903);
nand U995 (N_995,N_931,N_903);
nand U996 (N_996,N_938,N_952);
xor U997 (N_997,N_937,N_916);
or U998 (N_998,N_945,N_929);
xnor U999 (N_999,N_928,N_917);
nor U1000 (N_1000,N_930,N_932);
nor U1001 (N_1001,N_946,N_906);
or U1002 (N_1002,N_945,N_948);
nand U1003 (N_1003,N_920,N_952);
and U1004 (N_1004,N_900,N_931);
nand U1005 (N_1005,N_952,N_957);
or U1006 (N_1006,N_906,N_944);
xnor U1007 (N_1007,N_922,N_913);
and U1008 (N_1008,N_948,N_947);
xor U1009 (N_1009,N_917,N_948);
or U1010 (N_1010,N_929,N_933);
nor U1011 (N_1011,N_942,N_904);
or U1012 (N_1012,N_923,N_936);
or U1013 (N_1013,N_922,N_907);
xnor U1014 (N_1014,N_912,N_904);
xnor U1015 (N_1015,N_955,N_929);
or U1016 (N_1016,N_933,N_900);
and U1017 (N_1017,N_914,N_930);
nor U1018 (N_1018,N_939,N_943);
or U1019 (N_1019,N_931,N_926);
nand U1020 (N_1020,N_1011,N_982);
and U1021 (N_1021,N_990,N_1002);
nand U1022 (N_1022,N_973,N_967);
xor U1023 (N_1023,N_1006,N_983);
nand U1024 (N_1024,N_1015,N_988);
or U1025 (N_1025,N_1016,N_968);
nor U1026 (N_1026,N_992,N_1003);
xor U1027 (N_1027,N_972,N_994);
and U1028 (N_1028,N_999,N_975);
nand U1029 (N_1029,N_1012,N_1005);
nor U1030 (N_1030,N_980,N_985);
xor U1031 (N_1031,N_978,N_1008);
and U1032 (N_1032,N_993,N_979);
nand U1033 (N_1033,N_987,N_976);
xnor U1034 (N_1034,N_977,N_966);
and U1035 (N_1035,N_1019,N_1007);
or U1036 (N_1036,N_1000,N_984);
or U1037 (N_1037,N_995,N_991);
nand U1038 (N_1038,N_1018,N_998);
or U1039 (N_1039,N_965,N_986);
nand U1040 (N_1040,N_971,N_1004);
and U1041 (N_1041,N_989,N_960);
and U1042 (N_1042,N_963,N_1001);
nand U1043 (N_1043,N_981,N_962);
nor U1044 (N_1044,N_969,N_970);
and U1045 (N_1045,N_961,N_1010);
nand U1046 (N_1046,N_1009,N_1017);
or U1047 (N_1047,N_997,N_1013);
or U1048 (N_1048,N_974,N_996);
nor U1049 (N_1049,N_964,N_1014);
nand U1050 (N_1050,N_1013,N_971);
or U1051 (N_1051,N_990,N_1014);
and U1052 (N_1052,N_1006,N_982);
nand U1053 (N_1053,N_990,N_1003);
xnor U1054 (N_1054,N_975,N_991);
xor U1055 (N_1055,N_1013,N_999);
nor U1056 (N_1056,N_991,N_996);
nand U1057 (N_1057,N_962,N_966);
nand U1058 (N_1058,N_967,N_1018);
nand U1059 (N_1059,N_1012,N_988);
nor U1060 (N_1060,N_970,N_986);
and U1061 (N_1061,N_982,N_983);
xor U1062 (N_1062,N_981,N_1002);
nand U1063 (N_1063,N_1004,N_997);
or U1064 (N_1064,N_979,N_1019);
xor U1065 (N_1065,N_985,N_962);
and U1066 (N_1066,N_1013,N_978);
and U1067 (N_1067,N_990,N_995);
nor U1068 (N_1068,N_1012,N_972);
nand U1069 (N_1069,N_980,N_1006);
or U1070 (N_1070,N_998,N_984);
nand U1071 (N_1071,N_995,N_1017);
or U1072 (N_1072,N_995,N_970);
or U1073 (N_1073,N_1000,N_986);
and U1074 (N_1074,N_991,N_983);
nand U1075 (N_1075,N_973,N_1011);
nand U1076 (N_1076,N_1011,N_971);
nor U1077 (N_1077,N_1014,N_991);
and U1078 (N_1078,N_975,N_970);
or U1079 (N_1079,N_1012,N_993);
xor U1080 (N_1080,N_1048,N_1027);
nor U1081 (N_1081,N_1063,N_1033);
nor U1082 (N_1082,N_1072,N_1020);
nand U1083 (N_1083,N_1023,N_1079);
or U1084 (N_1084,N_1065,N_1057);
nand U1085 (N_1085,N_1066,N_1075);
and U1086 (N_1086,N_1024,N_1059);
or U1087 (N_1087,N_1045,N_1068);
and U1088 (N_1088,N_1032,N_1071);
nand U1089 (N_1089,N_1076,N_1038);
or U1090 (N_1090,N_1056,N_1021);
or U1091 (N_1091,N_1044,N_1025);
nor U1092 (N_1092,N_1036,N_1026);
and U1093 (N_1093,N_1047,N_1043);
and U1094 (N_1094,N_1050,N_1029);
or U1095 (N_1095,N_1028,N_1067);
and U1096 (N_1096,N_1060,N_1055);
and U1097 (N_1097,N_1074,N_1069);
nand U1098 (N_1098,N_1035,N_1052);
nor U1099 (N_1099,N_1037,N_1031);
nand U1100 (N_1100,N_1058,N_1046);
or U1101 (N_1101,N_1049,N_1040);
or U1102 (N_1102,N_1039,N_1051);
or U1103 (N_1103,N_1041,N_1034);
nand U1104 (N_1104,N_1054,N_1022);
and U1105 (N_1105,N_1053,N_1064);
nand U1106 (N_1106,N_1078,N_1073);
nor U1107 (N_1107,N_1062,N_1042);
nor U1108 (N_1108,N_1070,N_1077);
or U1109 (N_1109,N_1061,N_1030);
nor U1110 (N_1110,N_1034,N_1047);
and U1111 (N_1111,N_1049,N_1041);
or U1112 (N_1112,N_1034,N_1026);
nand U1113 (N_1113,N_1050,N_1043);
and U1114 (N_1114,N_1046,N_1068);
and U1115 (N_1115,N_1075,N_1034);
and U1116 (N_1116,N_1077,N_1044);
xnor U1117 (N_1117,N_1025,N_1056);
nor U1118 (N_1118,N_1075,N_1023);
or U1119 (N_1119,N_1052,N_1077);
nor U1120 (N_1120,N_1040,N_1059);
and U1121 (N_1121,N_1033,N_1040);
nand U1122 (N_1122,N_1040,N_1022);
nand U1123 (N_1123,N_1020,N_1077);
nor U1124 (N_1124,N_1044,N_1037);
and U1125 (N_1125,N_1026,N_1027);
and U1126 (N_1126,N_1052,N_1072);
nand U1127 (N_1127,N_1045,N_1042);
nand U1128 (N_1128,N_1023,N_1021);
and U1129 (N_1129,N_1069,N_1037);
xor U1130 (N_1130,N_1029,N_1068);
and U1131 (N_1131,N_1031,N_1034);
or U1132 (N_1132,N_1020,N_1065);
nor U1133 (N_1133,N_1022,N_1061);
and U1134 (N_1134,N_1050,N_1034);
nor U1135 (N_1135,N_1043,N_1046);
or U1136 (N_1136,N_1027,N_1063);
xor U1137 (N_1137,N_1028,N_1060);
and U1138 (N_1138,N_1062,N_1065);
and U1139 (N_1139,N_1076,N_1064);
nor U1140 (N_1140,N_1091,N_1114);
nor U1141 (N_1141,N_1122,N_1129);
nand U1142 (N_1142,N_1120,N_1093);
or U1143 (N_1143,N_1107,N_1090);
nor U1144 (N_1144,N_1104,N_1083);
and U1145 (N_1145,N_1130,N_1135);
xor U1146 (N_1146,N_1123,N_1136);
nand U1147 (N_1147,N_1099,N_1128);
nor U1148 (N_1148,N_1094,N_1121);
nor U1149 (N_1149,N_1097,N_1092);
and U1150 (N_1150,N_1084,N_1117);
nor U1151 (N_1151,N_1138,N_1087);
nand U1152 (N_1152,N_1081,N_1082);
or U1153 (N_1153,N_1111,N_1108);
nor U1154 (N_1154,N_1125,N_1118);
and U1155 (N_1155,N_1105,N_1109);
and U1156 (N_1156,N_1103,N_1132);
or U1157 (N_1157,N_1115,N_1112);
or U1158 (N_1158,N_1095,N_1110);
nand U1159 (N_1159,N_1127,N_1098);
nor U1160 (N_1160,N_1089,N_1100);
xnor U1161 (N_1161,N_1080,N_1113);
nor U1162 (N_1162,N_1106,N_1126);
or U1163 (N_1163,N_1101,N_1139);
nor U1164 (N_1164,N_1086,N_1102);
or U1165 (N_1165,N_1137,N_1119);
xor U1166 (N_1166,N_1088,N_1085);
nor U1167 (N_1167,N_1131,N_1116);
or U1168 (N_1168,N_1124,N_1096);
and U1169 (N_1169,N_1134,N_1133);
or U1170 (N_1170,N_1089,N_1125);
or U1171 (N_1171,N_1103,N_1134);
nand U1172 (N_1172,N_1107,N_1093);
and U1173 (N_1173,N_1110,N_1103);
nand U1174 (N_1174,N_1117,N_1122);
nor U1175 (N_1175,N_1096,N_1139);
and U1176 (N_1176,N_1085,N_1121);
xor U1177 (N_1177,N_1101,N_1120);
xor U1178 (N_1178,N_1109,N_1080);
or U1179 (N_1179,N_1136,N_1119);
nor U1180 (N_1180,N_1117,N_1094);
nor U1181 (N_1181,N_1108,N_1086);
nor U1182 (N_1182,N_1098,N_1112);
xor U1183 (N_1183,N_1130,N_1115);
nand U1184 (N_1184,N_1098,N_1086);
and U1185 (N_1185,N_1122,N_1134);
or U1186 (N_1186,N_1088,N_1127);
or U1187 (N_1187,N_1136,N_1131);
or U1188 (N_1188,N_1083,N_1116);
nand U1189 (N_1189,N_1111,N_1092);
or U1190 (N_1190,N_1112,N_1117);
and U1191 (N_1191,N_1081,N_1104);
xor U1192 (N_1192,N_1118,N_1116);
nand U1193 (N_1193,N_1084,N_1124);
nor U1194 (N_1194,N_1128,N_1085);
xor U1195 (N_1195,N_1085,N_1120);
or U1196 (N_1196,N_1130,N_1128);
nor U1197 (N_1197,N_1083,N_1125);
and U1198 (N_1198,N_1089,N_1130);
xnor U1199 (N_1199,N_1086,N_1110);
nand U1200 (N_1200,N_1192,N_1187);
or U1201 (N_1201,N_1197,N_1177);
xor U1202 (N_1202,N_1167,N_1199);
nand U1203 (N_1203,N_1194,N_1172);
xnor U1204 (N_1204,N_1176,N_1186);
or U1205 (N_1205,N_1196,N_1164);
nor U1206 (N_1206,N_1153,N_1174);
nand U1207 (N_1207,N_1159,N_1161);
nor U1208 (N_1208,N_1193,N_1181);
xnor U1209 (N_1209,N_1151,N_1155);
nor U1210 (N_1210,N_1145,N_1146);
xor U1211 (N_1211,N_1188,N_1173);
nor U1212 (N_1212,N_1184,N_1171);
nand U1213 (N_1213,N_1156,N_1178);
xnor U1214 (N_1214,N_1160,N_1180);
or U1215 (N_1215,N_1166,N_1142);
or U1216 (N_1216,N_1152,N_1158);
nand U1217 (N_1217,N_1163,N_1182);
nand U1218 (N_1218,N_1189,N_1169);
nor U1219 (N_1219,N_1165,N_1150);
nor U1220 (N_1220,N_1190,N_1140);
xnor U1221 (N_1221,N_1183,N_1148);
xnor U1222 (N_1222,N_1191,N_1149);
or U1223 (N_1223,N_1162,N_1195);
or U1224 (N_1224,N_1170,N_1157);
or U1225 (N_1225,N_1141,N_1198);
xor U1226 (N_1226,N_1185,N_1175);
and U1227 (N_1227,N_1144,N_1179);
nand U1228 (N_1228,N_1147,N_1168);
xor U1229 (N_1229,N_1154,N_1143);
or U1230 (N_1230,N_1153,N_1175);
or U1231 (N_1231,N_1172,N_1185);
or U1232 (N_1232,N_1193,N_1194);
nand U1233 (N_1233,N_1171,N_1193);
nor U1234 (N_1234,N_1169,N_1150);
nand U1235 (N_1235,N_1142,N_1143);
or U1236 (N_1236,N_1198,N_1192);
or U1237 (N_1237,N_1149,N_1177);
nor U1238 (N_1238,N_1158,N_1195);
or U1239 (N_1239,N_1187,N_1149);
xnor U1240 (N_1240,N_1160,N_1190);
nand U1241 (N_1241,N_1158,N_1165);
and U1242 (N_1242,N_1164,N_1171);
and U1243 (N_1243,N_1153,N_1196);
nand U1244 (N_1244,N_1167,N_1163);
nand U1245 (N_1245,N_1185,N_1186);
nor U1246 (N_1246,N_1169,N_1159);
and U1247 (N_1247,N_1189,N_1146);
and U1248 (N_1248,N_1164,N_1156);
xnor U1249 (N_1249,N_1151,N_1165);
nand U1250 (N_1250,N_1140,N_1184);
or U1251 (N_1251,N_1173,N_1141);
nand U1252 (N_1252,N_1159,N_1157);
nor U1253 (N_1253,N_1197,N_1181);
nand U1254 (N_1254,N_1157,N_1173);
nand U1255 (N_1255,N_1196,N_1147);
and U1256 (N_1256,N_1154,N_1169);
xor U1257 (N_1257,N_1152,N_1189);
nor U1258 (N_1258,N_1148,N_1159);
and U1259 (N_1259,N_1178,N_1186);
xor U1260 (N_1260,N_1251,N_1225);
nand U1261 (N_1261,N_1200,N_1236);
and U1262 (N_1262,N_1211,N_1232);
and U1263 (N_1263,N_1209,N_1219);
and U1264 (N_1264,N_1240,N_1206);
or U1265 (N_1265,N_1243,N_1217);
nand U1266 (N_1266,N_1215,N_1246);
nor U1267 (N_1267,N_1223,N_1252);
and U1268 (N_1268,N_1235,N_1230);
nor U1269 (N_1269,N_1242,N_1231);
and U1270 (N_1270,N_1229,N_1226);
nor U1271 (N_1271,N_1257,N_1221);
or U1272 (N_1272,N_1249,N_1205);
and U1273 (N_1273,N_1218,N_1212);
and U1274 (N_1274,N_1241,N_1204);
and U1275 (N_1275,N_1239,N_1250);
nand U1276 (N_1276,N_1247,N_1210);
and U1277 (N_1277,N_1227,N_1207);
or U1278 (N_1278,N_1220,N_1237);
or U1279 (N_1279,N_1238,N_1213);
or U1280 (N_1280,N_1253,N_1258);
and U1281 (N_1281,N_1234,N_1222);
or U1282 (N_1282,N_1259,N_1255);
xnor U1283 (N_1283,N_1256,N_1208);
nand U1284 (N_1284,N_1203,N_1245);
or U1285 (N_1285,N_1254,N_1224);
and U1286 (N_1286,N_1228,N_1201);
or U1287 (N_1287,N_1214,N_1248);
and U1288 (N_1288,N_1202,N_1233);
and U1289 (N_1289,N_1216,N_1244);
xor U1290 (N_1290,N_1254,N_1227);
and U1291 (N_1291,N_1212,N_1225);
and U1292 (N_1292,N_1234,N_1216);
nand U1293 (N_1293,N_1222,N_1223);
xnor U1294 (N_1294,N_1207,N_1216);
xnor U1295 (N_1295,N_1207,N_1205);
xnor U1296 (N_1296,N_1256,N_1209);
or U1297 (N_1297,N_1249,N_1256);
xor U1298 (N_1298,N_1240,N_1237);
or U1299 (N_1299,N_1203,N_1230);
xor U1300 (N_1300,N_1238,N_1236);
xor U1301 (N_1301,N_1255,N_1219);
xnor U1302 (N_1302,N_1234,N_1237);
nor U1303 (N_1303,N_1220,N_1251);
xor U1304 (N_1304,N_1248,N_1252);
nand U1305 (N_1305,N_1234,N_1235);
or U1306 (N_1306,N_1248,N_1203);
nand U1307 (N_1307,N_1237,N_1248);
nor U1308 (N_1308,N_1227,N_1245);
and U1309 (N_1309,N_1238,N_1214);
and U1310 (N_1310,N_1232,N_1220);
or U1311 (N_1311,N_1239,N_1258);
nor U1312 (N_1312,N_1213,N_1220);
xnor U1313 (N_1313,N_1239,N_1247);
nand U1314 (N_1314,N_1228,N_1219);
xnor U1315 (N_1315,N_1201,N_1218);
nor U1316 (N_1316,N_1200,N_1219);
and U1317 (N_1317,N_1250,N_1202);
or U1318 (N_1318,N_1259,N_1200);
and U1319 (N_1319,N_1233,N_1213);
nand U1320 (N_1320,N_1262,N_1276);
nand U1321 (N_1321,N_1311,N_1312);
nand U1322 (N_1322,N_1268,N_1300);
nor U1323 (N_1323,N_1318,N_1275);
or U1324 (N_1324,N_1310,N_1291);
nor U1325 (N_1325,N_1283,N_1274);
and U1326 (N_1326,N_1271,N_1277);
and U1327 (N_1327,N_1270,N_1263);
and U1328 (N_1328,N_1267,N_1316);
or U1329 (N_1329,N_1303,N_1319);
nor U1330 (N_1330,N_1296,N_1282);
or U1331 (N_1331,N_1293,N_1308);
xor U1332 (N_1332,N_1278,N_1313);
xor U1333 (N_1333,N_1314,N_1307);
nand U1334 (N_1334,N_1304,N_1317);
nand U1335 (N_1335,N_1286,N_1280);
or U1336 (N_1336,N_1284,N_1305);
xor U1337 (N_1337,N_1295,N_1261);
nand U1338 (N_1338,N_1272,N_1292);
and U1339 (N_1339,N_1260,N_1290);
nand U1340 (N_1340,N_1269,N_1301);
and U1341 (N_1341,N_1302,N_1297);
nor U1342 (N_1342,N_1287,N_1273);
nand U1343 (N_1343,N_1288,N_1266);
and U1344 (N_1344,N_1264,N_1265);
nor U1345 (N_1345,N_1279,N_1309);
nor U1346 (N_1346,N_1315,N_1306);
nand U1347 (N_1347,N_1281,N_1294);
nand U1348 (N_1348,N_1299,N_1285);
nand U1349 (N_1349,N_1289,N_1298);
nand U1350 (N_1350,N_1310,N_1313);
and U1351 (N_1351,N_1283,N_1286);
xnor U1352 (N_1352,N_1296,N_1314);
or U1353 (N_1353,N_1298,N_1279);
and U1354 (N_1354,N_1286,N_1291);
nor U1355 (N_1355,N_1271,N_1297);
nand U1356 (N_1356,N_1309,N_1312);
nor U1357 (N_1357,N_1311,N_1279);
or U1358 (N_1358,N_1272,N_1281);
xnor U1359 (N_1359,N_1268,N_1281);
nand U1360 (N_1360,N_1297,N_1301);
xnor U1361 (N_1361,N_1300,N_1281);
nand U1362 (N_1362,N_1265,N_1305);
nor U1363 (N_1363,N_1275,N_1283);
nor U1364 (N_1364,N_1318,N_1280);
nand U1365 (N_1365,N_1264,N_1267);
or U1366 (N_1366,N_1286,N_1271);
or U1367 (N_1367,N_1318,N_1284);
and U1368 (N_1368,N_1317,N_1282);
nand U1369 (N_1369,N_1290,N_1298);
nor U1370 (N_1370,N_1291,N_1292);
nand U1371 (N_1371,N_1291,N_1284);
xor U1372 (N_1372,N_1307,N_1268);
nand U1373 (N_1373,N_1315,N_1274);
or U1374 (N_1374,N_1300,N_1266);
nand U1375 (N_1375,N_1305,N_1282);
or U1376 (N_1376,N_1293,N_1314);
and U1377 (N_1377,N_1296,N_1300);
nand U1378 (N_1378,N_1279,N_1312);
or U1379 (N_1379,N_1301,N_1288);
xnor U1380 (N_1380,N_1327,N_1340);
and U1381 (N_1381,N_1366,N_1342);
xor U1382 (N_1382,N_1324,N_1323);
and U1383 (N_1383,N_1372,N_1351);
nand U1384 (N_1384,N_1345,N_1321);
or U1385 (N_1385,N_1322,N_1361);
and U1386 (N_1386,N_1373,N_1352);
or U1387 (N_1387,N_1320,N_1334);
nor U1388 (N_1388,N_1377,N_1326);
xor U1389 (N_1389,N_1325,N_1369);
and U1390 (N_1390,N_1335,N_1333);
nand U1391 (N_1391,N_1337,N_1365);
xor U1392 (N_1392,N_1353,N_1363);
xnor U1393 (N_1393,N_1338,N_1375);
or U1394 (N_1394,N_1341,N_1364);
nand U1395 (N_1395,N_1371,N_1379);
nor U1396 (N_1396,N_1330,N_1350);
nor U1397 (N_1397,N_1331,N_1348);
nand U1398 (N_1398,N_1370,N_1360);
and U1399 (N_1399,N_1368,N_1374);
or U1400 (N_1400,N_1346,N_1378);
or U1401 (N_1401,N_1343,N_1376);
nor U1402 (N_1402,N_1359,N_1357);
xnor U1403 (N_1403,N_1367,N_1329);
and U1404 (N_1404,N_1347,N_1362);
nand U1405 (N_1405,N_1332,N_1355);
or U1406 (N_1406,N_1336,N_1344);
xor U1407 (N_1407,N_1354,N_1358);
xor U1408 (N_1408,N_1356,N_1339);
nand U1409 (N_1409,N_1349,N_1328);
and U1410 (N_1410,N_1360,N_1349);
nand U1411 (N_1411,N_1355,N_1353);
nor U1412 (N_1412,N_1327,N_1366);
and U1413 (N_1413,N_1358,N_1360);
xor U1414 (N_1414,N_1349,N_1333);
nor U1415 (N_1415,N_1364,N_1365);
nor U1416 (N_1416,N_1359,N_1328);
nand U1417 (N_1417,N_1358,N_1327);
nand U1418 (N_1418,N_1326,N_1351);
nand U1419 (N_1419,N_1353,N_1368);
nand U1420 (N_1420,N_1365,N_1373);
or U1421 (N_1421,N_1323,N_1377);
xnor U1422 (N_1422,N_1332,N_1335);
xnor U1423 (N_1423,N_1356,N_1350);
nand U1424 (N_1424,N_1360,N_1367);
xnor U1425 (N_1425,N_1359,N_1325);
and U1426 (N_1426,N_1372,N_1334);
and U1427 (N_1427,N_1353,N_1345);
nand U1428 (N_1428,N_1351,N_1344);
and U1429 (N_1429,N_1338,N_1342);
nand U1430 (N_1430,N_1339,N_1351);
xor U1431 (N_1431,N_1328,N_1369);
and U1432 (N_1432,N_1375,N_1373);
nand U1433 (N_1433,N_1348,N_1343);
nand U1434 (N_1434,N_1355,N_1347);
nand U1435 (N_1435,N_1327,N_1373);
and U1436 (N_1436,N_1343,N_1333);
xor U1437 (N_1437,N_1347,N_1357);
nor U1438 (N_1438,N_1350,N_1370);
or U1439 (N_1439,N_1324,N_1369);
xnor U1440 (N_1440,N_1402,N_1437);
or U1441 (N_1441,N_1413,N_1389);
or U1442 (N_1442,N_1397,N_1399);
nor U1443 (N_1443,N_1395,N_1388);
xor U1444 (N_1444,N_1380,N_1439);
xor U1445 (N_1445,N_1421,N_1385);
or U1446 (N_1446,N_1411,N_1394);
nand U1447 (N_1447,N_1423,N_1426);
or U1448 (N_1448,N_1387,N_1431);
nor U1449 (N_1449,N_1432,N_1396);
nand U1450 (N_1450,N_1436,N_1408);
nor U1451 (N_1451,N_1418,N_1419);
and U1452 (N_1452,N_1386,N_1406);
nand U1453 (N_1453,N_1415,N_1424);
xnor U1454 (N_1454,N_1405,N_1409);
nand U1455 (N_1455,N_1400,N_1403);
xnor U1456 (N_1456,N_1430,N_1390);
and U1457 (N_1457,N_1429,N_1393);
xor U1458 (N_1458,N_1381,N_1428);
and U1459 (N_1459,N_1401,N_1391);
nor U1460 (N_1460,N_1435,N_1420);
and U1461 (N_1461,N_1410,N_1434);
and U1462 (N_1462,N_1416,N_1412);
nand U1463 (N_1463,N_1414,N_1425);
nor U1464 (N_1464,N_1384,N_1383);
nand U1465 (N_1465,N_1427,N_1438);
xnor U1466 (N_1466,N_1433,N_1417);
nor U1467 (N_1467,N_1392,N_1404);
nor U1468 (N_1468,N_1407,N_1398);
nand U1469 (N_1469,N_1382,N_1422);
and U1470 (N_1470,N_1422,N_1389);
nand U1471 (N_1471,N_1405,N_1435);
or U1472 (N_1472,N_1439,N_1431);
nand U1473 (N_1473,N_1432,N_1387);
or U1474 (N_1474,N_1394,N_1421);
nand U1475 (N_1475,N_1380,N_1382);
and U1476 (N_1476,N_1423,N_1389);
or U1477 (N_1477,N_1411,N_1428);
nand U1478 (N_1478,N_1401,N_1412);
xor U1479 (N_1479,N_1395,N_1413);
xor U1480 (N_1480,N_1423,N_1425);
nor U1481 (N_1481,N_1403,N_1430);
nand U1482 (N_1482,N_1406,N_1395);
nand U1483 (N_1483,N_1407,N_1403);
and U1484 (N_1484,N_1413,N_1436);
or U1485 (N_1485,N_1402,N_1429);
nand U1486 (N_1486,N_1391,N_1390);
nor U1487 (N_1487,N_1405,N_1402);
xnor U1488 (N_1488,N_1416,N_1387);
nor U1489 (N_1489,N_1427,N_1414);
or U1490 (N_1490,N_1391,N_1433);
or U1491 (N_1491,N_1405,N_1391);
and U1492 (N_1492,N_1420,N_1433);
or U1493 (N_1493,N_1405,N_1437);
nand U1494 (N_1494,N_1426,N_1386);
and U1495 (N_1495,N_1387,N_1397);
and U1496 (N_1496,N_1386,N_1389);
and U1497 (N_1497,N_1388,N_1421);
nand U1498 (N_1498,N_1392,N_1425);
and U1499 (N_1499,N_1385,N_1430);
nor U1500 (N_1500,N_1449,N_1482);
and U1501 (N_1501,N_1471,N_1458);
xnor U1502 (N_1502,N_1446,N_1499);
xnor U1503 (N_1503,N_1444,N_1465);
xnor U1504 (N_1504,N_1448,N_1452);
and U1505 (N_1505,N_1492,N_1489);
nor U1506 (N_1506,N_1457,N_1477);
nor U1507 (N_1507,N_1478,N_1455);
nand U1508 (N_1508,N_1466,N_1450);
or U1509 (N_1509,N_1447,N_1474);
xor U1510 (N_1510,N_1469,N_1440);
nand U1511 (N_1511,N_1494,N_1453);
xnor U1512 (N_1512,N_1473,N_1488);
and U1513 (N_1513,N_1493,N_1486);
and U1514 (N_1514,N_1491,N_1472);
or U1515 (N_1515,N_1464,N_1495);
xor U1516 (N_1516,N_1454,N_1456);
or U1517 (N_1517,N_1487,N_1476);
and U1518 (N_1518,N_1460,N_1445);
and U1519 (N_1519,N_1483,N_1496);
nor U1520 (N_1520,N_1451,N_1459);
xnor U1521 (N_1521,N_1467,N_1480);
or U1522 (N_1522,N_1485,N_1498);
nor U1523 (N_1523,N_1490,N_1441);
xor U1524 (N_1524,N_1475,N_1479);
xnor U1525 (N_1525,N_1443,N_1481);
nand U1526 (N_1526,N_1442,N_1470);
nor U1527 (N_1527,N_1462,N_1461);
nor U1528 (N_1528,N_1484,N_1468);
and U1529 (N_1529,N_1497,N_1463);
nor U1530 (N_1530,N_1496,N_1499);
nand U1531 (N_1531,N_1455,N_1444);
nand U1532 (N_1532,N_1443,N_1444);
and U1533 (N_1533,N_1496,N_1452);
xor U1534 (N_1534,N_1483,N_1443);
and U1535 (N_1535,N_1442,N_1494);
xnor U1536 (N_1536,N_1475,N_1462);
and U1537 (N_1537,N_1483,N_1469);
and U1538 (N_1538,N_1452,N_1480);
or U1539 (N_1539,N_1461,N_1494);
or U1540 (N_1540,N_1455,N_1462);
or U1541 (N_1541,N_1457,N_1493);
nand U1542 (N_1542,N_1443,N_1457);
xnor U1543 (N_1543,N_1476,N_1452);
or U1544 (N_1544,N_1458,N_1489);
nor U1545 (N_1545,N_1496,N_1458);
or U1546 (N_1546,N_1442,N_1467);
and U1547 (N_1547,N_1447,N_1499);
xor U1548 (N_1548,N_1442,N_1491);
nor U1549 (N_1549,N_1453,N_1486);
nor U1550 (N_1550,N_1465,N_1450);
nand U1551 (N_1551,N_1472,N_1458);
or U1552 (N_1552,N_1464,N_1469);
and U1553 (N_1553,N_1457,N_1467);
or U1554 (N_1554,N_1469,N_1441);
and U1555 (N_1555,N_1489,N_1465);
and U1556 (N_1556,N_1476,N_1444);
nor U1557 (N_1557,N_1476,N_1445);
nor U1558 (N_1558,N_1489,N_1454);
nor U1559 (N_1559,N_1459,N_1483);
nand U1560 (N_1560,N_1537,N_1513);
xor U1561 (N_1561,N_1538,N_1510);
or U1562 (N_1562,N_1501,N_1557);
or U1563 (N_1563,N_1507,N_1549);
xor U1564 (N_1564,N_1552,N_1512);
xor U1565 (N_1565,N_1550,N_1508);
nand U1566 (N_1566,N_1533,N_1520);
nor U1567 (N_1567,N_1555,N_1506);
nand U1568 (N_1568,N_1529,N_1516);
xor U1569 (N_1569,N_1551,N_1515);
or U1570 (N_1570,N_1502,N_1505);
nand U1571 (N_1571,N_1523,N_1554);
or U1572 (N_1572,N_1539,N_1556);
or U1573 (N_1573,N_1518,N_1548);
nand U1574 (N_1574,N_1503,N_1504);
or U1575 (N_1575,N_1541,N_1534);
nor U1576 (N_1576,N_1544,N_1530);
nand U1577 (N_1577,N_1528,N_1509);
or U1578 (N_1578,N_1527,N_1526);
xnor U1579 (N_1579,N_1522,N_1546);
xor U1580 (N_1580,N_1532,N_1559);
nor U1581 (N_1581,N_1545,N_1514);
xnor U1582 (N_1582,N_1540,N_1519);
and U1583 (N_1583,N_1543,N_1536);
xor U1584 (N_1584,N_1517,N_1542);
or U1585 (N_1585,N_1553,N_1521);
xnor U1586 (N_1586,N_1535,N_1525);
and U1587 (N_1587,N_1500,N_1558);
and U1588 (N_1588,N_1547,N_1511);
nor U1589 (N_1589,N_1524,N_1531);
xor U1590 (N_1590,N_1530,N_1543);
or U1591 (N_1591,N_1505,N_1536);
xnor U1592 (N_1592,N_1513,N_1542);
xnor U1593 (N_1593,N_1521,N_1534);
and U1594 (N_1594,N_1507,N_1505);
nor U1595 (N_1595,N_1539,N_1523);
nor U1596 (N_1596,N_1503,N_1547);
nand U1597 (N_1597,N_1501,N_1506);
nand U1598 (N_1598,N_1543,N_1526);
xor U1599 (N_1599,N_1521,N_1542);
nand U1600 (N_1600,N_1525,N_1523);
nand U1601 (N_1601,N_1529,N_1548);
and U1602 (N_1602,N_1549,N_1520);
xor U1603 (N_1603,N_1521,N_1556);
nor U1604 (N_1604,N_1510,N_1511);
xnor U1605 (N_1605,N_1516,N_1500);
and U1606 (N_1606,N_1555,N_1540);
or U1607 (N_1607,N_1552,N_1536);
and U1608 (N_1608,N_1514,N_1559);
or U1609 (N_1609,N_1526,N_1533);
xnor U1610 (N_1610,N_1500,N_1524);
xor U1611 (N_1611,N_1529,N_1523);
or U1612 (N_1612,N_1522,N_1513);
nand U1613 (N_1613,N_1525,N_1550);
nor U1614 (N_1614,N_1532,N_1553);
nor U1615 (N_1615,N_1533,N_1510);
nand U1616 (N_1616,N_1519,N_1512);
and U1617 (N_1617,N_1553,N_1549);
and U1618 (N_1618,N_1557,N_1521);
and U1619 (N_1619,N_1508,N_1540);
or U1620 (N_1620,N_1582,N_1591);
nand U1621 (N_1621,N_1587,N_1601);
or U1622 (N_1622,N_1599,N_1608);
and U1623 (N_1623,N_1618,N_1589);
nor U1624 (N_1624,N_1563,N_1600);
nand U1625 (N_1625,N_1598,N_1613);
xor U1626 (N_1626,N_1571,N_1584);
and U1627 (N_1627,N_1569,N_1568);
or U1628 (N_1628,N_1619,N_1606);
xnor U1629 (N_1629,N_1617,N_1588);
xnor U1630 (N_1630,N_1592,N_1576);
nand U1631 (N_1631,N_1604,N_1580);
nand U1632 (N_1632,N_1602,N_1597);
nor U1633 (N_1633,N_1614,N_1585);
xnor U1634 (N_1634,N_1575,N_1565);
and U1635 (N_1635,N_1578,N_1581);
and U1636 (N_1636,N_1564,N_1603);
xor U1637 (N_1637,N_1586,N_1610);
and U1638 (N_1638,N_1611,N_1594);
and U1639 (N_1639,N_1561,N_1560);
nor U1640 (N_1640,N_1616,N_1574);
nand U1641 (N_1641,N_1567,N_1607);
or U1642 (N_1642,N_1605,N_1583);
nand U1643 (N_1643,N_1562,N_1573);
nand U1644 (N_1644,N_1579,N_1612);
and U1645 (N_1645,N_1566,N_1572);
nor U1646 (N_1646,N_1595,N_1577);
nand U1647 (N_1647,N_1590,N_1593);
and U1648 (N_1648,N_1615,N_1609);
and U1649 (N_1649,N_1570,N_1596);
or U1650 (N_1650,N_1614,N_1601);
xor U1651 (N_1651,N_1617,N_1590);
nor U1652 (N_1652,N_1599,N_1612);
xor U1653 (N_1653,N_1606,N_1618);
xor U1654 (N_1654,N_1566,N_1589);
or U1655 (N_1655,N_1560,N_1584);
and U1656 (N_1656,N_1577,N_1615);
xor U1657 (N_1657,N_1578,N_1589);
xor U1658 (N_1658,N_1577,N_1571);
nor U1659 (N_1659,N_1590,N_1600);
or U1660 (N_1660,N_1569,N_1573);
nor U1661 (N_1661,N_1579,N_1574);
or U1662 (N_1662,N_1564,N_1560);
and U1663 (N_1663,N_1604,N_1567);
xnor U1664 (N_1664,N_1610,N_1584);
or U1665 (N_1665,N_1611,N_1581);
nor U1666 (N_1666,N_1599,N_1582);
nand U1667 (N_1667,N_1592,N_1574);
nand U1668 (N_1668,N_1578,N_1579);
or U1669 (N_1669,N_1569,N_1612);
nand U1670 (N_1670,N_1592,N_1588);
xor U1671 (N_1671,N_1606,N_1607);
or U1672 (N_1672,N_1588,N_1595);
nor U1673 (N_1673,N_1574,N_1569);
nor U1674 (N_1674,N_1560,N_1580);
nand U1675 (N_1675,N_1616,N_1618);
or U1676 (N_1676,N_1570,N_1617);
nor U1677 (N_1677,N_1560,N_1575);
xnor U1678 (N_1678,N_1584,N_1617);
nor U1679 (N_1679,N_1579,N_1591);
nor U1680 (N_1680,N_1646,N_1621);
nor U1681 (N_1681,N_1671,N_1669);
xor U1682 (N_1682,N_1641,N_1668);
nand U1683 (N_1683,N_1670,N_1630);
nand U1684 (N_1684,N_1667,N_1662);
nand U1685 (N_1685,N_1663,N_1653);
nand U1686 (N_1686,N_1650,N_1645);
and U1687 (N_1687,N_1655,N_1626);
and U1688 (N_1688,N_1660,N_1627);
or U1689 (N_1689,N_1673,N_1675);
nand U1690 (N_1690,N_1664,N_1623);
nor U1691 (N_1691,N_1629,N_1659);
nor U1692 (N_1692,N_1622,N_1679);
and U1693 (N_1693,N_1634,N_1628);
xnor U1694 (N_1694,N_1656,N_1636);
nor U1695 (N_1695,N_1649,N_1639);
nor U1696 (N_1696,N_1674,N_1644);
nand U1697 (N_1697,N_1637,N_1648);
and U1698 (N_1698,N_1620,N_1678);
nor U1699 (N_1699,N_1642,N_1657);
or U1700 (N_1700,N_1632,N_1635);
and U1701 (N_1701,N_1638,N_1665);
nor U1702 (N_1702,N_1643,N_1647);
or U1703 (N_1703,N_1640,N_1666);
or U1704 (N_1704,N_1661,N_1652);
xor U1705 (N_1705,N_1658,N_1677);
or U1706 (N_1706,N_1651,N_1625);
xnor U1707 (N_1707,N_1676,N_1624);
and U1708 (N_1708,N_1672,N_1631);
nand U1709 (N_1709,N_1633,N_1654);
and U1710 (N_1710,N_1668,N_1644);
nor U1711 (N_1711,N_1633,N_1665);
and U1712 (N_1712,N_1628,N_1678);
xor U1713 (N_1713,N_1659,N_1632);
or U1714 (N_1714,N_1667,N_1639);
nor U1715 (N_1715,N_1649,N_1661);
nand U1716 (N_1716,N_1676,N_1626);
or U1717 (N_1717,N_1649,N_1655);
xnor U1718 (N_1718,N_1676,N_1634);
nor U1719 (N_1719,N_1651,N_1639);
xnor U1720 (N_1720,N_1634,N_1663);
nor U1721 (N_1721,N_1630,N_1651);
nand U1722 (N_1722,N_1645,N_1641);
nor U1723 (N_1723,N_1675,N_1663);
xor U1724 (N_1724,N_1647,N_1662);
and U1725 (N_1725,N_1666,N_1675);
nand U1726 (N_1726,N_1679,N_1671);
or U1727 (N_1727,N_1643,N_1651);
nand U1728 (N_1728,N_1650,N_1633);
xnor U1729 (N_1729,N_1657,N_1656);
xnor U1730 (N_1730,N_1675,N_1636);
or U1731 (N_1731,N_1658,N_1671);
xnor U1732 (N_1732,N_1628,N_1679);
and U1733 (N_1733,N_1672,N_1678);
nand U1734 (N_1734,N_1630,N_1679);
and U1735 (N_1735,N_1640,N_1630);
nor U1736 (N_1736,N_1630,N_1646);
nor U1737 (N_1737,N_1637,N_1643);
nand U1738 (N_1738,N_1664,N_1674);
nand U1739 (N_1739,N_1658,N_1668);
xor U1740 (N_1740,N_1691,N_1724);
or U1741 (N_1741,N_1697,N_1723);
xor U1742 (N_1742,N_1739,N_1719);
and U1743 (N_1743,N_1716,N_1727);
xnor U1744 (N_1744,N_1689,N_1738);
and U1745 (N_1745,N_1690,N_1737);
and U1746 (N_1746,N_1682,N_1709);
xnor U1747 (N_1747,N_1711,N_1692);
nor U1748 (N_1748,N_1681,N_1736);
xnor U1749 (N_1749,N_1732,N_1698);
xor U1750 (N_1750,N_1717,N_1725);
xnor U1751 (N_1751,N_1695,N_1718);
nor U1752 (N_1752,N_1706,N_1702);
nor U1753 (N_1753,N_1730,N_1708);
nor U1754 (N_1754,N_1731,N_1703);
nor U1755 (N_1755,N_1712,N_1710);
xor U1756 (N_1756,N_1699,N_1685);
and U1757 (N_1757,N_1696,N_1701);
xor U1758 (N_1758,N_1726,N_1722);
and U1759 (N_1759,N_1733,N_1734);
nor U1760 (N_1760,N_1735,N_1713);
xnor U1761 (N_1761,N_1720,N_1729);
xnor U1762 (N_1762,N_1687,N_1700);
nor U1763 (N_1763,N_1721,N_1686);
and U1764 (N_1764,N_1683,N_1704);
and U1765 (N_1765,N_1680,N_1693);
nor U1766 (N_1766,N_1705,N_1728);
and U1767 (N_1767,N_1707,N_1688);
and U1768 (N_1768,N_1684,N_1714);
xnor U1769 (N_1769,N_1715,N_1694);
nor U1770 (N_1770,N_1711,N_1703);
nand U1771 (N_1771,N_1732,N_1708);
xnor U1772 (N_1772,N_1713,N_1723);
nand U1773 (N_1773,N_1680,N_1728);
nand U1774 (N_1774,N_1735,N_1711);
nor U1775 (N_1775,N_1730,N_1723);
xnor U1776 (N_1776,N_1703,N_1688);
xor U1777 (N_1777,N_1696,N_1689);
nor U1778 (N_1778,N_1712,N_1718);
and U1779 (N_1779,N_1689,N_1716);
nand U1780 (N_1780,N_1693,N_1703);
and U1781 (N_1781,N_1703,N_1698);
xor U1782 (N_1782,N_1708,N_1690);
and U1783 (N_1783,N_1728,N_1703);
and U1784 (N_1784,N_1729,N_1688);
nor U1785 (N_1785,N_1686,N_1680);
xor U1786 (N_1786,N_1687,N_1698);
and U1787 (N_1787,N_1689,N_1704);
nor U1788 (N_1788,N_1689,N_1718);
or U1789 (N_1789,N_1681,N_1727);
and U1790 (N_1790,N_1703,N_1680);
and U1791 (N_1791,N_1708,N_1724);
nor U1792 (N_1792,N_1720,N_1699);
xor U1793 (N_1793,N_1703,N_1694);
nor U1794 (N_1794,N_1681,N_1709);
xnor U1795 (N_1795,N_1695,N_1737);
or U1796 (N_1796,N_1711,N_1698);
or U1797 (N_1797,N_1680,N_1691);
and U1798 (N_1798,N_1695,N_1729);
xor U1799 (N_1799,N_1710,N_1732);
and U1800 (N_1800,N_1782,N_1760);
nand U1801 (N_1801,N_1771,N_1747);
or U1802 (N_1802,N_1792,N_1797);
and U1803 (N_1803,N_1776,N_1783);
and U1804 (N_1804,N_1762,N_1790);
nand U1805 (N_1805,N_1780,N_1746);
nand U1806 (N_1806,N_1787,N_1794);
nor U1807 (N_1807,N_1784,N_1781);
nand U1808 (N_1808,N_1785,N_1769);
xnor U1809 (N_1809,N_1755,N_1754);
xor U1810 (N_1810,N_1750,N_1761);
xnor U1811 (N_1811,N_1768,N_1774);
nand U1812 (N_1812,N_1748,N_1743);
nand U1813 (N_1813,N_1751,N_1767);
xnor U1814 (N_1814,N_1796,N_1777);
xnor U1815 (N_1815,N_1740,N_1799);
and U1816 (N_1816,N_1752,N_1789);
nor U1817 (N_1817,N_1765,N_1753);
or U1818 (N_1818,N_1744,N_1798);
nand U1819 (N_1819,N_1779,N_1742);
xnor U1820 (N_1820,N_1793,N_1759);
xnor U1821 (N_1821,N_1775,N_1772);
nor U1822 (N_1822,N_1764,N_1770);
nand U1823 (N_1823,N_1745,N_1788);
nand U1824 (N_1824,N_1773,N_1757);
nor U1825 (N_1825,N_1741,N_1758);
nor U1826 (N_1826,N_1766,N_1791);
xor U1827 (N_1827,N_1756,N_1749);
nor U1828 (N_1828,N_1795,N_1763);
xor U1829 (N_1829,N_1786,N_1778);
xor U1830 (N_1830,N_1764,N_1771);
and U1831 (N_1831,N_1744,N_1768);
nand U1832 (N_1832,N_1749,N_1750);
and U1833 (N_1833,N_1782,N_1788);
nand U1834 (N_1834,N_1792,N_1796);
and U1835 (N_1835,N_1765,N_1762);
or U1836 (N_1836,N_1741,N_1743);
nand U1837 (N_1837,N_1773,N_1784);
xor U1838 (N_1838,N_1785,N_1744);
xor U1839 (N_1839,N_1749,N_1744);
xor U1840 (N_1840,N_1794,N_1749);
nand U1841 (N_1841,N_1770,N_1758);
xnor U1842 (N_1842,N_1755,N_1749);
xnor U1843 (N_1843,N_1798,N_1791);
and U1844 (N_1844,N_1759,N_1772);
or U1845 (N_1845,N_1751,N_1744);
xnor U1846 (N_1846,N_1776,N_1782);
nor U1847 (N_1847,N_1775,N_1788);
nor U1848 (N_1848,N_1769,N_1795);
nand U1849 (N_1849,N_1786,N_1744);
and U1850 (N_1850,N_1757,N_1795);
nand U1851 (N_1851,N_1792,N_1774);
xor U1852 (N_1852,N_1755,N_1769);
nand U1853 (N_1853,N_1792,N_1750);
and U1854 (N_1854,N_1749,N_1774);
xor U1855 (N_1855,N_1750,N_1784);
nor U1856 (N_1856,N_1779,N_1769);
nand U1857 (N_1857,N_1794,N_1784);
and U1858 (N_1858,N_1765,N_1766);
nand U1859 (N_1859,N_1795,N_1742);
xor U1860 (N_1860,N_1851,N_1807);
xnor U1861 (N_1861,N_1837,N_1850);
xor U1862 (N_1862,N_1804,N_1858);
nor U1863 (N_1863,N_1835,N_1821);
xnor U1864 (N_1864,N_1802,N_1831);
or U1865 (N_1865,N_1823,N_1853);
and U1866 (N_1866,N_1833,N_1852);
and U1867 (N_1867,N_1834,N_1813);
or U1868 (N_1868,N_1845,N_1839);
xor U1869 (N_1869,N_1838,N_1815);
nand U1870 (N_1870,N_1808,N_1803);
nor U1871 (N_1871,N_1827,N_1846);
nor U1872 (N_1872,N_1805,N_1849);
and U1873 (N_1873,N_1842,N_1857);
or U1874 (N_1874,N_1830,N_1856);
or U1875 (N_1875,N_1814,N_1819);
or U1876 (N_1876,N_1848,N_1847);
nand U1877 (N_1877,N_1844,N_1855);
and U1878 (N_1878,N_1810,N_1859);
xnor U1879 (N_1879,N_1806,N_1826);
xor U1880 (N_1880,N_1822,N_1825);
and U1881 (N_1881,N_1801,N_1811);
and U1882 (N_1882,N_1854,N_1843);
or U1883 (N_1883,N_1817,N_1809);
nor U1884 (N_1884,N_1820,N_1816);
xnor U1885 (N_1885,N_1832,N_1841);
and U1886 (N_1886,N_1812,N_1824);
xor U1887 (N_1887,N_1818,N_1828);
or U1888 (N_1888,N_1829,N_1836);
or U1889 (N_1889,N_1800,N_1840);
nand U1890 (N_1890,N_1859,N_1831);
or U1891 (N_1891,N_1853,N_1802);
nor U1892 (N_1892,N_1831,N_1848);
nand U1893 (N_1893,N_1848,N_1840);
nor U1894 (N_1894,N_1810,N_1843);
nand U1895 (N_1895,N_1819,N_1804);
nand U1896 (N_1896,N_1823,N_1842);
and U1897 (N_1897,N_1844,N_1835);
nor U1898 (N_1898,N_1812,N_1856);
nor U1899 (N_1899,N_1840,N_1841);
and U1900 (N_1900,N_1850,N_1820);
or U1901 (N_1901,N_1844,N_1845);
nor U1902 (N_1902,N_1830,N_1800);
nor U1903 (N_1903,N_1840,N_1834);
xnor U1904 (N_1904,N_1838,N_1812);
xnor U1905 (N_1905,N_1805,N_1855);
xnor U1906 (N_1906,N_1835,N_1849);
nor U1907 (N_1907,N_1817,N_1826);
nand U1908 (N_1908,N_1839,N_1819);
or U1909 (N_1909,N_1819,N_1857);
xor U1910 (N_1910,N_1802,N_1854);
and U1911 (N_1911,N_1806,N_1833);
nand U1912 (N_1912,N_1812,N_1818);
xnor U1913 (N_1913,N_1831,N_1854);
nor U1914 (N_1914,N_1839,N_1841);
nor U1915 (N_1915,N_1821,N_1837);
or U1916 (N_1916,N_1828,N_1858);
xor U1917 (N_1917,N_1855,N_1846);
and U1918 (N_1918,N_1855,N_1806);
nor U1919 (N_1919,N_1835,N_1841);
nand U1920 (N_1920,N_1862,N_1880);
xor U1921 (N_1921,N_1866,N_1894);
and U1922 (N_1922,N_1873,N_1863);
nand U1923 (N_1923,N_1882,N_1870);
and U1924 (N_1924,N_1879,N_1919);
nor U1925 (N_1925,N_1913,N_1915);
nor U1926 (N_1926,N_1878,N_1907);
nand U1927 (N_1927,N_1892,N_1872);
and U1928 (N_1928,N_1902,N_1898);
nand U1929 (N_1929,N_1917,N_1876);
nand U1930 (N_1930,N_1884,N_1916);
nor U1931 (N_1931,N_1891,N_1867);
nand U1932 (N_1932,N_1893,N_1910);
nand U1933 (N_1933,N_1908,N_1912);
nand U1934 (N_1934,N_1909,N_1885);
nand U1935 (N_1935,N_1904,N_1911);
xnor U1936 (N_1936,N_1861,N_1914);
or U1937 (N_1937,N_1869,N_1888);
nand U1938 (N_1938,N_1889,N_1864);
or U1939 (N_1939,N_1865,N_1874);
and U1940 (N_1940,N_1886,N_1905);
nand U1941 (N_1941,N_1875,N_1906);
xor U1942 (N_1942,N_1881,N_1900);
or U1943 (N_1943,N_1887,N_1896);
or U1944 (N_1944,N_1918,N_1890);
nor U1945 (N_1945,N_1895,N_1871);
nand U1946 (N_1946,N_1883,N_1901);
or U1947 (N_1947,N_1868,N_1877);
xor U1948 (N_1948,N_1897,N_1903);
and U1949 (N_1949,N_1860,N_1899);
or U1950 (N_1950,N_1903,N_1899);
or U1951 (N_1951,N_1882,N_1901);
nand U1952 (N_1952,N_1912,N_1906);
xor U1953 (N_1953,N_1909,N_1913);
xnor U1954 (N_1954,N_1918,N_1884);
and U1955 (N_1955,N_1874,N_1913);
nand U1956 (N_1956,N_1902,N_1909);
and U1957 (N_1957,N_1882,N_1881);
nor U1958 (N_1958,N_1887,N_1907);
nor U1959 (N_1959,N_1915,N_1902);
xnor U1960 (N_1960,N_1887,N_1917);
nor U1961 (N_1961,N_1917,N_1877);
or U1962 (N_1962,N_1880,N_1872);
xor U1963 (N_1963,N_1860,N_1917);
or U1964 (N_1964,N_1903,N_1865);
nor U1965 (N_1965,N_1894,N_1873);
and U1966 (N_1966,N_1873,N_1883);
nand U1967 (N_1967,N_1881,N_1883);
and U1968 (N_1968,N_1891,N_1864);
nor U1969 (N_1969,N_1906,N_1862);
nand U1970 (N_1970,N_1902,N_1918);
and U1971 (N_1971,N_1888,N_1904);
nand U1972 (N_1972,N_1910,N_1873);
nor U1973 (N_1973,N_1900,N_1869);
nor U1974 (N_1974,N_1880,N_1860);
xor U1975 (N_1975,N_1886,N_1916);
nand U1976 (N_1976,N_1903,N_1898);
and U1977 (N_1977,N_1910,N_1911);
xnor U1978 (N_1978,N_1907,N_1918);
or U1979 (N_1979,N_1891,N_1863);
or U1980 (N_1980,N_1974,N_1972);
nand U1981 (N_1981,N_1957,N_1941);
xnor U1982 (N_1982,N_1979,N_1938);
or U1983 (N_1983,N_1936,N_1970);
nor U1984 (N_1984,N_1920,N_1930);
and U1985 (N_1985,N_1944,N_1964);
and U1986 (N_1986,N_1942,N_1962);
nor U1987 (N_1987,N_1955,N_1969);
xnor U1988 (N_1988,N_1978,N_1924);
and U1989 (N_1989,N_1929,N_1965);
xnor U1990 (N_1990,N_1943,N_1939);
or U1991 (N_1991,N_1968,N_1960);
and U1992 (N_1992,N_1958,N_1946);
xor U1993 (N_1993,N_1947,N_1976);
or U1994 (N_1994,N_1954,N_1948);
xor U1995 (N_1995,N_1975,N_1926);
and U1996 (N_1996,N_1923,N_1927);
nand U1997 (N_1997,N_1934,N_1956);
and U1998 (N_1998,N_1971,N_1977);
and U1999 (N_1999,N_1950,N_1953);
nor U2000 (N_2000,N_1922,N_1961);
and U2001 (N_2001,N_1945,N_1931);
or U2002 (N_2002,N_1963,N_1959);
nor U2003 (N_2003,N_1932,N_1966);
xnor U2004 (N_2004,N_1935,N_1928);
and U2005 (N_2005,N_1925,N_1933);
xor U2006 (N_2006,N_1973,N_1921);
nor U2007 (N_2007,N_1949,N_1940);
nand U2008 (N_2008,N_1937,N_1951);
xor U2009 (N_2009,N_1967,N_1952);
nand U2010 (N_2010,N_1976,N_1941);
and U2011 (N_2011,N_1974,N_1959);
or U2012 (N_2012,N_1933,N_1939);
nor U2013 (N_2013,N_1972,N_1944);
nand U2014 (N_2014,N_1970,N_1940);
xnor U2015 (N_2015,N_1924,N_1933);
and U2016 (N_2016,N_1929,N_1948);
xor U2017 (N_2017,N_1938,N_1966);
or U2018 (N_2018,N_1969,N_1956);
nand U2019 (N_2019,N_1954,N_1953);
nand U2020 (N_2020,N_1971,N_1936);
nor U2021 (N_2021,N_1931,N_1946);
or U2022 (N_2022,N_1974,N_1943);
and U2023 (N_2023,N_1977,N_1974);
or U2024 (N_2024,N_1934,N_1970);
nand U2025 (N_2025,N_1966,N_1933);
or U2026 (N_2026,N_1939,N_1938);
xor U2027 (N_2027,N_1945,N_1974);
xor U2028 (N_2028,N_1958,N_1932);
or U2029 (N_2029,N_1954,N_1965);
or U2030 (N_2030,N_1957,N_1943);
nor U2031 (N_2031,N_1978,N_1930);
nor U2032 (N_2032,N_1931,N_1935);
and U2033 (N_2033,N_1978,N_1960);
and U2034 (N_2034,N_1943,N_1940);
or U2035 (N_2035,N_1956,N_1950);
or U2036 (N_2036,N_1957,N_1964);
or U2037 (N_2037,N_1958,N_1944);
nor U2038 (N_2038,N_1966,N_1970);
or U2039 (N_2039,N_1927,N_1974);
xor U2040 (N_2040,N_2001,N_2030);
or U2041 (N_2041,N_2021,N_2000);
nand U2042 (N_2042,N_2033,N_2026);
xnor U2043 (N_2043,N_1982,N_2011);
xnor U2044 (N_2044,N_2018,N_2019);
xor U2045 (N_2045,N_1998,N_1996);
nand U2046 (N_2046,N_2013,N_2032);
nand U2047 (N_2047,N_2022,N_1987);
or U2048 (N_2048,N_1980,N_2023);
or U2049 (N_2049,N_1992,N_2028);
nor U2050 (N_2050,N_1997,N_2015);
xor U2051 (N_2051,N_1999,N_2039);
and U2052 (N_2052,N_2031,N_2008);
nand U2053 (N_2053,N_2027,N_2029);
nor U2054 (N_2054,N_2034,N_2037);
xor U2055 (N_2055,N_2010,N_1984);
and U2056 (N_2056,N_1995,N_2038);
nor U2057 (N_2057,N_2017,N_1985);
nand U2058 (N_2058,N_1989,N_2014);
or U2059 (N_2059,N_2009,N_1991);
nand U2060 (N_2060,N_2004,N_1983);
nor U2061 (N_2061,N_1988,N_2035);
xor U2062 (N_2062,N_1994,N_2024);
xor U2063 (N_2063,N_2012,N_1993);
and U2064 (N_2064,N_2006,N_1981);
nor U2065 (N_2065,N_1990,N_1986);
xnor U2066 (N_2066,N_2003,N_2020);
or U2067 (N_2067,N_2025,N_2005);
nand U2068 (N_2068,N_2007,N_2002);
and U2069 (N_2069,N_2016,N_2036);
xnor U2070 (N_2070,N_2001,N_2023);
nand U2071 (N_2071,N_1992,N_2026);
or U2072 (N_2072,N_2025,N_2015);
nor U2073 (N_2073,N_2004,N_1980);
and U2074 (N_2074,N_2008,N_2012);
nand U2075 (N_2075,N_1980,N_2016);
nand U2076 (N_2076,N_2038,N_1987);
or U2077 (N_2077,N_2017,N_2033);
nand U2078 (N_2078,N_2039,N_1987);
and U2079 (N_2079,N_2029,N_2003);
or U2080 (N_2080,N_2024,N_1998);
or U2081 (N_2081,N_2021,N_1991);
and U2082 (N_2082,N_2038,N_2001);
nand U2083 (N_2083,N_2021,N_2018);
nor U2084 (N_2084,N_2015,N_2038);
nand U2085 (N_2085,N_2031,N_1990);
or U2086 (N_2086,N_2035,N_2039);
and U2087 (N_2087,N_2002,N_1988);
nor U2088 (N_2088,N_2016,N_1985);
nand U2089 (N_2089,N_2003,N_1988);
and U2090 (N_2090,N_2004,N_1986);
xnor U2091 (N_2091,N_1989,N_2031);
and U2092 (N_2092,N_2029,N_2036);
nor U2093 (N_2093,N_2000,N_2017);
xor U2094 (N_2094,N_2015,N_2020);
and U2095 (N_2095,N_2015,N_2032);
xor U2096 (N_2096,N_2012,N_2017);
nand U2097 (N_2097,N_1994,N_2038);
or U2098 (N_2098,N_2013,N_2017);
nor U2099 (N_2099,N_2030,N_1999);
and U2100 (N_2100,N_2069,N_2055);
nor U2101 (N_2101,N_2095,N_2094);
or U2102 (N_2102,N_2090,N_2080);
xnor U2103 (N_2103,N_2053,N_2056);
xor U2104 (N_2104,N_2076,N_2040);
or U2105 (N_2105,N_2081,N_2078);
nand U2106 (N_2106,N_2070,N_2082);
nand U2107 (N_2107,N_2065,N_2072);
and U2108 (N_2108,N_2099,N_2071);
nand U2109 (N_2109,N_2073,N_2077);
nand U2110 (N_2110,N_2074,N_2085);
nand U2111 (N_2111,N_2096,N_2050);
nand U2112 (N_2112,N_2097,N_2062);
nor U2113 (N_2113,N_2079,N_2052);
nor U2114 (N_2114,N_2054,N_2042);
or U2115 (N_2115,N_2087,N_2058);
nand U2116 (N_2116,N_2048,N_2088);
nor U2117 (N_2117,N_2046,N_2084);
nor U2118 (N_2118,N_2075,N_2093);
or U2119 (N_2119,N_2045,N_2057);
or U2120 (N_2120,N_2067,N_2063);
xnor U2121 (N_2121,N_2049,N_2089);
or U2122 (N_2122,N_2051,N_2041);
and U2123 (N_2123,N_2068,N_2044);
xnor U2124 (N_2124,N_2083,N_2086);
and U2125 (N_2125,N_2047,N_2066);
xor U2126 (N_2126,N_2091,N_2064);
and U2127 (N_2127,N_2059,N_2060);
nor U2128 (N_2128,N_2061,N_2043);
and U2129 (N_2129,N_2098,N_2092);
nor U2130 (N_2130,N_2069,N_2077);
or U2131 (N_2131,N_2066,N_2078);
or U2132 (N_2132,N_2099,N_2095);
xnor U2133 (N_2133,N_2069,N_2060);
or U2134 (N_2134,N_2064,N_2052);
nor U2135 (N_2135,N_2054,N_2074);
or U2136 (N_2136,N_2060,N_2094);
nand U2137 (N_2137,N_2049,N_2085);
nor U2138 (N_2138,N_2040,N_2065);
nand U2139 (N_2139,N_2078,N_2091);
xnor U2140 (N_2140,N_2081,N_2044);
nand U2141 (N_2141,N_2096,N_2040);
or U2142 (N_2142,N_2058,N_2051);
and U2143 (N_2143,N_2062,N_2092);
and U2144 (N_2144,N_2079,N_2084);
nor U2145 (N_2145,N_2094,N_2055);
nor U2146 (N_2146,N_2068,N_2050);
nand U2147 (N_2147,N_2052,N_2043);
and U2148 (N_2148,N_2061,N_2089);
nor U2149 (N_2149,N_2061,N_2082);
and U2150 (N_2150,N_2073,N_2046);
nor U2151 (N_2151,N_2056,N_2040);
nor U2152 (N_2152,N_2081,N_2084);
and U2153 (N_2153,N_2043,N_2060);
nand U2154 (N_2154,N_2087,N_2067);
xnor U2155 (N_2155,N_2089,N_2076);
or U2156 (N_2156,N_2052,N_2055);
xnor U2157 (N_2157,N_2051,N_2057);
nor U2158 (N_2158,N_2095,N_2059);
xor U2159 (N_2159,N_2096,N_2053);
nor U2160 (N_2160,N_2113,N_2124);
xor U2161 (N_2161,N_2128,N_2130);
nand U2162 (N_2162,N_2146,N_2108);
nand U2163 (N_2163,N_2112,N_2103);
and U2164 (N_2164,N_2137,N_2117);
or U2165 (N_2165,N_2102,N_2155);
or U2166 (N_2166,N_2123,N_2119);
nand U2167 (N_2167,N_2133,N_2144);
nor U2168 (N_2168,N_2142,N_2140);
nor U2169 (N_2169,N_2118,N_2121);
and U2170 (N_2170,N_2159,N_2106);
and U2171 (N_2171,N_2135,N_2158);
xor U2172 (N_2172,N_2139,N_2148);
or U2173 (N_2173,N_2105,N_2151);
nor U2174 (N_2174,N_2157,N_2126);
nand U2175 (N_2175,N_2145,N_2132);
xor U2176 (N_2176,N_2101,N_2125);
nand U2177 (N_2177,N_2152,N_2122);
or U2178 (N_2178,N_2136,N_2100);
xor U2179 (N_2179,N_2116,N_2111);
xor U2180 (N_2180,N_2115,N_2156);
or U2181 (N_2181,N_2153,N_2154);
xnor U2182 (N_2182,N_2104,N_2129);
nor U2183 (N_2183,N_2149,N_2141);
xor U2184 (N_2184,N_2107,N_2110);
nand U2185 (N_2185,N_2114,N_2109);
nand U2186 (N_2186,N_2138,N_2134);
nand U2187 (N_2187,N_2127,N_2143);
and U2188 (N_2188,N_2150,N_2131);
nand U2189 (N_2189,N_2120,N_2147);
xor U2190 (N_2190,N_2159,N_2136);
and U2191 (N_2191,N_2135,N_2142);
nand U2192 (N_2192,N_2106,N_2105);
nand U2193 (N_2193,N_2148,N_2112);
nor U2194 (N_2194,N_2131,N_2151);
or U2195 (N_2195,N_2100,N_2147);
xnor U2196 (N_2196,N_2155,N_2141);
or U2197 (N_2197,N_2142,N_2141);
or U2198 (N_2198,N_2142,N_2122);
or U2199 (N_2199,N_2124,N_2111);
or U2200 (N_2200,N_2149,N_2154);
and U2201 (N_2201,N_2126,N_2116);
xnor U2202 (N_2202,N_2141,N_2138);
nand U2203 (N_2203,N_2135,N_2111);
or U2204 (N_2204,N_2141,N_2156);
nor U2205 (N_2205,N_2105,N_2126);
or U2206 (N_2206,N_2104,N_2124);
or U2207 (N_2207,N_2123,N_2139);
xnor U2208 (N_2208,N_2105,N_2142);
nand U2209 (N_2209,N_2147,N_2138);
or U2210 (N_2210,N_2101,N_2103);
nor U2211 (N_2211,N_2100,N_2115);
xnor U2212 (N_2212,N_2158,N_2113);
or U2213 (N_2213,N_2159,N_2124);
or U2214 (N_2214,N_2107,N_2143);
xnor U2215 (N_2215,N_2119,N_2149);
or U2216 (N_2216,N_2122,N_2117);
xor U2217 (N_2217,N_2127,N_2150);
nand U2218 (N_2218,N_2154,N_2152);
xnor U2219 (N_2219,N_2151,N_2149);
or U2220 (N_2220,N_2215,N_2185);
and U2221 (N_2221,N_2162,N_2187);
nor U2222 (N_2222,N_2204,N_2200);
nand U2223 (N_2223,N_2163,N_2195);
xor U2224 (N_2224,N_2219,N_2205);
nor U2225 (N_2225,N_2184,N_2206);
and U2226 (N_2226,N_2161,N_2172);
nand U2227 (N_2227,N_2176,N_2193);
and U2228 (N_2228,N_2173,N_2191);
or U2229 (N_2229,N_2192,N_2214);
and U2230 (N_2230,N_2216,N_2198);
nand U2231 (N_2231,N_2186,N_2208);
and U2232 (N_2232,N_2197,N_2211);
nor U2233 (N_2233,N_2170,N_2171);
and U2234 (N_2234,N_2203,N_2181);
nand U2235 (N_2235,N_2177,N_2210);
nor U2236 (N_2236,N_2194,N_2178);
xnor U2237 (N_2237,N_2207,N_2180);
and U2238 (N_2238,N_2212,N_2218);
or U2239 (N_2239,N_2188,N_2183);
nor U2240 (N_2240,N_2166,N_2167);
nand U2241 (N_2241,N_2182,N_2160);
or U2242 (N_2242,N_2209,N_2190);
nand U2243 (N_2243,N_2217,N_2202);
or U2244 (N_2244,N_2196,N_2168);
nand U2245 (N_2245,N_2165,N_2199);
xor U2246 (N_2246,N_2174,N_2164);
and U2247 (N_2247,N_2189,N_2169);
nor U2248 (N_2248,N_2213,N_2201);
nor U2249 (N_2249,N_2175,N_2179);
nand U2250 (N_2250,N_2190,N_2208);
nor U2251 (N_2251,N_2218,N_2164);
xnor U2252 (N_2252,N_2160,N_2219);
nor U2253 (N_2253,N_2188,N_2208);
and U2254 (N_2254,N_2205,N_2160);
nand U2255 (N_2255,N_2169,N_2178);
and U2256 (N_2256,N_2216,N_2163);
xnor U2257 (N_2257,N_2164,N_2190);
nor U2258 (N_2258,N_2215,N_2189);
nor U2259 (N_2259,N_2162,N_2165);
nor U2260 (N_2260,N_2166,N_2216);
xor U2261 (N_2261,N_2168,N_2191);
nor U2262 (N_2262,N_2169,N_2179);
or U2263 (N_2263,N_2198,N_2185);
nand U2264 (N_2264,N_2188,N_2203);
or U2265 (N_2265,N_2180,N_2219);
and U2266 (N_2266,N_2162,N_2161);
or U2267 (N_2267,N_2161,N_2178);
nor U2268 (N_2268,N_2205,N_2172);
and U2269 (N_2269,N_2216,N_2171);
nor U2270 (N_2270,N_2185,N_2164);
nor U2271 (N_2271,N_2192,N_2179);
and U2272 (N_2272,N_2167,N_2189);
and U2273 (N_2273,N_2207,N_2210);
xnor U2274 (N_2274,N_2172,N_2198);
or U2275 (N_2275,N_2219,N_2208);
nor U2276 (N_2276,N_2205,N_2184);
nor U2277 (N_2277,N_2178,N_2160);
xor U2278 (N_2278,N_2201,N_2185);
nor U2279 (N_2279,N_2197,N_2176);
xor U2280 (N_2280,N_2262,N_2236);
and U2281 (N_2281,N_2275,N_2249);
and U2282 (N_2282,N_2263,N_2279);
nand U2283 (N_2283,N_2222,N_2226);
xor U2284 (N_2284,N_2235,N_2239);
nor U2285 (N_2285,N_2243,N_2278);
and U2286 (N_2286,N_2265,N_2264);
or U2287 (N_2287,N_2257,N_2224);
xor U2288 (N_2288,N_2229,N_2227);
nor U2289 (N_2289,N_2241,N_2261);
nand U2290 (N_2290,N_2271,N_2255);
or U2291 (N_2291,N_2245,N_2274);
and U2292 (N_2292,N_2260,N_2270);
nand U2293 (N_2293,N_2221,N_2266);
or U2294 (N_2294,N_2228,N_2277);
nor U2295 (N_2295,N_2272,N_2269);
or U2296 (N_2296,N_2256,N_2220);
nand U2297 (N_2297,N_2233,N_2231);
nor U2298 (N_2298,N_2248,N_2247);
or U2299 (N_2299,N_2276,N_2251);
nand U2300 (N_2300,N_2240,N_2232);
xnor U2301 (N_2301,N_2230,N_2252);
and U2302 (N_2302,N_2254,N_2223);
nand U2303 (N_2303,N_2268,N_2238);
nand U2304 (N_2304,N_2234,N_2253);
and U2305 (N_2305,N_2242,N_2267);
and U2306 (N_2306,N_2237,N_2258);
xor U2307 (N_2307,N_2246,N_2273);
or U2308 (N_2308,N_2225,N_2244);
and U2309 (N_2309,N_2250,N_2259);
xnor U2310 (N_2310,N_2248,N_2259);
nor U2311 (N_2311,N_2235,N_2266);
xnor U2312 (N_2312,N_2270,N_2252);
and U2313 (N_2313,N_2261,N_2228);
nand U2314 (N_2314,N_2264,N_2255);
nand U2315 (N_2315,N_2271,N_2228);
nor U2316 (N_2316,N_2220,N_2230);
nor U2317 (N_2317,N_2258,N_2234);
xor U2318 (N_2318,N_2227,N_2220);
nor U2319 (N_2319,N_2279,N_2271);
or U2320 (N_2320,N_2234,N_2266);
xnor U2321 (N_2321,N_2242,N_2274);
nand U2322 (N_2322,N_2264,N_2222);
nand U2323 (N_2323,N_2279,N_2254);
nand U2324 (N_2324,N_2249,N_2258);
or U2325 (N_2325,N_2252,N_2256);
nand U2326 (N_2326,N_2244,N_2222);
and U2327 (N_2327,N_2224,N_2252);
nor U2328 (N_2328,N_2229,N_2259);
or U2329 (N_2329,N_2252,N_2267);
or U2330 (N_2330,N_2228,N_2233);
xnor U2331 (N_2331,N_2270,N_2222);
and U2332 (N_2332,N_2279,N_2241);
nor U2333 (N_2333,N_2262,N_2276);
nor U2334 (N_2334,N_2258,N_2224);
or U2335 (N_2335,N_2231,N_2238);
and U2336 (N_2336,N_2222,N_2256);
or U2337 (N_2337,N_2249,N_2270);
nand U2338 (N_2338,N_2254,N_2249);
nand U2339 (N_2339,N_2248,N_2249);
nor U2340 (N_2340,N_2295,N_2311);
xnor U2341 (N_2341,N_2334,N_2280);
nand U2342 (N_2342,N_2327,N_2332);
and U2343 (N_2343,N_2296,N_2310);
nor U2344 (N_2344,N_2305,N_2323);
and U2345 (N_2345,N_2307,N_2281);
nor U2346 (N_2346,N_2330,N_2335);
nand U2347 (N_2347,N_2285,N_2338);
or U2348 (N_2348,N_2326,N_2293);
and U2349 (N_2349,N_2325,N_2319);
nand U2350 (N_2350,N_2292,N_2304);
or U2351 (N_2351,N_2312,N_2282);
or U2352 (N_2352,N_2317,N_2289);
and U2353 (N_2353,N_2333,N_2300);
or U2354 (N_2354,N_2320,N_2337);
or U2355 (N_2355,N_2336,N_2314);
xor U2356 (N_2356,N_2297,N_2313);
nand U2357 (N_2357,N_2284,N_2287);
nor U2358 (N_2358,N_2315,N_2316);
xor U2359 (N_2359,N_2324,N_2294);
or U2360 (N_2360,N_2288,N_2299);
nor U2361 (N_2361,N_2309,N_2302);
nand U2362 (N_2362,N_2301,N_2339);
and U2363 (N_2363,N_2283,N_2291);
nand U2364 (N_2364,N_2329,N_2298);
xnor U2365 (N_2365,N_2286,N_2308);
nand U2366 (N_2366,N_2328,N_2321);
and U2367 (N_2367,N_2303,N_2331);
nand U2368 (N_2368,N_2290,N_2318);
nor U2369 (N_2369,N_2322,N_2306);
and U2370 (N_2370,N_2285,N_2314);
and U2371 (N_2371,N_2324,N_2319);
nand U2372 (N_2372,N_2295,N_2312);
or U2373 (N_2373,N_2328,N_2282);
nand U2374 (N_2374,N_2282,N_2329);
nand U2375 (N_2375,N_2309,N_2310);
xnor U2376 (N_2376,N_2294,N_2291);
nand U2377 (N_2377,N_2318,N_2306);
and U2378 (N_2378,N_2328,N_2296);
nand U2379 (N_2379,N_2324,N_2292);
nor U2380 (N_2380,N_2330,N_2327);
xor U2381 (N_2381,N_2318,N_2304);
xnor U2382 (N_2382,N_2336,N_2297);
xor U2383 (N_2383,N_2326,N_2305);
or U2384 (N_2384,N_2298,N_2304);
or U2385 (N_2385,N_2285,N_2311);
and U2386 (N_2386,N_2290,N_2306);
and U2387 (N_2387,N_2303,N_2293);
nand U2388 (N_2388,N_2304,N_2306);
or U2389 (N_2389,N_2298,N_2305);
nor U2390 (N_2390,N_2311,N_2300);
nor U2391 (N_2391,N_2309,N_2315);
or U2392 (N_2392,N_2291,N_2286);
xor U2393 (N_2393,N_2316,N_2330);
or U2394 (N_2394,N_2333,N_2307);
and U2395 (N_2395,N_2282,N_2292);
nor U2396 (N_2396,N_2309,N_2295);
and U2397 (N_2397,N_2305,N_2330);
or U2398 (N_2398,N_2314,N_2299);
nor U2399 (N_2399,N_2313,N_2306);
nand U2400 (N_2400,N_2395,N_2386);
xor U2401 (N_2401,N_2380,N_2344);
nand U2402 (N_2402,N_2371,N_2364);
nand U2403 (N_2403,N_2373,N_2341);
or U2404 (N_2404,N_2399,N_2357);
xor U2405 (N_2405,N_2394,N_2393);
nor U2406 (N_2406,N_2388,N_2392);
nand U2407 (N_2407,N_2366,N_2363);
xnor U2408 (N_2408,N_2375,N_2355);
nand U2409 (N_2409,N_2384,N_2389);
xor U2410 (N_2410,N_2359,N_2346);
nand U2411 (N_2411,N_2352,N_2374);
nand U2412 (N_2412,N_2387,N_2390);
and U2413 (N_2413,N_2368,N_2396);
nand U2414 (N_2414,N_2376,N_2377);
or U2415 (N_2415,N_2351,N_2360);
or U2416 (N_2416,N_2361,N_2340);
nand U2417 (N_2417,N_2342,N_2369);
xor U2418 (N_2418,N_2354,N_2349);
nor U2419 (N_2419,N_2348,N_2383);
and U2420 (N_2420,N_2358,N_2378);
xor U2421 (N_2421,N_2353,N_2391);
nor U2422 (N_2422,N_2382,N_2367);
nor U2423 (N_2423,N_2362,N_2398);
and U2424 (N_2424,N_2350,N_2365);
nand U2425 (N_2425,N_2397,N_2379);
and U2426 (N_2426,N_2370,N_2356);
nand U2427 (N_2427,N_2372,N_2345);
and U2428 (N_2428,N_2381,N_2385);
nand U2429 (N_2429,N_2347,N_2343);
or U2430 (N_2430,N_2383,N_2373);
or U2431 (N_2431,N_2385,N_2386);
nor U2432 (N_2432,N_2393,N_2366);
nand U2433 (N_2433,N_2355,N_2365);
nor U2434 (N_2434,N_2366,N_2388);
nand U2435 (N_2435,N_2376,N_2374);
nand U2436 (N_2436,N_2392,N_2354);
nor U2437 (N_2437,N_2372,N_2354);
and U2438 (N_2438,N_2342,N_2370);
nand U2439 (N_2439,N_2340,N_2351);
nor U2440 (N_2440,N_2354,N_2389);
xnor U2441 (N_2441,N_2390,N_2378);
or U2442 (N_2442,N_2387,N_2399);
nor U2443 (N_2443,N_2353,N_2358);
or U2444 (N_2444,N_2386,N_2382);
xor U2445 (N_2445,N_2377,N_2396);
xnor U2446 (N_2446,N_2362,N_2397);
and U2447 (N_2447,N_2354,N_2365);
xor U2448 (N_2448,N_2380,N_2341);
xor U2449 (N_2449,N_2397,N_2356);
or U2450 (N_2450,N_2345,N_2377);
and U2451 (N_2451,N_2397,N_2349);
nor U2452 (N_2452,N_2357,N_2366);
and U2453 (N_2453,N_2361,N_2398);
and U2454 (N_2454,N_2387,N_2382);
nor U2455 (N_2455,N_2364,N_2342);
and U2456 (N_2456,N_2355,N_2374);
xor U2457 (N_2457,N_2364,N_2368);
nor U2458 (N_2458,N_2372,N_2357);
or U2459 (N_2459,N_2371,N_2362);
nor U2460 (N_2460,N_2458,N_2436);
nand U2461 (N_2461,N_2421,N_2404);
nand U2462 (N_2462,N_2418,N_2427);
xor U2463 (N_2463,N_2405,N_2417);
nand U2464 (N_2464,N_2434,N_2401);
nand U2465 (N_2465,N_2438,N_2420);
or U2466 (N_2466,N_2450,N_2451);
or U2467 (N_2467,N_2416,N_2412);
nand U2468 (N_2468,N_2435,N_2407);
nor U2469 (N_2469,N_2400,N_2430);
and U2470 (N_2470,N_2449,N_2459);
and U2471 (N_2471,N_2456,N_2415);
nor U2472 (N_2472,N_2428,N_2419);
and U2473 (N_2473,N_2432,N_2442);
nor U2474 (N_2474,N_2444,N_2409);
and U2475 (N_2475,N_2424,N_2455);
and U2476 (N_2476,N_2410,N_2423);
nand U2477 (N_2477,N_2403,N_2452);
nand U2478 (N_2478,N_2446,N_2457);
nor U2479 (N_2479,N_2441,N_2439);
or U2480 (N_2480,N_2413,N_2411);
and U2481 (N_2481,N_2453,N_2408);
or U2482 (N_2482,N_2454,N_2447);
nor U2483 (N_2483,N_2433,N_2443);
and U2484 (N_2484,N_2431,N_2445);
and U2485 (N_2485,N_2429,N_2425);
nand U2486 (N_2486,N_2422,N_2448);
xor U2487 (N_2487,N_2437,N_2440);
and U2488 (N_2488,N_2426,N_2406);
or U2489 (N_2489,N_2402,N_2414);
or U2490 (N_2490,N_2403,N_2455);
nor U2491 (N_2491,N_2402,N_2444);
nor U2492 (N_2492,N_2444,N_2411);
nor U2493 (N_2493,N_2414,N_2415);
or U2494 (N_2494,N_2427,N_2404);
or U2495 (N_2495,N_2402,N_2423);
or U2496 (N_2496,N_2437,N_2425);
nand U2497 (N_2497,N_2436,N_2445);
or U2498 (N_2498,N_2452,N_2432);
and U2499 (N_2499,N_2428,N_2410);
or U2500 (N_2500,N_2444,N_2450);
xnor U2501 (N_2501,N_2445,N_2435);
and U2502 (N_2502,N_2415,N_2453);
or U2503 (N_2503,N_2411,N_2441);
and U2504 (N_2504,N_2414,N_2435);
nor U2505 (N_2505,N_2443,N_2441);
or U2506 (N_2506,N_2434,N_2435);
or U2507 (N_2507,N_2448,N_2441);
nor U2508 (N_2508,N_2400,N_2428);
xor U2509 (N_2509,N_2444,N_2400);
xnor U2510 (N_2510,N_2413,N_2424);
and U2511 (N_2511,N_2408,N_2450);
xnor U2512 (N_2512,N_2439,N_2416);
nand U2513 (N_2513,N_2412,N_2444);
nand U2514 (N_2514,N_2404,N_2432);
or U2515 (N_2515,N_2436,N_2434);
or U2516 (N_2516,N_2425,N_2413);
xnor U2517 (N_2517,N_2413,N_2435);
nand U2518 (N_2518,N_2410,N_2417);
or U2519 (N_2519,N_2454,N_2435);
xnor U2520 (N_2520,N_2486,N_2496);
and U2521 (N_2521,N_2485,N_2519);
and U2522 (N_2522,N_2503,N_2494);
and U2523 (N_2523,N_2472,N_2488);
nor U2524 (N_2524,N_2492,N_2468);
nor U2525 (N_2525,N_2465,N_2506);
and U2526 (N_2526,N_2510,N_2463);
and U2527 (N_2527,N_2516,N_2469);
xor U2528 (N_2528,N_2489,N_2514);
and U2529 (N_2529,N_2493,N_2475);
nor U2530 (N_2530,N_2499,N_2467);
nand U2531 (N_2531,N_2481,N_2495);
nand U2532 (N_2532,N_2487,N_2515);
or U2533 (N_2533,N_2464,N_2476);
and U2534 (N_2534,N_2474,N_2471);
nand U2535 (N_2535,N_2482,N_2484);
xnor U2536 (N_2536,N_2466,N_2505);
xor U2537 (N_2537,N_2498,N_2517);
nor U2538 (N_2538,N_2508,N_2507);
nor U2539 (N_2539,N_2461,N_2483);
and U2540 (N_2540,N_2518,N_2460);
xnor U2541 (N_2541,N_2497,N_2513);
or U2542 (N_2542,N_2480,N_2470);
and U2543 (N_2543,N_2509,N_2462);
and U2544 (N_2544,N_2479,N_2478);
and U2545 (N_2545,N_2500,N_2477);
nand U2546 (N_2546,N_2511,N_2473);
xor U2547 (N_2547,N_2504,N_2502);
xor U2548 (N_2548,N_2491,N_2490);
nand U2549 (N_2549,N_2512,N_2501);
or U2550 (N_2550,N_2486,N_2507);
nor U2551 (N_2551,N_2519,N_2505);
xor U2552 (N_2552,N_2503,N_2511);
or U2553 (N_2553,N_2484,N_2479);
nor U2554 (N_2554,N_2482,N_2492);
or U2555 (N_2555,N_2465,N_2482);
nor U2556 (N_2556,N_2477,N_2470);
and U2557 (N_2557,N_2511,N_2501);
nor U2558 (N_2558,N_2509,N_2506);
and U2559 (N_2559,N_2515,N_2519);
nor U2560 (N_2560,N_2515,N_2509);
or U2561 (N_2561,N_2492,N_2504);
nand U2562 (N_2562,N_2482,N_2503);
and U2563 (N_2563,N_2474,N_2502);
xnor U2564 (N_2564,N_2486,N_2470);
nand U2565 (N_2565,N_2517,N_2495);
xnor U2566 (N_2566,N_2506,N_2494);
nand U2567 (N_2567,N_2479,N_2477);
and U2568 (N_2568,N_2503,N_2502);
or U2569 (N_2569,N_2484,N_2519);
xor U2570 (N_2570,N_2462,N_2470);
nand U2571 (N_2571,N_2494,N_2478);
xnor U2572 (N_2572,N_2495,N_2484);
nand U2573 (N_2573,N_2500,N_2513);
xor U2574 (N_2574,N_2491,N_2512);
nor U2575 (N_2575,N_2481,N_2486);
or U2576 (N_2576,N_2490,N_2478);
nor U2577 (N_2577,N_2464,N_2500);
nor U2578 (N_2578,N_2460,N_2515);
nand U2579 (N_2579,N_2491,N_2466);
and U2580 (N_2580,N_2535,N_2547);
and U2581 (N_2581,N_2534,N_2540);
or U2582 (N_2582,N_2541,N_2528);
nor U2583 (N_2583,N_2543,N_2556);
nand U2584 (N_2584,N_2521,N_2529);
nor U2585 (N_2585,N_2539,N_2560);
xor U2586 (N_2586,N_2527,N_2525);
or U2587 (N_2587,N_2526,N_2571);
or U2588 (N_2588,N_2559,N_2533);
xor U2589 (N_2589,N_2537,N_2562);
xnor U2590 (N_2590,N_2548,N_2564);
or U2591 (N_2591,N_2531,N_2553);
or U2592 (N_2592,N_2542,N_2552);
nor U2593 (N_2593,N_2563,N_2549);
xnor U2594 (N_2594,N_2575,N_2523);
and U2595 (N_2595,N_2522,N_2578);
or U2596 (N_2596,N_2530,N_2546);
nor U2597 (N_2597,N_2576,N_2550);
nand U2598 (N_2598,N_2558,N_2579);
nor U2599 (N_2599,N_2566,N_2545);
xor U2600 (N_2600,N_2572,N_2561);
or U2601 (N_2601,N_2524,N_2573);
and U2602 (N_2602,N_2551,N_2536);
and U2603 (N_2603,N_2538,N_2520);
and U2604 (N_2604,N_2570,N_2557);
xnor U2605 (N_2605,N_2568,N_2554);
or U2606 (N_2606,N_2544,N_2567);
or U2607 (N_2607,N_2565,N_2577);
nor U2608 (N_2608,N_2569,N_2555);
or U2609 (N_2609,N_2532,N_2574);
nand U2610 (N_2610,N_2578,N_2527);
xor U2611 (N_2611,N_2566,N_2528);
xnor U2612 (N_2612,N_2549,N_2523);
or U2613 (N_2613,N_2572,N_2527);
xnor U2614 (N_2614,N_2579,N_2532);
nand U2615 (N_2615,N_2549,N_2537);
nand U2616 (N_2616,N_2557,N_2556);
xnor U2617 (N_2617,N_2544,N_2537);
nand U2618 (N_2618,N_2531,N_2533);
nand U2619 (N_2619,N_2521,N_2574);
nor U2620 (N_2620,N_2540,N_2571);
nand U2621 (N_2621,N_2564,N_2532);
xnor U2622 (N_2622,N_2523,N_2551);
xor U2623 (N_2623,N_2539,N_2570);
nor U2624 (N_2624,N_2579,N_2522);
xnor U2625 (N_2625,N_2535,N_2558);
or U2626 (N_2626,N_2523,N_2569);
xnor U2627 (N_2627,N_2529,N_2558);
nor U2628 (N_2628,N_2576,N_2524);
xnor U2629 (N_2629,N_2573,N_2544);
or U2630 (N_2630,N_2566,N_2546);
and U2631 (N_2631,N_2572,N_2533);
xor U2632 (N_2632,N_2553,N_2560);
and U2633 (N_2633,N_2563,N_2569);
nand U2634 (N_2634,N_2558,N_2563);
or U2635 (N_2635,N_2570,N_2524);
nand U2636 (N_2636,N_2551,N_2571);
nand U2637 (N_2637,N_2532,N_2573);
xor U2638 (N_2638,N_2522,N_2577);
and U2639 (N_2639,N_2523,N_2527);
xnor U2640 (N_2640,N_2607,N_2615);
or U2641 (N_2641,N_2604,N_2608);
nand U2642 (N_2642,N_2601,N_2613);
xnor U2643 (N_2643,N_2597,N_2585);
nor U2644 (N_2644,N_2587,N_2583);
nor U2645 (N_2645,N_2639,N_2606);
and U2646 (N_2646,N_2588,N_2632);
xor U2647 (N_2647,N_2610,N_2628);
nor U2648 (N_2648,N_2635,N_2581);
xnor U2649 (N_2649,N_2631,N_2586);
and U2650 (N_2650,N_2638,N_2605);
xnor U2651 (N_2651,N_2584,N_2633);
or U2652 (N_2652,N_2629,N_2617);
nor U2653 (N_2653,N_2598,N_2609);
nor U2654 (N_2654,N_2591,N_2618);
xor U2655 (N_2655,N_2616,N_2634);
nand U2656 (N_2656,N_2612,N_2625);
xnor U2657 (N_2657,N_2630,N_2592);
or U2658 (N_2658,N_2619,N_2582);
xor U2659 (N_2659,N_2602,N_2611);
nand U2660 (N_2660,N_2620,N_2594);
xnor U2661 (N_2661,N_2603,N_2590);
nand U2662 (N_2662,N_2636,N_2600);
nand U2663 (N_2663,N_2621,N_2593);
and U2664 (N_2664,N_2627,N_2637);
nand U2665 (N_2665,N_2580,N_2596);
and U2666 (N_2666,N_2624,N_2589);
nor U2667 (N_2667,N_2626,N_2599);
xnor U2668 (N_2668,N_2623,N_2622);
nand U2669 (N_2669,N_2595,N_2614);
nand U2670 (N_2670,N_2585,N_2624);
or U2671 (N_2671,N_2633,N_2624);
or U2672 (N_2672,N_2638,N_2613);
and U2673 (N_2673,N_2601,N_2623);
nor U2674 (N_2674,N_2592,N_2606);
xnor U2675 (N_2675,N_2602,N_2589);
and U2676 (N_2676,N_2632,N_2612);
or U2677 (N_2677,N_2601,N_2584);
nor U2678 (N_2678,N_2608,N_2595);
nor U2679 (N_2679,N_2633,N_2609);
nor U2680 (N_2680,N_2635,N_2624);
xnor U2681 (N_2681,N_2608,N_2594);
and U2682 (N_2682,N_2639,N_2599);
nor U2683 (N_2683,N_2633,N_2636);
or U2684 (N_2684,N_2583,N_2594);
and U2685 (N_2685,N_2592,N_2638);
xor U2686 (N_2686,N_2615,N_2595);
or U2687 (N_2687,N_2605,N_2618);
and U2688 (N_2688,N_2585,N_2609);
nand U2689 (N_2689,N_2625,N_2596);
or U2690 (N_2690,N_2634,N_2609);
nor U2691 (N_2691,N_2605,N_2606);
nand U2692 (N_2692,N_2611,N_2631);
xnor U2693 (N_2693,N_2606,N_2614);
nand U2694 (N_2694,N_2614,N_2620);
or U2695 (N_2695,N_2587,N_2585);
and U2696 (N_2696,N_2601,N_2585);
and U2697 (N_2697,N_2617,N_2636);
xnor U2698 (N_2698,N_2600,N_2584);
or U2699 (N_2699,N_2622,N_2620);
and U2700 (N_2700,N_2646,N_2667);
or U2701 (N_2701,N_2696,N_2676);
xor U2702 (N_2702,N_2643,N_2660);
or U2703 (N_2703,N_2679,N_2693);
xnor U2704 (N_2704,N_2653,N_2678);
or U2705 (N_2705,N_2692,N_2661);
or U2706 (N_2706,N_2658,N_2684);
xor U2707 (N_2707,N_2657,N_2683);
nand U2708 (N_2708,N_2694,N_2649);
and U2709 (N_2709,N_2647,N_2670);
xor U2710 (N_2710,N_2698,N_2640);
nor U2711 (N_2711,N_2675,N_2677);
xnor U2712 (N_2712,N_2674,N_2672);
and U2713 (N_2713,N_2664,N_2685);
nor U2714 (N_2714,N_2697,N_2689);
xnor U2715 (N_2715,N_2665,N_2662);
nor U2716 (N_2716,N_2682,N_2680);
and U2717 (N_2717,N_2687,N_2656);
and U2718 (N_2718,N_2659,N_2669);
nor U2719 (N_2719,N_2663,N_2668);
or U2720 (N_2720,N_2699,N_2655);
xor U2721 (N_2721,N_2686,N_2688);
nand U2722 (N_2722,N_2666,N_2644);
nand U2723 (N_2723,N_2645,N_2671);
xnor U2724 (N_2724,N_2641,N_2652);
nor U2725 (N_2725,N_2673,N_2650);
xnor U2726 (N_2726,N_2648,N_2651);
nor U2727 (N_2727,N_2691,N_2654);
nand U2728 (N_2728,N_2642,N_2695);
and U2729 (N_2729,N_2690,N_2681);
nor U2730 (N_2730,N_2651,N_2669);
xor U2731 (N_2731,N_2660,N_2645);
nand U2732 (N_2732,N_2670,N_2693);
nor U2733 (N_2733,N_2650,N_2657);
nor U2734 (N_2734,N_2654,N_2645);
or U2735 (N_2735,N_2654,N_2651);
nor U2736 (N_2736,N_2688,N_2643);
and U2737 (N_2737,N_2682,N_2675);
nor U2738 (N_2738,N_2688,N_2654);
xnor U2739 (N_2739,N_2691,N_2668);
nand U2740 (N_2740,N_2687,N_2693);
and U2741 (N_2741,N_2672,N_2661);
xnor U2742 (N_2742,N_2646,N_2692);
nand U2743 (N_2743,N_2665,N_2664);
or U2744 (N_2744,N_2653,N_2669);
and U2745 (N_2745,N_2661,N_2649);
or U2746 (N_2746,N_2678,N_2688);
xnor U2747 (N_2747,N_2688,N_2684);
or U2748 (N_2748,N_2642,N_2684);
nand U2749 (N_2749,N_2691,N_2671);
nor U2750 (N_2750,N_2684,N_2689);
and U2751 (N_2751,N_2659,N_2691);
nand U2752 (N_2752,N_2666,N_2659);
and U2753 (N_2753,N_2668,N_2645);
nand U2754 (N_2754,N_2672,N_2668);
and U2755 (N_2755,N_2662,N_2658);
nor U2756 (N_2756,N_2668,N_2693);
nand U2757 (N_2757,N_2677,N_2685);
nand U2758 (N_2758,N_2697,N_2672);
xnor U2759 (N_2759,N_2685,N_2687);
xor U2760 (N_2760,N_2702,N_2757);
nor U2761 (N_2761,N_2759,N_2758);
or U2762 (N_2762,N_2739,N_2710);
xnor U2763 (N_2763,N_2704,N_2746);
xor U2764 (N_2764,N_2736,N_2705);
or U2765 (N_2765,N_2738,N_2719);
or U2766 (N_2766,N_2714,N_2703);
and U2767 (N_2767,N_2700,N_2755);
nand U2768 (N_2768,N_2753,N_2747);
nand U2769 (N_2769,N_2731,N_2751);
and U2770 (N_2770,N_2722,N_2727);
nor U2771 (N_2771,N_2752,N_2749);
nor U2772 (N_2772,N_2754,N_2708);
nor U2773 (N_2773,N_2706,N_2717);
or U2774 (N_2774,N_2732,N_2756);
nor U2775 (N_2775,N_2715,N_2734);
nor U2776 (N_2776,N_2712,N_2745);
or U2777 (N_2777,N_2716,N_2748);
and U2778 (N_2778,N_2723,N_2711);
nor U2779 (N_2779,N_2726,N_2729);
xnor U2780 (N_2780,N_2721,N_2701);
nor U2781 (N_2781,N_2737,N_2718);
or U2782 (N_2782,N_2735,N_2733);
or U2783 (N_2783,N_2740,N_2724);
or U2784 (N_2784,N_2744,N_2707);
or U2785 (N_2785,N_2720,N_2728);
or U2786 (N_2786,N_2743,N_2725);
xnor U2787 (N_2787,N_2750,N_2713);
and U2788 (N_2788,N_2742,N_2709);
or U2789 (N_2789,N_2741,N_2730);
and U2790 (N_2790,N_2719,N_2740);
xor U2791 (N_2791,N_2726,N_2752);
or U2792 (N_2792,N_2754,N_2747);
nor U2793 (N_2793,N_2755,N_2724);
and U2794 (N_2794,N_2712,N_2717);
nand U2795 (N_2795,N_2741,N_2745);
and U2796 (N_2796,N_2742,N_2731);
nand U2797 (N_2797,N_2704,N_2734);
or U2798 (N_2798,N_2725,N_2709);
nor U2799 (N_2799,N_2713,N_2749);
nor U2800 (N_2800,N_2753,N_2727);
nor U2801 (N_2801,N_2758,N_2730);
nor U2802 (N_2802,N_2752,N_2751);
xnor U2803 (N_2803,N_2751,N_2720);
or U2804 (N_2804,N_2708,N_2726);
xor U2805 (N_2805,N_2712,N_2749);
nand U2806 (N_2806,N_2708,N_2723);
xor U2807 (N_2807,N_2708,N_2725);
and U2808 (N_2808,N_2719,N_2710);
nor U2809 (N_2809,N_2758,N_2733);
xor U2810 (N_2810,N_2700,N_2729);
and U2811 (N_2811,N_2759,N_2757);
nor U2812 (N_2812,N_2759,N_2752);
xor U2813 (N_2813,N_2728,N_2712);
nor U2814 (N_2814,N_2706,N_2718);
nor U2815 (N_2815,N_2730,N_2712);
nand U2816 (N_2816,N_2734,N_2749);
and U2817 (N_2817,N_2720,N_2758);
nor U2818 (N_2818,N_2729,N_2754);
nand U2819 (N_2819,N_2704,N_2725);
and U2820 (N_2820,N_2817,N_2774);
and U2821 (N_2821,N_2772,N_2783);
nand U2822 (N_2822,N_2761,N_2788);
nand U2823 (N_2823,N_2775,N_2765);
and U2824 (N_2824,N_2789,N_2810);
nand U2825 (N_2825,N_2787,N_2807);
and U2826 (N_2826,N_2764,N_2791);
nand U2827 (N_2827,N_2805,N_2762);
xnor U2828 (N_2828,N_2806,N_2763);
and U2829 (N_2829,N_2792,N_2814);
xor U2830 (N_2830,N_2813,N_2816);
nand U2831 (N_2831,N_2785,N_2794);
nor U2832 (N_2832,N_2767,N_2782);
xnor U2833 (N_2833,N_2804,N_2780);
or U2834 (N_2834,N_2786,N_2790);
xnor U2835 (N_2835,N_2798,N_2769);
or U2836 (N_2836,N_2803,N_2815);
and U2837 (N_2837,N_2771,N_2796);
nand U2838 (N_2838,N_2760,N_2781);
and U2839 (N_2839,N_2808,N_2779);
and U2840 (N_2840,N_2818,N_2784);
nand U2841 (N_2841,N_2802,N_2795);
or U2842 (N_2842,N_2778,N_2819);
nor U2843 (N_2843,N_2776,N_2777);
or U2844 (N_2844,N_2768,N_2801);
nand U2845 (N_2845,N_2770,N_2811);
xor U2846 (N_2846,N_2812,N_2809);
and U2847 (N_2847,N_2793,N_2797);
nor U2848 (N_2848,N_2799,N_2800);
nor U2849 (N_2849,N_2773,N_2766);
nor U2850 (N_2850,N_2760,N_2810);
nand U2851 (N_2851,N_2783,N_2801);
or U2852 (N_2852,N_2799,N_2809);
or U2853 (N_2853,N_2804,N_2811);
and U2854 (N_2854,N_2778,N_2786);
xnor U2855 (N_2855,N_2774,N_2810);
or U2856 (N_2856,N_2763,N_2815);
and U2857 (N_2857,N_2807,N_2766);
and U2858 (N_2858,N_2770,N_2819);
nand U2859 (N_2859,N_2810,N_2786);
and U2860 (N_2860,N_2816,N_2794);
and U2861 (N_2861,N_2778,N_2782);
xor U2862 (N_2862,N_2768,N_2762);
nor U2863 (N_2863,N_2772,N_2811);
nand U2864 (N_2864,N_2796,N_2789);
or U2865 (N_2865,N_2781,N_2818);
nand U2866 (N_2866,N_2800,N_2775);
xnor U2867 (N_2867,N_2765,N_2814);
nand U2868 (N_2868,N_2794,N_2815);
or U2869 (N_2869,N_2798,N_2776);
and U2870 (N_2870,N_2804,N_2776);
and U2871 (N_2871,N_2799,N_2768);
nand U2872 (N_2872,N_2760,N_2818);
and U2873 (N_2873,N_2766,N_2782);
xnor U2874 (N_2874,N_2784,N_2769);
xor U2875 (N_2875,N_2818,N_2772);
nand U2876 (N_2876,N_2796,N_2817);
xor U2877 (N_2877,N_2777,N_2771);
nor U2878 (N_2878,N_2815,N_2788);
and U2879 (N_2879,N_2806,N_2775);
nor U2880 (N_2880,N_2879,N_2833);
nand U2881 (N_2881,N_2823,N_2834);
and U2882 (N_2882,N_2855,N_2868);
xnor U2883 (N_2883,N_2842,N_2852);
nor U2884 (N_2884,N_2847,N_2874);
xor U2885 (N_2885,N_2858,N_2837);
nor U2886 (N_2886,N_2829,N_2867);
nor U2887 (N_2887,N_2865,N_2835);
or U2888 (N_2888,N_2878,N_2846);
xnor U2889 (N_2889,N_2827,N_2822);
and U2890 (N_2890,N_2843,N_2832);
xor U2891 (N_2891,N_2838,N_2824);
nand U2892 (N_2892,N_2826,N_2856);
xor U2893 (N_2893,N_2875,N_2866);
xnor U2894 (N_2894,N_2828,N_2839);
xor U2895 (N_2895,N_2825,N_2872);
nor U2896 (N_2896,N_2851,N_2850);
and U2897 (N_2897,N_2848,N_2821);
nor U2898 (N_2898,N_2863,N_2831);
xnor U2899 (N_2899,N_2830,N_2877);
xor U2900 (N_2900,N_2845,N_2844);
nor U2901 (N_2901,N_2864,N_2861);
or U2902 (N_2902,N_2840,N_2857);
xor U2903 (N_2903,N_2871,N_2870);
and U2904 (N_2904,N_2836,N_2841);
nor U2905 (N_2905,N_2869,N_2876);
xor U2906 (N_2906,N_2862,N_2860);
nand U2907 (N_2907,N_2849,N_2873);
or U2908 (N_2908,N_2859,N_2853);
nand U2909 (N_2909,N_2854,N_2820);
and U2910 (N_2910,N_2879,N_2867);
and U2911 (N_2911,N_2831,N_2854);
nor U2912 (N_2912,N_2868,N_2874);
xnor U2913 (N_2913,N_2829,N_2872);
xor U2914 (N_2914,N_2859,N_2851);
and U2915 (N_2915,N_2870,N_2859);
nand U2916 (N_2916,N_2876,N_2870);
xnor U2917 (N_2917,N_2872,N_2838);
xnor U2918 (N_2918,N_2828,N_2851);
xor U2919 (N_2919,N_2843,N_2865);
and U2920 (N_2920,N_2866,N_2871);
xor U2921 (N_2921,N_2847,N_2863);
xor U2922 (N_2922,N_2850,N_2823);
nor U2923 (N_2923,N_2863,N_2861);
xnor U2924 (N_2924,N_2877,N_2872);
nor U2925 (N_2925,N_2867,N_2866);
or U2926 (N_2926,N_2875,N_2827);
nand U2927 (N_2927,N_2827,N_2834);
and U2928 (N_2928,N_2871,N_2878);
or U2929 (N_2929,N_2852,N_2878);
nor U2930 (N_2930,N_2877,N_2854);
nand U2931 (N_2931,N_2847,N_2869);
and U2932 (N_2932,N_2876,N_2877);
nand U2933 (N_2933,N_2850,N_2843);
and U2934 (N_2934,N_2835,N_2830);
or U2935 (N_2935,N_2847,N_2864);
or U2936 (N_2936,N_2877,N_2860);
xor U2937 (N_2937,N_2874,N_2845);
and U2938 (N_2938,N_2860,N_2879);
xnor U2939 (N_2939,N_2863,N_2850);
xor U2940 (N_2940,N_2896,N_2893);
nor U2941 (N_2941,N_2925,N_2928);
nand U2942 (N_2942,N_2880,N_2913);
nor U2943 (N_2943,N_2919,N_2926);
and U2944 (N_2944,N_2900,N_2901);
nor U2945 (N_2945,N_2921,N_2936);
and U2946 (N_2946,N_2897,N_2932);
nand U2947 (N_2947,N_2912,N_2917);
or U2948 (N_2948,N_2908,N_2891);
and U2949 (N_2949,N_2914,N_2882);
xnor U2950 (N_2950,N_2937,N_2927);
xor U2951 (N_2951,N_2920,N_2884);
or U2952 (N_2952,N_2933,N_2885);
nand U2953 (N_2953,N_2910,N_2907);
nand U2954 (N_2954,N_2887,N_2918);
nor U2955 (N_2955,N_2899,N_2930);
xnor U2956 (N_2956,N_2892,N_2924);
xnor U2957 (N_2957,N_2931,N_2886);
or U2958 (N_2958,N_2894,N_2923);
or U2959 (N_2959,N_2909,N_2889);
nand U2960 (N_2960,N_2929,N_2938);
nor U2961 (N_2961,N_2890,N_2902);
and U2962 (N_2962,N_2905,N_2935);
and U2963 (N_2963,N_2904,N_2915);
nor U2964 (N_2964,N_2895,N_2922);
nand U2965 (N_2965,N_2888,N_2916);
nand U2966 (N_2966,N_2939,N_2903);
xnor U2967 (N_2967,N_2906,N_2911);
xnor U2968 (N_2968,N_2883,N_2898);
and U2969 (N_2969,N_2934,N_2881);
nand U2970 (N_2970,N_2913,N_2885);
or U2971 (N_2971,N_2911,N_2890);
xnor U2972 (N_2972,N_2910,N_2896);
xnor U2973 (N_2973,N_2916,N_2937);
nor U2974 (N_2974,N_2896,N_2916);
and U2975 (N_2975,N_2896,N_2928);
and U2976 (N_2976,N_2930,N_2918);
xor U2977 (N_2977,N_2891,N_2907);
and U2978 (N_2978,N_2914,N_2930);
or U2979 (N_2979,N_2897,N_2896);
nor U2980 (N_2980,N_2893,N_2905);
or U2981 (N_2981,N_2921,N_2922);
xnor U2982 (N_2982,N_2907,N_2900);
xnor U2983 (N_2983,N_2911,N_2910);
and U2984 (N_2984,N_2908,N_2904);
xor U2985 (N_2985,N_2910,N_2887);
xor U2986 (N_2986,N_2921,N_2894);
or U2987 (N_2987,N_2918,N_2907);
or U2988 (N_2988,N_2931,N_2922);
nor U2989 (N_2989,N_2889,N_2933);
or U2990 (N_2990,N_2928,N_2921);
xnor U2991 (N_2991,N_2906,N_2907);
and U2992 (N_2992,N_2891,N_2917);
and U2993 (N_2993,N_2887,N_2899);
xnor U2994 (N_2994,N_2909,N_2918);
nor U2995 (N_2995,N_2885,N_2897);
nor U2996 (N_2996,N_2934,N_2907);
nand U2997 (N_2997,N_2884,N_2895);
xnor U2998 (N_2998,N_2888,N_2899);
or U2999 (N_2999,N_2883,N_2904);
or UO_0 (O_0,N_2984,N_2967);
and UO_1 (O_1,N_2998,N_2941);
and UO_2 (O_2,N_2988,N_2976);
and UO_3 (O_3,N_2954,N_2983);
xor UO_4 (O_4,N_2965,N_2971);
nor UO_5 (O_5,N_2968,N_2962);
and UO_6 (O_6,N_2959,N_2989);
nand UO_7 (O_7,N_2985,N_2973);
nand UO_8 (O_8,N_2981,N_2940);
and UO_9 (O_9,N_2969,N_2995);
nor UO_10 (O_10,N_2999,N_2992);
and UO_11 (O_11,N_2980,N_2996);
nor UO_12 (O_12,N_2960,N_2972);
or UO_13 (O_13,N_2957,N_2944);
xnor UO_14 (O_14,N_2970,N_2952);
and UO_15 (O_15,N_2982,N_2955);
and UO_16 (O_16,N_2994,N_2943);
or UO_17 (O_17,N_2978,N_2986);
and UO_18 (O_18,N_2950,N_2964);
xnor UO_19 (O_19,N_2979,N_2958);
or UO_20 (O_20,N_2949,N_2974);
nor UO_21 (O_21,N_2993,N_2953);
nand UO_22 (O_22,N_2956,N_2990);
and UO_23 (O_23,N_2946,N_2977);
nand UO_24 (O_24,N_2997,N_2951);
and UO_25 (O_25,N_2966,N_2948);
and UO_26 (O_26,N_2963,N_2987);
or UO_27 (O_27,N_2961,N_2947);
nor UO_28 (O_28,N_2991,N_2945);
or UO_29 (O_29,N_2975,N_2942);
xnor UO_30 (O_30,N_2984,N_2978);
and UO_31 (O_31,N_2984,N_2980);
xor UO_32 (O_32,N_2991,N_2970);
xnor UO_33 (O_33,N_2993,N_2988);
or UO_34 (O_34,N_2976,N_2954);
nor UO_35 (O_35,N_2965,N_2951);
xnor UO_36 (O_36,N_2953,N_2948);
and UO_37 (O_37,N_2988,N_2991);
nand UO_38 (O_38,N_2968,N_2957);
or UO_39 (O_39,N_2978,N_2962);
and UO_40 (O_40,N_2980,N_2995);
or UO_41 (O_41,N_2993,N_2974);
nor UO_42 (O_42,N_2965,N_2960);
nor UO_43 (O_43,N_2950,N_2987);
and UO_44 (O_44,N_2954,N_2979);
and UO_45 (O_45,N_2953,N_2947);
nor UO_46 (O_46,N_2974,N_2997);
nand UO_47 (O_47,N_2955,N_2945);
nand UO_48 (O_48,N_2950,N_2955);
xnor UO_49 (O_49,N_2945,N_2944);
nor UO_50 (O_50,N_2997,N_2944);
xor UO_51 (O_51,N_2974,N_2945);
or UO_52 (O_52,N_2997,N_2968);
or UO_53 (O_53,N_2957,N_2943);
nor UO_54 (O_54,N_2977,N_2966);
xnor UO_55 (O_55,N_2958,N_2957);
nor UO_56 (O_56,N_2975,N_2948);
xnor UO_57 (O_57,N_2961,N_2970);
xnor UO_58 (O_58,N_2980,N_2949);
nor UO_59 (O_59,N_2953,N_2978);
and UO_60 (O_60,N_2959,N_2977);
nand UO_61 (O_61,N_2964,N_2974);
xnor UO_62 (O_62,N_2978,N_2973);
and UO_63 (O_63,N_2952,N_2961);
or UO_64 (O_64,N_2985,N_2955);
xnor UO_65 (O_65,N_2946,N_2955);
nor UO_66 (O_66,N_2967,N_2982);
nor UO_67 (O_67,N_2975,N_2940);
and UO_68 (O_68,N_2997,N_2971);
or UO_69 (O_69,N_2943,N_2940);
nand UO_70 (O_70,N_2996,N_2977);
or UO_71 (O_71,N_2944,N_2999);
nor UO_72 (O_72,N_2944,N_2965);
and UO_73 (O_73,N_2940,N_2942);
and UO_74 (O_74,N_2996,N_2987);
nor UO_75 (O_75,N_2977,N_2972);
or UO_76 (O_76,N_2963,N_2979);
and UO_77 (O_77,N_2971,N_2943);
and UO_78 (O_78,N_2985,N_2950);
nand UO_79 (O_79,N_2952,N_2968);
nor UO_80 (O_80,N_2988,N_2985);
nor UO_81 (O_81,N_2973,N_2946);
and UO_82 (O_82,N_2943,N_2978);
and UO_83 (O_83,N_2945,N_2949);
nor UO_84 (O_84,N_2966,N_2960);
or UO_85 (O_85,N_2940,N_2985);
or UO_86 (O_86,N_2991,N_2980);
or UO_87 (O_87,N_2993,N_2979);
or UO_88 (O_88,N_2967,N_2992);
or UO_89 (O_89,N_2961,N_2998);
nand UO_90 (O_90,N_2975,N_2950);
nor UO_91 (O_91,N_2942,N_2961);
nand UO_92 (O_92,N_2993,N_2984);
or UO_93 (O_93,N_2983,N_2942);
nor UO_94 (O_94,N_2980,N_2971);
xor UO_95 (O_95,N_2963,N_2998);
nor UO_96 (O_96,N_2971,N_2967);
nor UO_97 (O_97,N_2950,N_2971);
and UO_98 (O_98,N_2967,N_2997);
or UO_99 (O_99,N_2962,N_2982);
or UO_100 (O_100,N_2995,N_2972);
and UO_101 (O_101,N_2949,N_2964);
and UO_102 (O_102,N_2947,N_2943);
xnor UO_103 (O_103,N_2980,N_2988);
nand UO_104 (O_104,N_2962,N_2991);
or UO_105 (O_105,N_2988,N_2961);
nand UO_106 (O_106,N_2960,N_2951);
nor UO_107 (O_107,N_2961,N_2968);
nor UO_108 (O_108,N_2982,N_2957);
and UO_109 (O_109,N_2976,N_2992);
nor UO_110 (O_110,N_2991,N_2954);
or UO_111 (O_111,N_2948,N_2974);
xnor UO_112 (O_112,N_2974,N_2940);
nor UO_113 (O_113,N_2981,N_2990);
or UO_114 (O_114,N_2966,N_2964);
nor UO_115 (O_115,N_2949,N_2965);
and UO_116 (O_116,N_2985,N_2945);
xnor UO_117 (O_117,N_2988,N_2972);
nand UO_118 (O_118,N_2983,N_2970);
nand UO_119 (O_119,N_2997,N_2987);
or UO_120 (O_120,N_2964,N_2985);
nor UO_121 (O_121,N_2960,N_2992);
xor UO_122 (O_122,N_2964,N_2972);
xnor UO_123 (O_123,N_2984,N_2954);
and UO_124 (O_124,N_2969,N_2970);
nand UO_125 (O_125,N_2983,N_2969);
nor UO_126 (O_126,N_2968,N_2967);
xor UO_127 (O_127,N_2979,N_2988);
xor UO_128 (O_128,N_2969,N_2942);
nand UO_129 (O_129,N_2969,N_2941);
nor UO_130 (O_130,N_2983,N_2975);
xnor UO_131 (O_131,N_2998,N_2992);
xnor UO_132 (O_132,N_2953,N_2941);
nor UO_133 (O_133,N_2947,N_2999);
or UO_134 (O_134,N_2995,N_2975);
or UO_135 (O_135,N_2975,N_2966);
and UO_136 (O_136,N_2967,N_2983);
and UO_137 (O_137,N_2944,N_2985);
nand UO_138 (O_138,N_2947,N_2956);
or UO_139 (O_139,N_2940,N_2995);
xnor UO_140 (O_140,N_2959,N_2946);
nand UO_141 (O_141,N_2975,N_2955);
nor UO_142 (O_142,N_2957,N_2980);
xor UO_143 (O_143,N_2973,N_2963);
or UO_144 (O_144,N_2965,N_2988);
nor UO_145 (O_145,N_2961,N_2976);
nand UO_146 (O_146,N_2940,N_2993);
and UO_147 (O_147,N_2942,N_2974);
xor UO_148 (O_148,N_2952,N_2949);
nand UO_149 (O_149,N_2948,N_2971);
nand UO_150 (O_150,N_2999,N_2955);
xnor UO_151 (O_151,N_2999,N_2950);
xnor UO_152 (O_152,N_2978,N_2980);
and UO_153 (O_153,N_2989,N_2977);
or UO_154 (O_154,N_2970,N_2948);
or UO_155 (O_155,N_2995,N_2968);
nor UO_156 (O_156,N_2963,N_2967);
and UO_157 (O_157,N_2948,N_2957);
or UO_158 (O_158,N_2965,N_2957);
or UO_159 (O_159,N_2957,N_2955);
or UO_160 (O_160,N_2969,N_2963);
or UO_161 (O_161,N_2970,N_2973);
and UO_162 (O_162,N_2961,N_2948);
nor UO_163 (O_163,N_2994,N_2983);
nor UO_164 (O_164,N_2945,N_2984);
nor UO_165 (O_165,N_2979,N_2967);
or UO_166 (O_166,N_2941,N_2972);
and UO_167 (O_167,N_2963,N_2982);
and UO_168 (O_168,N_2967,N_2952);
xnor UO_169 (O_169,N_2978,N_2966);
nor UO_170 (O_170,N_2947,N_2981);
or UO_171 (O_171,N_2980,N_2946);
and UO_172 (O_172,N_2940,N_2984);
xor UO_173 (O_173,N_2999,N_2941);
nand UO_174 (O_174,N_2941,N_2942);
nand UO_175 (O_175,N_2953,N_2976);
nand UO_176 (O_176,N_2961,N_2946);
or UO_177 (O_177,N_2967,N_2976);
nand UO_178 (O_178,N_2947,N_2959);
or UO_179 (O_179,N_2987,N_2940);
nand UO_180 (O_180,N_2956,N_2961);
or UO_181 (O_181,N_2959,N_2985);
nor UO_182 (O_182,N_2997,N_2945);
or UO_183 (O_183,N_2948,N_2996);
and UO_184 (O_184,N_2992,N_2968);
nand UO_185 (O_185,N_2976,N_2964);
and UO_186 (O_186,N_2970,N_2967);
nor UO_187 (O_187,N_2976,N_2969);
and UO_188 (O_188,N_2971,N_2963);
nor UO_189 (O_189,N_2977,N_2958);
or UO_190 (O_190,N_2991,N_2957);
nor UO_191 (O_191,N_2955,N_2952);
xnor UO_192 (O_192,N_2957,N_2997);
or UO_193 (O_193,N_2988,N_2959);
or UO_194 (O_194,N_2976,N_2946);
nand UO_195 (O_195,N_2972,N_2954);
or UO_196 (O_196,N_2942,N_2965);
nor UO_197 (O_197,N_2965,N_2954);
and UO_198 (O_198,N_2985,N_2953);
nor UO_199 (O_199,N_2971,N_2969);
nand UO_200 (O_200,N_2959,N_2994);
xnor UO_201 (O_201,N_2967,N_2961);
nor UO_202 (O_202,N_2977,N_2943);
nand UO_203 (O_203,N_2970,N_2954);
xor UO_204 (O_204,N_2993,N_2976);
xor UO_205 (O_205,N_2982,N_2975);
and UO_206 (O_206,N_2948,N_2993);
xnor UO_207 (O_207,N_2998,N_2974);
nand UO_208 (O_208,N_2953,N_2954);
nor UO_209 (O_209,N_2956,N_2960);
nor UO_210 (O_210,N_2940,N_2956);
and UO_211 (O_211,N_2953,N_2973);
and UO_212 (O_212,N_2993,N_2985);
and UO_213 (O_213,N_2989,N_2995);
and UO_214 (O_214,N_2940,N_2953);
xor UO_215 (O_215,N_2998,N_2970);
and UO_216 (O_216,N_2974,N_2954);
nand UO_217 (O_217,N_2942,N_2979);
xor UO_218 (O_218,N_2941,N_2943);
and UO_219 (O_219,N_2981,N_2964);
nor UO_220 (O_220,N_2977,N_2944);
xor UO_221 (O_221,N_2979,N_2986);
and UO_222 (O_222,N_2949,N_2971);
xnor UO_223 (O_223,N_2992,N_2985);
and UO_224 (O_224,N_2951,N_2981);
nor UO_225 (O_225,N_2948,N_2977);
and UO_226 (O_226,N_2990,N_2964);
and UO_227 (O_227,N_2960,N_2997);
nand UO_228 (O_228,N_2997,N_2981);
and UO_229 (O_229,N_2981,N_2985);
and UO_230 (O_230,N_2957,N_2956);
xnor UO_231 (O_231,N_2948,N_2960);
nor UO_232 (O_232,N_2994,N_2999);
nor UO_233 (O_233,N_2964,N_2948);
nand UO_234 (O_234,N_2951,N_2999);
nor UO_235 (O_235,N_2962,N_2997);
or UO_236 (O_236,N_2974,N_2967);
and UO_237 (O_237,N_2986,N_2942);
or UO_238 (O_238,N_2956,N_2997);
or UO_239 (O_239,N_2943,N_2946);
nor UO_240 (O_240,N_2975,N_2976);
nand UO_241 (O_241,N_2947,N_2998);
nand UO_242 (O_242,N_2944,N_2962);
and UO_243 (O_243,N_2975,N_2952);
and UO_244 (O_244,N_2973,N_2980);
xor UO_245 (O_245,N_2998,N_2956);
and UO_246 (O_246,N_2959,N_2982);
and UO_247 (O_247,N_2954,N_2973);
and UO_248 (O_248,N_2972,N_2962);
nor UO_249 (O_249,N_2963,N_2943);
nor UO_250 (O_250,N_2953,N_2945);
nand UO_251 (O_251,N_2961,N_2994);
nor UO_252 (O_252,N_2947,N_2978);
nand UO_253 (O_253,N_2951,N_2947);
or UO_254 (O_254,N_2962,N_2965);
nand UO_255 (O_255,N_2962,N_2966);
or UO_256 (O_256,N_2981,N_2952);
or UO_257 (O_257,N_2989,N_2955);
nand UO_258 (O_258,N_2949,N_2970);
xor UO_259 (O_259,N_2942,N_2992);
xnor UO_260 (O_260,N_2949,N_2986);
or UO_261 (O_261,N_2960,N_2976);
nand UO_262 (O_262,N_2966,N_2957);
nor UO_263 (O_263,N_2996,N_2974);
nand UO_264 (O_264,N_2985,N_2963);
or UO_265 (O_265,N_2963,N_2962);
xor UO_266 (O_266,N_2973,N_2969);
or UO_267 (O_267,N_2986,N_2992);
xor UO_268 (O_268,N_2963,N_2978);
nor UO_269 (O_269,N_2953,N_2966);
xor UO_270 (O_270,N_2964,N_2944);
or UO_271 (O_271,N_2964,N_2965);
nand UO_272 (O_272,N_2992,N_2952);
or UO_273 (O_273,N_2983,N_2966);
and UO_274 (O_274,N_2977,N_2960);
or UO_275 (O_275,N_2995,N_2999);
nand UO_276 (O_276,N_2977,N_2945);
and UO_277 (O_277,N_2943,N_2967);
nand UO_278 (O_278,N_2986,N_2973);
nor UO_279 (O_279,N_2956,N_2954);
xor UO_280 (O_280,N_2987,N_2967);
nor UO_281 (O_281,N_2970,N_2987);
nor UO_282 (O_282,N_2956,N_2995);
xnor UO_283 (O_283,N_2972,N_2982);
nand UO_284 (O_284,N_2951,N_2969);
xor UO_285 (O_285,N_2984,N_2994);
or UO_286 (O_286,N_2944,N_2971);
nand UO_287 (O_287,N_2997,N_2946);
xnor UO_288 (O_288,N_2965,N_2994);
and UO_289 (O_289,N_2993,N_2978);
and UO_290 (O_290,N_2987,N_2978);
nor UO_291 (O_291,N_2967,N_2996);
or UO_292 (O_292,N_2978,N_2985);
nor UO_293 (O_293,N_2945,N_2951);
nor UO_294 (O_294,N_2947,N_2989);
nor UO_295 (O_295,N_2947,N_2941);
nand UO_296 (O_296,N_2963,N_2974);
xnor UO_297 (O_297,N_2982,N_2964);
nand UO_298 (O_298,N_2987,N_2956);
or UO_299 (O_299,N_2940,N_2963);
nand UO_300 (O_300,N_2987,N_2966);
or UO_301 (O_301,N_2961,N_2951);
or UO_302 (O_302,N_2977,N_2978);
nor UO_303 (O_303,N_2960,N_2987);
nor UO_304 (O_304,N_2969,N_2999);
nor UO_305 (O_305,N_2948,N_2951);
and UO_306 (O_306,N_2979,N_2972);
nor UO_307 (O_307,N_2998,N_2975);
nand UO_308 (O_308,N_2973,N_2991);
nor UO_309 (O_309,N_2999,N_2984);
and UO_310 (O_310,N_2981,N_2958);
xor UO_311 (O_311,N_2954,N_2942);
xnor UO_312 (O_312,N_2989,N_2979);
and UO_313 (O_313,N_2961,N_2943);
nor UO_314 (O_314,N_2987,N_2991);
nand UO_315 (O_315,N_2970,N_2941);
and UO_316 (O_316,N_2954,N_2962);
nor UO_317 (O_317,N_2963,N_2948);
xor UO_318 (O_318,N_2990,N_2945);
and UO_319 (O_319,N_2993,N_2987);
xnor UO_320 (O_320,N_2957,N_2962);
nand UO_321 (O_321,N_2958,N_2996);
nor UO_322 (O_322,N_2968,N_2941);
xor UO_323 (O_323,N_2969,N_2950);
and UO_324 (O_324,N_2974,N_2991);
nor UO_325 (O_325,N_2960,N_2994);
xor UO_326 (O_326,N_2997,N_2972);
xnor UO_327 (O_327,N_2989,N_2968);
xor UO_328 (O_328,N_2976,N_2958);
nor UO_329 (O_329,N_2954,N_2944);
and UO_330 (O_330,N_2969,N_2994);
and UO_331 (O_331,N_2941,N_2960);
nor UO_332 (O_332,N_2984,N_2968);
nand UO_333 (O_333,N_2992,N_2948);
and UO_334 (O_334,N_2987,N_2959);
and UO_335 (O_335,N_2992,N_2979);
or UO_336 (O_336,N_2982,N_2995);
nor UO_337 (O_337,N_2952,N_2980);
nand UO_338 (O_338,N_2968,N_2973);
nand UO_339 (O_339,N_2962,N_2974);
xor UO_340 (O_340,N_2983,N_2986);
nand UO_341 (O_341,N_2970,N_2974);
or UO_342 (O_342,N_2981,N_2996);
xor UO_343 (O_343,N_2962,N_2988);
nand UO_344 (O_344,N_2941,N_2955);
nor UO_345 (O_345,N_2957,N_2963);
nand UO_346 (O_346,N_2964,N_2998);
or UO_347 (O_347,N_2978,N_2968);
and UO_348 (O_348,N_2975,N_2951);
nor UO_349 (O_349,N_2986,N_2943);
xnor UO_350 (O_350,N_2984,N_2964);
and UO_351 (O_351,N_2986,N_2984);
or UO_352 (O_352,N_2978,N_2988);
or UO_353 (O_353,N_2966,N_2970);
or UO_354 (O_354,N_2962,N_2977);
or UO_355 (O_355,N_2944,N_2968);
or UO_356 (O_356,N_2991,N_2946);
or UO_357 (O_357,N_2973,N_2966);
nand UO_358 (O_358,N_2962,N_2985);
or UO_359 (O_359,N_2987,N_2944);
or UO_360 (O_360,N_2975,N_2991);
and UO_361 (O_361,N_2999,N_2993);
or UO_362 (O_362,N_2980,N_2940);
or UO_363 (O_363,N_2978,N_2961);
nor UO_364 (O_364,N_2970,N_2976);
or UO_365 (O_365,N_2986,N_2959);
and UO_366 (O_366,N_2945,N_2970);
nand UO_367 (O_367,N_2978,N_2972);
nand UO_368 (O_368,N_2947,N_2993);
xnor UO_369 (O_369,N_2974,N_2961);
xor UO_370 (O_370,N_2965,N_2993);
nor UO_371 (O_371,N_2949,N_2989);
and UO_372 (O_372,N_2980,N_2993);
and UO_373 (O_373,N_2964,N_2988);
xnor UO_374 (O_374,N_2970,N_2965);
nand UO_375 (O_375,N_2951,N_2955);
nor UO_376 (O_376,N_2974,N_2969);
and UO_377 (O_377,N_2990,N_2940);
and UO_378 (O_378,N_2996,N_2976);
nor UO_379 (O_379,N_2978,N_2974);
nand UO_380 (O_380,N_2989,N_2944);
nor UO_381 (O_381,N_2995,N_2962);
and UO_382 (O_382,N_2958,N_2993);
xnor UO_383 (O_383,N_2973,N_2984);
nor UO_384 (O_384,N_2956,N_2943);
and UO_385 (O_385,N_2987,N_2957);
nand UO_386 (O_386,N_2980,N_2950);
nor UO_387 (O_387,N_2974,N_2977);
or UO_388 (O_388,N_2954,N_2990);
nand UO_389 (O_389,N_2958,N_2988);
or UO_390 (O_390,N_2977,N_2942);
or UO_391 (O_391,N_2950,N_2953);
and UO_392 (O_392,N_2949,N_2944);
nor UO_393 (O_393,N_2968,N_2949);
or UO_394 (O_394,N_2995,N_2974);
xnor UO_395 (O_395,N_2959,N_2990);
nor UO_396 (O_396,N_2950,N_2993);
nor UO_397 (O_397,N_2954,N_2977);
nor UO_398 (O_398,N_2973,N_2982);
xor UO_399 (O_399,N_2976,N_2973);
xnor UO_400 (O_400,N_2955,N_2944);
nor UO_401 (O_401,N_2974,N_2989);
nor UO_402 (O_402,N_2969,N_2975);
or UO_403 (O_403,N_2942,N_2997);
and UO_404 (O_404,N_2957,N_2994);
nand UO_405 (O_405,N_2995,N_2943);
or UO_406 (O_406,N_2963,N_2966);
xor UO_407 (O_407,N_2951,N_2976);
nand UO_408 (O_408,N_2978,N_2971);
xnor UO_409 (O_409,N_2950,N_2952);
nor UO_410 (O_410,N_2973,N_2959);
nand UO_411 (O_411,N_2949,N_2983);
or UO_412 (O_412,N_2956,N_2963);
xor UO_413 (O_413,N_2999,N_2960);
nor UO_414 (O_414,N_2989,N_2991);
xor UO_415 (O_415,N_2946,N_2953);
nand UO_416 (O_416,N_2948,N_2952);
or UO_417 (O_417,N_2943,N_2982);
nor UO_418 (O_418,N_2965,N_2940);
nand UO_419 (O_419,N_2978,N_2995);
or UO_420 (O_420,N_2998,N_2944);
and UO_421 (O_421,N_2993,N_2986);
xor UO_422 (O_422,N_2985,N_2990);
or UO_423 (O_423,N_2941,N_2944);
xnor UO_424 (O_424,N_2977,N_2971);
or UO_425 (O_425,N_2948,N_2981);
nor UO_426 (O_426,N_2967,N_2969);
and UO_427 (O_427,N_2964,N_2978);
nand UO_428 (O_428,N_2999,N_2942);
nand UO_429 (O_429,N_2981,N_2965);
nor UO_430 (O_430,N_2992,N_2940);
or UO_431 (O_431,N_2976,N_2942);
xnor UO_432 (O_432,N_2986,N_2963);
nor UO_433 (O_433,N_2969,N_2962);
or UO_434 (O_434,N_2952,N_2997);
nor UO_435 (O_435,N_2980,N_2986);
xnor UO_436 (O_436,N_2966,N_2996);
and UO_437 (O_437,N_2973,N_2955);
nand UO_438 (O_438,N_2966,N_2993);
nor UO_439 (O_439,N_2963,N_2999);
and UO_440 (O_440,N_2997,N_2964);
or UO_441 (O_441,N_2996,N_2986);
xor UO_442 (O_442,N_2982,N_2991);
nand UO_443 (O_443,N_2958,N_2944);
xor UO_444 (O_444,N_2943,N_2964);
xor UO_445 (O_445,N_2949,N_2976);
nor UO_446 (O_446,N_2961,N_2950);
and UO_447 (O_447,N_2954,N_2949);
nor UO_448 (O_448,N_2961,N_2940);
xor UO_449 (O_449,N_2992,N_2951);
and UO_450 (O_450,N_2981,N_2968);
or UO_451 (O_451,N_2963,N_2981);
xor UO_452 (O_452,N_2948,N_2989);
xor UO_453 (O_453,N_2995,N_2966);
nand UO_454 (O_454,N_2945,N_2967);
xor UO_455 (O_455,N_2949,N_2956);
xnor UO_456 (O_456,N_2982,N_2965);
or UO_457 (O_457,N_2980,N_2945);
nand UO_458 (O_458,N_2963,N_2949);
nand UO_459 (O_459,N_2954,N_2997);
nor UO_460 (O_460,N_2948,N_2973);
and UO_461 (O_461,N_2949,N_2977);
nor UO_462 (O_462,N_2942,N_2962);
xor UO_463 (O_463,N_2940,N_2947);
or UO_464 (O_464,N_2999,N_2973);
nand UO_465 (O_465,N_2984,N_2957);
nor UO_466 (O_466,N_2940,N_2950);
or UO_467 (O_467,N_2945,N_2978);
nor UO_468 (O_468,N_2962,N_2994);
nor UO_469 (O_469,N_2944,N_2960);
or UO_470 (O_470,N_2994,N_2942);
and UO_471 (O_471,N_2944,N_2983);
xnor UO_472 (O_472,N_2973,N_2994);
or UO_473 (O_473,N_2966,N_2979);
and UO_474 (O_474,N_2997,N_2940);
or UO_475 (O_475,N_2989,N_2990);
and UO_476 (O_476,N_2969,N_2948);
xor UO_477 (O_477,N_2984,N_2966);
or UO_478 (O_478,N_2957,N_2951);
or UO_479 (O_479,N_2964,N_2961);
xor UO_480 (O_480,N_2961,N_2959);
or UO_481 (O_481,N_2961,N_2955);
or UO_482 (O_482,N_2960,N_2969);
nor UO_483 (O_483,N_2992,N_2987);
xor UO_484 (O_484,N_2946,N_2981);
and UO_485 (O_485,N_2994,N_2997);
and UO_486 (O_486,N_2970,N_2962);
xor UO_487 (O_487,N_2971,N_2947);
or UO_488 (O_488,N_2975,N_2954);
or UO_489 (O_489,N_2956,N_2972);
nand UO_490 (O_490,N_2964,N_2995);
or UO_491 (O_491,N_2951,N_2970);
xnor UO_492 (O_492,N_2954,N_2981);
or UO_493 (O_493,N_2982,N_2954);
or UO_494 (O_494,N_2957,N_2959);
xor UO_495 (O_495,N_2982,N_2949);
or UO_496 (O_496,N_2954,N_2989);
nor UO_497 (O_497,N_2985,N_2976);
xnor UO_498 (O_498,N_2955,N_2974);
xnor UO_499 (O_499,N_2988,N_2973);
endmodule