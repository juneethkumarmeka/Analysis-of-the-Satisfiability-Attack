module basic_1000_10000_1500_50_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_470,In_588);
or U1 (N_1,In_806,In_957);
nand U2 (N_2,In_492,In_722);
nand U3 (N_3,In_691,In_598);
nor U4 (N_4,In_522,In_425);
or U5 (N_5,In_201,In_919);
and U6 (N_6,In_413,In_79);
and U7 (N_7,In_737,In_213);
nand U8 (N_8,In_874,In_973);
xor U9 (N_9,In_170,In_904);
xor U10 (N_10,In_929,In_310);
nor U11 (N_11,In_19,In_85);
nand U12 (N_12,In_117,In_840);
and U13 (N_13,In_134,In_266);
nand U14 (N_14,In_547,In_561);
nand U15 (N_15,In_426,In_686);
and U16 (N_16,In_819,In_464);
nor U17 (N_17,In_37,In_485);
or U18 (N_18,In_195,In_996);
nor U19 (N_19,In_750,In_854);
nor U20 (N_20,In_497,In_967);
and U21 (N_21,In_365,In_924);
nand U22 (N_22,In_931,In_409);
nor U23 (N_23,In_900,In_476);
and U24 (N_24,In_120,In_294);
and U25 (N_25,In_226,In_937);
nor U26 (N_26,In_38,In_752);
nor U27 (N_27,In_742,In_692);
nor U28 (N_28,In_3,In_200);
or U29 (N_29,In_495,In_756);
nand U30 (N_30,In_728,In_110);
nor U31 (N_31,In_999,In_24);
xor U32 (N_32,In_979,In_76);
or U33 (N_33,In_263,In_576);
nor U34 (N_34,In_600,In_143);
nand U35 (N_35,In_34,In_23);
or U36 (N_36,In_718,In_455);
nand U37 (N_37,In_100,In_665);
nand U38 (N_38,In_368,In_80);
nor U39 (N_39,In_594,In_624);
or U40 (N_40,In_214,In_968);
xnor U41 (N_41,In_963,In_389);
xor U42 (N_42,In_606,In_644);
nor U43 (N_43,In_813,In_658);
and U44 (N_44,In_474,In_468);
and U45 (N_45,In_460,In_851);
xnor U46 (N_46,In_156,In_866);
nor U47 (N_47,In_596,In_798);
nand U48 (N_48,In_613,In_735);
and U49 (N_49,In_843,In_431);
and U50 (N_50,In_281,In_630);
nor U51 (N_51,In_52,In_99);
xor U52 (N_52,In_188,In_885);
nand U53 (N_53,In_231,In_387);
or U54 (N_54,In_295,In_577);
nand U55 (N_55,In_567,In_941);
xnor U56 (N_56,In_933,In_140);
or U57 (N_57,In_126,In_340);
nor U58 (N_58,In_660,In_792);
and U59 (N_59,In_706,In_308);
xnor U60 (N_60,In_595,In_920);
nand U61 (N_61,In_357,In_720);
xnor U62 (N_62,In_636,In_564);
nand U63 (N_63,In_709,In_884);
or U64 (N_64,In_590,In_190);
or U65 (N_65,In_865,In_732);
or U66 (N_66,In_825,In_557);
or U67 (N_67,In_956,In_939);
xnor U68 (N_68,In_17,In_58);
nor U69 (N_69,In_786,In_127);
nor U70 (N_70,In_723,In_647);
or U71 (N_71,In_318,In_898);
or U72 (N_72,In_44,In_662);
nand U73 (N_73,In_244,In_30);
nor U74 (N_74,In_301,In_314);
nor U75 (N_75,In_95,In_404);
xnor U76 (N_76,In_254,In_291);
nor U77 (N_77,In_240,In_418);
nand U78 (N_78,In_589,In_882);
nor U79 (N_79,In_947,In_66);
and U80 (N_80,In_118,In_356);
nand U81 (N_81,In_493,In_326);
xnor U82 (N_82,In_207,In_70);
nand U83 (N_83,In_237,In_247);
xor U84 (N_84,In_142,In_345);
xor U85 (N_85,In_976,In_73);
xor U86 (N_86,In_498,In_333);
nor U87 (N_87,In_611,In_63);
nand U88 (N_88,In_778,In_75);
or U89 (N_89,In_123,In_27);
or U90 (N_90,In_727,In_958);
or U91 (N_91,In_151,In_678);
nand U92 (N_92,In_661,In_158);
and U93 (N_93,In_65,In_128);
and U94 (N_94,In_500,In_11);
nand U95 (N_95,In_946,In_991);
or U96 (N_96,In_646,In_265);
or U97 (N_97,In_508,In_290);
xor U98 (N_98,In_275,In_969);
nor U99 (N_99,In_154,In_36);
nand U100 (N_100,In_91,In_125);
nand U101 (N_101,In_452,In_930);
or U102 (N_102,In_615,In_812);
nor U103 (N_103,In_233,In_109);
nor U104 (N_104,In_67,In_679);
xnor U105 (N_105,In_415,In_952);
or U106 (N_106,In_530,In_748);
and U107 (N_107,In_248,In_55);
nor U108 (N_108,In_824,In_815);
or U109 (N_109,In_563,In_965);
or U110 (N_110,In_139,In_372);
and U111 (N_111,In_451,In_446);
nand U112 (N_112,In_483,In_977);
or U113 (N_113,In_381,In_971);
and U114 (N_114,In_124,In_717);
nor U115 (N_115,In_593,In_829);
xnor U116 (N_116,In_434,In_499);
nor U117 (N_117,In_922,In_512);
xnor U118 (N_118,In_478,In_974);
or U119 (N_119,In_699,In_166);
nor U120 (N_120,In_932,In_582);
and U121 (N_121,In_986,In_719);
or U122 (N_122,In_241,In_890);
nor U123 (N_123,In_227,In_304);
xnor U124 (N_124,In_463,In_774);
or U125 (N_125,In_726,In_799);
and U126 (N_126,In_74,In_521);
nor U127 (N_127,In_934,In_373);
xor U128 (N_128,In_320,In_927);
xor U129 (N_129,In_211,In_776);
xnor U130 (N_130,In_664,In_212);
xnor U131 (N_131,In_670,In_849);
nor U132 (N_132,In_654,In_566);
nand U133 (N_133,In_641,In_48);
nand U134 (N_134,In_453,In_697);
nand U135 (N_135,In_961,In_22);
and U136 (N_136,In_584,In_210);
nand U137 (N_137,In_773,In_349);
or U138 (N_138,In_362,In_808);
nand U139 (N_139,In_449,In_358);
nand U140 (N_140,In_571,In_2);
and U141 (N_141,In_4,In_185);
nand U142 (N_142,In_954,In_271);
and U143 (N_143,In_714,In_666);
nor U144 (N_144,In_873,In_323);
or U145 (N_145,In_758,In_383);
xor U146 (N_146,In_385,In_674);
and U147 (N_147,In_183,In_89);
xnor U148 (N_148,In_42,In_917);
and U149 (N_149,In_7,In_995);
nor U150 (N_150,In_804,In_159);
and U151 (N_151,In_867,In_307);
and U152 (N_152,In_472,In_380);
nand U153 (N_153,In_779,In_793);
xor U154 (N_154,In_155,In_861);
and U155 (N_155,In_940,In_57);
nor U156 (N_156,In_671,In_517);
and U157 (N_157,In_948,In_132);
xnor U158 (N_158,In_410,In_157);
nand U159 (N_159,In_620,In_520);
nor U160 (N_160,In_342,In_878);
and U161 (N_161,In_261,In_13);
and U162 (N_162,In_545,In_273);
or U163 (N_163,In_423,In_788);
or U164 (N_164,In_894,In_928);
nand U165 (N_165,In_145,In_574);
nor U166 (N_166,In_264,In_762);
nand U167 (N_167,In_315,In_831);
nand U168 (N_168,In_311,In_419);
or U169 (N_169,In_256,In_760);
and U170 (N_170,In_18,In_649);
nand U171 (N_171,In_822,In_568);
or U172 (N_172,In_909,In_397);
nor U173 (N_173,In_411,In_570);
and U174 (N_174,In_113,In_82);
xnor U175 (N_175,In_1,In_562);
nand U176 (N_176,In_329,In_970);
xnor U177 (N_177,In_586,In_502);
or U178 (N_178,In_33,In_627);
xor U179 (N_179,In_787,In_121);
xor U180 (N_180,In_703,In_442);
nor U181 (N_181,In_989,In_285);
nor U182 (N_182,In_889,In_730);
and U183 (N_183,In_833,In_81);
or U184 (N_184,In_313,In_436);
nand U185 (N_185,In_114,In_300);
or U186 (N_186,In_685,In_303);
and U187 (N_187,In_642,In_191);
nand U188 (N_188,In_777,In_847);
nor U189 (N_189,In_603,In_921);
or U190 (N_190,In_529,In_949);
nor U191 (N_191,In_136,In_165);
xor U192 (N_192,In_6,In_386);
nand U193 (N_193,In_287,In_454);
or U194 (N_194,In_108,In_111);
and U195 (N_195,In_267,In_149);
or U196 (N_196,In_344,In_797);
and U197 (N_197,In_86,In_407);
xnor U198 (N_198,In_655,In_236);
or U199 (N_199,In_913,In_115);
nand U200 (N_200,N_183,N_103);
xor U201 (N_201,In_177,In_651);
nand U202 (N_202,In_626,In_169);
and U203 (N_203,N_113,N_187);
xnor U204 (N_204,In_791,N_88);
xnor U205 (N_205,In_14,In_775);
nor U206 (N_206,In_993,In_648);
nor U207 (N_207,In_461,In_417);
and U208 (N_208,In_68,In_339);
nor U209 (N_209,In_650,In_559);
nand U210 (N_210,In_994,In_286);
or U211 (N_211,In_288,N_142);
and U212 (N_212,In_980,In_49);
or U213 (N_213,N_49,In_72);
and U214 (N_214,In_950,In_260);
nand U215 (N_215,In_908,In_440);
xor U216 (N_216,N_163,In_435);
nand U217 (N_217,N_145,In_875);
nand U218 (N_218,In_886,In_533);
and U219 (N_219,In_428,In_604);
nand U220 (N_220,In_635,In_987);
nand U221 (N_221,In_540,N_8);
nor U222 (N_222,N_140,In_332);
or U223 (N_223,N_62,N_84);
nor U224 (N_224,In_197,In_811);
nor U225 (N_225,N_128,In_633);
nor U226 (N_226,In_964,In_814);
nand U227 (N_227,In_462,In_607);
xnor U228 (N_228,N_19,In_97);
nand U229 (N_229,In_997,In_141);
nand U230 (N_230,N_6,N_148);
and U231 (N_231,N_52,N_139);
or U232 (N_232,In_284,N_4);
nand U233 (N_233,In_59,In_205);
or U234 (N_234,In_712,In_312);
nand U235 (N_235,In_809,N_144);
nand U236 (N_236,In_915,N_149);
and U237 (N_237,In_219,In_579);
nor U238 (N_238,N_21,In_768);
or U239 (N_239,In_251,In_269);
nand U240 (N_240,In_743,In_724);
nand U241 (N_241,In_370,In_807);
or U242 (N_242,In_837,In_926);
xor U243 (N_243,In_558,N_189);
or U244 (N_244,N_66,In_252);
nor U245 (N_245,In_523,N_196);
xnor U246 (N_246,In_892,In_278);
nand U247 (N_247,N_43,In_507);
nor U248 (N_248,In_783,In_374);
xnor U249 (N_249,In_751,In_622);
nor U250 (N_250,In_580,N_94);
nor U251 (N_251,In_21,In_710);
nor U252 (N_252,In_222,In_178);
and U253 (N_253,In_769,N_178);
nor U254 (N_254,In_176,N_61);
or U255 (N_255,In_863,In_62);
nor U256 (N_256,In_475,N_73);
and U257 (N_257,In_322,In_221);
nand U258 (N_258,In_872,In_518);
xor U259 (N_259,In_84,N_25);
nor U260 (N_260,In_309,N_10);
nand U261 (N_261,In_810,In_47);
nand U262 (N_262,N_86,In_198);
or U263 (N_263,In_560,In_489);
or U264 (N_264,In_317,N_87);
nand U265 (N_265,N_117,N_132);
nand U266 (N_266,In_179,In_782);
or U267 (N_267,In_232,In_511);
xor U268 (N_268,In_652,In_700);
xnor U269 (N_269,In_781,In_150);
nor U270 (N_270,In_384,N_146);
or U271 (N_271,In_458,In_516);
and U272 (N_272,In_43,N_18);
nand U273 (N_273,In_695,In_282);
and U274 (N_274,In_98,In_54);
or U275 (N_275,N_158,N_157);
nor U276 (N_276,N_192,In_868);
or U277 (N_277,N_64,N_194);
nand U278 (N_278,In_45,In_618);
xor U279 (N_279,In_803,In_167);
nor U280 (N_280,In_293,N_55);
xor U281 (N_281,In_888,In_864);
or U282 (N_282,N_155,N_81);
xor U283 (N_283,In_350,In_616);
and U284 (N_284,In_443,N_124);
or U285 (N_285,In_850,In_28);
xor U286 (N_286,N_170,In_550);
and U287 (N_287,N_95,In_8);
and U288 (N_288,In_245,In_9);
xor U289 (N_289,In_754,N_102);
nor U290 (N_290,In_32,N_36);
and U291 (N_291,In_677,In_536);
and U292 (N_292,In_733,In_524);
nand U293 (N_293,In_747,In_257);
nor U294 (N_294,N_177,In_528);
nor U295 (N_295,In_355,In_77);
nand U296 (N_296,In_610,In_535);
xor U297 (N_297,In_725,In_501);
or U298 (N_298,In_399,N_114);
nand U299 (N_299,In_130,In_916);
nor U300 (N_300,In_601,In_160);
and U301 (N_301,In_148,In_643);
xnor U302 (N_302,In_820,In_862);
xnor U303 (N_303,N_26,N_184);
or U304 (N_304,N_17,In_10);
nor U305 (N_305,In_541,In_279);
xor U306 (N_306,In_41,In_897);
nand U307 (N_307,N_160,In_334);
or U308 (N_308,In_194,In_767);
and U309 (N_309,In_795,In_962);
nor U310 (N_310,In_430,In_336);
or U311 (N_311,In_390,In_164);
xor U312 (N_312,In_481,N_59);
xnor U313 (N_313,In_623,In_983);
xor U314 (N_314,In_78,N_7);
nand U315 (N_315,N_180,N_93);
and U316 (N_316,N_159,In_942);
or U317 (N_317,In_484,In_467);
or U318 (N_318,N_186,In_94);
or U319 (N_319,In_966,In_450);
nand U320 (N_320,In_363,In_346);
and U321 (N_321,In_551,In_585);
nand U322 (N_322,N_16,N_51);
nor U323 (N_323,In_944,N_154);
or U324 (N_324,In_180,In_96);
xnor U325 (N_325,In_640,In_348);
nor U326 (N_326,In_659,In_525);
nand U327 (N_327,In_527,In_734);
nand U328 (N_328,In_899,In_532);
nand U329 (N_329,In_255,N_0);
and U330 (N_330,N_137,In_208);
nor U331 (N_331,In_869,In_746);
xor U332 (N_332,In_376,In_53);
and U333 (N_333,N_190,N_1);
nand U334 (N_334,N_127,N_150);
nor U335 (N_335,In_539,In_327);
and U336 (N_336,In_513,N_133);
nand U337 (N_337,In_144,N_22);
or U338 (N_338,In_675,In_494);
and U339 (N_339,In_519,In_785);
nand U340 (N_340,In_341,N_120);
nor U341 (N_341,N_75,In_138);
nand U342 (N_342,In_534,In_935);
xor U343 (N_343,In_716,In_510);
or U344 (N_344,N_90,In_135);
and U345 (N_345,In_87,N_104);
or U346 (N_346,In_592,In_509);
and U347 (N_347,In_337,In_552);
or U348 (N_348,N_72,In_223);
xor U349 (N_349,In_262,In_92);
xor U350 (N_350,In_910,In_591);
nand U351 (N_351,In_229,In_998);
nand U352 (N_352,In_29,In_230);
and U353 (N_353,In_347,In_631);
xor U354 (N_354,In_801,In_441);
xor U355 (N_355,In_444,In_871);
or U356 (N_356,N_134,In_876);
and U357 (N_357,N_83,In_653);
nand U358 (N_358,In_181,In_209);
and U359 (N_359,In_107,In_259);
xor U360 (N_360,In_147,In_672);
nand U361 (N_361,N_176,In_161);
or U362 (N_362,N_67,In_629);
nor U363 (N_363,In_856,N_168);
xor U364 (N_364,N_31,In_555);
nand U365 (N_365,In_408,In_395);
nand U366 (N_366,In_238,N_33);
nor U367 (N_367,In_25,In_152);
or U368 (N_368,N_98,In_466);
and U369 (N_369,In_826,In_16);
nor U370 (N_370,In_985,In_137);
and U371 (N_371,In_951,In_400);
xnor U372 (N_372,N_27,N_14);
and U373 (N_373,In_901,N_53);
or U374 (N_374,In_857,In_189);
or U375 (N_375,In_770,In_292);
nor U376 (N_376,In_575,In_503);
and U377 (N_377,N_136,In_379);
nor U378 (N_378,In_371,In_828);
or U379 (N_379,In_548,In_272);
and U380 (N_380,In_903,N_165);
xor U381 (N_381,In_172,In_701);
nor U382 (N_382,In_845,In_682);
nand U383 (N_383,N_101,In_26);
or U384 (N_384,In_71,In_634);
nor U385 (N_385,In_538,In_496);
and U386 (N_386,N_123,N_5);
nand U387 (N_387,N_23,In_39);
or U388 (N_388,N_96,N_112);
xor U389 (N_389,In_184,In_122);
nand U390 (N_390,In_578,In_784);
nor U391 (N_391,In_681,In_447);
or U392 (N_392,In_193,In_708);
xor U393 (N_393,In_855,In_736);
or U394 (N_394,In_852,In_978);
and U395 (N_395,In_242,In_702);
nand U396 (N_396,In_473,In_0);
and U397 (N_397,N_105,N_15);
or U398 (N_398,In_325,In_583);
xnor U399 (N_399,N_11,N_169);
xnor U400 (N_400,In_945,In_249);
nand U401 (N_401,N_244,In_883);
nand U402 (N_402,In_422,N_349);
and U403 (N_403,N_37,N_201);
nor U404 (N_404,In_343,N_272);
or U405 (N_405,N_256,In_597);
nor U406 (N_406,In_763,In_187);
and U407 (N_407,In_805,In_173);
nand U408 (N_408,N_230,N_269);
or U409 (N_409,In_895,N_388);
and U410 (N_410,N_34,N_40);
and U411 (N_411,N_250,In_705);
and U412 (N_412,In_234,In_554);
and U413 (N_413,In_253,In_186);
nor U414 (N_414,N_339,In_12);
xnor U415 (N_415,In_953,N_351);
and U416 (N_416,N_239,N_391);
xor U417 (N_417,In_960,In_764);
xor U418 (N_418,In_599,N_381);
and U419 (N_419,N_32,N_108);
or U420 (N_420,N_397,N_205);
and U421 (N_421,In_490,In_835);
xnor U422 (N_422,In_739,N_131);
nor U423 (N_423,In_424,In_761);
nand U424 (N_424,N_212,N_130);
nand U425 (N_425,N_82,In_324);
or U426 (N_426,N_213,In_90);
or U427 (N_427,N_312,In_738);
or U428 (N_428,N_232,In_394);
or U429 (N_429,In_907,In_696);
or U430 (N_430,N_358,In_684);
nor U431 (N_431,N_209,In_438);
xor U432 (N_432,N_365,N_368);
or U433 (N_433,In_657,N_100);
or U434 (N_434,N_153,In_354);
nand U435 (N_435,N_185,N_370);
and U436 (N_436,In_638,N_47);
or U437 (N_437,In_830,N_276);
nor U438 (N_438,N_389,N_92);
nand U439 (N_439,N_291,N_226);
nor U440 (N_440,N_138,N_208);
nand U441 (N_441,N_362,In_405);
nor U442 (N_442,In_800,In_352);
or U443 (N_443,N_227,N_204);
or U444 (N_444,N_387,In_608);
and U445 (N_445,In_975,N_390);
nor U446 (N_446,N_344,N_299);
nand U447 (N_447,In_171,N_333);
or U448 (N_448,N_392,N_3);
or U449 (N_449,N_12,In_549);
xor U450 (N_450,N_216,In_639);
or U451 (N_451,In_765,In_881);
nor U452 (N_452,N_316,N_210);
nand U453 (N_453,N_340,In_217);
or U454 (N_454,N_287,In_715);
nor U455 (N_455,In_687,N_374);
and U456 (N_456,N_314,N_89);
or U457 (N_457,N_273,In_250);
and U458 (N_458,In_133,N_39);
and U459 (N_459,In_988,N_69);
or U460 (N_460,N_279,N_218);
nor U461 (N_461,N_313,In_106);
or U462 (N_462,In_429,In_297);
and U463 (N_463,In_388,N_231);
or U464 (N_464,N_296,In_393);
xnor U465 (N_465,In_375,In_199);
nor U466 (N_466,N_41,In_556);
xor U467 (N_467,In_572,N_56);
xnor U468 (N_468,In_543,In_235);
nand U469 (N_469,In_328,N_282);
nor U470 (N_470,N_293,In_880);
nand U471 (N_471,In_175,N_164);
nand U472 (N_472,N_193,N_175);
nand U473 (N_473,N_307,In_69);
xor U474 (N_474,N_382,In_335);
nand U475 (N_475,In_224,In_617);
or U476 (N_476,In_925,In_602);
nand U477 (N_477,In_471,N_295);
nand U478 (N_478,In_174,N_331);
nor U479 (N_479,In_46,N_118);
and U480 (N_480,In_858,In_353);
nor U481 (N_481,In_305,In_64);
or U482 (N_482,N_236,N_320);
or U483 (N_483,In_515,In_704);
nor U484 (N_484,In_162,N_30);
xnor U485 (N_485,In_351,N_181);
and U486 (N_486,In_20,N_42);
xnor U487 (N_487,N_294,In_711);
or U488 (N_488,N_115,N_199);
nand U489 (N_489,In_105,N_283);
nor U490 (N_490,N_57,In_749);
or U491 (N_491,N_161,In_359);
nor U492 (N_492,N_45,N_305);
or U493 (N_493,In_280,In_406);
nand U494 (N_494,In_296,In_816);
nor U495 (N_495,In_656,In_319);
and U496 (N_496,In_955,In_731);
nand U497 (N_497,N_359,N_277);
and U498 (N_498,N_174,In_215);
xor U499 (N_499,N_135,N_308);
and U500 (N_500,In_729,In_488);
and U501 (N_501,N_197,In_378);
nand U502 (N_502,N_259,In_243);
nand U503 (N_503,In_565,In_771);
xnor U504 (N_504,N_9,In_621);
nor U505 (N_505,In_839,N_321);
nand U506 (N_506,In_887,In_605);
xor U507 (N_507,In_984,In_896);
nand U508 (N_508,N_311,N_342);
xor U509 (N_509,In_836,N_267);
or U510 (N_510,In_412,In_506);
nor U511 (N_511,N_97,N_166);
nor U512 (N_512,N_361,In_859);
xnor U513 (N_513,N_182,N_309);
nor U514 (N_514,N_111,N_71);
nor U515 (N_515,In_270,N_372);
xor U516 (N_516,In_218,In_698);
nand U517 (N_517,N_355,In_790);
nor U518 (N_518,In_302,In_741);
or U519 (N_519,N_345,In_401);
nor U520 (N_520,In_83,N_141);
and U521 (N_521,In_131,N_380);
xor U522 (N_522,N_375,In_316);
nand U523 (N_523,In_283,N_384);
or U524 (N_524,In_146,In_690);
nand U525 (N_525,N_325,In_338);
nor U526 (N_526,In_990,In_817);
and U527 (N_527,N_29,N_284);
nor U528 (N_528,N_237,In_766);
or U529 (N_529,In_673,N_38);
xnor U530 (N_530,N_386,N_206);
nand U531 (N_531,In_35,In_504);
nor U532 (N_532,N_242,In_537);
nor U533 (N_533,In_669,N_247);
nor U534 (N_534,In_289,In_459);
nand U535 (N_535,N_255,N_352);
and U536 (N_536,In_182,In_693);
nor U537 (N_537,In_361,In_204);
xor U538 (N_538,In_914,N_122);
nor U539 (N_539,In_683,In_694);
or U540 (N_540,In_5,In_821);
nand U541 (N_541,In_268,N_246);
xnor U542 (N_542,In_688,In_391);
nor U543 (N_543,N_233,N_65);
xnor U544 (N_544,In_905,In_40);
or U545 (N_545,N_13,In_796);
xnor U546 (N_546,N_211,In_206);
nor U547 (N_547,N_195,In_220);
and U548 (N_548,In_860,N_110);
and U549 (N_549,In_482,N_106);
and U550 (N_550,N_35,N_357);
nor U551 (N_551,In_542,In_366);
and U552 (N_552,N_58,In_276);
or U553 (N_553,In_433,N_290);
or U554 (N_554,N_376,In_938);
nand U555 (N_555,N_300,N_215);
and U556 (N_556,N_371,N_77);
xnor U557 (N_557,N_281,In_581);
and U558 (N_558,In_246,N_297);
or U559 (N_559,In_663,N_254);
and U560 (N_560,N_366,In_129);
and U561 (N_561,N_346,In_403);
or U562 (N_562,In_239,In_757);
nor U563 (N_563,In_56,N_332);
nor U564 (N_564,N_200,N_398);
nand U565 (N_565,In_367,In_546);
nand U566 (N_566,In_486,In_959);
xnor U567 (N_567,N_235,N_234);
xnor U568 (N_568,N_315,In_587);
nor U569 (N_569,In_680,N_151);
nand U570 (N_570,In_465,N_63);
or U571 (N_571,N_379,In_420);
nand U572 (N_572,N_78,In_753);
and U573 (N_573,In_870,In_360);
xor U574 (N_574,In_31,In_982);
nor U575 (N_575,N_119,In_637);
nor U576 (N_576,In_844,In_823);
nor U577 (N_577,N_243,In_645);
xor U578 (N_578,In_479,N_179);
and U579 (N_579,N_44,N_356);
nand U580 (N_580,N_394,N_280);
and U581 (N_581,N_167,In_612);
and U582 (N_582,N_173,N_129);
nand U583 (N_583,N_275,In_573);
nand U584 (N_584,N_348,In_553);
xnor U585 (N_585,In_102,In_258);
nand U586 (N_586,In_364,N_24);
nor U587 (N_587,In_330,N_306);
nand U588 (N_588,In_619,N_202);
or U589 (N_589,N_198,N_109);
xnor U590 (N_590,N_285,N_220);
nand U591 (N_591,N_360,N_260);
nor U592 (N_592,N_341,In_912);
nor U593 (N_593,N_147,In_972);
xor U594 (N_594,In_848,In_981);
nor U595 (N_595,In_203,N_328);
or U596 (N_596,In_755,N_322);
nand U597 (N_597,N_229,N_369);
and U598 (N_598,N_262,N_347);
or U599 (N_599,In_392,N_60);
xnor U600 (N_600,N_444,N_405);
and U601 (N_601,N_495,N_511);
and U602 (N_602,N_461,N_538);
or U603 (N_603,N_418,N_427);
nand U604 (N_604,N_578,N_403);
xor U605 (N_605,N_472,N_432);
xnor U606 (N_606,N_518,N_425);
or U607 (N_607,N_579,N_546);
and U608 (N_608,N_459,N_191);
nor U609 (N_609,N_583,N_363);
nand U610 (N_610,In_891,N_270);
nor U611 (N_611,N_261,N_457);
nand U612 (N_612,In_456,N_171);
and U613 (N_613,N_404,N_525);
xnor U614 (N_614,N_527,N_493);
xnor U615 (N_615,In_744,In_491);
nor U616 (N_616,In_877,In_842);
nand U617 (N_617,N_485,N_480);
nand U618 (N_618,N_594,N_523);
or U619 (N_619,N_467,N_248);
or U620 (N_620,In_936,N_324);
and U621 (N_621,In_923,In_846);
xnor U622 (N_622,N_458,N_593);
or U623 (N_623,N_524,N_488);
nand U624 (N_624,N_557,N_599);
nor U625 (N_625,N_529,In_772);
xor U626 (N_626,In_625,N_519);
nor U627 (N_627,In_228,N_268);
nor U628 (N_628,N_559,N_568);
nand U629 (N_629,N_564,In_480);
xor U630 (N_630,N_249,In_526);
and U631 (N_631,N_415,In_382);
nor U632 (N_632,In_101,N_449);
xor U633 (N_633,N_595,N_534);
xor U634 (N_634,N_503,N_500);
xor U635 (N_635,N_482,N_402);
nand U636 (N_636,N_567,In_609);
xor U637 (N_637,N_552,In_745);
and U638 (N_638,N_532,N_50);
nor U639 (N_639,N_126,N_207);
and U640 (N_640,N_162,N_121);
nor U641 (N_641,N_494,N_399);
nor U642 (N_642,N_264,N_413);
or U643 (N_643,N_514,N_188);
and U644 (N_644,In_396,N_228);
or U645 (N_645,N_253,N_396);
and U646 (N_646,N_116,In_51);
and U647 (N_647,N_240,In_369);
nand U648 (N_648,N_489,N_490);
nor U649 (N_649,In_841,N_597);
nor U650 (N_650,In_759,N_589);
nor U651 (N_651,In_632,N_452);
or U652 (N_652,N_301,N_563);
nor U653 (N_653,In_414,N_419);
and U654 (N_654,In_216,N_414);
nor U655 (N_655,N_421,In_906);
nor U656 (N_656,In_104,In_196);
or U657 (N_657,N_393,N_203);
nor U658 (N_658,N_302,N_492);
xor U659 (N_659,N_571,In_918);
and U660 (N_660,In_437,N_542);
xnor U661 (N_661,N_79,N_501);
or U662 (N_662,N_411,N_28);
or U663 (N_663,N_453,N_70);
nor U664 (N_664,N_225,N_515);
and U665 (N_665,N_326,N_505);
nor U666 (N_666,N_550,N_378);
or U667 (N_667,N_412,N_545);
and U668 (N_668,N_558,N_156);
nor U669 (N_669,In_119,In_879);
or U670 (N_670,In_544,N_516);
xnor U671 (N_671,N_318,N_541);
nor U672 (N_672,N_330,N_469);
and U673 (N_673,N_274,N_576);
or U674 (N_674,N_245,In_448);
or U675 (N_675,In_116,In_445);
and U676 (N_676,N_329,N_540);
xnor U677 (N_677,In_487,N_286);
nor U678 (N_678,N_241,In_153);
nor U679 (N_679,N_460,N_426);
nand U680 (N_680,N_553,In_277);
or U681 (N_681,N_303,In_911);
xnor U682 (N_682,N_441,N_46);
xor U683 (N_683,N_508,N_581);
xor U684 (N_684,N_451,N_338);
and U685 (N_685,In_838,In_439);
or U686 (N_686,N_420,N_475);
nor U687 (N_687,In_274,N_507);
xnor U688 (N_688,N_454,N_548);
nor U689 (N_689,N_543,N_172);
nor U690 (N_690,In_15,N_437);
nor U691 (N_691,N_510,N_439);
nand U692 (N_692,N_377,N_539);
and U693 (N_693,N_544,N_336);
nor U694 (N_694,N_463,In_943);
nor U695 (N_695,In_88,N_468);
or U696 (N_696,N_478,In_202);
and U697 (N_697,N_400,N_434);
or U698 (N_698,N_504,N_143);
or U699 (N_699,N_520,N_590);
or U700 (N_700,In_377,In_168);
xnor U701 (N_701,N_217,N_592);
or U702 (N_702,N_317,In_794);
and U703 (N_703,N_423,N_481);
nor U704 (N_704,N_68,In_818);
nor U705 (N_705,N_2,N_20);
nand U706 (N_706,N_431,N_555);
nor U707 (N_707,N_223,N_450);
xor U708 (N_708,N_319,N_438);
xor U709 (N_709,In_902,N_486);
or U710 (N_710,N_577,N_512);
nand U711 (N_711,N_526,N_584);
nor U712 (N_712,N_288,N_497);
or U713 (N_713,N_513,N_566);
xor U714 (N_714,N_487,N_407);
or U715 (N_715,N_424,N_263);
or U716 (N_716,In_628,N_266);
and U717 (N_717,In_469,N_591);
xor U718 (N_718,N_278,N_477);
and U719 (N_719,In_721,N_74);
and U720 (N_720,N_572,N_334);
and U721 (N_721,N_440,N_354);
nor U722 (N_722,N_416,N_80);
or U723 (N_723,N_221,In_834);
nor U724 (N_724,N_238,N_343);
xor U725 (N_725,N_473,In_298);
nand U726 (N_726,N_385,N_353);
nor U727 (N_727,N_547,N_446);
xor U728 (N_728,N_502,In_61);
or U729 (N_729,N_289,N_335);
nand U730 (N_730,N_556,In_505);
or U731 (N_731,In_427,N_466);
nor U732 (N_732,N_470,N_409);
or U733 (N_733,N_456,N_430);
or U734 (N_734,N_462,N_588);
nand U735 (N_735,N_565,N_417);
or U736 (N_736,N_498,In_416);
or U737 (N_737,N_530,In_331);
and U738 (N_738,N_484,N_443);
or U739 (N_739,N_265,In_306);
nand U740 (N_740,In_802,N_435);
nor U741 (N_741,N_222,N_465);
nand U742 (N_742,In_780,N_491);
or U743 (N_743,N_561,In_992);
and U744 (N_744,N_506,N_533);
xor U745 (N_745,N_251,N_521);
nand U746 (N_746,N_496,N_570);
xnor U747 (N_747,N_476,N_323);
nand U748 (N_748,N_401,In_668);
or U749 (N_749,N_367,N_499);
xnor U750 (N_750,N_522,N_587);
nand U751 (N_751,N_509,N_535);
or U752 (N_752,N_350,N_536);
nor U753 (N_753,N_447,N_573);
or U754 (N_754,N_528,N_76);
nor U755 (N_755,In_514,N_125);
and U756 (N_756,In_853,N_455);
or U757 (N_757,N_436,N_531);
nand U758 (N_758,N_410,N_214);
xor U759 (N_759,N_85,In_667);
nand U760 (N_760,N_364,In_225);
nand U761 (N_761,N_445,N_337);
nor U762 (N_762,N_224,N_598);
and U763 (N_763,N_48,N_574);
nor U764 (N_764,In_421,N_91);
nand U765 (N_765,N_551,N_483);
xnor U766 (N_766,N_152,N_537);
xnor U767 (N_767,N_99,N_586);
nor U768 (N_768,N_479,N_429);
and U769 (N_769,N_554,In_60);
nand U770 (N_770,N_252,In_689);
or U771 (N_771,N_471,In_707);
and U772 (N_772,N_271,In_789);
or U773 (N_773,N_580,In_93);
or U774 (N_774,In_112,In_893);
xor U775 (N_775,N_569,In_321);
nand U776 (N_776,N_433,N_292);
xor U777 (N_777,N_408,N_582);
and U778 (N_778,N_448,N_383);
nand U779 (N_779,In_432,In_832);
nor U780 (N_780,In_569,In_457);
nor U781 (N_781,N_442,In_827);
nand U782 (N_782,In_50,N_258);
nor U783 (N_783,N_428,N_257);
nor U784 (N_784,In_676,N_575);
or U785 (N_785,N_310,N_560);
and U786 (N_786,N_474,N_406);
xor U787 (N_787,N_298,In_477);
nand U788 (N_788,N_373,In_299);
xor U789 (N_789,N_395,In_531);
xnor U790 (N_790,N_549,N_54);
xor U791 (N_791,In_614,N_596);
xor U792 (N_792,N_304,In_740);
and U793 (N_793,N_422,N_327);
xor U794 (N_794,In_192,In_402);
nor U795 (N_795,N_107,In_398);
nand U796 (N_796,N_585,In_103);
or U797 (N_797,In_713,In_163);
nand U798 (N_798,N_219,N_517);
nor U799 (N_799,N_562,N_464);
xnor U800 (N_800,N_730,N_774);
xnor U801 (N_801,N_748,N_636);
or U802 (N_802,N_680,N_699);
and U803 (N_803,N_610,N_734);
and U804 (N_804,N_754,N_652);
or U805 (N_805,N_724,N_667);
nand U806 (N_806,N_720,N_693);
xnor U807 (N_807,N_723,N_691);
nand U808 (N_808,N_687,N_784);
or U809 (N_809,N_726,N_778);
nand U810 (N_810,N_702,N_744);
nand U811 (N_811,N_722,N_738);
or U812 (N_812,N_780,N_753);
xor U813 (N_813,N_655,N_740);
nand U814 (N_814,N_609,N_616);
and U815 (N_815,N_706,N_612);
nor U816 (N_816,N_653,N_679);
xor U817 (N_817,N_683,N_617);
nor U818 (N_818,N_697,N_786);
and U819 (N_819,N_606,N_641);
nor U820 (N_820,N_710,N_767);
nand U821 (N_821,N_619,N_764);
and U822 (N_822,N_659,N_692);
and U823 (N_823,N_631,N_777);
nand U824 (N_824,N_731,N_634);
and U825 (N_825,N_625,N_694);
nor U826 (N_826,N_672,N_678);
xnor U827 (N_827,N_732,N_714);
xor U828 (N_828,N_628,N_637);
and U829 (N_829,N_765,N_772);
and U830 (N_830,N_638,N_799);
xor U831 (N_831,N_763,N_604);
or U832 (N_832,N_712,N_709);
or U833 (N_833,N_622,N_645);
xor U834 (N_834,N_749,N_623);
nand U835 (N_835,N_707,N_776);
or U836 (N_836,N_658,N_607);
xor U837 (N_837,N_755,N_721);
nand U838 (N_838,N_790,N_686);
or U839 (N_839,N_635,N_779);
and U840 (N_840,N_698,N_627);
nor U841 (N_841,N_770,N_789);
and U842 (N_842,N_781,N_798);
or U843 (N_843,N_758,N_689);
and U844 (N_844,N_797,N_639);
and U845 (N_845,N_752,N_751);
or U846 (N_846,N_768,N_633);
and U847 (N_847,N_727,N_671);
and U848 (N_848,N_773,N_685);
and U849 (N_849,N_743,N_759);
or U850 (N_850,N_665,N_771);
xnor U851 (N_851,N_651,N_642);
nor U852 (N_852,N_795,N_729);
nor U853 (N_853,N_716,N_626);
nand U854 (N_854,N_794,N_646);
xnor U855 (N_855,N_737,N_708);
xor U856 (N_856,N_696,N_673);
and U857 (N_857,N_717,N_647);
xnor U858 (N_858,N_654,N_664);
xnor U859 (N_859,N_669,N_701);
nand U860 (N_860,N_747,N_757);
and U861 (N_861,N_640,N_736);
nand U862 (N_862,N_677,N_787);
and U863 (N_863,N_766,N_661);
nor U864 (N_864,N_618,N_621);
and U865 (N_865,N_785,N_613);
nand U866 (N_866,N_704,N_644);
xor U867 (N_867,N_733,N_614);
or U868 (N_868,N_674,N_602);
xnor U869 (N_869,N_741,N_695);
or U870 (N_870,N_608,N_656);
or U871 (N_871,N_760,N_684);
or U872 (N_872,N_670,N_601);
or U873 (N_873,N_775,N_713);
nand U874 (N_874,N_682,N_746);
or U875 (N_875,N_650,N_681);
xor U876 (N_876,N_796,N_648);
nand U877 (N_877,N_761,N_600);
nor U878 (N_878,N_762,N_611);
nand U879 (N_879,N_630,N_783);
nor U880 (N_880,N_792,N_660);
xnor U881 (N_881,N_718,N_649);
xor U882 (N_882,N_725,N_769);
nand U883 (N_883,N_705,N_615);
nor U884 (N_884,N_629,N_793);
nand U885 (N_885,N_620,N_782);
nor U886 (N_886,N_690,N_715);
xor U887 (N_887,N_791,N_742);
nor U888 (N_888,N_728,N_750);
xor U889 (N_889,N_605,N_666);
and U890 (N_890,N_711,N_663);
or U891 (N_891,N_700,N_624);
nand U892 (N_892,N_719,N_739);
nand U893 (N_893,N_735,N_668);
nand U894 (N_894,N_632,N_688);
or U895 (N_895,N_676,N_603);
and U896 (N_896,N_662,N_643);
xnor U897 (N_897,N_788,N_657);
xor U898 (N_898,N_675,N_745);
nand U899 (N_899,N_703,N_756);
xnor U900 (N_900,N_762,N_694);
or U901 (N_901,N_621,N_654);
and U902 (N_902,N_791,N_776);
and U903 (N_903,N_753,N_606);
and U904 (N_904,N_757,N_671);
or U905 (N_905,N_785,N_643);
xnor U906 (N_906,N_716,N_622);
nand U907 (N_907,N_756,N_761);
and U908 (N_908,N_692,N_649);
and U909 (N_909,N_618,N_629);
or U910 (N_910,N_712,N_646);
xor U911 (N_911,N_670,N_660);
nor U912 (N_912,N_650,N_765);
and U913 (N_913,N_710,N_714);
nor U914 (N_914,N_748,N_791);
or U915 (N_915,N_686,N_784);
and U916 (N_916,N_648,N_605);
nand U917 (N_917,N_633,N_696);
or U918 (N_918,N_731,N_769);
nor U919 (N_919,N_627,N_787);
or U920 (N_920,N_707,N_779);
nor U921 (N_921,N_630,N_653);
and U922 (N_922,N_780,N_718);
xor U923 (N_923,N_618,N_714);
nor U924 (N_924,N_698,N_784);
nand U925 (N_925,N_760,N_793);
xor U926 (N_926,N_782,N_601);
xnor U927 (N_927,N_708,N_752);
and U928 (N_928,N_647,N_658);
nand U929 (N_929,N_700,N_762);
nor U930 (N_930,N_755,N_725);
nor U931 (N_931,N_716,N_627);
nor U932 (N_932,N_790,N_669);
or U933 (N_933,N_724,N_606);
nand U934 (N_934,N_698,N_791);
and U935 (N_935,N_648,N_677);
and U936 (N_936,N_765,N_694);
or U937 (N_937,N_704,N_639);
nor U938 (N_938,N_722,N_613);
or U939 (N_939,N_741,N_715);
or U940 (N_940,N_653,N_762);
or U941 (N_941,N_693,N_635);
and U942 (N_942,N_706,N_721);
nand U943 (N_943,N_765,N_674);
xor U944 (N_944,N_799,N_747);
and U945 (N_945,N_610,N_674);
xor U946 (N_946,N_708,N_689);
and U947 (N_947,N_789,N_643);
nor U948 (N_948,N_760,N_634);
xor U949 (N_949,N_787,N_600);
and U950 (N_950,N_687,N_718);
xor U951 (N_951,N_642,N_731);
nor U952 (N_952,N_734,N_617);
nand U953 (N_953,N_650,N_791);
or U954 (N_954,N_762,N_663);
nor U955 (N_955,N_659,N_622);
nand U956 (N_956,N_743,N_790);
and U957 (N_957,N_736,N_676);
nand U958 (N_958,N_725,N_742);
and U959 (N_959,N_751,N_601);
or U960 (N_960,N_646,N_736);
nor U961 (N_961,N_683,N_701);
nand U962 (N_962,N_621,N_652);
nor U963 (N_963,N_662,N_756);
xor U964 (N_964,N_700,N_638);
xnor U965 (N_965,N_731,N_775);
nor U966 (N_966,N_602,N_777);
or U967 (N_967,N_711,N_791);
and U968 (N_968,N_752,N_700);
and U969 (N_969,N_796,N_697);
nand U970 (N_970,N_668,N_673);
xor U971 (N_971,N_657,N_713);
nor U972 (N_972,N_724,N_668);
nand U973 (N_973,N_799,N_647);
nor U974 (N_974,N_727,N_612);
nand U975 (N_975,N_781,N_690);
or U976 (N_976,N_643,N_758);
and U977 (N_977,N_627,N_794);
and U978 (N_978,N_734,N_678);
nor U979 (N_979,N_621,N_689);
or U980 (N_980,N_635,N_761);
and U981 (N_981,N_781,N_642);
nor U982 (N_982,N_619,N_702);
or U983 (N_983,N_741,N_671);
and U984 (N_984,N_663,N_695);
and U985 (N_985,N_605,N_698);
nand U986 (N_986,N_656,N_767);
xnor U987 (N_987,N_644,N_739);
nand U988 (N_988,N_689,N_616);
and U989 (N_989,N_740,N_650);
or U990 (N_990,N_727,N_797);
nand U991 (N_991,N_678,N_783);
and U992 (N_992,N_679,N_706);
or U993 (N_993,N_798,N_776);
and U994 (N_994,N_736,N_719);
nand U995 (N_995,N_653,N_664);
xor U996 (N_996,N_667,N_793);
xor U997 (N_997,N_776,N_631);
and U998 (N_998,N_613,N_696);
and U999 (N_999,N_671,N_679);
nand U1000 (N_1000,N_854,N_987);
or U1001 (N_1001,N_984,N_909);
nand U1002 (N_1002,N_800,N_975);
and U1003 (N_1003,N_934,N_836);
nand U1004 (N_1004,N_940,N_872);
or U1005 (N_1005,N_873,N_811);
xnor U1006 (N_1006,N_885,N_847);
xnor U1007 (N_1007,N_851,N_804);
xor U1008 (N_1008,N_979,N_924);
and U1009 (N_1009,N_818,N_995);
or U1010 (N_1010,N_939,N_802);
and U1011 (N_1011,N_982,N_961);
or U1012 (N_1012,N_805,N_861);
xor U1013 (N_1013,N_834,N_897);
or U1014 (N_1014,N_911,N_892);
and U1015 (N_1015,N_853,N_833);
nor U1016 (N_1016,N_823,N_910);
nor U1017 (N_1017,N_827,N_916);
and U1018 (N_1018,N_843,N_868);
and U1019 (N_1019,N_822,N_908);
xnor U1020 (N_1020,N_947,N_957);
nand U1021 (N_1021,N_922,N_944);
nand U1022 (N_1022,N_881,N_876);
nand U1023 (N_1023,N_973,N_849);
nor U1024 (N_1024,N_869,N_878);
nor U1025 (N_1025,N_978,N_974);
nand U1026 (N_1026,N_866,N_801);
or U1027 (N_1027,N_965,N_955);
xnor U1028 (N_1028,N_862,N_942);
nand U1029 (N_1029,N_859,N_882);
or U1030 (N_1030,N_956,N_980);
xnor U1031 (N_1031,N_929,N_837);
and U1032 (N_1032,N_863,N_923);
nor U1033 (N_1033,N_994,N_893);
nor U1034 (N_1034,N_831,N_858);
nor U1035 (N_1035,N_913,N_846);
nand U1036 (N_1036,N_814,N_932);
or U1037 (N_1037,N_951,N_945);
and U1038 (N_1038,N_954,N_865);
nor U1039 (N_1039,N_819,N_884);
xor U1040 (N_1040,N_890,N_825);
nand U1041 (N_1041,N_920,N_960);
nor U1042 (N_1042,N_894,N_915);
xor U1043 (N_1043,N_842,N_998);
and U1044 (N_1044,N_952,N_966);
xnor U1045 (N_1045,N_983,N_815);
and U1046 (N_1046,N_864,N_953);
or U1047 (N_1047,N_935,N_826);
xnor U1048 (N_1048,N_990,N_900);
nand U1049 (N_1049,N_883,N_963);
and U1050 (N_1050,N_964,N_852);
nor U1051 (N_1051,N_879,N_810);
nand U1052 (N_1052,N_970,N_928);
and U1053 (N_1053,N_898,N_968);
nand U1054 (N_1054,N_938,N_976);
and U1055 (N_1055,N_830,N_871);
or U1056 (N_1056,N_848,N_835);
nand U1057 (N_1057,N_850,N_941);
and U1058 (N_1058,N_971,N_914);
nand U1059 (N_1059,N_905,N_997);
nand U1060 (N_1060,N_839,N_989);
nand U1061 (N_1061,N_959,N_886);
nand U1062 (N_1062,N_840,N_902);
nor U1063 (N_1063,N_903,N_933);
xnor U1064 (N_1064,N_917,N_889);
xor U1065 (N_1065,N_808,N_930);
nand U1066 (N_1066,N_949,N_918);
nand U1067 (N_1067,N_860,N_829);
or U1068 (N_1068,N_943,N_999);
or U1069 (N_1069,N_907,N_996);
and U1070 (N_1070,N_950,N_906);
nand U1071 (N_1071,N_888,N_946);
xor U1072 (N_1072,N_832,N_958);
nor U1073 (N_1073,N_972,N_856);
nor U1074 (N_1074,N_967,N_919);
nand U1075 (N_1075,N_936,N_981);
and U1076 (N_1076,N_838,N_845);
xor U1077 (N_1077,N_896,N_912);
nor U1078 (N_1078,N_986,N_991);
nor U1079 (N_1079,N_841,N_844);
nor U1080 (N_1080,N_874,N_817);
nand U1081 (N_1081,N_867,N_812);
xor U1082 (N_1082,N_895,N_937);
or U1083 (N_1083,N_985,N_969);
and U1084 (N_1084,N_931,N_948);
and U1085 (N_1085,N_988,N_821);
nor U1086 (N_1086,N_803,N_824);
xor U1087 (N_1087,N_901,N_870);
xor U1088 (N_1088,N_925,N_899);
nand U1089 (N_1089,N_809,N_877);
or U1090 (N_1090,N_816,N_880);
and U1091 (N_1091,N_887,N_904);
nor U1092 (N_1092,N_813,N_806);
or U1093 (N_1093,N_857,N_962);
and U1094 (N_1094,N_807,N_828);
nor U1095 (N_1095,N_977,N_855);
and U1096 (N_1096,N_927,N_875);
nand U1097 (N_1097,N_820,N_992);
xnor U1098 (N_1098,N_926,N_921);
xnor U1099 (N_1099,N_993,N_891);
nor U1100 (N_1100,N_887,N_957);
and U1101 (N_1101,N_921,N_844);
xor U1102 (N_1102,N_991,N_973);
and U1103 (N_1103,N_856,N_921);
xnor U1104 (N_1104,N_949,N_823);
nand U1105 (N_1105,N_943,N_957);
nor U1106 (N_1106,N_837,N_823);
nor U1107 (N_1107,N_871,N_926);
and U1108 (N_1108,N_888,N_972);
xor U1109 (N_1109,N_921,N_987);
nand U1110 (N_1110,N_906,N_863);
nand U1111 (N_1111,N_965,N_859);
nor U1112 (N_1112,N_849,N_952);
nand U1113 (N_1113,N_928,N_978);
xnor U1114 (N_1114,N_840,N_909);
or U1115 (N_1115,N_900,N_915);
and U1116 (N_1116,N_977,N_976);
and U1117 (N_1117,N_890,N_826);
or U1118 (N_1118,N_925,N_877);
xor U1119 (N_1119,N_859,N_983);
nor U1120 (N_1120,N_930,N_962);
or U1121 (N_1121,N_993,N_871);
and U1122 (N_1122,N_929,N_919);
and U1123 (N_1123,N_919,N_811);
and U1124 (N_1124,N_939,N_838);
and U1125 (N_1125,N_990,N_932);
nand U1126 (N_1126,N_806,N_987);
and U1127 (N_1127,N_884,N_980);
or U1128 (N_1128,N_888,N_843);
nand U1129 (N_1129,N_946,N_992);
xor U1130 (N_1130,N_990,N_903);
or U1131 (N_1131,N_870,N_814);
xnor U1132 (N_1132,N_848,N_982);
nor U1133 (N_1133,N_979,N_922);
or U1134 (N_1134,N_949,N_914);
nand U1135 (N_1135,N_857,N_977);
nor U1136 (N_1136,N_813,N_947);
and U1137 (N_1137,N_944,N_896);
and U1138 (N_1138,N_901,N_970);
xor U1139 (N_1139,N_906,N_959);
and U1140 (N_1140,N_802,N_892);
nor U1141 (N_1141,N_942,N_816);
and U1142 (N_1142,N_911,N_900);
and U1143 (N_1143,N_807,N_883);
xnor U1144 (N_1144,N_998,N_800);
and U1145 (N_1145,N_846,N_995);
xnor U1146 (N_1146,N_921,N_885);
nor U1147 (N_1147,N_869,N_972);
or U1148 (N_1148,N_928,N_965);
or U1149 (N_1149,N_919,N_996);
or U1150 (N_1150,N_941,N_834);
nor U1151 (N_1151,N_858,N_847);
nor U1152 (N_1152,N_821,N_945);
nor U1153 (N_1153,N_934,N_971);
nor U1154 (N_1154,N_820,N_846);
or U1155 (N_1155,N_997,N_948);
nor U1156 (N_1156,N_899,N_956);
nand U1157 (N_1157,N_980,N_972);
or U1158 (N_1158,N_883,N_929);
nand U1159 (N_1159,N_899,N_886);
or U1160 (N_1160,N_927,N_967);
or U1161 (N_1161,N_876,N_974);
xor U1162 (N_1162,N_980,N_886);
nand U1163 (N_1163,N_902,N_963);
and U1164 (N_1164,N_982,N_932);
and U1165 (N_1165,N_966,N_867);
nand U1166 (N_1166,N_895,N_813);
nand U1167 (N_1167,N_993,N_872);
and U1168 (N_1168,N_810,N_979);
or U1169 (N_1169,N_990,N_872);
nand U1170 (N_1170,N_920,N_939);
and U1171 (N_1171,N_933,N_810);
nor U1172 (N_1172,N_961,N_866);
nor U1173 (N_1173,N_837,N_824);
nand U1174 (N_1174,N_987,N_932);
nand U1175 (N_1175,N_973,N_917);
nand U1176 (N_1176,N_941,N_983);
and U1177 (N_1177,N_885,N_932);
nor U1178 (N_1178,N_871,N_880);
nor U1179 (N_1179,N_830,N_850);
and U1180 (N_1180,N_946,N_877);
xor U1181 (N_1181,N_911,N_852);
or U1182 (N_1182,N_897,N_901);
and U1183 (N_1183,N_829,N_954);
xnor U1184 (N_1184,N_804,N_854);
xnor U1185 (N_1185,N_802,N_991);
and U1186 (N_1186,N_833,N_900);
and U1187 (N_1187,N_963,N_956);
and U1188 (N_1188,N_938,N_837);
and U1189 (N_1189,N_801,N_804);
nand U1190 (N_1190,N_987,N_976);
xor U1191 (N_1191,N_877,N_943);
nand U1192 (N_1192,N_958,N_809);
nand U1193 (N_1193,N_806,N_852);
nor U1194 (N_1194,N_805,N_802);
or U1195 (N_1195,N_938,N_974);
or U1196 (N_1196,N_867,N_945);
and U1197 (N_1197,N_865,N_887);
nand U1198 (N_1198,N_962,N_861);
nand U1199 (N_1199,N_968,N_821);
nand U1200 (N_1200,N_1067,N_1009);
xor U1201 (N_1201,N_1141,N_1037);
or U1202 (N_1202,N_1072,N_1137);
nand U1203 (N_1203,N_1020,N_1046);
xnor U1204 (N_1204,N_1051,N_1171);
xor U1205 (N_1205,N_1085,N_1138);
nor U1206 (N_1206,N_1173,N_1021);
and U1207 (N_1207,N_1157,N_1189);
or U1208 (N_1208,N_1101,N_1090);
nand U1209 (N_1209,N_1008,N_1047);
and U1210 (N_1210,N_1055,N_1011);
xor U1211 (N_1211,N_1073,N_1110);
nand U1212 (N_1212,N_1103,N_1054);
or U1213 (N_1213,N_1043,N_1148);
xnor U1214 (N_1214,N_1019,N_1163);
and U1215 (N_1215,N_1109,N_1078);
and U1216 (N_1216,N_1079,N_1015);
and U1217 (N_1217,N_1113,N_1169);
xnor U1218 (N_1218,N_1188,N_1036);
nor U1219 (N_1219,N_1121,N_1029);
and U1220 (N_1220,N_1147,N_1197);
or U1221 (N_1221,N_1187,N_1108);
nor U1222 (N_1222,N_1002,N_1177);
or U1223 (N_1223,N_1026,N_1151);
and U1224 (N_1224,N_1013,N_1125);
nor U1225 (N_1225,N_1032,N_1003);
or U1226 (N_1226,N_1070,N_1166);
nor U1227 (N_1227,N_1153,N_1099);
nand U1228 (N_1228,N_1024,N_1144);
or U1229 (N_1229,N_1028,N_1058);
and U1230 (N_1230,N_1066,N_1164);
nand U1231 (N_1231,N_1034,N_1194);
nand U1232 (N_1232,N_1087,N_1143);
or U1233 (N_1233,N_1042,N_1154);
nor U1234 (N_1234,N_1084,N_1118);
nand U1235 (N_1235,N_1033,N_1035);
xor U1236 (N_1236,N_1074,N_1105);
nor U1237 (N_1237,N_1162,N_1077);
and U1238 (N_1238,N_1129,N_1114);
nand U1239 (N_1239,N_1007,N_1132);
xnor U1240 (N_1240,N_1191,N_1175);
or U1241 (N_1241,N_1061,N_1181);
or U1242 (N_1242,N_1117,N_1075);
nand U1243 (N_1243,N_1041,N_1119);
xnor U1244 (N_1244,N_1112,N_1089);
nand U1245 (N_1245,N_1102,N_1111);
and U1246 (N_1246,N_1196,N_1053);
and U1247 (N_1247,N_1165,N_1150);
or U1248 (N_1248,N_1180,N_1185);
and U1249 (N_1249,N_1128,N_1023);
or U1250 (N_1250,N_1134,N_1104);
nor U1251 (N_1251,N_1081,N_1178);
and U1252 (N_1252,N_1159,N_1062);
xor U1253 (N_1253,N_1063,N_1065);
nand U1254 (N_1254,N_1155,N_1017);
nand U1255 (N_1255,N_1006,N_1038);
and U1256 (N_1256,N_1176,N_1198);
and U1257 (N_1257,N_1136,N_1146);
and U1258 (N_1258,N_1004,N_1122);
nor U1259 (N_1259,N_1131,N_1071);
or U1260 (N_1260,N_1027,N_1001);
and U1261 (N_1261,N_1091,N_1167);
nand U1262 (N_1262,N_1127,N_1082);
xnor U1263 (N_1263,N_1096,N_1039);
nand U1264 (N_1264,N_1133,N_1098);
xor U1265 (N_1265,N_1135,N_1040);
xor U1266 (N_1266,N_1184,N_1179);
xor U1267 (N_1267,N_1064,N_1161);
nor U1268 (N_1268,N_1022,N_1048);
and U1269 (N_1269,N_1130,N_1076);
or U1270 (N_1270,N_1142,N_1192);
and U1271 (N_1271,N_1156,N_1140);
and U1272 (N_1272,N_1195,N_1095);
and U1273 (N_1273,N_1083,N_1107);
xor U1274 (N_1274,N_1050,N_1031);
xor U1275 (N_1275,N_1094,N_1174);
or U1276 (N_1276,N_1049,N_1193);
nor U1277 (N_1277,N_1116,N_1152);
xor U1278 (N_1278,N_1052,N_1186);
or U1279 (N_1279,N_1160,N_1059);
and U1280 (N_1280,N_1030,N_1123);
xor U1281 (N_1281,N_1000,N_1018);
nor U1282 (N_1282,N_1126,N_1182);
or U1283 (N_1283,N_1080,N_1005);
nand U1284 (N_1284,N_1045,N_1158);
nand U1285 (N_1285,N_1100,N_1106);
xnor U1286 (N_1286,N_1149,N_1139);
or U1287 (N_1287,N_1057,N_1088);
nor U1288 (N_1288,N_1172,N_1115);
nand U1289 (N_1289,N_1093,N_1199);
nor U1290 (N_1290,N_1120,N_1016);
nor U1291 (N_1291,N_1124,N_1170);
nand U1292 (N_1292,N_1097,N_1183);
or U1293 (N_1293,N_1060,N_1044);
nand U1294 (N_1294,N_1012,N_1014);
nand U1295 (N_1295,N_1068,N_1069);
nor U1296 (N_1296,N_1056,N_1190);
and U1297 (N_1297,N_1025,N_1145);
xnor U1298 (N_1298,N_1168,N_1010);
or U1299 (N_1299,N_1092,N_1086);
and U1300 (N_1300,N_1094,N_1044);
nand U1301 (N_1301,N_1164,N_1006);
xnor U1302 (N_1302,N_1142,N_1143);
xor U1303 (N_1303,N_1032,N_1006);
nand U1304 (N_1304,N_1137,N_1107);
or U1305 (N_1305,N_1003,N_1072);
xor U1306 (N_1306,N_1111,N_1109);
nor U1307 (N_1307,N_1124,N_1015);
xnor U1308 (N_1308,N_1055,N_1072);
or U1309 (N_1309,N_1023,N_1178);
nor U1310 (N_1310,N_1100,N_1165);
or U1311 (N_1311,N_1069,N_1008);
or U1312 (N_1312,N_1001,N_1089);
and U1313 (N_1313,N_1130,N_1007);
nand U1314 (N_1314,N_1101,N_1003);
nor U1315 (N_1315,N_1182,N_1005);
nor U1316 (N_1316,N_1002,N_1091);
nor U1317 (N_1317,N_1197,N_1112);
and U1318 (N_1318,N_1161,N_1058);
nand U1319 (N_1319,N_1072,N_1040);
and U1320 (N_1320,N_1010,N_1179);
nand U1321 (N_1321,N_1116,N_1076);
nand U1322 (N_1322,N_1147,N_1026);
nor U1323 (N_1323,N_1039,N_1042);
and U1324 (N_1324,N_1096,N_1132);
or U1325 (N_1325,N_1085,N_1087);
xnor U1326 (N_1326,N_1157,N_1003);
nand U1327 (N_1327,N_1177,N_1166);
nand U1328 (N_1328,N_1146,N_1079);
nand U1329 (N_1329,N_1132,N_1072);
xor U1330 (N_1330,N_1039,N_1098);
and U1331 (N_1331,N_1135,N_1193);
xor U1332 (N_1332,N_1149,N_1039);
xor U1333 (N_1333,N_1008,N_1048);
or U1334 (N_1334,N_1145,N_1190);
nand U1335 (N_1335,N_1198,N_1022);
nor U1336 (N_1336,N_1050,N_1090);
xnor U1337 (N_1337,N_1130,N_1148);
nand U1338 (N_1338,N_1025,N_1028);
or U1339 (N_1339,N_1118,N_1074);
nand U1340 (N_1340,N_1144,N_1034);
nand U1341 (N_1341,N_1174,N_1153);
or U1342 (N_1342,N_1059,N_1002);
xor U1343 (N_1343,N_1137,N_1038);
or U1344 (N_1344,N_1006,N_1119);
and U1345 (N_1345,N_1060,N_1186);
or U1346 (N_1346,N_1156,N_1090);
nand U1347 (N_1347,N_1123,N_1067);
nor U1348 (N_1348,N_1019,N_1199);
nor U1349 (N_1349,N_1000,N_1062);
or U1350 (N_1350,N_1120,N_1085);
xnor U1351 (N_1351,N_1114,N_1023);
or U1352 (N_1352,N_1018,N_1050);
nand U1353 (N_1353,N_1132,N_1102);
and U1354 (N_1354,N_1043,N_1161);
nor U1355 (N_1355,N_1165,N_1020);
or U1356 (N_1356,N_1193,N_1059);
nor U1357 (N_1357,N_1138,N_1173);
nor U1358 (N_1358,N_1037,N_1000);
and U1359 (N_1359,N_1136,N_1009);
xnor U1360 (N_1360,N_1193,N_1027);
nor U1361 (N_1361,N_1145,N_1051);
nor U1362 (N_1362,N_1184,N_1120);
nor U1363 (N_1363,N_1065,N_1194);
nand U1364 (N_1364,N_1011,N_1005);
nand U1365 (N_1365,N_1018,N_1023);
xor U1366 (N_1366,N_1000,N_1133);
xnor U1367 (N_1367,N_1000,N_1088);
and U1368 (N_1368,N_1182,N_1089);
xor U1369 (N_1369,N_1073,N_1054);
nand U1370 (N_1370,N_1010,N_1046);
xor U1371 (N_1371,N_1171,N_1121);
nand U1372 (N_1372,N_1144,N_1110);
nor U1373 (N_1373,N_1056,N_1055);
and U1374 (N_1374,N_1073,N_1079);
xnor U1375 (N_1375,N_1160,N_1134);
nand U1376 (N_1376,N_1000,N_1058);
nor U1377 (N_1377,N_1145,N_1171);
xor U1378 (N_1378,N_1172,N_1067);
or U1379 (N_1379,N_1064,N_1184);
nand U1380 (N_1380,N_1132,N_1014);
nand U1381 (N_1381,N_1163,N_1127);
and U1382 (N_1382,N_1058,N_1151);
and U1383 (N_1383,N_1191,N_1180);
xnor U1384 (N_1384,N_1055,N_1171);
nor U1385 (N_1385,N_1019,N_1116);
nand U1386 (N_1386,N_1084,N_1100);
nand U1387 (N_1387,N_1145,N_1111);
nor U1388 (N_1388,N_1103,N_1097);
xor U1389 (N_1389,N_1004,N_1042);
and U1390 (N_1390,N_1195,N_1116);
xor U1391 (N_1391,N_1190,N_1194);
nand U1392 (N_1392,N_1062,N_1164);
nor U1393 (N_1393,N_1014,N_1006);
nor U1394 (N_1394,N_1087,N_1124);
or U1395 (N_1395,N_1130,N_1093);
nand U1396 (N_1396,N_1131,N_1015);
or U1397 (N_1397,N_1057,N_1140);
nand U1398 (N_1398,N_1022,N_1096);
or U1399 (N_1399,N_1051,N_1097);
nor U1400 (N_1400,N_1264,N_1297);
or U1401 (N_1401,N_1273,N_1373);
and U1402 (N_1402,N_1222,N_1368);
and U1403 (N_1403,N_1309,N_1259);
nor U1404 (N_1404,N_1200,N_1208);
xor U1405 (N_1405,N_1382,N_1263);
or U1406 (N_1406,N_1251,N_1293);
nand U1407 (N_1407,N_1262,N_1385);
nor U1408 (N_1408,N_1355,N_1363);
nor U1409 (N_1409,N_1324,N_1244);
nor U1410 (N_1410,N_1289,N_1321);
nor U1411 (N_1411,N_1322,N_1336);
nor U1412 (N_1412,N_1284,N_1371);
or U1413 (N_1413,N_1234,N_1299);
or U1414 (N_1414,N_1215,N_1378);
nand U1415 (N_1415,N_1316,N_1246);
or U1416 (N_1416,N_1218,N_1384);
and U1417 (N_1417,N_1361,N_1372);
nor U1418 (N_1418,N_1365,N_1317);
xor U1419 (N_1419,N_1353,N_1364);
nand U1420 (N_1420,N_1216,N_1390);
xor U1421 (N_1421,N_1279,N_1315);
and U1422 (N_1422,N_1210,N_1287);
xnor U1423 (N_1423,N_1277,N_1255);
or U1424 (N_1424,N_1313,N_1204);
or U1425 (N_1425,N_1359,N_1338);
and U1426 (N_1426,N_1312,N_1270);
or U1427 (N_1427,N_1213,N_1349);
xor U1428 (N_1428,N_1254,N_1394);
xnor U1429 (N_1429,N_1351,N_1203);
xor U1430 (N_1430,N_1265,N_1374);
and U1431 (N_1431,N_1212,N_1228);
xor U1432 (N_1432,N_1221,N_1250);
nor U1433 (N_1433,N_1360,N_1340);
and U1434 (N_1434,N_1295,N_1240);
or U1435 (N_1435,N_1326,N_1375);
and U1436 (N_1436,N_1387,N_1268);
nand U1437 (N_1437,N_1343,N_1391);
or U1438 (N_1438,N_1288,N_1386);
or U1439 (N_1439,N_1245,N_1337);
and U1440 (N_1440,N_1260,N_1211);
nor U1441 (N_1441,N_1292,N_1307);
or U1442 (N_1442,N_1381,N_1318);
xor U1443 (N_1443,N_1267,N_1226);
nor U1444 (N_1444,N_1370,N_1231);
and U1445 (N_1445,N_1329,N_1223);
nor U1446 (N_1446,N_1306,N_1206);
xor U1447 (N_1447,N_1207,N_1201);
or U1448 (N_1448,N_1333,N_1367);
nor U1449 (N_1449,N_1271,N_1300);
or U1450 (N_1450,N_1393,N_1369);
nand U1451 (N_1451,N_1323,N_1352);
or U1452 (N_1452,N_1274,N_1238);
nand U1453 (N_1453,N_1296,N_1357);
and U1454 (N_1454,N_1217,N_1236);
or U1455 (N_1455,N_1302,N_1269);
xor U1456 (N_1456,N_1311,N_1278);
xnor U1457 (N_1457,N_1304,N_1258);
or U1458 (N_1458,N_1358,N_1275);
or U1459 (N_1459,N_1332,N_1227);
or U1460 (N_1460,N_1339,N_1319);
nand U1461 (N_1461,N_1376,N_1243);
nand U1462 (N_1462,N_1314,N_1354);
xnor U1463 (N_1463,N_1272,N_1350);
nand U1464 (N_1464,N_1392,N_1341);
and U1465 (N_1465,N_1253,N_1248);
nand U1466 (N_1466,N_1256,N_1230);
and U1467 (N_1467,N_1325,N_1396);
nor U1468 (N_1468,N_1291,N_1280);
xnor U1469 (N_1469,N_1219,N_1366);
nor U1470 (N_1470,N_1335,N_1282);
or U1471 (N_1471,N_1290,N_1225);
nand U1472 (N_1472,N_1383,N_1249);
and U1473 (N_1473,N_1362,N_1379);
and U1474 (N_1474,N_1389,N_1239);
and U1475 (N_1475,N_1202,N_1345);
and U1476 (N_1476,N_1346,N_1214);
nor U1477 (N_1477,N_1235,N_1397);
and U1478 (N_1478,N_1294,N_1233);
or U1479 (N_1479,N_1310,N_1220);
nor U1480 (N_1480,N_1266,N_1320);
xnor U1481 (N_1481,N_1257,N_1308);
nor U1482 (N_1482,N_1348,N_1347);
or U1483 (N_1483,N_1388,N_1229);
nor U1484 (N_1484,N_1330,N_1224);
xor U1485 (N_1485,N_1285,N_1237);
or U1486 (N_1486,N_1303,N_1344);
nor U1487 (N_1487,N_1298,N_1398);
xor U1488 (N_1488,N_1380,N_1305);
nor U1489 (N_1489,N_1241,N_1209);
or U1490 (N_1490,N_1276,N_1328);
and U1491 (N_1491,N_1395,N_1286);
nand U1492 (N_1492,N_1242,N_1301);
and U1493 (N_1493,N_1247,N_1252);
xnor U1494 (N_1494,N_1399,N_1205);
xnor U1495 (N_1495,N_1261,N_1356);
nor U1496 (N_1496,N_1377,N_1327);
nand U1497 (N_1497,N_1331,N_1283);
or U1498 (N_1498,N_1232,N_1342);
nor U1499 (N_1499,N_1281,N_1334);
nand U1500 (N_1500,N_1369,N_1365);
and U1501 (N_1501,N_1387,N_1330);
xor U1502 (N_1502,N_1276,N_1312);
nor U1503 (N_1503,N_1324,N_1335);
xnor U1504 (N_1504,N_1220,N_1267);
nand U1505 (N_1505,N_1359,N_1221);
and U1506 (N_1506,N_1287,N_1281);
nand U1507 (N_1507,N_1202,N_1311);
xor U1508 (N_1508,N_1217,N_1357);
and U1509 (N_1509,N_1303,N_1208);
nor U1510 (N_1510,N_1375,N_1264);
and U1511 (N_1511,N_1379,N_1334);
or U1512 (N_1512,N_1266,N_1241);
or U1513 (N_1513,N_1385,N_1209);
and U1514 (N_1514,N_1207,N_1345);
or U1515 (N_1515,N_1240,N_1321);
nor U1516 (N_1516,N_1358,N_1264);
nor U1517 (N_1517,N_1271,N_1252);
xor U1518 (N_1518,N_1351,N_1329);
or U1519 (N_1519,N_1394,N_1304);
and U1520 (N_1520,N_1276,N_1351);
or U1521 (N_1521,N_1214,N_1349);
nand U1522 (N_1522,N_1357,N_1343);
xnor U1523 (N_1523,N_1390,N_1214);
xnor U1524 (N_1524,N_1368,N_1326);
nand U1525 (N_1525,N_1380,N_1343);
xnor U1526 (N_1526,N_1256,N_1314);
xor U1527 (N_1527,N_1247,N_1329);
or U1528 (N_1528,N_1330,N_1351);
and U1529 (N_1529,N_1236,N_1392);
nand U1530 (N_1530,N_1252,N_1378);
or U1531 (N_1531,N_1292,N_1336);
nand U1532 (N_1532,N_1260,N_1352);
nor U1533 (N_1533,N_1259,N_1206);
xnor U1534 (N_1534,N_1211,N_1275);
nor U1535 (N_1535,N_1351,N_1224);
nand U1536 (N_1536,N_1266,N_1291);
xnor U1537 (N_1537,N_1298,N_1227);
nor U1538 (N_1538,N_1204,N_1231);
xnor U1539 (N_1539,N_1359,N_1330);
and U1540 (N_1540,N_1236,N_1208);
nor U1541 (N_1541,N_1331,N_1372);
xor U1542 (N_1542,N_1258,N_1260);
nand U1543 (N_1543,N_1356,N_1311);
or U1544 (N_1544,N_1311,N_1352);
nand U1545 (N_1545,N_1260,N_1360);
and U1546 (N_1546,N_1246,N_1213);
or U1547 (N_1547,N_1370,N_1222);
nor U1548 (N_1548,N_1287,N_1248);
xor U1549 (N_1549,N_1251,N_1349);
nand U1550 (N_1550,N_1344,N_1371);
or U1551 (N_1551,N_1300,N_1287);
nor U1552 (N_1552,N_1269,N_1287);
xnor U1553 (N_1553,N_1217,N_1200);
nor U1554 (N_1554,N_1299,N_1295);
xnor U1555 (N_1555,N_1304,N_1243);
nand U1556 (N_1556,N_1304,N_1308);
nor U1557 (N_1557,N_1239,N_1326);
or U1558 (N_1558,N_1245,N_1280);
nor U1559 (N_1559,N_1270,N_1367);
xnor U1560 (N_1560,N_1381,N_1379);
and U1561 (N_1561,N_1390,N_1230);
or U1562 (N_1562,N_1208,N_1355);
nor U1563 (N_1563,N_1201,N_1292);
and U1564 (N_1564,N_1397,N_1203);
or U1565 (N_1565,N_1331,N_1337);
or U1566 (N_1566,N_1239,N_1365);
nand U1567 (N_1567,N_1222,N_1226);
and U1568 (N_1568,N_1259,N_1253);
nand U1569 (N_1569,N_1235,N_1228);
nor U1570 (N_1570,N_1222,N_1318);
and U1571 (N_1571,N_1330,N_1274);
or U1572 (N_1572,N_1347,N_1231);
nand U1573 (N_1573,N_1392,N_1208);
and U1574 (N_1574,N_1353,N_1228);
nor U1575 (N_1575,N_1366,N_1333);
and U1576 (N_1576,N_1285,N_1281);
and U1577 (N_1577,N_1252,N_1219);
nor U1578 (N_1578,N_1292,N_1355);
xnor U1579 (N_1579,N_1272,N_1241);
or U1580 (N_1580,N_1239,N_1385);
and U1581 (N_1581,N_1324,N_1371);
nand U1582 (N_1582,N_1221,N_1347);
nand U1583 (N_1583,N_1233,N_1247);
nor U1584 (N_1584,N_1201,N_1390);
xnor U1585 (N_1585,N_1357,N_1260);
xor U1586 (N_1586,N_1223,N_1353);
or U1587 (N_1587,N_1280,N_1307);
xnor U1588 (N_1588,N_1283,N_1221);
or U1589 (N_1589,N_1275,N_1383);
or U1590 (N_1590,N_1226,N_1275);
xnor U1591 (N_1591,N_1333,N_1314);
and U1592 (N_1592,N_1334,N_1319);
nor U1593 (N_1593,N_1334,N_1376);
nor U1594 (N_1594,N_1229,N_1397);
nor U1595 (N_1595,N_1203,N_1350);
nand U1596 (N_1596,N_1252,N_1295);
nand U1597 (N_1597,N_1356,N_1390);
nor U1598 (N_1598,N_1257,N_1232);
nand U1599 (N_1599,N_1313,N_1257);
and U1600 (N_1600,N_1423,N_1561);
nand U1601 (N_1601,N_1491,N_1574);
nor U1602 (N_1602,N_1540,N_1573);
xnor U1603 (N_1603,N_1509,N_1485);
nor U1604 (N_1604,N_1546,N_1437);
nor U1605 (N_1605,N_1487,N_1403);
or U1606 (N_1606,N_1468,N_1440);
nor U1607 (N_1607,N_1500,N_1590);
or U1608 (N_1608,N_1415,N_1518);
xor U1609 (N_1609,N_1476,N_1554);
xor U1610 (N_1610,N_1421,N_1410);
nor U1611 (N_1611,N_1532,N_1568);
and U1612 (N_1612,N_1585,N_1531);
xor U1613 (N_1613,N_1458,N_1427);
or U1614 (N_1614,N_1513,N_1482);
nand U1615 (N_1615,N_1588,N_1508);
xor U1616 (N_1616,N_1497,N_1582);
or U1617 (N_1617,N_1455,N_1489);
nor U1618 (N_1618,N_1412,N_1417);
nand U1619 (N_1619,N_1526,N_1443);
nor U1620 (N_1620,N_1511,N_1597);
nand U1621 (N_1621,N_1529,N_1569);
or U1622 (N_1622,N_1404,N_1406);
or U1623 (N_1623,N_1408,N_1555);
nor U1624 (N_1624,N_1436,N_1571);
or U1625 (N_1625,N_1547,N_1589);
and U1626 (N_1626,N_1549,N_1539);
or U1627 (N_1627,N_1467,N_1535);
and U1628 (N_1628,N_1504,N_1542);
nand U1629 (N_1629,N_1405,N_1472);
xnor U1630 (N_1630,N_1543,N_1557);
and U1631 (N_1631,N_1441,N_1591);
nand U1632 (N_1632,N_1495,N_1420);
nor U1633 (N_1633,N_1550,N_1515);
nor U1634 (N_1634,N_1502,N_1469);
nor U1635 (N_1635,N_1541,N_1435);
nand U1636 (N_1636,N_1537,N_1481);
and U1637 (N_1637,N_1488,N_1471);
nor U1638 (N_1638,N_1456,N_1570);
nor U1639 (N_1639,N_1560,N_1538);
nand U1640 (N_1640,N_1490,N_1466);
and U1641 (N_1641,N_1496,N_1521);
nand U1642 (N_1642,N_1516,N_1517);
nand U1643 (N_1643,N_1473,N_1401);
and U1644 (N_1644,N_1477,N_1510);
xor U1645 (N_1645,N_1434,N_1501);
nand U1646 (N_1646,N_1483,N_1586);
and U1647 (N_1647,N_1494,N_1565);
or U1648 (N_1648,N_1411,N_1407);
nor U1649 (N_1649,N_1583,N_1450);
or U1650 (N_1650,N_1463,N_1428);
xor U1651 (N_1651,N_1492,N_1593);
nand U1652 (N_1652,N_1442,N_1562);
nor U1653 (N_1653,N_1548,N_1594);
or U1654 (N_1654,N_1451,N_1556);
or U1655 (N_1655,N_1519,N_1584);
or U1656 (N_1656,N_1478,N_1544);
nor U1657 (N_1657,N_1457,N_1452);
xnor U1658 (N_1658,N_1567,N_1430);
and U1659 (N_1659,N_1553,N_1470);
nand U1660 (N_1660,N_1465,N_1413);
xnor U1661 (N_1661,N_1460,N_1576);
nor U1662 (N_1662,N_1425,N_1580);
nor U1663 (N_1663,N_1462,N_1429);
or U1664 (N_1664,N_1480,N_1464);
nor U1665 (N_1665,N_1559,N_1474);
nor U1666 (N_1666,N_1432,N_1524);
or U1667 (N_1667,N_1445,N_1577);
or U1668 (N_1668,N_1534,N_1479);
nor U1669 (N_1669,N_1447,N_1475);
nand U1670 (N_1670,N_1424,N_1505);
and U1671 (N_1671,N_1564,N_1461);
nor U1672 (N_1672,N_1545,N_1595);
and U1673 (N_1673,N_1431,N_1409);
or U1674 (N_1674,N_1506,N_1599);
nor U1675 (N_1675,N_1551,N_1575);
nor U1676 (N_1676,N_1438,N_1530);
xor U1677 (N_1677,N_1418,N_1528);
and U1678 (N_1678,N_1414,N_1454);
and U1679 (N_1679,N_1499,N_1433);
and U1680 (N_1680,N_1453,N_1444);
xor U1681 (N_1681,N_1572,N_1592);
and U1682 (N_1682,N_1449,N_1579);
nor U1683 (N_1683,N_1536,N_1422);
and U1684 (N_1684,N_1446,N_1566);
xnor U1685 (N_1685,N_1514,N_1426);
and U1686 (N_1686,N_1493,N_1507);
nor U1687 (N_1687,N_1527,N_1587);
and U1688 (N_1688,N_1448,N_1486);
nand U1689 (N_1689,N_1416,N_1484);
nand U1690 (N_1690,N_1596,N_1533);
and U1691 (N_1691,N_1512,N_1525);
nor U1692 (N_1692,N_1523,N_1552);
nor U1693 (N_1693,N_1439,N_1400);
xnor U1694 (N_1694,N_1503,N_1522);
nand U1695 (N_1695,N_1578,N_1498);
nand U1696 (N_1696,N_1402,N_1558);
or U1697 (N_1697,N_1598,N_1459);
nor U1698 (N_1698,N_1581,N_1563);
or U1699 (N_1699,N_1419,N_1520);
and U1700 (N_1700,N_1525,N_1402);
nor U1701 (N_1701,N_1514,N_1454);
nor U1702 (N_1702,N_1525,N_1442);
xnor U1703 (N_1703,N_1517,N_1593);
nor U1704 (N_1704,N_1402,N_1580);
nand U1705 (N_1705,N_1565,N_1514);
or U1706 (N_1706,N_1534,N_1451);
xnor U1707 (N_1707,N_1540,N_1570);
xor U1708 (N_1708,N_1562,N_1519);
or U1709 (N_1709,N_1431,N_1536);
and U1710 (N_1710,N_1431,N_1564);
nor U1711 (N_1711,N_1522,N_1565);
nand U1712 (N_1712,N_1432,N_1585);
and U1713 (N_1713,N_1515,N_1443);
and U1714 (N_1714,N_1592,N_1560);
and U1715 (N_1715,N_1467,N_1468);
or U1716 (N_1716,N_1519,N_1508);
nor U1717 (N_1717,N_1499,N_1494);
nand U1718 (N_1718,N_1428,N_1527);
or U1719 (N_1719,N_1596,N_1419);
nor U1720 (N_1720,N_1493,N_1531);
nand U1721 (N_1721,N_1595,N_1505);
xor U1722 (N_1722,N_1583,N_1500);
and U1723 (N_1723,N_1438,N_1419);
or U1724 (N_1724,N_1497,N_1537);
nor U1725 (N_1725,N_1589,N_1586);
nor U1726 (N_1726,N_1458,N_1461);
nor U1727 (N_1727,N_1510,N_1595);
and U1728 (N_1728,N_1523,N_1477);
and U1729 (N_1729,N_1414,N_1578);
nor U1730 (N_1730,N_1422,N_1453);
and U1731 (N_1731,N_1570,N_1496);
and U1732 (N_1732,N_1468,N_1422);
nor U1733 (N_1733,N_1520,N_1435);
and U1734 (N_1734,N_1459,N_1422);
and U1735 (N_1735,N_1406,N_1493);
xnor U1736 (N_1736,N_1498,N_1449);
nor U1737 (N_1737,N_1459,N_1558);
xnor U1738 (N_1738,N_1527,N_1583);
xor U1739 (N_1739,N_1520,N_1595);
and U1740 (N_1740,N_1446,N_1562);
xor U1741 (N_1741,N_1504,N_1416);
nor U1742 (N_1742,N_1469,N_1474);
nand U1743 (N_1743,N_1598,N_1513);
xnor U1744 (N_1744,N_1548,N_1584);
and U1745 (N_1745,N_1496,N_1490);
and U1746 (N_1746,N_1547,N_1585);
or U1747 (N_1747,N_1460,N_1596);
and U1748 (N_1748,N_1468,N_1471);
or U1749 (N_1749,N_1506,N_1571);
nand U1750 (N_1750,N_1542,N_1526);
nand U1751 (N_1751,N_1508,N_1587);
nand U1752 (N_1752,N_1559,N_1563);
nor U1753 (N_1753,N_1422,N_1560);
nor U1754 (N_1754,N_1569,N_1528);
xnor U1755 (N_1755,N_1483,N_1404);
nand U1756 (N_1756,N_1572,N_1568);
xor U1757 (N_1757,N_1429,N_1482);
xor U1758 (N_1758,N_1490,N_1571);
nand U1759 (N_1759,N_1419,N_1427);
or U1760 (N_1760,N_1557,N_1523);
xor U1761 (N_1761,N_1487,N_1407);
and U1762 (N_1762,N_1582,N_1409);
or U1763 (N_1763,N_1476,N_1412);
or U1764 (N_1764,N_1517,N_1592);
xor U1765 (N_1765,N_1589,N_1475);
nand U1766 (N_1766,N_1488,N_1538);
nor U1767 (N_1767,N_1424,N_1488);
or U1768 (N_1768,N_1555,N_1534);
or U1769 (N_1769,N_1412,N_1474);
nor U1770 (N_1770,N_1597,N_1500);
and U1771 (N_1771,N_1536,N_1537);
or U1772 (N_1772,N_1527,N_1586);
and U1773 (N_1773,N_1586,N_1551);
or U1774 (N_1774,N_1539,N_1444);
nand U1775 (N_1775,N_1573,N_1529);
nor U1776 (N_1776,N_1415,N_1424);
nand U1777 (N_1777,N_1571,N_1497);
xor U1778 (N_1778,N_1404,N_1482);
and U1779 (N_1779,N_1573,N_1409);
and U1780 (N_1780,N_1549,N_1546);
or U1781 (N_1781,N_1549,N_1556);
xnor U1782 (N_1782,N_1403,N_1437);
xnor U1783 (N_1783,N_1524,N_1474);
or U1784 (N_1784,N_1563,N_1497);
xor U1785 (N_1785,N_1541,N_1549);
nand U1786 (N_1786,N_1576,N_1495);
or U1787 (N_1787,N_1466,N_1547);
or U1788 (N_1788,N_1542,N_1575);
or U1789 (N_1789,N_1438,N_1599);
and U1790 (N_1790,N_1530,N_1415);
or U1791 (N_1791,N_1510,N_1562);
xnor U1792 (N_1792,N_1566,N_1421);
or U1793 (N_1793,N_1429,N_1448);
and U1794 (N_1794,N_1469,N_1562);
xor U1795 (N_1795,N_1581,N_1485);
nor U1796 (N_1796,N_1589,N_1410);
xnor U1797 (N_1797,N_1451,N_1426);
nor U1798 (N_1798,N_1472,N_1468);
nor U1799 (N_1799,N_1479,N_1520);
nand U1800 (N_1800,N_1632,N_1734);
xnor U1801 (N_1801,N_1767,N_1640);
xor U1802 (N_1802,N_1624,N_1675);
nor U1803 (N_1803,N_1631,N_1704);
xnor U1804 (N_1804,N_1647,N_1664);
and U1805 (N_1805,N_1783,N_1680);
and U1806 (N_1806,N_1738,N_1743);
or U1807 (N_1807,N_1777,N_1623);
nand U1808 (N_1808,N_1699,N_1622);
nor U1809 (N_1809,N_1672,N_1733);
and U1810 (N_1810,N_1790,N_1719);
nand U1811 (N_1811,N_1685,N_1628);
nor U1812 (N_1812,N_1627,N_1762);
nor U1813 (N_1813,N_1797,N_1779);
nor U1814 (N_1814,N_1639,N_1755);
nor U1815 (N_1815,N_1774,N_1731);
nor U1816 (N_1816,N_1683,N_1727);
and U1817 (N_1817,N_1608,N_1748);
xnor U1818 (N_1818,N_1674,N_1619);
or U1819 (N_1819,N_1785,N_1725);
nor U1820 (N_1820,N_1669,N_1626);
nand U1821 (N_1821,N_1605,N_1614);
nand U1822 (N_1822,N_1718,N_1667);
or U1823 (N_1823,N_1645,N_1659);
or U1824 (N_1824,N_1687,N_1751);
nor U1825 (N_1825,N_1766,N_1764);
nand U1826 (N_1826,N_1749,N_1752);
or U1827 (N_1827,N_1660,N_1700);
and U1828 (N_1828,N_1646,N_1671);
or U1829 (N_1829,N_1713,N_1601);
or U1830 (N_1830,N_1653,N_1726);
or U1831 (N_1831,N_1791,N_1656);
nand U1832 (N_1832,N_1615,N_1682);
and U1833 (N_1833,N_1651,N_1698);
nand U1834 (N_1834,N_1650,N_1701);
nor U1835 (N_1835,N_1720,N_1729);
and U1836 (N_1836,N_1668,N_1629);
or U1837 (N_1837,N_1696,N_1786);
nand U1838 (N_1838,N_1691,N_1717);
nor U1839 (N_1839,N_1689,N_1746);
and U1840 (N_1840,N_1678,N_1728);
and U1841 (N_1841,N_1613,N_1692);
nand U1842 (N_1842,N_1787,N_1711);
nor U1843 (N_1843,N_1756,N_1759);
xor U1844 (N_1844,N_1775,N_1600);
nor U1845 (N_1845,N_1611,N_1679);
and U1846 (N_1846,N_1604,N_1636);
nor U1847 (N_1847,N_1633,N_1773);
nand U1848 (N_1848,N_1754,N_1655);
or U1849 (N_1849,N_1799,N_1630);
xor U1850 (N_1850,N_1771,N_1770);
nand U1851 (N_1851,N_1657,N_1673);
xor U1852 (N_1852,N_1607,N_1686);
xor U1853 (N_1853,N_1643,N_1693);
nor U1854 (N_1854,N_1694,N_1765);
nor U1855 (N_1855,N_1781,N_1690);
xnor U1856 (N_1856,N_1760,N_1745);
nand U1857 (N_1857,N_1708,N_1753);
and U1858 (N_1858,N_1665,N_1737);
nand U1859 (N_1859,N_1684,N_1714);
or U1860 (N_1860,N_1741,N_1663);
xnor U1861 (N_1861,N_1792,N_1677);
nor U1862 (N_1862,N_1635,N_1634);
nand U1863 (N_1863,N_1795,N_1722);
and U1864 (N_1864,N_1681,N_1747);
nand U1865 (N_1865,N_1723,N_1620);
and U1866 (N_1866,N_1610,N_1606);
and U1867 (N_1867,N_1621,N_1763);
or U1868 (N_1868,N_1789,N_1716);
or U1869 (N_1869,N_1715,N_1778);
nand U1870 (N_1870,N_1617,N_1648);
nand U1871 (N_1871,N_1744,N_1794);
or U1872 (N_1872,N_1772,N_1649);
and U1873 (N_1873,N_1768,N_1782);
nand U1874 (N_1874,N_1769,N_1654);
or U1875 (N_1875,N_1658,N_1724);
or U1876 (N_1876,N_1784,N_1641);
and U1877 (N_1877,N_1712,N_1788);
or U1878 (N_1878,N_1742,N_1676);
xnor U1879 (N_1879,N_1703,N_1798);
and U1880 (N_1880,N_1618,N_1642);
and U1881 (N_1881,N_1793,N_1730);
or U1882 (N_1882,N_1688,N_1603);
or U1883 (N_1883,N_1625,N_1710);
or U1884 (N_1884,N_1609,N_1740);
xnor U1885 (N_1885,N_1796,N_1638);
nand U1886 (N_1886,N_1721,N_1637);
xor U1887 (N_1887,N_1757,N_1758);
nor U1888 (N_1888,N_1706,N_1666);
nand U1889 (N_1889,N_1644,N_1612);
nand U1890 (N_1890,N_1776,N_1736);
and U1891 (N_1891,N_1616,N_1697);
xor U1892 (N_1892,N_1707,N_1732);
xor U1893 (N_1893,N_1602,N_1661);
xor U1894 (N_1894,N_1739,N_1709);
nand U1895 (N_1895,N_1670,N_1652);
nand U1896 (N_1896,N_1705,N_1735);
nand U1897 (N_1897,N_1780,N_1702);
or U1898 (N_1898,N_1761,N_1695);
nand U1899 (N_1899,N_1662,N_1750);
nand U1900 (N_1900,N_1721,N_1731);
nand U1901 (N_1901,N_1651,N_1685);
and U1902 (N_1902,N_1665,N_1688);
xor U1903 (N_1903,N_1733,N_1744);
nand U1904 (N_1904,N_1619,N_1652);
nor U1905 (N_1905,N_1695,N_1678);
nand U1906 (N_1906,N_1701,N_1647);
and U1907 (N_1907,N_1717,N_1618);
nor U1908 (N_1908,N_1638,N_1776);
nand U1909 (N_1909,N_1708,N_1608);
nand U1910 (N_1910,N_1646,N_1602);
nand U1911 (N_1911,N_1796,N_1797);
xor U1912 (N_1912,N_1681,N_1744);
and U1913 (N_1913,N_1659,N_1781);
xnor U1914 (N_1914,N_1748,N_1714);
nor U1915 (N_1915,N_1673,N_1712);
or U1916 (N_1916,N_1655,N_1767);
and U1917 (N_1917,N_1726,N_1646);
nand U1918 (N_1918,N_1682,N_1724);
xor U1919 (N_1919,N_1698,N_1704);
or U1920 (N_1920,N_1754,N_1700);
nand U1921 (N_1921,N_1698,N_1779);
nor U1922 (N_1922,N_1753,N_1681);
or U1923 (N_1923,N_1689,N_1745);
or U1924 (N_1924,N_1792,N_1609);
and U1925 (N_1925,N_1781,N_1798);
nor U1926 (N_1926,N_1630,N_1700);
and U1927 (N_1927,N_1700,N_1710);
xnor U1928 (N_1928,N_1641,N_1604);
and U1929 (N_1929,N_1733,N_1657);
and U1930 (N_1930,N_1771,N_1617);
and U1931 (N_1931,N_1621,N_1759);
and U1932 (N_1932,N_1796,N_1641);
and U1933 (N_1933,N_1674,N_1784);
and U1934 (N_1934,N_1681,N_1616);
nand U1935 (N_1935,N_1681,N_1760);
xnor U1936 (N_1936,N_1778,N_1659);
nand U1937 (N_1937,N_1741,N_1717);
and U1938 (N_1938,N_1771,N_1705);
xnor U1939 (N_1939,N_1724,N_1648);
nor U1940 (N_1940,N_1609,N_1622);
and U1941 (N_1941,N_1693,N_1649);
nand U1942 (N_1942,N_1772,N_1783);
or U1943 (N_1943,N_1715,N_1695);
nand U1944 (N_1944,N_1735,N_1671);
nand U1945 (N_1945,N_1684,N_1695);
or U1946 (N_1946,N_1759,N_1632);
and U1947 (N_1947,N_1775,N_1642);
nand U1948 (N_1948,N_1753,N_1688);
or U1949 (N_1949,N_1705,N_1667);
and U1950 (N_1950,N_1761,N_1671);
and U1951 (N_1951,N_1684,N_1755);
or U1952 (N_1952,N_1618,N_1600);
nand U1953 (N_1953,N_1761,N_1757);
xor U1954 (N_1954,N_1647,N_1627);
or U1955 (N_1955,N_1661,N_1798);
nor U1956 (N_1956,N_1776,N_1645);
and U1957 (N_1957,N_1799,N_1615);
xor U1958 (N_1958,N_1639,N_1722);
nand U1959 (N_1959,N_1751,N_1756);
nand U1960 (N_1960,N_1698,N_1617);
xnor U1961 (N_1961,N_1766,N_1732);
xnor U1962 (N_1962,N_1643,N_1676);
xor U1963 (N_1963,N_1759,N_1773);
nor U1964 (N_1964,N_1648,N_1669);
and U1965 (N_1965,N_1734,N_1605);
and U1966 (N_1966,N_1751,N_1626);
nand U1967 (N_1967,N_1749,N_1784);
nand U1968 (N_1968,N_1736,N_1637);
nand U1969 (N_1969,N_1680,N_1757);
nor U1970 (N_1970,N_1734,N_1600);
nor U1971 (N_1971,N_1743,N_1633);
xnor U1972 (N_1972,N_1619,N_1780);
and U1973 (N_1973,N_1681,N_1745);
or U1974 (N_1974,N_1745,N_1618);
and U1975 (N_1975,N_1646,N_1611);
xnor U1976 (N_1976,N_1699,N_1634);
and U1977 (N_1977,N_1645,N_1696);
and U1978 (N_1978,N_1767,N_1642);
xnor U1979 (N_1979,N_1712,N_1774);
or U1980 (N_1980,N_1757,N_1617);
nor U1981 (N_1981,N_1682,N_1786);
nand U1982 (N_1982,N_1713,N_1607);
nor U1983 (N_1983,N_1686,N_1789);
nor U1984 (N_1984,N_1782,N_1630);
nand U1985 (N_1985,N_1702,N_1707);
and U1986 (N_1986,N_1701,N_1645);
or U1987 (N_1987,N_1751,N_1704);
and U1988 (N_1988,N_1744,N_1628);
nand U1989 (N_1989,N_1751,N_1707);
and U1990 (N_1990,N_1606,N_1726);
nor U1991 (N_1991,N_1736,N_1636);
xor U1992 (N_1992,N_1684,N_1793);
or U1993 (N_1993,N_1764,N_1752);
nand U1994 (N_1994,N_1710,N_1662);
xnor U1995 (N_1995,N_1716,N_1650);
xnor U1996 (N_1996,N_1739,N_1723);
nor U1997 (N_1997,N_1609,N_1783);
nor U1998 (N_1998,N_1793,N_1757);
nor U1999 (N_1999,N_1668,N_1707);
and U2000 (N_2000,N_1819,N_1837);
or U2001 (N_2001,N_1957,N_1824);
nand U2002 (N_2002,N_1909,N_1835);
nand U2003 (N_2003,N_1942,N_1915);
nor U2004 (N_2004,N_1864,N_1876);
nand U2005 (N_2005,N_1826,N_1847);
nand U2006 (N_2006,N_1963,N_1857);
nand U2007 (N_2007,N_1984,N_1865);
or U2008 (N_2008,N_1883,N_1889);
nand U2009 (N_2009,N_1801,N_1822);
or U2010 (N_2010,N_1871,N_1992);
nand U2011 (N_2011,N_1813,N_1874);
xnor U2012 (N_2012,N_1914,N_1922);
nor U2013 (N_2013,N_1939,N_1917);
and U2014 (N_2014,N_1959,N_1867);
and U2015 (N_2015,N_1800,N_1825);
nand U2016 (N_2016,N_1806,N_1869);
xnor U2017 (N_2017,N_1958,N_1892);
and U2018 (N_2018,N_1817,N_1993);
and U2019 (N_2019,N_1821,N_1997);
nand U2020 (N_2020,N_1863,N_1870);
and U2021 (N_2021,N_1833,N_1930);
or U2022 (N_2022,N_1947,N_1980);
nor U2023 (N_2023,N_1814,N_1991);
nand U2024 (N_2024,N_1938,N_1972);
xor U2025 (N_2025,N_1954,N_1907);
nand U2026 (N_2026,N_1851,N_1898);
and U2027 (N_2027,N_1921,N_1969);
or U2028 (N_2028,N_1836,N_1998);
and U2029 (N_2029,N_1919,N_1977);
nor U2030 (N_2030,N_1924,N_1975);
or U2031 (N_2031,N_1941,N_1890);
nor U2032 (N_2032,N_1880,N_1846);
xor U2033 (N_2033,N_1911,N_1931);
and U2034 (N_2034,N_1979,N_1920);
nand U2035 (N_2035,N_1987,N_1809);
xnor U2036 (N_2036,N_1950,N_1970);
nor U2037 (N_2037,N_1965,N_1861);
xnor U2038 (N_2038,N_1960,N_1808);
xnor U2039 (N_2039,N_1912,N_1897);
and U2040 (N_2040,N_1974,N_1905);
nand U2041 (N_2041,N_1816,N_1955);
nand U2042 (N_2042,N_1860,N_1881);
xnor U2043 (N_2043,N_1953,N_1815);
and U2044 (N_2044,N_1810,N_1926);
or U2045 (N_2045,N_1873,N_1886);
and U2046 (N_2046,N_1976,N_1859);
xnor U2047 (N_2047,N_1830,N_1916);
xor U2048 (N_2048,N_1850,N_1988);
nor U2049 (N_2049,N_1981,N_1811);
xnor U2050 (N_2050,N_1862,N_1834);
nor U2051 (N_2051,N_1854,N_1841);
and U2052 (N_2052,N_1840,N_1994);
xnor U2053 (N_2053,N_1936,N_1875);
and U2054 (N_2054,N_1927,N_1985);
or U2055 (N_2055,N_1807,N_1966);
and U2056 (N_2056,N_1956,N_1858);
and U2057 (N_2057,N_1843,N_1868);
and U2058 (N_2058,N_1804,N_1934);
xnor U2059 (N_2059,N_1946,N_1802);
or U2060 (N_2060,N_1853,N_1933);
or U2061 (N_2061,N_1838,N_1973);
nand U2062 (N_2062,N_1918,N_1849);
and U2063 (N_2063,N_1805,N_1894);
and U2064 (N_2064,N_1884,N_1823);
nor U2065 (N_2065,N_1989,N_1866);
or U2066 (N_2066,N_1856,N_1820);
and U2067 (N_2067,N_1845,N_1902);
nand U2068 (N_2068,N_1827,N_1879);
and U2069 (N_2069,N_1872,N_1948);
and U2070 (N_2070,N_1803,N_1896);
or U2071 (N_2071,N_1925,N_1962);
or U2072 (N_2072,N_1913,N_1910);
nor U2073 (N_2073,N_1929,N_1852);
or U2074 (N_2074,N_1887,N_1828);
or U2075 (N_2075,N_1831,N_1945);
nand U2076 (N_2076,N_1971,N_1900);
xor U2077 (N_2077,N_1903,N_1932);
nor U2078 (N_2078,N_1848,N_1995);
or U2079 (N_2079,N_1983,N_1949);
or U2080 (N_2080,N_1967,N_1943);
or U2081 (N_2081,N_1935,N_1982);
or U2082 (N_2082,N_1891,N_1878);
or U2083 (N_2083,N_1888,N_1855);
xor U2084 (N_2084,N_1842,N_1906);
xor U2085 (N_2085,N_1968,N_1996);
or U2086 (N_2086,N_1978,N_1901);
nor U2087 (N_2087,N_1986,N_1937);
nand U2088 (N_2088,N_1885,N_1829);
or U2089 (N_2089,N_1832,N_1844);
xnor U2090 (N_2090,N_1818,N_1904);
nand U2091 (N_2091,N_1839,N_1951);
or U2092 (N_2092,N_1944,N_1952);
or U2093 (N_2093,N_1893,N_1899);
nand U2094 (N_2094,N_1908,N_1895);
nand U2095 (N_2095,N_1877,N_1812);
or U2096 (N_2096,N_1964,N_1940);
or U2097 (N_2097,N_1928,N_1961);
nor U2098 (N_2098,N_1923,N_1999);
nand U2099 (N_2099,N_1882,N_1990);
and U2100 (N_2100,N_1864,N_1857);
or U2101 (N_2101,N_1923,N_1843);
xor U2102 (N_2102,N_1824,N_1989);
nand U2103 (N_2103,N_1842,N_1964);
xnor U2104 (N_2104,N_1949,N_1893);
or U2105 (N_2105,N_1991,N_1876);
and U2106 (N_2106,N_1975,N_1955);
or U2107 (N_2107,N_1929,N_1944);
nor U2108 (N_2108,N_1851,N_1824);
nor U2109 (N_2109,N_1860,N_1886);
nand U2110 (N_2110,N_1878,N_1851);
nor U2111 (N_2111,N_1924,N_1884);
xnor U2112 (N_2112,N_1940,N_1825);
or U2113 (N_2113,N_1825,N_1965);
or U2114 (N_2114,N_1907,N_1912);
or U2115 (N_2115,N_1951,N_1942);
and U2116 (N_2116,N_1836,N_1835);
nand U2117 (N_2117,N_1959,N_1920);
xnor U2118 (N_2118,N_1864,N_1878);
and U2119 (N_2119,N_1910,N_1829);
nor U2120 (N_2120,N_1928,N_1964);
and U2121 (N_2121,N_1926,N_1824);
xnor U2122 (N_2122,N_1815,N_1882);
xor U2123 (N_2123,N_1914,N_1805);
nor U2124 (N_2124,N_1951,N_1804);
xnor U2125 (N_2125,N_1806,N_1846);
xnor U2126 (N_2126,N_1998,N_1940);
xor U2127 (N_2127,N_1814,N_1904);
nand U2128 (N_2128,N_1955,N_1872);
and U2129 (N_2129,N_1876,N_1913);
nand U2130 (N_2130,N_1954,N_1951);
or U2131 (N_2131,N_1955,N_1997);
or U2132 (N_2132,N_1846,N_1938);
xnor U2133 (N_2133,N_1905,N_1892);
or U2134 (N_2134,N_1880,N_1943);
or U2135 (N_2135,N_1872,N_1867);
or U2136 (N_2136,N_1815,N_1843);
nand U2137 (N_2137,N_1836,N_1825);
nand U2138 (N_2138,N_1901,N_1950);
nor U2139 (N_2139,N_1844,N_1860);
or U2140 (N_2140,N_1894,N_1911);
nor U2141 (N_2141,N_1926,N_1843);
and U2142 (N_2142,N_1803,N_1816);
or U2143 (N_2143,N_1944,N_1853);
xnor U2144 (N_2144,N_1993,N_1867);
nand U2145 (N_2145,N_1977,N_1943);
nor U2146 (N_2146,N_1881,N_1813);
and U2147 (N_2147,N_1846,N_1811);
and U2148 (N_2148,N_1946,N_1840);
and U2149 (N_2149,N_1993,N_1900);
or U2150 (N_2150,N_1941,N_1948);
nor U2151 (N_2151,N_1800,N_1955);
nor U2152 (N_2152,N_1969,N_1800);
xnor U2153 (N_2153,N_1861,N_1995);
xnor U2154 (N_2154,N_1934,N_1920);
xnor U2155 (N_2155,N_1837,N_1875);
or U2156 (N_2156,N_1948,N_1909);
or U2157 (N_2157,N_1847,N_1956);
and U2158 (N_2158,N_1971,N_1973);
or U2159 (N_2159,N_1862,N_1853);
xnor U2160 (N_2160,N_1945,N_1813);
and U2161 (N_2161,N_1861,N_1823);
or U2162 (N_2162,N_1837,N_1873);
or U2163 (N_2163,N_1987,N_1858);
nand U2164 (N_2164,N_1862,N_1967);
xnor U2165 (N_2165,N_1826,N_1837);
and U2166 (N_2166,N_1818,N_1907);
and U2167 (N_2167,N_1998,N_1903);
nor U2168 (N_2168,N_1908,N_1953);
nor U2169 (N_2169,N_1893,N_1848);
xor U2170 (N_2170,N_1921,N_1886);
nand U2171 (N_2171,N_1873,N_1878);
xnor U2172 (N_2172,N_1911,N_1848);
or U2173 (N_2173,N_1980,N_1978);
or U2174 (N_2174,N_1922,N_1906);
nand U2175 (N_2175,N_1887,N_1972);
and U2176 (N_2176,N_1936,N_1990);
nor U2177 (N_2177,N_1886,N_1845);
or U2178 (N_2178,N_1916,N_1829);
nor U2179 (N_2179,N_1985,N_1952);
nand U2180 (N_2180,N_1899,N_1808);
nand U2181 (N_2181,N_1874,N_1867);
and U2182 (N_2182,N_1810,N_1869);
nor U2183 (N_2183,N_1965,N_1987);
nand U2184 (N_2184,N_1977,N_1855);
and U2185 (N_2185,N_1902,N_1947);
or U2186 (N_2186,N_1975,N_1825);
xnor U2187 (N_2187,N_1982,N_1813);
nand U2188 (N_2188,N_1979,N_1928);
nand U2189 (N_2189,N_1829,N_1989);
and U2190 (N_2190,N_1875,N_1862);
and U2191 (N_2191,N_1900,N_1824);
xnor U2192 (N_2192,N_1883,N_1933);
and U2193 (N_2193,N_1959,N_1859);
nand U2194 (N_2194,N_1975,N_1993);
xor U2195 (N_2195,N_1936,N_1923);
and U2196 (N_2196,N_1961,N_1858);
and U2197 (N_2197,N_1804,N_1941);
or U2198 (N_2198,N_1903,N_1836);
nand U2199 (N_2199,N_1916,N_1963);
xor U2200 (N_2200,N_2135,N_2067);
xor U2201 (N_2201,N_2052,N_2133);
or U2202 (N_2202,N_2169,N_2022);
nor U2203 (N_2203,N_2080,N_2175);
nand U2204 (N_2204,N_2004,N_2179);
or U2205 (N_2205,N_2060,N_2159);
xnor U2206 (N_2206,N_2103,N_2180);
and U2207 (N_2207,N_2125,N_2116);
or U2208 (N_2208,N_2074,N_2010);
nor U2209 (N_2209,N_2153,N_2195);
nand U2210 (N_2210,N_2113,N_2143);
nor U2211 (N_2211,N_2163,N_2014);
nor U2212 (N_2212,N_2005,N_2138);
and U2213 (N_2213,N_2006,N_2114);
or U2214 (N_2214,N_2025,N_2155);
nand U2215 (N_2215,N_2099,N_2156);
and U2216 (N_2216,N_2036,N_2019);
and U2217 (N_2217,N_2146,N_2012);
and U2218 (N_2218,N_2024,N_2164);
nor U2219 (N_2219,N_2101,N_2105);
nand U2220 (N_2220,N_2154,N_2192);
and U2221 (N_2221,N_2127,N_2176);
nor U2222 (N_2222,N_2097,N_2062);
nand U2223 (N_2223,N_2166,N_2087);
and U2224 (N_2224,N_2042,N_2131);
and U2225 (N_2225,N_2196,N_2044);
or U2226 (N_2226,N_2041,N_2003);
or U2227 (N_2227,N_2043,N_2034);
xor U2228 (N_2228,N_2017,N_2057);
nand U2229 (N_2229,N_2158,N_2089);
or U2230 (N_2230,N_2141,N_2077);
and U2231 (N_2231,N_2157,N_2094);
nor U2232 (N_2232,N_2035,N_2130);
xnor U2233 (N_2233,N_2132,N_2096);
and U2234 (N_2234,N_2072,N_2183);
nor U2235 (N_2235,N_2013,N_2174);
nor U2236 (N_2236,N_2108,N_2149);
or U2237 (N_2237,N_2191,N_2063);
nand U2238 (N_2238,N_2082,N_2121);
xor U2239 (N_2239,N_2048,N_2136);
nand U2240 (N_2240,N_2151,N_2181);
nand U2241 (N_2241,N_2173,N_2083);
and U2242 (N_2242,N_2002,N_2061);
or U2243 (N_2243,N_2055,N_2129);
nor U2244 (N_2244,N_2126,N_2148);
nand U2245 (N_2245,N_2177,N_2020);
nand U2246 (N_2246,N_2168,N_2115);
xor U2247 (N_2247,N_2053,N_2095);
and U2248 (N_2248,N_2160,N_2039);
nor U2249 (N_2249,N_2018,N_2139);
nor U2250 (N_2250,N_2104,N_2142);
and U2251 (N_2251,N_2015,N_2075);
xor U2252 (N_2252,N_2051,N_2147);
and U2253 (N_2253,N_2100,N_2137);
nand U2254 (N_2254,N_2172,N_2198);
xor U2255 (N_2255,N_2056,N_2008);
nor U2256 (N_2256,N_2190,N_2186);
xor U2257 (N_2257,N_2066,N_2079);
and U2258 (N_2258,N_2011,N_2187);
xnor U2259 (N_2259,N_2118,N_2152);
and U2260 (N_2260,N_2110,N_2009);
or U2261 (N_2261,N_2167,N_2016);
nor U2262 (N_2262,N_2047,N_2161);
and U2263 (N_2263,N_2049,N_2124);
xnor U2264 (N_2264,N_2054,N_2162);
and U2265 (N_2265,N_2026,N_2050);
nand U2266 (N_2266,N_2111,N_2064);
nand U2267 (N_2267,N_2093,N_2182);
xnor U2268 (N_2268,N_2032,N_2001);
nor U2269 (N_2269,N_2178,N_2029);
and U2270 (N_2270,N_2038,N_2033);
nand U2271 (N_2271,N_2122,N_2091);
xnor U2272 (N_2272,N_2046,N_2098);
nor U2273 (N_2273,N_2134,N_2081);
nor U2274 (N_2274,N_2102,N_2058);
or U2275 (N_2275,N_2184,N_2076);
nor U2276 (N_2276,N_2194,N_2199);
xnor U2277 (N_2277,N_2150,N_2107);
and U2278 (N_2278,N_2085,N_2092);
nor U2279 (N_2279,N_2073,N_2170);
nand U2280 (N_2280,N_2065,N_2145);
and U2281 (N_2281,N_2069,N_2068);
xnor U2282 (N_2282,N_2023,N_2059);
nor U2283 (N_2283,N_2071,N_2090);
or U2284 (N_2284,N_2021,N_2165);
nand U2285 (N_2285,N_2084,N_2027);
or U2286 (N_2286,N_2189,N_2031);
nand U2287 (N_2287,N_2070,N_2123);
or U2288 (N_2288,N_2112,N_2078);
xor U2289 (N_2289,N_2045,N_2040);
and U2290 (N_2290,N_2000,N_2193);
nor U2291 (N_2291,N_2144,N_2197);
and U2292 (N_2292,N_2007,N_2119);
or U2293 (N_2293,N_2188,N_2086);
nor U2294 (N_2294,N_2171,N_2030);
or U2295 (N_2295,N_2028,N_2037);
and U2296 (N_2296,N_2140,N_2120);
xnor U2297 (N_2297,N_2106,N_2185);
and U2298 (N_2298,N_2117,N_2088);
or U2299 (N_2299,N_2109,N_2128);
or U2300 (N_2300,N_2093,N_2172);
nand U2301 (N_2301,N_2083,N_2104);
nor U2302 (N_2302,N_2167,N_2020);
nand U2303 (N_2303,N_2103,N_2167);
nor U2304 (N_2304,N_2121,N_2086);
xnor U2305 (N_2305,N_2183,N_2130);
and U2306 (N_2306,N_2126,N_2002);
nand U2307 (N_2307,N_2156,N_2187);
xnor U2308 (N_2308,N_2180,N_2068);
or U2309 (N_2309,N_2004,N_2033);
nor U2310 (N_2310,N_2166,N_2110);
xnor U2311 (N_2311,N_2139,N_2126);
nor U2312 (N_2312,N_2150,N_2027);
xnor U2313 (N_2313,N_2044,N_2129);
or U2314 (N_2314,N_2107,N_2171);
xor U2315 (N_2315,N_2197,N_2011);
and U2316 (N_2316,N_2138,N_2043);
nand U2317 (N_2317,N_2104,N_2031);
xnor U2318 (N_2318,N_2133,N_2032);
xnor U2319 (N_2319,N_2114,N_2062);
xnor U2320 (N_2320,N_2151,N_2030);
nand U2321 (N_2321,N_2033,N_2055);
and U2322 (N_2322,N_2042,N_2123);
nor U2323 (N_2323,N_2178,N_2063);
and U2324 (N_2324,N_2092,N_2173);
xnor U2325 (N_2325,N_2061,N_2058);
or U2326 (N_2326,N_2119,N_2135);
nand U2327 (N_2327,N_2002,N_2179);
or U2328 (N_2328,N_2010,N_2067);
xnor U2329 (N_2329,N_2195,N_2162);
nor U2330 (N_2330,N_2176,N_2152);
or U2331 (N_2331,N_2003,N_2070);
nor U2332 (N_2332,N_2109,N_2168);
nor U2333 (N_2333,N_2059,N_2183);
nand U2334 (N_2334,N_2117,N_2175);
or U2335 (N_2335,N_2002,N_2088);
xor U2336 (N_2336,N_2030,N_2115);
xor U2337 (N_2337,N_2187,N_2112);
nand U2338 (N_2338,N_2163,N_2181);
and U2339 (N_2339,N_2171,N_2031);
and U2340 (N_2340,N_2112,N_2000);
and U2341 (N_2341,N_2029,N_2082);
xnor U2342 (N_2342,N_2119,N_2014);
xor U2343 (N_2343,N_2159,N_2098);
nor U2344 (N_2344,N_2027,N_2136);
xor U2345 (N_2345,N_2178,N_2173);
xnor U2346 (N_2346,N_2059,N_2076);
nand U2347 (N_2347,N_2049,N_2100);
nor U2348 (N_2348,N_2150,N_2189);
nand U2349 (N_2349,N_2131,N_2100);
or U2350 (N_2350,N_2017,N_2043);
nand U2351 (N_2351,N_2132,N_2167);
nor U2352 (N_2352,N_2013,N_2049);
nand U2353 (N_2353,N_2107,N_2083);
nand U2354 (N_2354,N_2125,N_2128);
xor U2355 (N_2355,N_2024,N_2135);
nand U2356 (N_2356,N_2120,N_2150);
nor U2357 (N_2357,N_2036,N_2140);
or U2358 (N_2358,N_2110,N_2070);
nor U2359 (N_2359,N_2077,N_2185);
or U2360 (N_2360,N_2136,N_2101);
xor U2361 (N_2361,N_2163,N_2185);
xnor U2362 (N_2362,N_2171,N_2175);
xnor U2363 (N_2363,N_2046,N_2070);
or U2364 (N_2364,N_2020,N_2192);
or U2365 (N_2365,N_2163,N_2157);
xor U2366 (N_2366,N_2120,N_2094);
nor U2367 (N_2367,N_2094,N_2026);
nor U2368 (N_2368,N_2098,N_2026);
nand U2369 (N_2369,N_2109,N_2050);
nand U2370 (N_2370,N_2164,N_2114);
or U2371 (N_2371,N_2059,N_2081);
and U2372 (N_2372,N_2050,N_2022);
or U2373 (N_2373,N_2017,N_2091);
or U2374 (N_2374,N_2192,N_2170);
nand U2375 (N_2375,N_2186,N_2162);
nor U2376 (N_2376,N_2111,N_2047);
and U2377 (N_2377,N_2188,N_2037);
nand U2378 (N_2378,N_2131,N_2041);
or U2379 (N_2379,N_2114,N_2028);
nand U2380 (N_2380,N_2127,N_2198);
nand U2381 (N_2381,N_2160,N_2165);
xnor U2382 (N_2382,N_2170,N_2018);
xnor U2383 (N_2383,N_2135,N_2007);
nand U2384 (N_2384,N_2035,N_2031);
nand U2385 (N_2385,N_2080,N_2147);
or U2386 (N_2386,N_2175,N_2159);
xnor U2387 (N_2387,N_2161,N_2079);
or U2388 (N_2388,N_2184,N_2183);
or U2389 (N_2389,N_2004,N_2197);
xor U2390 (N_2390,N_2002,N_2110);
nor U2391 (N_2391,N_2134,N_2097);
xor U2392 (N_2392,N_2009,N_2147);
nand U2393 (N_2393,N_2196,N_2096);
and U2394 (N_2394,N_2196,N_2105);
xnor U2395 (N_2395,N_2110,N_2150);
nor U2396 (N_2396,N_2128,N_2009);
nand U2397 (N_2397,N_2153,N_2159);
or U2398 (N_2398,N_2111,N_2115);
and U2399 (N_2399,N_2080,N_2179);
or U2400 (N_2400,N_2335,N_2261);
nor U2401 (N_2401,N_2205,N_2249);
and U2402 (N_2402,N_2328,N_2283);
xnor U2403 (N_2403,N_2372,N_2343);
and U2404 (N_2404,N_2342,N_2236);
xor U2405 (N_2405,N_2221,N_2332);
and U2406 (N_2406,N_2351,N_2256);
nand U2407 (N_2407,N_2290,N_2211);
or U2408 (N_2408,N_2257,N_2223);
xor U2409 (N_2409,N_2299,N_2248);
xor U2410 (N_2410,N_2293,N_2271);
or U2411 (N_2411,N_2207,N_2219);
and U2412 (N_2412,N_2339,N_2309);
nor U2413 (N_2413,N_2352,N_2364);
or U2414 (N_2414,N_2302,N_2275);
xnor U2415 (N_2415,N_2241,N_2289);
nor U2416 (N_2416,N_2220,N_2312);
and U2417 (N_2417,N_2315,N_2370);
xnor U2418 (N_2418,N_2329,N_2297);
and U2419 (N_2419,N_2396,N_2310);
and U2420 (N_2420,N_2233,N_2318);
and U2421 (N_2421,N_2252,N_2284);
or U2422 (N_2422,N_2327,N_2239);
xnor U2423 (N_2423,N_2334,N_2345);
and U2424 (N_2424,N_2368,N_2308);
or U2425 (N_2425,N_2273,N_2388);
nand U2426 (N_2426,N_2350,N_2262);
or U2427 (N_2427,N_2304,N_2287);
xnor U2428 (N_2428,N_2242,N_2353);
or U2429 (N_2429,N_2206,N_2369);
xnor U2430 (N_2430,N_2266,N_2210);
or U2431 (N_2431,N_2389,N_2348);
or U2432 (N_2432,N_2244,N_2208);
nand U2433 (N_2433,N_2373,N_2215);
nand U2434 (N_2434,N_2323,N_2386);
nand U2435 (N_2435,N_2243,N_2213);
nand U2436 (N_2436,N_2317,N_2379);
xor U2437 (N_2437,N_2203,N_2321);
nand U2438 (N_2438,N_2240,N_2381);
nand U2439 (N_2439,N_2232,N_2229);
and U2440 (N_2440,N_2225,N_2295);
nand U2441 (N_2441,N_2286,N_2399);
xor U2442 (N_2442,N_2365,N_2292);
and U2443 (N_2443,N_2383,N_2263);
xnor U2444 (N_2444,N_2288,N_2260);
nand U2445 (N_2445,N_2347,N_2235);
xor U2446 (N_2446,N_2360,N_2255);
and U2447 (N_2447,N_2227,N_2326);
or U2448 (N_2448,N_2333,N_2387);
nor U2449 (N_2449,N_2307,N_2270);
and U2450 (N_2450,N_2361,N_2354);
nor U2451 (N_2451,N_2325,N_2204);
nor U2452 (N_2452,N_2395,N_2313);
xor U2453 (N_2453,N_2214,N_2280);
nand U2454 (N_2454,N_2322,N_2294);
xnor U2455 (N_2455,N_2269,N_2316);
nor U2456 (N_2456,N_2397,N_2259);
xor U2457 (N_2457,N_2380,N_2382);
nand U2458 (N_2458,N_2366,N_2391);
and U2459 (N_2459,N_2222,N_2282);
nand U2460 (N_2460,N_2362,N_2247);
nand U2461 (N_2461,N_2238,N_2226);
or U2462 (N_2462,N_2224,N_2200);
nand U2463 (N_2463,N_2338,N_2245);
nor U2464 (N_2464,N_2279,N_2276);
xnor U2465 (N_2465,N_2230,N_2331);
nor U2466 (N_2466,N_2250,N_2392);
and U2467 (N_2467,N_2390,N_2394);
nor U2468 (N_2468,N_2201,N_2385);
and U2469 (N_2469,N_2336,N_2377);
and U2470 (N_2470,N_2349,N_2251);
nor U2471 (N_2471,N_2384,N_2371);
or U2472 (N_2472,N_2376,N_2231);
nor U2473 (N_2473,N_2356,N_2254);
xor U2474 (N_2474,N_2264,N_2202);
nand U2475 (N_2475,N_2357,N_2209);
nand U2476 (N_2476,N_2278,N_2306);
nand U2477 (N_2477,N_2355,N_2367);
and U2478 (N_2478,N_2359,N_2344);
nor U2479 (N_2479,N_2281,N_2305);
or U2480 (N_2480,N_2237,N_2246);
nor U2481 (N_2481,N_2311,N_2340);
nand U2482 (N_2482,N_2324,N_2253);
nand U2483 (N_2483,N_2303,N_2267);
and U2484 (N_2484,N_2285,N_2218);
nand U2485 (N_2485,N_2300,N_2298);
nand U2486 (N_2486,N_2319,N_2330);
nor U2487 (N_2487,N_2398,N_2393);
xor U2488 (N_2488,N_2320,N_2277);
nor U2489 (N_2489,N_2234,N_2217);
nand U2490 (N_2490,N_2212,N_2375);
xor U2491 (N_2491,N_2374,N_2228);
and U2492 (N_2492,N_2274,N_2301);
or U2493 (N_2493,N_2314,N_2291);
nand U2494 (N_2494,N_2268,N_2346);
nand U2495 (N_2495,N_2341,N_2296);
or U2496 (N_2496,N_2265,N_2272);
xor U2497 (N_2497,N_2216,N_2378);
and U2498 (N_2498,N_2337,N_2358);
nor U2499 (N_2499,N_2258,N_2363);
nand U2500 (N_2500,N_2222,N_2373);
nor U2501 (N_2501,N_2233,N_2320);
nand U2502 (N_2502,N_2276,N_2370);
nand U2503 (N_2503,N_2304,N_2396);
or U2504 (N_2504,N_2367,N_2210);
xnor U2505 (N_2505,N_2253,N_2322);
nand U2506 (N_2506,N_2292,N_2228);
or U2507 (N_2507,N_2249,N_2348);
xor U2508 (N_2508,N_2303,N_2255);
nor U2509 (N_2509,N_2256,N_2397);
nand U2510 (N_2510,N_2390,N_2367);
nor U2511 (N_2511,N_2297,N_2243);
and U2512 (N_2512,N_2341,N_2294);
xnor U2513 (N_2513,N_2316,N_2324);
nor U2514 (N_2514,N_2320,N_2310);
xnor U2515 (N_2515,N_2254,N_2333);
and U2516 (N_2516,N_2395,N_2311);
or U2517 (N_2517,N_2379,N_2232);
xor U2518 (N_2518,N_2355,N_2393);
xnor U2519 (N_2519,N_2385,N_2200);
and U2520 (N_2520,N_2354,N_2282);
nand U2521 (N_2521,N_2293,N_2203);
nand U2522 (N_2522,N_2226,N_2320);
nand U2523 (N_2523,N_2335,N_2318);
nand U2524 (N_2524,N_2259,N_2246);
or U2525 (N_2525,N_2323,N_2396);
xor U2526 (N_2526,N_2352,N_2304);
and U2527 (N_2527,N_2399,N_2394);
nor U2528 (N_2528,N_2281,N_2391);
or U2529 (N_2529,N_2399,N_2309);
or U2530 (N_2530,N_2291,N_2387);
nor U2531 (N_2531,N_2322,N_2332);
and U2532 (N_2532,N_2225,N_2206);
nand U2533 (N_2533,N_2318,N_2280);
nand U2534 (N_2534,N_2378,N_2315);
xnor U2535 (N_2535,N_2245,N_2239);
nand U2536 (N_2536,N_2368,N_2274);
nor U2537 (N_2537,N_2396,N_2379);
or U2538 (N_2538,N_2239,N_2360);
xor U2539 (N_2539,N_2229,N_2307);
or U2540 (N_2540,N_2382,N_2232);
or U2541 (N_2541,N_2333,N_2347);
or U2542 (N_2542,N_2293,N_2330);
or U2543 (N_2543,N_2202,N_2222);
and U2544 (N_2544,N_2287,N_2345);
or U2545 (N_2545,N_2201,N_2262);
and U2546 (N_2546,N_2392,N_2229);
xnor U2547 (N_2547,N_2307,N_2248);
nor U2548 (N_2548,N_2277,N_2351);
and U2549 (N_2549,N_2224,N_2253);
or U2550 (N_2550,N_2254,N_2201);
or U2551 (N_2551,N_2203,N_2357);
nand U2552 (N_2552,N_2325,N_2364);
xor U2553 (N_2553,N_2356,N_2248);
and U2554 (N_2554,N_2281,N_2392);
nand U2555 (N_2555,N_2333,N_2367);
and U2556 (N_2556,N_2387,N_2318);
nand U2557 (N_2557,N_2304,N_2318);
or U2558 (N_2558,N_2202,N_2336);
xnor U2559 (N_2559,N_2314,N_2303);
nor U2560 (N_2560,N_2244,N_2292);
nor U2561 (N_2561,N_2357,N_2355);
xor U2562 (N_2562,N_2262,N_2364);
nor U2563 (N_2563,N_2297,N_2322);
xnor U2564 (N_2564,N_2257,N_2294);
or U2565 (N_2565,N_2296,N_2380);
xor U2566 (N_2566,N_2227,N_2301);
xnor U2567 (N_2567,N_2397,N_2393);
xor U2568 (N_2568,N_2227,N_2309);
or U2569 (N_2569,N_2249,N_2251);
xor U2570 (N_2570,N_2364,N_2317);
nand U2571 (N_2571,N_2377,N_2315);
xnor U2572 (N_2572,N_2319,N_2235);
nand U2573 (N_2573,N_2244,N_2210);
nand U2574 (N_2574,N_2353,N_2346);
nor U2575 (N_2575,N_2363,N_2261);
nor U2576 (N_2576,N_2222,N_2316);
xor U2577 (N_2577,N_2399,N_2244);
nor U2578 (N_2578,N_2333,N_2354);
nand U2579 (N_2579,N_2346,N_2270);
nor U2580 (N_2580,N_2356,N_2290);
and U2581 (N_2581,N_2382,N_2318);
and U2582 (N_2582,N_2203,N_2209);
xnor U2583 (N_2583,N_2219,N_2280);
nor U2584 (N_2584,N_2343,N_2266);
or U2585 (N_2585,N_2383,N_2308);
xnor U2586 (N_2586,N_2262,N_2254);
and U2587 (N_2587,N_2266,N_2301);
or U2588 (N_2588,N_2290,N_2379);
nand U2589 (N_2589,N_2388,N_2200);
xnor U2590 (N_2590,N_2306,N_2285);
nor U2591 (N_2591,N_2283,N_2302);
xor U2592 (N_2592,N_2388,N_2267);
and U2593 (N_2593,N_2254,N_2267);
nand U2594 (N_2594,N_2247,N_2360);
or U2595 (N_2595,N_2387,N_2247);
and U2596 (N_2596,N_2305,N_2319);
or U2597 (N_2597,N_2247,N_2286);
and U2598 (N_2598,N_2381,N_2396);
or U2599 (N_2599,N_2242,N_2364);
or U2600 (N_2600,N_2554,N_2481);
xor U2601 (N_2601,N_2423,N_2430);
xnor U2602 (N_2602,N_2522,N_2446);
nor U2603 (N_2603,N_2424,N_2445);
and U2604 (N_2604,N_2418,N_2487);
or U2605 (N_2605,N_2587,N_2441);
or U2606 (N_2606,N_2502,N_2553);
and U2607 (N_2607,N_2503,N_2412);
or U2608 (N_2608,N_2457,N_2484);
xnor U2609 (N_2609,N_2540,N_2595);
nand U2610 (N_2610,N_2547,N_2570);
and U2611 (N_2611,N_2546,N_2574);
and U2612 (N_2612,N_2401,N_2597);
and U2613 (N_2613,N_2551,N_2447);
nand U2614 (N_2614,N_2590,N_2488);
xor U2615 (N_2615,N_2460,N_2432);
nor U2616 (N_2616,N_2500,N_2405);
nand U2617 (N_2617,N_2462,N_2419);
nand U2618 (N_2618,N_2489,N_2542);
and U2619 (N_2619,N_2429,N_2596);
nor U2620 (N_2620,N_2579,N_2582);
nand U2621 (N_2621,N_2584,N_2544);
nand U2622 (N_2622,N_2598,N_2518);
xor U2623 (N_2623,N_2491,N_2404);
and U2624 (N_2624,N_2478,N_2559);
or U2625 (N_2625,N_2538,N_2564);
xnor U2626 (N_2626,N_2480,N_2434);
nand U2627 (N_2627,N_2586,N_2466);
or U2628 (N_2628,N_2433,N_2519);
nand U2629 (N_2629,N_2452,N_2558);
or U2630 (N_2630,N_2575,N_2515);
nor U2631 (N_2631,N_2509,N_2413);
nor U2632 (N_2632,N_2409,N_2456);
nor U2633 (N_2633,N_2567,N_2490);
nand U2634 (N_2634,N_2520,N_2465);
xor U2635 (N_2635,N_2511,N_2531);
nor U2636 (N_2636,N_2536,N_2562);
and U2637 (N_2637,N_2420,N_2422);
and U2638 (N_2638,N_2534,N_2400);
nor U2639 (N_2639,N_2474,N_2557);
and U2640 (N_2640,N_2499,N_2594);
xnor U2641 (N_2641,N_2498,N_2449);
and U2642 (N_2642,N_2569,N_2578);
nor U2643 (N_2643,N_2440,N_2463);
nand U2644 (N_2644,N_2427,N_2439);
nand U2645 (N_2645,N_2532,N_2537);
and U2646 (N_2646,N_2591,N_2479);
xor U2647 (N_2647,N_2402,N_2572);
or U2648 (N_2648,N_2568,N_2437);
and U2649 (N_2649,N_2451,N_2548);
xor U2650 (N_2650,N_2493,N_2485);
nor U2651 (N_2651,N_2461,N_2468);
or U2652 (N_2652,N_2425,N_2549);
or U2653 (N_2653,N_2443,N_2450);
nor U2654 (N_2654,N_2428,N_2406);
nor U2655 (N_2655,N_2454,N_2593);
nor U2656 (N_2656,N_2426,N_2482);
and U2657 (N_2657,N_2475,N_2560);
nand U2658 (N_2658,N_2469,N_2588);
nor U2659 (N_2659,N_2566,N_2455);
and U2660 (N_2660,N_2528,N_2486);
or U2661 (N_2661,N_2471,N_2444);
or U2662 (N_2662,N_2526,N_2431);
nor U2663 (N_2663,N_2525,N_2507);
and U2664 (N_2664,N_2472,N_2506);
xnor U2665 (N_2665,N_2508,N_2417);
or U2666 (N_2666,N_2513,N_2421);
or U2667 (N_2667,N_2581,N_2573);
or U2668 (N_2668,N_2415,N_2563);
nand U2669 (N_2669,N_2521,N_2448);
nor U2670 (N_2670,N_2533,N_2556);
nand U2671 (N_2671,N_2545,N_2414);
xor U2672 (N_2672,N_2523,N_2577);
or U2673 (N_2673,N_2517,N_2530);
and U2674 (N_2674,N_2416,N_2483);
nand U2675 (N_2675,N_2410,N_2550);
or U2676 (N_2676,N_2516,N_2497);
nor U2677 (N_2677,N_2505,N_2408);
nand U2678 (N_2678,N_2496,N_2552);
nor U2679 (N_2679,N_2583,N_2473);
nand U2680 (N_2680,N_2411,N_2599);
or U2681 (N_2681,N_2501,N_2561);
or U2682 (N_2682,N_2529,N_2476);
or U2683 (N_2683,N_2592,N_2495);
or U2684 (N_2684,N_2535,N_2555);
and U2685 (N_2685,N_2470,N_2580);
nor U2686 (N_2686,N_2543,N_2492);
nand U2687 (N_2687,N_2438,N_2453);
or U2688 (N_2688,N_2403,N_2459);
nand U2689 (N_2689,N_2477,N_2494);
nand U2690 (N_2690,N_2589,N_2436);
nor U2691 (N_2691,N_2442,N_2539);
nor U2692 (N_2692,N_2407,N_2458);
nor U2693 (N_2693,N_2464,N_2541);
or U2694 (N_2694,N_2571,N_2565);
nand U2695 (N_2695,N_2510,N_2585);
or U2696 (N_2696,N_2467,N_2524);
xor U2697 (N_2697,N_2512,N_2435);
or U2698 (N_2698,N_2576,N_2504);
nor U2699 (N_2699,N_2514,N_2527);
or U2700 (N_2700,N_2550,N_2541);
xor U2701 (N_2701,N_2496,N_2491);
or U2702 (N_2702,N_2451,N_2522);
nor U2703 (N_2703,N_2483,N_2547);
nor U2704 (N_2704,N_2548,N_2538);
nor U2705 (N_2705,N_2429,N_2489);
xor U2706 (N_2706,N_2488,N_2423);
nand U2707 (N_2707,N_2562,N_2461);
xnor U2708 (N_2708,N_2547,N_2497);
xnor U2709 (N_2709,N_2453,N_2481);
and U2710 (N_2710,N_2558,N_2556);
nor U2711 (N_2711,N_2450,N_2469);
nand U2712 (N_2712,N_2475,N_2520);
nor U2713 (N_2713,N_2561,N_2530);
or U2714 (N_2714,N_2446,N_2444);
nor U2715 (N_2715,N_2555,N_2406);
nand U2716 (N_2716,N_2584,N_2534);
nand U2717 (N_2717,N_2405,N_2430);
and U2718 (N_2718,N_2509,N_2506);
or U2719 (N_2719,N_2443,N_2469);
nor U2720 (N_2720,N_2497,N_2423);
xor U2721 (N_2721,N_2494,N_2577);
nand U2722 (N_2722,N_2593,N_2404);
nor U2723 (N_2723,N_2485,N_2518);
and U2724 (N_2724,N_2446,N_2573);
or U2725 (N_2725,N_2459,N_2439);
nand U2726 (N_2726,N_2483,N_2529);
nand U2727 (N_2727,N_2492,N_2413);
nand U2728 (N_2728,N_2467,N_2409);
or U2729 (N_2729,N_2464,N_2506);
and U2730 (N_2730,N_2471,N_2561);
nand U2731 (N_2731,N_2492,N_2441);
nand U2732 (N_2732,N_2513,N_2475);
nand U2733 (N_2733,N_2566,N_2523);
and U2734 (N_2734,N_2480,N_2576);
xnor U2735 (N_2735,N_2570,N_2583);
nand U2736 (N_2736,N_2472,N_2463);
or U2737 (N_2737,N_2510,N_2465);
xor U2738 (N_2738,N_2596,N_2595);
nand U2739 (N_2739,N_2588,N_2507);
nand U2740 (N_2740,N_2448,N_2587);
nand U2741 (N_2741,N_2430,N_2468);
or U2742 (N_2742,N_2519,N_2530);
nand U2743 (N_2743,N_2515,N_2479);
nor U2744 (N_2744,N_2517,N_2595);
or U2745 (N_2745,N_2463,N_2568);
xnor U2746 (N_2746,N_2511,N_2525);
or U2747 (N_2747,N_2403,N_2426);
nand U2748 (N_2748,N_2540,N_2542);
nor U2749 (N_2749,N_2409,N_2562);
or U2750 (N_2750,N_2424,N_2410);
nand U2751 (N_2751,N_2530,N_2449);
and U2752 (N_2752,N_2586,N_2405);
xor U2753 (N_2753,N_2531,N_2403);
xor U2754 (N_2754,N_2490,N_2527);
and U2755 (N_2755,N_2523,N_2551);
or U2756 (N_2756,N_2446,N_2578);
and U2757 (N_2757,N_2404,N_2585);
or U2758 (N_2758,N_2491,N_2401);
xnor U2759 (N_2759,N_2412,N_2592);
nand U2760 (N_2760,N_2526,N_2529);
nor U2761 (N_2761,N_2497,N_2539);
and U2762 (N_2762,N_2470,N_2512);
xnor U2763 (N_2763,N_2411,N_2440);
nor U2764 (N_2764,N_2580,N_2485);
nand U2765 (N_2765,N_2496,N_2489);
or U2766 (N_2766,N_2523,N_2418);
nand U2767 (N_2767,N_2512,N_2408);
xnor U2768 (N_2768,N_2535,N_2417);
nand U2769 (N_2769,N_2544,N_2511);
nand U2770 (N_2770,N_2538,N_2595);
xor U2771 (N_2771,N_2547,N_2493);
and U2772 (N_2772,N_2486,N_2578);
nor U2773 (N_2773,N_2579,N_2520);
and U2774 (N_2774,N_2599,N_2557);
or U2775 (N_2775,N_2479,N_2439);
nand U2776 (N_2776,N_2478,N_2429);
nor U2777 (N_2777,N_2543,N_2588);
nor U2778 (N_2778,N_2501,N_2472);
nand U2779 (N_2779,N_2403,N_2566);
xor U2780 (N_2780,N_2549,N_2570);
nand U2781 (N_2781,N_2534,N_2593);
or U2782 (N_2782,N_2450,N_2557);
xor U2783 (N_2783,N_2559,N_2441);
nand U2784 (N_2784,N_2404,N_2590);
nor U2785 (N_2785,N_2461,N_2483);
or U2786 (N_2786,N_2415,N_2512);
nor U2787 (N_2787,N_2571,N_2519);
and U2788 (N_2788,N_2501,N_2546);
nand U2789 (N_2789,N_2477,N_2530);
nand U2790 (N_2790,N_2509,N_2420);
xor U2791 (N_2791,N_2453,N_2504);
nand U2792 (N_2792,N_2538,N_2516);
or U2793 (N_2793,N_2591,N_2516);
xor U2794 (N_2794,N_2556,N_2469);
or U2795 (N_2795,N_2558,N_2536);
and U2796 (N_2796,N_2571,N_2441);
xor U2797 (N_2797,N_2512,N_2419);
or U2798 (N_2798,N_2590,N_2424);
and U2799 (N_2799,N_2496,N_2430);
and U2800 (N_2800,N_2635,N_2694);
or U2801 (N_2801,N_2678,N_2703);
or U2802 (N_2802,N_2711,N_2627);
and U2803 (N_2803,N_2710,N_2672);
or U2804 (N_2804,N_2731,N_2713);
xnor U2805 (N_2805,N_2773,N_2641);
or U2806 (N_2806,N_2708,N_2698);
xor U2807 (N_2807,N_2646,N_2718);
nor U2808 (N_2808,N_2729,N_2722);
nand U2809 (N_2809,N_2670,N_2676);
or U2810 (N_2810,N_2606,N_2648);
xnor U2811 (N_2811,N_2747,N_2687);
and U2812 (N_2812,N_2787,N_2780);
nor U2813 (N_2813,N_2732,N_2782);
and U2814 (N_2814,N_2629,N_2727);
nor U2815 (N_2815,N_2626,N_2684);
nor U2816 (N_2816,N_2734,N_2697);
and U2817 (N_2817,N_2612,N_2602);
nor U2818 (N_2818,N_2701,N_2771);
or U2819 (N_2819,N_2749,N_2705);
or U2820 (N_2820,N_2737,N_2762);
xnor U2821 (N_2821,N_2791,N_2797);
nand U2822 (N_2822,N_2743,N_2784);
and U2823 (N_2823,N_2746,N_2764);
or U2824 (N_2824,N_2654,N_2742);
and U2825 (N_2825,N_2643,N_2664);
and U2826 (N_2826,N_2666,N_2733);
nand U2827 (N_2827,N_2653,N_2618);
xnor U2828 (N_2828,N_2695,N_2691);
xnor U2829 (N_2829,N_2735,N_2677);
or U2830 (N_2830,N_2604,N_2645);
and U2831 (N_2831,N_2686,N_2603);
xor U2832 (N_2832,N_2615,N_2776);
xor U2833 (N_2833,N_2652,N_2725);
nor U2834 (N_2834,N_2685,N_2779);
or U2835 (N_2835,N_2763,N_2706);
xor U2836 (N_2836,N_2611,N_2744);
or U2837 (N_2837,N_2667,N_2794);
xnor U2838 (N_2838,N_2623,N_2638);
nor U2839 (N_2839,N_2688,N_2689);
xnor U2840 (N_2840,N_2739,N_2690);
or U2841 (N_2841,N_2683,N_2620);
or U2842 (N_2842,N_2745,N_2757);
nor U2843 (N_2843,N_2616,N_2799);
and U2844 (N_2844,N_2783,N_2786);
nand U2845 (N_2845,N_2637,N_2750);
or U2846 (N_2846,N_2658,N_2649);
or U2847 (N_2847,N_2702,N_2723);
and U2848 (N_2848,N_2753,N_2625);
and U2849 (N_2849,N_2761,N_2659);
or U2850 (N_2850,N_2774,N_2600);
nor U2851 (N_2851,N_2741,N_2639);
nor U2852 (N_2852,N_2704,N_2700);
nor U2853 (N_2853,N_2693,N_2751);
nor U2854 (N_2854,N_2756,N_2696);
xor U2855 (N_2855,N_2699,N_2647);
and U2856 (N_2856,N_2714,N_2798);
xor U2857 (N_2857,N_2709,N_2631);
xor U2858 (N_2858,N_2622,N_2657);
and U2859 (N_2859,N_2665,N_2765);
xor U2860 (N_2860,N_2717,N_2621);
and U2861 (N_2861,N_2632,N_2758);
or U2862 (N_2862,N_2682,N_2795);
xor U2863 (N_2863,N_2719,N_2777);
nor U2864 (N_2864,N_2755,N_2634);
nor U2865 (N_2865,N_2721,N_2679);
xor U2866 (N_2866,N_2692,N_2644);
nor U2867 (N_2867,N_2778,N_2740);
and U2868 (N_2868,N_2720,N_2673);
or U2869 (N_2869,N_2605,N_2770);
nor U2870 (N_2870,N_2661,N_2716);
nand U2871 (N_2871,N_2788,N_2752);
xor U2872 (N_2872,N_2608,N_2663);
nand U2873 (N_2873,N_2650,N_2681);
xnor U2874 (N_2874,N_2724,N_2772);
and U2875 (N_2875,N_2712,N_2607);
nor U2876 (N_2876,N_2748,N_2789);
nor U2877 (N_2877,N_2726,N_2660);
nand U2878 (N_2878,N_2617,N_2760);
or U2879 (N_2879,N_2640,N_2736);
xor U2880 (N_2880,N_2636,N_2781);
or U2881 (N_2881,N_2609,N_2668);
or U2882 (N_2882,N_2790,N_2680);
nand U2883 (N_2883,N_2796,N_2651);
or U2884 (N_2884,N_2759,N_2766);
nand U2885 (N_2885,N_2793,N_2610);
or U2886 (N_2886,N_2662,N_2754);
xor U2887 (N_2887,N_2669,N_2728);
xor U2888 (N_2888,N_2630,N_2785);
xor U2889 (N_2889,N_2613,N_2671);
or U2890 (N_2890,N_2619,N_2642);
nand U2891 (N_2891,N_2675,N_2768);
nand U2892 (N_2892,N_2775,N_2769);
nor U2893 (N_2893,N_2601,N_2633);
or U2894 (N_2894,N_2715,N_2707);
nor U2895 (N_2895,N_2674,N_2730);
xnor U2896 (N_2896,N_2614,N_2656);
xnor U2897 (N_2897,N_2655,N_2624);
nand U2898 (N_2898,N_2738,N_2792);
or U2899 (N_2899,N_2767,N_2628);
xnor U2900 (N_2900,N_2653,N_2644);
or U2901 (N_2901,N_2799,N_2679);
nor U2902 (N_2902,N_2661,N_2756);
and U2903 (N_2903,N_2695,N_2733);
and U2904 (N_2904,N_2629,N_2736);
nand U2905 (N_2905,N_2728,N_2726);
or U2906 (N_2906,N_2620,N_2759);
xor U2907 (N_2907,N_2754,N_2674);
xor U2908 (N_2908,N_2716,N_2671);
and U2909 (N_2909,N_2771,N_2601);
nand U2910 (N_2910,N_2635,N_2748);
nor U2911 (N_2911,N_2626,N_2672);
xnor U2912 (N_2912,N_2698,N_2783);
nor U2913 (N_2913,N_2635,N_2711);
and U2914 (N_2914,N_2732,N_2747);
nor U2915 (N_2915,N_2766,N_2661);
nor U2916 (N_2916,N_2710,N_2740);
xor U2917 (N_2917,N_2602,N_2730);
nor U2918 (N_2918,N_2611,N_2764);
and U2919 (N_2919,N_2799,N_2625);
nor U2920 (N_2920,N_2648,N_2708);
and U2921 (N_2921,N_2710,N_2605);
or U2922 (N_2922,N_2792,N_2747);
xor U2923 (N_2923,N_2797,N_2793);
and U2924 (N_2924,N_2688,N_2626);
and U2925 (N_2925,N_2705,N_2771);
or U2926 (N_2926,N_2740,N_2763);
or U2927 (N_2927,N_2691,N_2655);
nand U2928 (N_2928,N_2631,N_2645);
or U2929 (N_2929,N_2753,N_2794);
nor U2930 (N_2930,N_2601,N_2647);
and U2931 (N_2931,N_2663,N_2777);
nand U2932 (N_2932,N_2766,N_2648);
nand U2933 (N_2933,N_2735,N_2682);
nand U2934 (N_2934,N_2602,N_2760);
nor U2935 (N_2935,N_2713,N_2657);
or U2936 (N_2936,N_2692,N_2610);
or U2937 (N_2937,N_2616,N_2694);
xnor U2938 (N_2938,N_2677,N_2624);
or U2939 (N_2939,N_2640,N_2606);
and U2940 (N_2940,N_2777,N_2781);
or U2941 (N_2941,N_2713,N_2649);
xor U2942 (N_2942,N_2670,N_2799);
nand U2943 (N_2943,N_2753,N_2680);
and U2944 (N_2944,N_2673,N_2674);
or U2945 (N_2945,N_2689,N_2728);
and U2946 (N_2946,N_2677,N_2784);
nor U2947 (N_2947,N_2698,N_2735);
nor U2948 (N_2948,N_2772,N_2710);
and U2949 (N_2949,N_2660,N_2667);
xor U2950 (N_2950,N_2728,N_2655);
nor U2951 (N_2951,N_2616,N_2747);
xor U2952 (N_2952,N_2642,N_2624);
nor U2953 (N_2953,N_2602,N_2790);
and U2954 (N_2954,N_2712,N_2794);
and U2955 (N_2955,N_2735,N_2762);
nor U2956 (N_2956,N_2675,N_2645);
nor U2957 (N_2957,N_2727,N_2631);
and U2958 (N_2958,N_2771,N_2653);
nor U2959 (N_2959,N_2625,N_2722);
or U2960 (N_2960,N_2795,N_2670);
nor U2961 (N_2961,N_2643,N_2750);
or U2962 (N_2962,N_2640,N_2783);
or U2963 (N_2963,N_2698,N_2764);
xnor U2964 (N_2964,N_2706,N_2653);
and U2965 (N_2965,N_2657,N_2681);
xor U2966 (N_2966,N_2760,N_2750);
nor U2967 (N_2967,N_2699,N_2687);
nand U2968 (N_2968,N_2679,N_2739);
or U2969 (N_2969,N_2747,N_2607);
and U2970 (N_2970,N_2720,N_2614);
nand U2971 (N_2971,N_2625,N_2796);
and U2972 (N_2972,N_2661,N_2767);
nor U2973 (N_2973,N_2625,N_2789);
nand U2974 (N_2974,N_2761,N_2781);
nor U2975 (N_2975,N_2633,N_2670);
xnor U2976 (N_2976,N_2640,N_2684);
and U2977 (N_2977,N_2690,N_2651);
and U2978 (N_2978,N_2673,N_2614);
nand U2979 (N_2979,N_2706,N_2643);
nand U2980 (N_2980,N_2764,N_2657);
xor U2981 (N_2981,N_2694,N_2649);
and U2982 (N_2982,N_2705,N_2737);
nand U2983 (N_2983,N_2713,N_2703);
nor U2984 (N_2984,N_2628,N_2649);
or U2985 (N_2985,N_2764,N_2629);
nand U2986 (N_2986,N_2761,N_2758);
or U2987 (N_2987,N_2784,N_2645);
or U2988 (N_2988,N_2777,N_2718);
xor U2989 (N_2989,N_2734,N_2648);
and U2990 (N_2990,N_2656,N_2658);
nor U2991 (N_2991,N_2739,N_2719);
or U2992 (N_2992,N_2773,N_2795);
or U2993 (N_2993,N_2694,N_2626);
nand U2994 (N_2994,N_2693,N_2625);
xor U2995 (N_2995,N_2727,N_2630);
nand U2996 (N_2996,N_2604,N_2630);
xor U2997 (N_2997,N_2648,N_2730);
nor U2998 (N_2998,N_2784,N_2793);
and U2999 (N_2999,N_2789,N_2774);
nand U3000 (N_3000,N_2909,N_2817);
nor U3001 (N_3001,N_2904,N_2920);
and U3002 (N_3002,N_2905,N_2981);
nand U3003 (N_3003,N_2808,N_2853);
xnor U3004 (N_3004,N_2991,N_2851);
and U3005 (N_3005,N_2875,N_2941);
nor U3006 (N_3006,N_2839,N_2939);
nand U3007 (N_3007,N_2840,N_2878);
and U3008 (N_3008,N_2935,N_2982);
or U3009 (N_3009,N_2956,N_2934);
nor U3010 (N_3010,N_2940,N_2830);
nand U3011 (N_3011,N_2859,N_2983);
nor U3012 (N_3012,N_2881,N_2845);
and U3013 (N_3013,N_2907,N_2973);
xnor U3014 (N_3014,N_2911,N_2959);
or U3015 (N_3015,N_2996,N_2919);
or U3016 (N_3016,N_2899,N_2971);
and U3017 (N_3017,N_2949,N_2995);
xnor U3018 (N_3018,N_2962,N_2898);
and U3019 (N_3019,N_2832,N_2879);
nand U3020 (N_3020,N_2882,N_2812);
or U3021 (N_3021,N_2821,N_2979);
and U3022 (N_3022,N_2886,N_2809);
nor U3023 (N_3023,N_2970,N_2855);
or U3024 (N_3024,N_2997,N_2837);
nand U3025 (N_3025,N_2813,N_2807);
or U3026 (N_3026,N_2926,N_2893);
and U3027 (N_3027,N_2819,N_2924);
and U3028 (N_3028,N_2804,N_2923);
xnor U3029 (N_3029,N_2922,N_2987);
or U3030 (N_3030,N_2890,N_2968);
or U3031 (N_3031,N_2884,N_2969);
xor U3032 (N_3032,N_2883,N_2810);
xnor U3033 (N_3033,N_2918,N_2960);
or U3034 (N_3034,N_2906,N_2929);
xnor U3035 (N_3035,N_2823,N_2865);
xnor U3036 (N_3036,N_2989,N_2877);
nand U3037 (N_3037,N_2897,N_2966);
or U3038 (N_3038,N_2938,N_2847);
nor U3039 (N_3039,N_2901,N_2867);
or U3040 (N_3040,N_2834,N_2955);
and U3041 (N_3041,N_2892,N_2931);
nor U3042 (N_3042,N_2836,N_2951);
and U3043 (N_3043,N_2833,N_2914);
or U3044 (N_3044,N_2858,N_2930);
nand U3045 (N_3045,N_2888,N_2862);
xnor U3046 (N_3046,N_2903,N_2999);
xor U3047 (N_3047,N_2811,N_2988);
nand U3048 (N_3048,N_2975,N_2946);
xnor U3049 (N_3049,N_2976,N_2835);
or U3050 (N_3050,N_2844,N_2826);
nand U3051 (N_3051,N_2933,N_2871);
xnor U3052 (N_3052,N_2803,N_2885);
xor U3053 (N_3053,N_2985,N_2992);
nand U3054 (N_3054,N_2829,N_2891);
nor U3055 (N_3055,N_2980,N_2954);
xor U3056 (N_3056,N_2876,N_2921);
or U3057 (N_3057,N_2814,N_2852);
nand U3058 (N_3058,N_2986,N_2850);
nand U3059 (N_3059,N_2869,N_2972);
or U3060 (N_3060,N_2942,N_2843);
nor U3061 (N_3061,N_2947,N_2857);
or U3062 (N_3062,N_2902,N_2831);
or U3063 (N_3063,N_2964,N_2896);
xnor U3064 (N_3064,N_2838,N_2864);
or U3065 (N_3065,N_2846,N_2894);
or U3066 (N_3066,N_2863,N_2880);
nor U3067 (N_3067,N_2910,N_2873);
nand U3068 (N_3068,N_2827,N_2945);
xnor U3069 (N_3069,N_2990,N_2872);
nor U3070 (N_3070,N_2856,N_2908);
and U3071 (N_3071,N_2870,N_2801);
and U3072 (N_3072,N_2825,N_2944);
and U3073 (N_3073,N_2822,N_2861);
nand U3074 (N_3074,N_2828,N_2913);
nor U3075 (N_3075,N_2974,N_2800);
nand U3076 (N_3076,N_2977,N_2937);
nor U3077 (N_3077,N_2965,N_2887);
xnor U3078 (N_3078,N_2915,N_2998);
and U3079 (N_3079,N_2841,N_2818);
nand U3080 (N_3080,N_2994,N_2805);
or U3081 (N_3081,N_2860,N_2993);
or U3082 (N_3082,N_2868,N_2932);
nand U3083 (N_3083,N_2889,N_2820);
or U3084 (N_3084,N_2963,N_2948);
or U3085 (N_3085,N_2806,N_2928);
and U3086 (N_3086,N_2936,N_2815);
xnor U3087 (N_3087,N_2950,N_2900);
and U3088 (N_3088,N_2957,N_2925);
and U3089 (N_3089,N_2953,N_2816);
and U3090 (N_3090,N_2961,N_2848);
and U3091 (N_3091,N_2895,N_2916);
xor U3092 (N_3092,N_2967,N_2912);
nand U3093 (N_3093,N_2866,N_2824);
nand U3094 (N_3094,N_2917,N_2802);
or U3095 (N_3095,N_2952,N_2874);
and U3096 (N_3096,N_2842,N_2854);
xnor U3097 (N_3097,N_2927,N_2849);
xor U3098 (N_3098,N_2958,N_2978);
and U3099 (N_3099,N_2943,N_2984);
nor U3100 (N_3100,N_2980,N_2905);
and U3101 (N_3101,N_2809,N_2926);
nand U3102 (N_3102,N_2874,N_2842);
xnor U3103 (N_3103,N_2844,N_2813);
xnor U3104 (N_3104,N_2961,N_2922);
and U3105 (N_3105,N_2944,N_2853);
and U3106 (N_3106,N_2849,N_2923);
xor U3107 (N_3107,N_2965,N_2828);
or U3108 (N_3108,N_2990,N_2976);
nor U3109 (N_3109,N_2985,N_2957);
xor U3110 (N_3110,N_2874,N_2959);
nand U3111 (N_3111,N_2825,N_2935);
nor U3112 (N_3112,N_2960,N_2943);
or U3113 (N_3113,N_2865,N_2857);
xor U3114 (N_3114,N_2818,N_2927);
or U3115 (N_3115,N_2828,N_2807);
xnor U3116 (N_3116,N_2919,N_2807);
xor U3117 (N_3117,N_2908,N_2900);
and U3118 (N_3118,N_2924,N_2874);
nand U3119 (N_3119,N_2842,N_2815);
nor U3120 (N_3120,N_2960,N_2908);
xor U3121 (N_3121,N_2967,N_2959);
xor U3122 (N_3122,N_2921,N_2843);
xnor U3123 (N_3123,N_2874,N_2906);
nand U3124 (N_3124,N_2802,N_2850);
nand U3125 (N_3125,N_2813,N_2949);
and U3126 (N_3126,N_2884,N_2831);
and U3127 (N_3127,N_2808,N_2809);
or U3128 (N_3128,N_2847,N_2876);
nor U3129 (N_3129,N_2896,N_2971);
and U3130 (N_3130,N_2971,N_2815);
nor U3131 (N_3131,N_2884,N_2995);
nand U3132 (N_3132,N_2873,N_2822);
nor U3133 (N_3133,N_2835,N_2944);
nor U3134 (N_3134,N_2809,N_2876);
xor U3135 (N_3135,N_2984,N_2877);
nor U3136 (N_3136,N_2974,N_2888);
nor U3137 (N_3137,N_2817,N_2807);
xnor U3138 (N_3138,N_2941,N_2988);
nand U3139 (N_3139,N_2827,N_2927);
or U3140 (N_3140,N_2900,N_2833);
xnor U3141 (N_3141,N_2928,N_2955);
nor U3142 (N_3142,N_2881,N_2926);
nand U3143 (N_3143,N_2976,N_2937);
xnor U3144 (N_3144,N_2889,N_2864);
and U3145 (N_3145,N_2968,N_2964);
xnor U3146 (N_3146,N_2915,N_2954);
nor U3147 (N_3147,N_2920,N_2964);
and U3148 (N_3148,N_2834,N_2858);
nand U3149 (N_3149,N_2952,N_2811);
and U3150 (N_3150,N_2915,N_2860);
or U3151 (N_3151,N_2974,N_2928);
and U3152 (N_3152,N_2987,N_2911);
nand U3153 (N_3153,N_2903,N_2828);
or U3154 (N_3154,N_2800,N_2828);
or U3155 (N_3155,N_2928,N_2850);
or U3156 (N_3156,N_2940,N_2833);
nand U3157 (N_3157,N_2969,N_2979);
or U3158 (N_3158,N_2928,N_2914);
nor U3159 (N_3159,N_2887,N_2801);
and U3160 (N_3160,N_2810,N_2966);
or U3161 (N_3161,N_2867,N_2845);
nor U3162 (N_3162,N_2956,N_2936);
nor U3163 (N_3163,N_2834,N_2992);
nor U3164 (N_3164,N_2951,N_2835);
xnor U3165 (N_3165,N_2927,N_2931);
or U3166 (N_3166,N_2951,N_2863);
and U3167 (N_3167,N_2900,N_2841);
or U3168 (N_3168,N_2956,N_2969);
or U3169 (N_3169,N_2800,N_2872);
and U3170 (N_3170,N_2901,N_2829);
nor U3171 (N_3171,N_2970,N_2954);
nand U3172 (N_3172,N_2844,N_2881);
nand U3173 (N_3173,N_2817,N_2955);
or U3174 (N_3174,N_2986,N_2985);
or U3175 (N_3175,N_2875,N_2912);
nor U3176 (N_3176,N_2838,N_2960);
nand U3177 (N_3177,N_2912,N_2897);
or U3178 (N_3178,N_2909,N_2807);
and U3179 (N_3179,N_2822,N_2836);
nand U3180 (N_3180,N_2940,N_2818);
and U3181 (N_3181,N_2907,N_2919);
xor U3182 (N_3182,N_2888,N_2928);
and U3183 (N_3183,N_2956,N_2913);
nand U3184 (N_3184,N_2932,N_2897);
or U3185 (N_3185,N_2948,N_2804);
xor U3186 (N_3186,N_2858,N_2964);
and U3187 (N_3187,N_2962,N_2952);
and U3188 (N_3188,N_2921,N_2989);
or U3189 (N_3189,N_2801,N_2989);
nor U3190 (N_3190,N_2807,N_2816);
and U3191 (N_3191,N_2962,N_2817);
nor U3192 (N_3192,N_2871,N_2824);
nand U3193 (N_3193,N_2956,N_2945);
or U3194 (N_3194,N_2804,N_2906);
and U3195 (N_3195,N_2928,N_2962);
xor U3196 (N_3196,N_2825,N_2889);
nor U3197 (N_3197,N_2899,N_2993);
and U3198 (N_3198,N_2939,N_2942);
nand U3199 (N_3199,N_2848,N_2947);
and U3200 (N_3200,N_3085,N_3147);
nor U3201 (N_3201,N_3014,N_3083);
nand U3202 (N_3202,N_3159,N_3132);
nand U3203 (N_3203,N_3035,N_3011);
xnor U3204 (N_3204,N_3045,N_3198);
and U3205 (N_3205,N_3195,N_3025);
nor U3206 (N_3206,N_3193,N_3057);
or U3207 (N_3207,N_3197,N_3016);
or U3208 (N_3208,N_3033,N_3115);
xor U3209 (N_3209,N_3126,N_3114);
and U3210 (N_3210,N_3120,N_3130);
and U3211 (N_3211,N_3189,N_3020);
nand U3212 (N_3212,N_3070,N_3122);
nor U3213 (N_3213,N_3173,N_3190);
nand U3214 (N_3214,N_3111,N_3178);
or U3215 (N_3215,N_3087,N_3041);
xnor U3216 (N_3216,N_3116,N_3082);
nand U3217 (N_3217,N_3187,N_3047);
nor U3218 (N_3218,N_3053,N_3103);
nor U3219 (N_3219,N_3007,N_3001);
xnor U3220 (N_3220,N_3167,N_3142);
or U3221 (N_3221,N_3086,N_3068);
nand U3222 (N_3222,N_3042,N_3181);
nand U3223 (N_3223,N_3049,N_3029);
and U3224 (N_3224,N_3145,N_3133);
xnor U3225 (N_3225,N_3196,N_3139);
or U3226 (N_3226,N_3165,N_3146);
and U3227 (N_3227,N_3191,N_3008);
nor U3228 (N_3228,N_3121,N_3168);
xnor U3229 (N_3229,N_3162,N_3136);
nor U3230 (N_3230,N_3158,N_3022);
or U3231 (N_3231,N_3100,N_3038);
nor U3232 (N_3232,N_3170,N_3063);
xor U3233 (N_3233,N_3036,N_3096);
or U3234 (N_3234,N_3175,N_3177);
xnor U3235 (N_3235,N_3051,N_3043);
or U3236 (N_3236,N_3023,N_3015);
and U3237 (N_3237,N_3027,N_3194);
and U3238 (N_3238,N_3021,N_3060);
and U3239 (N_3239,N_3143,N_3140);
nor U3240 (N_3240,N_3095,N_3090);
nor U3241 (N_3241,N_3138,N_3163);
xnor U3242 (N_3242,N_3006,N_3108);
or U3243 (N_3243,N_3172,N_3135);
or U3244 (N_3244,N_3056,N_3012);
and U3245 (N_3245,N_3066,N_3048);
and U3246 (N_3246,N_3094,N_3032);
nor U3247 (N_3247,N_3131,N_3176);
or U3248 (N_3248,N_3149,N_3064);
or U3249 (N_3249,N_3185,N_3044);
nand U3250 (N_3250,N_3153,N_3157);
or U3251 (N_3251,N_3052,N_3169);
and U3252 (N_3252,N_3099,N_3156);
xnor U3253 (N_3253,N_3166,N_3039);
or U3254 (N_3254,N_3088,N_3151);
xor U3255 (N_3255,N_3071,N_3091);
xnor U3256 (N_3256,N_3188,N_3124);
xor U3257 (N_3257,N_3125,N_3005);
nand U3258 (N_3258,N_3002,N_3079);
nor U3259 (N_3259,N_3019,N_3192);
or U3260 (N_3260,N_3065,N_3104);
and U3261 (N_3261,N_3127,N_3113);
nand U3262 (N_3262,N_3102,N_3031);
or U3263 (N_3263,N_3017,N_3141);
nor U3264 (N_3264,N_3078,N_3093);
nand U3265 (N_3265,N_3034,N_3073);
xnor U3266 (N_3266,N_3069,N_3046);
and U3267 (N_3267,N_3084,N_3098);
nand U3268 (N_3268,N_3128,N_3097);
nand U3269 (N_3269,N_3199,N_3081);
or U3270 (N_3270,N_3186,N_3129);
nand U3271 (N_3271,N_3101,N_3003);
nand U3272 (N_3272,N_3160,N_3010);
and U3273 (N_3273,N_3055,N_3054);
and U3274 (N_3274,N_3004,N_3144);
or U3275 (N_3275,N_3164,N_3092);
xor U3276 (N_3276,N_3076,N_3174);
nor U3277 (N_3277,N_3182,N_3062);
and U3278 (N_3278,N_3150,N_3080);
nand U3279 (N_3279,N_3154,N_3067);
and U3280 (N_3280,N_3118,N_3119);
and U3281 (N_3281,N_3018,N_3161);
nand U3282 (N_3282,N_3180,N_3171);
nand U3283 (N_3283,N_3037,N_3106);
nor U3284 (N_3284,N_3028,N_3179);
xnor U3285 (N_3285,N_3109,N_3077);
xor U3286 (N_3286,N_3026,N_3112);
nand U3287 (N_3287,N_3030,N_3058);
nor U3288 (N_3288,N_3013,N_3024);
nand U3289 (N_3289,N_3183,N_3075);
nor U3290 (N_3290,N_3123,N_3155);
xor U3291 (N_3291,N_3009,N_3110);
xnor U3292 (N_3292,N_3000,N_3152);
nor U3293 (N_3293,N_3107,N_3184);
nor U3294 (N_3294,N_3148,N_3089);
nand U3295 (N_3295,N_3059,N_3105);
nor U3296 (N_3296,N_3074,N_3072);
and U3297 (N_3297,N_3134,N_3050);
nand U3298 (N_3298,N_3040,N_3061);
xnor U3299 (N_3299,N_3137,N_3117);
and U3300 (N_3300,N_3143,N_3106);
nor U3301 (N_3301,N_3028,N_3052);
and U3302 (N_3302,N_3006,N_3067);
or U3303 (N_3303,N_3011,N_3184);
nand U3304 (N_3304,N_3005,N_3175);
and U3305 (N_3305,N_3149,N_3061);
nor U3306 (N_3306,N_3151,N_3067);
or U3307 (N_3307,N_3107,N_3049);
or U3308 (N_3308,N_3041,N_3006);
or U3309 (N_3309,N_3184,N_3052);
xor U3310 (N_3310,N_3185,N_3193);
and U3311 (N_3311,N_3020,N_3103);
nor U3312 (N_3312,N_3056,N_3045);
and U3313 (N_3313,N_3058,N_3089);
xnor U3314 (N_3314,N_3193,N_3067);
xor U3315 (N_3315,N_3035,N_3191);
or U3316 (N_3316,N_3031,N_3054);
or U3317 (N_3317,N_3192,N_3197);
and U3318 (N_3318,N_3178,N_3108);
and U3319 (N_3319,N_3125,N_3046);
nand U3320 (N_3320,N_3064,N_3116);
and U3321 (N_3321,N_3009,N_3096);
and U3322 (N_3322,N_3068,N_3083);
and U3323 (N_3323,N_3143,N_3074);
xnor U3324 (N_3324,N_3134,N_3017);
nand U3325 (N_3325,N_3093,N_3161);
nor U3326 (N_3326,N_3118,N_3022);
nor U3327 (N_3327,N_3123,N_3050);
nor U3328 (N_3328,N_3069,N_3120);
or U3329 (N_3329,N_3130,N_3189);
or U3330 (N_3330,N_3087,N_3069);
nand U3331 (N_3331,N_3194,N_3010);
xnor U3332 (N_3332,N_3060,N_3026);
or U3333 (N_3333,N_3107,N_3094);
xnor U3334 (N_3334,N_3039,N_3170);
and U3335 (N_3335,N_3105,N_3129);
nor U3336 (N_3336,N_3157,N_3180);
or U3337 (N_3337,N_3183,N_3005);
or U3338 (N_3338,N_3136,N_3053);
nand U3339 (N_3339,N_3169,N_3144);
xor U3340 (N_3340,N_3150,N_3033);
xor U3341 (N_3341,N_3098,N_3036);
nand U3342 (N_3342,N_3032,N_3055);
nor U3343 (N_3343,N_3066,N_3108);
or U3344 (N_3344,N_3108,N_3198);
xor U3345 (N_3345,N_3112,N_3151);
nand U3346 (N_3346,N_3003,N_3039);
xor U3347 (N_3347,N_3161,N_3198);
xor U3348 (N_3348,N_3012,N_3136);
nor U3349 (N_3349,N_3160,N_3167);
xnor U3350 (N_3350,N_3016,N_3012);
nor U3351 (N_3351,N_3033,N_3139);
and U3352 (N_3352,N_3030,N_3187);
xnor U3353 (N_3353,N_3135,N_3125);
nor U3354 (N_3354,N_3105,N_3048);
and U3355 (N_3355,N_3154,N_3095);
and U3356 (N_3356,N_3192,N_3070);
nand U3357 (N_3357,N_3125,N_3025);
and U3358 (N_3358,N_3057,N_3157);
and U3359 (N_3359,N_3181,N_3066);
nand U3360 (N_3360,N_3141,N_3142);
xnor U3361 (N_3361,N_3141,N_3008);
nor U3362 (N_3362,N_3052,N_3199);
xnor U3363 (N_3363,N_3033,N_3198);
or U3364 (N_3364,N_3174,N_3170);
xor U3365 (N_3365,N_3177,N_3032);
and U3366 (N_3366,N_3168,N_3056);
xnor U3367 (N_3367,N_3108,N_3186);
xnor U3368 (N_3368,N_3028,N_3043);
and U3369 (N_3369,N_3113,N_3002);
or U3370 (N_3370,N_3157,N_3058);
xor U3371 (N_3371,N_3112,N_3196);
or U3372 (N_3372,N_3163,N_3151);
or U3373 (N_3373,N_3154,N_3016);
nand U3374 (N_3374,N_3186,N_3029);
xor U3375 (N_3375,N_3094,N_3133);
and U3376 (N_3376,N_3065,N_3055);
nand U3377 (N_3377,N_3122,N_3199);
nor U3378 (N_3378,N_3099,N_3072);
xnor U3379 (N_3379,N_3015,N_3003);
or U3380 (N_3380,N_3182,N_3024);
and U3381 (N_3381,N_3106,N_3183);
nor U3382 (N_3382,N_3058,N_3135);
nor U3383 (N_3383,N_3010,N_3018);
nor U3384 (N_3384,N_3008,N_3046);
nor U3385 (N_3385,N_3028,N_3198);
nor U3386 (N_3386,N_3054,N_3165);
and U3387 (N_3387,N_3038,N_3181);
and U3388 (N_3388,N_3166,N_3005);
or U3389 (N_3389,N_3198,N_3012);
and U3390 (N_3390,N_3066,N_3018);
and U3391 (N_3391,N_3189,N_3137);
nor U3392 (N_3392,N_3157,N_3085);
nand U3393 (N_3393,N_3148,N_3191);
or U3394 (N_3394,N_3063,N_3000);
nand U3395 (N_3395,N_3005,N_3143);
xnor U3396 (N_3396,N_3198,N_3169);
and U3397 (N_3397,N_3188,N_3119);
and U3398 (N_3398,N_3136,N_3154);
nor U3399 (N_3399,N_3086,N_3158);
nand U3400 (N_3400,N_3300,N_3238);
nor U3401 (N_3401,N_3389,N_3381);
nand U3402 (N_3402,N_3379,N_3334);
and U3403 (N_3403,N_3348,N_3222);
and U3404 (N_3404,N_3245,N_3362);
or U3405 (N_3405,N_3296,N_3380);
nand U3406 (N_3406,N_3292,N_3359);
or U3407 (N_3407,N_3237,N_3270);
nor U3408 (N_3408,N_3304,N_3263);
xnor U3409 (N_3409,N_3282,N_3204);
nand U3410 (N_3410,N_3347,N_3374);
or U3411 (N_3411,N_3322,N_3349);
nor U3412 (N_3412,N_3303,N_3258);
and U3413 (N_3413,N_3345,N_3317);
and U3414 (N_3414,N_3257,N_3360);
xor U3415 (N_3415,N_3249,N_3235);
xor U3416 (N_3416,N_3221,N_3210);
or U3417 (N_3417,N_3329,N_3307);
nand U3418 (N_3418,N_3243,N_3261);
or U3419 (N_3419,N_3295,N_3248);
nor U3420 (N_3420,N_3352,N_3276);
nor U3421 (N_3421,N_3217,N_3285);
and U3422 (N_3422,N_3337,N_3393);
xor U3423 (N_3423,N_3355,N_3211);
or U3424 (N_3424,N_3284,N_3223);
xor U3425 (N_3425,N_3364,N_3318);
nand U3426 (N_3426,N_3226,N_3251);
nand U3427 (N_3427,N_3325,N_3346);
nand U3428 (N_3428,N_3290,N_3373);
nand U3429 (N_3429,N_3395,N_3240);
nor U3430 (N_3430,N_3225,N_3365);
or U3431 (N_3431,N_3377,N_3326);
xor U3432 (N_3432,N_3394,N_3219);
nor U3433 (N_3433,N_3302,N_3305);
or U3434 (N_3434,N_3202,N_3227);
xnor U3435 (N_3435,N_3336,N_3330);
xor U3436 (N_3436,N_3264,N_3387);
or U3437 (N_3437,N_3321,N_3333);
nand U3438 (N_3438,N_3340,N_3378);
and U3439 (N_3439,N_3372,N_3254);
nand U3440 (N_3440,N_3200,N_3239);
nand U3441 (N_3441,N_3272,N_3324);
nand U3442 (N_3442,N_3207,N_3370);
nand U3443 (N_3443,N_3286,N_3242);
nor U3444 (N_3444,N_3259,N_3354);
nand U3445 (N_3445,N_3338,N_3383);
nor U3446 (N_3446,N_3265,N_3301);
and U3447 (N_3447,N_3241,N_3375);
and U3448 (N_3448,N_3320,N_3234);
or U3449 (N_3449,N_3312,N_3368);
or U3450 (N_3450,N_3294,N_3201);
or U3451 (N_3451,N_3203,N_3213);
nand U3452 (N_3452,N_3246,N_3310);
and U3453 (N_3453,N_3319,N_3357);
nor U3454 (N_3454,N_3311,N_3356);
and U3455 (N_3455,N_3262,N_3371);
and U3456 (N_3456,N_3343,N_3396);
nand U3457 (N_3457,N_3367,N_3232);
nor U3458 (N_3458,N_3332,N_3266);
and U3459 (N_3459,N_3275,N_3293);
xnor U3460 (N_3460,N_3268,N_3398);
nand U3461 (N_3461,N_3280,N_3218);
nor U3462 (N_3462,N_3236,N_3391);
or U3463 (N_3463,N_3271,N_3224);
and U3464 (N_3464,N_3289,N_3358);
and U3465 (N_3465,N_3327,N_3366);
and U3466 (N_3466,N_3328,N_3350);
nand U3467 (N_3467,N_3388,N_3369);
and U3468 (N_3468,N_3287,N_3313);
nor U3469 (N_3469,N_3291,N_3376);
nand U3470 (N_3470,N_3212,N_3386);
nor U3471 (N_3471,N_3206,N_3215);
xor U3472 (N_3472,N_3309,N_3397);
and U3473 (N_3473,N_3274,N_3230);
and U3474 (N_3474,N_3382,N_3255);
and U3475 (N_3475,N_3233,N_3385);
or U3476 (N_3476,N_3256,N_3344);
xnor U3477 (N_3477,N_3278,N_3273);
nand U3478 (N_3478,N_3253,N_3269);
xor U3479 (N_3479,N_3353,N_3315);
xor U3480 (N_3480,N_3316,N_3247);
and U3481 (N_3481,N_3323,N_3351);
nand U3482 (N_3482,N_3384,N_3214);
nand U3483 (N_3483,N_3229,N_3341);
nand U3484 (N_3484,N_3361,N_3209);
xor U3485 (N_3485,N_3308,N_3390);
nor U3486 (N_3486,N_3216,N_3342);
nor U3487 (N_3487,N_3231,N_3339);
nand U3488 (N_3488,N_3399,N_3306);
and U3489 (N_3489,N_3281,N_3260);
xnor U3490 (N_3490,N_3279,N_3250);
xor U3491 (N_3491,N_3363,N_3205);
nor U3492 (N_3492,N_3392,N_3331);
nand U3493 (N_3493,N_3252,N_3220);
and U3494 (N_3494,N_3208,N_3314);
and U3495 (N_3495,N_3277,N_3267);
nor U3496 (N_3496,N_3244,N_3283);
nand U3497 (N_3497,N_3288,N_3298);
nand U3498 (N_3498,N_3335,N_3228);
nand U3499 (N_3499,N_3297,N_3299);
nand U3500 (N_3500,N_3326,N_3256);
and U3501 (N_3501,N_3371,N_3335);
or U3502 (N_3502,N_3324,N_3323);
xnor U3503 (N_3503,N_3309,N_3286);
nor U3504 (N_3504,N_3329,N_3259);
nor U3505 (N_3505,N_3375,N_3263);
xnor U3506 (N_3506,N_3360,N_3391);
and U3507 (N_3507,N_3303,N_3326);
and U3508 (N_3508,N_3272,N_3347);
nor U3509 (N_3509,N_3321,N_3205);
nand U3510 (N_3510,N_3202,N_3387);
or U3511 (N_3511,N_3338,N_3280);
nand U3512 (N_3512,N_3209,N_3212);
or U3513 (N_3513,N_3305,N_3399);
nand U3514 (N_3514,N_3202,N_3327);
xnor U3515 (N_3515,N_3273,N_3368);
nand U3516 (N_3516,N_3233,N_3286);
nor U3517 (N_3517,N_3347,N_3201);
and U3518 (N_3518,N_3214,N_3299);
and U3519 (N_3519,N_3329,N_3234);
nor U3520 (N_3520,N_3210,N_3376);
xnor U3521 (N_3521,N_3215,N_3246);
xor U3522 (N_3522,N_3203,N_3299);
xor U3523 (N_3523,N_3202,N_3226);
or U3524 (N_3524,N_3355,N_3207);
and U3525 (N_3525,N_3319,N_3343);
xnor U3526 (N_3526,N_3318,N_3289);
xor U3527 (N_3527,N_3224,N_3233);
xor U3528 (N_3528,N_3265,N_3331);
xor U3529 (N_3529,N_3329,N_3380);
nor U3530 (N_3530,N_3247,N_3259);
nand U3531 (N_3531,N_3292,N_3331);
xor U3532 (N_3532,N_3374,N_3244);
nand U3533 (N_3533,N_3319,N_3387);
and U3534 (N_3534,N_3397,N_3222);
nor U3535 (N_3535,N_3303,N_3363);
and U3536 (N_3536,N_3386,N_3246);
and U3537 (N_3537,N_3397,N_3317);
or U3538 (N_3538,N_3238,N_3298);
xor U3539 (N_3539,N_3293,N_3325);
and U3540 (N_3540,N_3386,N_3342);
and U3541 (N_3541,N_3285,N_3208);
nand U3542 (N_3542,N_3372,N_3313);
nor U3543 (N_3543,N_3382,N_3387);
or U3544 (N_3544,N_3225,N_3311);
nand U3545 (N_3545,N_3383,N_3250);
or U3546 (N_3546,N_3367,N_3255);
or U3547 (N_3547,N_3300,N_3365);
nor U3548 (N_3548,N_3266,N_3371);
or U3549 (N_3549,N_3286,N_3331);
nor U3550 (N_3550,N_3276,N_3241);
nand U3551 (N_3551,N_3261,N_3225);
nor U3552 (N_3552,N_3379,N_3319);
or U3553 (N_3553,N_3296,N_3302);
nand U3554 (N_3554,N_3315,N_3324);
xor U3555 (N_3555,N_3236,N_3228);
or U3556 (N_3556,N_3212,N_3326);
or U3557 (N_3557,N_3384,N_3342);
nand U3558 (N_3558,N_3397,N_3242);
nor U3559 (N_3559,N_3238,N_3378);
and U3560 (N_3560,N_3363,N_3228);
nand U3561 (N_3561,N_3268,N_3332);
nand U3562 (N_3562,N_3222,N_3327);
xor U3563 (N_3563,N_3205,N_3314);
nor U3564 (N_3564,N_3340,N_3253);
nor U3565 (N_3565,N_3330,N_3343);
nand U3566 (N_3566,N_3326,N_3209);
nand U3567 (N_3567,N_3387,N_3388);
or U3568 (N_3568,N_3306,N_3272);
or U3569 (N_3569,N_3380,N_3227);
nand U3570 (N_3570,N_3229,N_3238);
nor U3571 (N_3571,N_3346,N_3280);
nor U3572 (N_3572,N_3370,N_3321);
or U3573 (N_3573,N_3366,N_3281);
and U3574 (N_3574,N_3367,N_3294);
or U3575 (N_3575,N_3349,N_3218);
nand U3576 (N_3576,N_3332,N_3390);
nor U3577 (N_3577,N_3224,N_3268);
and U3578 (N_3578,N_3241,N_3253);
nor U3579 (N_3579,N_3236,N_3384);
nor U3580 (N_3580,N_3350,N_3213);
nor U3581 (N_3581,N_3322,N_3260);
nand U3582 (N_3582,N_3383,N_3270);
nor U3583 (N_3583,N_3238,N_3379);
and U3584 (N_3584,N_3244,N_3270);
nand U3585 (N_3585,N_3333,N_3266);
nor U3586 (N_3586,N_3256,N_3279);
or U3587 (N_3587,N_3355,N_3381);
and U3588 (N_3588,N_3344,N_3209);
nor U3589 (N_3589,N_3305,N_3380);
xnor U3590 (N_3590,N_3382,N_3235);
xor U3591 (N_3591,N_3208,N_3366);
nor U3592 (N_3592,N_3222,N_3341);
nor U3593 (N_3593,N_3216,N_3287);
or U3594 (N_3594,N_3322,N_3356);
or U3595 (N_3595,N_3201,N_3383);
or U3596 (N_3596,N_3217,N_3339);
xnor U3597 (N_3597,N_3365,N_3330);
xor U3598 (N_3598,N_3368,N_3257);
nor U3599 (N_3599,N_3353,N_3285);
or U3600 (N_3600,N_3448,N_3460);
or U3601 (N_3601,N_3569,N_3582);
and U3602 (N_3602,N_3566,N_3400);
xor U3603 (N_3603,N_3482,N_3465);
and U3604 (N_3604,N_3459,N_3499);
nor U3605 (N_3605,N_3521,N_3562);
or U3606 (N_3606,N_3526,N_3542);
nand U3607 (N_3607,N_3440,N_3513);
nor U3608 (N_3608,N_3584,N_3596);
and U3609 (N_3609,N_3401,N_3473);
xnor U3610 (N_3610,N_3544,N_3451);
nor U3611 (N_3611,N_3445,N_3579);
and U3612 (N_3612,N_3510,N_3593);
nand U3613 (N_3613,N_3549,N_3547);
nand U3614 (N_3614,N_3444,N_3421);
nor U3615 (N_3615,N_3537,N_3560);
and U3616 (N_3616,N_3597,N_3552);
or U3617 (N_3617,N_3412,N_3518);
or U3618 (N_3618,N_3423,N_3551);
or U3619 (N_3619,N_3527,N_3458);
xor U3620 (N_3620,N_3590,N_3457);
nand U3621 (N_3621,N_3468,N_3425);
nand U3622 (N_3622,N_3419,N_3557);
and U3623 (N_3623,N_3453,N_3567);
nand U3624 (N_3624,N_3464,N_3452);
nand U3625 (N_3625,N_3483,N_3558);
or U3626 (N_3626,N_3503,N_3563);
nand U3627 (N_3627,N_3591,N_3575);
nand U3628 (N_3628,N_3406,N_3493);
and U3629 (N_3629,N_3443,N_3507);
nor U3630 (N_3630,N_3446,N_3508);
xnor U3631 (N_3631,N_3422,N_3413);
nor U3632 (N_3632,N_3427,N_3494);
nor U3633 (N_3633,N_3462,N_3441);
xnor U3634 (N_3634,N_3496,N_3501);
nor U3635 (N_3635,N_3592,N_3583);
nand U3636 (N_3636,N_3486,N_3478);
nor U3637 (N_3637,N_3484,N_3403);
xor U3638 (N_3638,N_3594,N_3571);
nand U3639 (N_3639,N_3565,N_3580);
or U3640 (N_3640,N_3587,N_3532);
nor U3641 (N_3641,N_3574,N_3429);
nor U3642 (N_3642,N_3442,N_3463);
nor U3643 (N_3643,N_3439,N_3469);
or U3644 (N_3644,N_3489,N_3530);
nor U3645 (N_3645,N_3511,N_3472);
xnor U3646 (N_3646,N_3498,N_3519);
nor U3647 (N_3647,N_3430,N_3540);
nand U3648 (N_3648,N_3553,N_3481);
nor U3649 (N_3649,N_3598,N_3417);
or U3650 (N_3650,N_3432,N_3546);
and U3651 (N_3651,N_3585,N_3586);
nand U3652 (N_3652,N_3520,N_3477);
and U3653 (N_3653,N_3467,N_3536);
or U3654 (N_3654,N_3599,N_3595);
nor U3655 (N_3655,N_3435,N_3576);
nand U3656 (N_3656,N_3466,N_3506);
xnor U3657 (N_3657,N_3411,N_3538);
and U3658 (N_3658,N_3455,N_3415);
nand U3659 (N_3659,N_3500,N_3561);
or U3660 (N_3660,N_3479,N_3447);
nor U3661 (N_3661,N_3414,N_3438);
nor U3662 (N_3662,N_3539,N_3535);
xnor U3663 (N_3663,N_3424,N_3504);
xnor U3664 (N_3664,N_3426,N_3497);
xnor U3665 (N_3665,N_3517,N_3556);
xor U3666 (N_3666,N_3408,N_3509);
or U3667 (N_3667,N_3487,N_3528);
or U3668 (N_3668,N_3515,N_3437);
xnor U3669 (N_3669,N_3525,N_3434);
nor U3670 (N_3670,N_3485,N_3454);
nor U3671 (N_3671,N_3531,N_3545);
xnor U3672 (N_3672,N_3490,N_3431);
xor U3673 (N_3673,N_3554,N_3502);
or U3674 (N_3674,N_3450,N_3541);
nor U3675 (N_3675,N_3409,N_3449);
and U3676 (N_3676,N_3550,N_3461);
or U3677 (N_3677,N_3588,N_3420);
and U3678 (N_3678,N_3410,N_3578);
and U3679 (N_3679,N_3470,N_3512);
xor U3680 (N_3680,N_3529,N_3488);
nor U3681 (N_3681,N_3573,N_3524);
and U3682 (N_3682,N_3402,N_3492);
xor U3683 (N_3683,N_3416,N_3505);
and U3684 (N_3684,N_3568,N_3533);
nor U3685 (N_3685,N_3559,N_3581);
nor U3686 (N_3686,N_3534,N_3564);
nor U3687 (N_3687,N_3548,N_3572);
nor U3688 (N_3688,N_3570,N_3522);
or U3689 (N_3689,N_3474,N_3471);
xnor U3690 (N_3690,N_3418,N_3555);
nand U3691 (N_3691,N_3577,N_3407);
xnor U3692 (N_3692,N_3405,N_3589);
or U3693 (N_3693,N_3543,N_3475);
nand U3694 (N_3694,N_3516,N_3491);
xor U3695 (N_3695,N_3433,N_3456);
or U3696 (N_3696,N_3480,N_3428);
and U3697 (N_3697,N_3436,N_3514);
and U3698 (N_3698,N_3495,N_3476);
nand U3699 (N_3699,N_3523,N_3404);
and U3700 (N_3700,N_3436,N_3402);
or U3701 (N_3701,N_3558,N_3407);
nor U3702 (N_3702,N_3454,N_3594);
xnor U3703 (N_3703,N_3422,N_3562);
xnor U3704 (N_3704,N_3533,N_3549);
and U3705 (N_3705,N_3511,N_3486);
nor U3706 (N_3706,N_3425,N_3540);
and U3707 (N_3707,N_3557,N_3482);
and U3708 (N_3708,N_3586,N_3448);
xnor U3709 (N_3709,N_3490,N_3442);
and U3710 (N_3710,N_3440,N_3410);
nor U3711 (N_3711,N_3416,N_3572);
xnor U3712 (N_3712,N_3596,N_3500);
and U3713 (N_3713,N_3423,N_3471);
xor U3714 (N_3714,N_3555,N_3459);
and U3715 (N_3715,N_3551,N_3532);
nor U3716 (N_3716,N_3524,N_3514);
xor U3717 (N_3717,N_3404,N_3498);
nand U3718 (N_3718,N_3496,N_3408);
xnor U3719 (N_3719,N_3549,N_3417);
and U3720 (N_3720,N_3489,N_3585);
or U3721 (N_3721,N_3417,N_3573);
or U3722 (N_3722,N_3429,N_3533);
xor U3723 (N_3723,N_3508,N_3553);
xor U3724 (N_3724,N_3595,N_3562);
nor U3725 (N_3725,N_3473,N_3469);
and U3726 (N_3726,N_3419,N_3484);
and U3727 (N_3727,N_3420,N_3522);
or U3728 (N_3728,N_3565,N_3416);
nor U3729 (N_3729,N_3458,N_3488);
or U3730 (N_3730,N_3533,N_3405);
nor U3731 (N_3731,N_3472,N_3572);
nand U3732 (N_3732,N_3563,N_3552);
or U3733 (N_3733,N_3531,N_3534);
nor U3734 (N_3734,N_3488,N_3546);
or U3735 (N_3735,N_3567,N_3435);
or U3736 (N_3736,N_3516,N_3584);
or U3737 (N_3737,N_3495,N_3493);
xor U3738 (N_3738,N_3580,N_3412);
or U3739 (N_3739,N_3426,N_3452);
nand U3740 (N_3740,N_3597,N_3509);
nor U3741 (N_3741,N_3554,N_3490);
xor U3742 (N_3742,N_3481,N_3502);
and U3743 (N_3743,N_3503,N_3529);
nor U3744 (N_3744,N_3594,N_3524);
xnor U3745 (N_3745,N_3587,N_3475);
and U3746 (N_3746,N_3401,N_3419);
nor U3747 (N_3747,N_3595,N_3429);
or U3748 (N_3748,N_3587,N_3489);
xnor U3749 (N_3749,N_3472,N_3598);
xnor U3750 (N_3750,N_3441,N_3487);
nor U3751 (N_3751,N_3566,N_3573);
nand U3752 (N_3752,N_3442,N_3521);
and U3753 (N_3753,N_3461,N_3495);
nand U3754 (N_3754,N_3402,N_3545);
and U3755 (N_3755,N_3479,N_3451);
nor U3756 (N_3756,N_3498,N_3495);
or U3757 (N_3757,N_3417,N_3447);
or U3758 (N_3758,N_3436,N_3580);
nand U3759 (N_3759,N_3568,N_3546);
or U3760 (N_3760,N_3599,N_3478);
and U3761 (N_3761,N_3522,N_3406);
xor U3762 (N_3762,N_3402,N_3507);
nand U3763 (N_3763,N_3416,N_3519);
nand U3764 (N_3764,N_3458,N_3502);
xnor U3765 (N_3765,N_3472,N_3469);
or U3766 (N_3766,N_3542,N_3583);
or U3767 (N_3767,N_3517,N_3515);
and U3768 (N_3768,N_3410,N_3468);
or U3769 (N_3769,N_3574,N_3586);
xor U3770 (N_3770,N_3403,N_3429);
nor U3771 (N_3771,N_3509,N_3582);
xor U3772 (N_3772,N_3508,N_3484);
nand U3773 (N_3773,N_3567,N_3470);
nand U3774 (N_3774,N_3460,N_3586);
or U3775 (N_3775,N_3448,N_3481);
or U3776 (N_3776,N_3513,N_3421);
or U3777 (N_3777,N_3437,N_3401);
and U3778 (N_3778,N_3405,N_3571);
nor U3779 (N_3779,N_3450,N_3537);
nand U3780 (N_3780,N_3546,N_3541);
and U3781 (N_3781,N_3546,N_3565);
or U3782 (N_3782,N_3408,N_3527);
xor U3783 (N_3783,N_3486,N_3438);
xnor U3784 (N_3784,N_3429,N_3576);
nor U3785 (N_3785,N_3503,N_3516);
nand U3786 (N_3786,N_3531,N_3413);
nor U3787 (N_3787,N_3471,N_3547);
xnor U3788 (N_3788,N_3591,N_3574);
and U3789 (N_3789,N_3587,N_3406);
or U3790 (N_3790,N_3531,N_3580);
and U3791 (N_3791,N_3577,N_3566);
nand U3792 (N_3792,N_3468,N_3583);
and U3793 (N_3793,N_3555,N_3596);
nor U3794 (N_3794,N_3489,N_3425);
or U3795 (N_3795,N_3444,N_3585);
nand U3796 (N_3796,N_3415,N_3523);
nand U3797 (N_3797,N_3545,N_3587);
and U3798 (N_3798,N_3459,N_3441);
and U3799 (N_3799,N_3560,N_3435);
nor U3800 (N_3800,N_3621,N_3661);
and U3801 (N_3801,N_3749,N_3697);
and U3802 (N_3802,N_3716,N_3788);
or U3803 (N_3803,N_3771,N_3724);
and U3804 (N_3804,N_3732,N_3746);
or U3805 (N_3805,N_3617,N_3758);
nand U3806 (N_3806,N_3734,N_3708);
xor U3807 (N_3807,N_3774,N_3640);
or U3808 (N_3808,N_3632,N_3789);
xnor U3809 (N_3809,N_3768,N_3750);
nand U3810 (N_3810,N_3764,N_3616);
and U3811 (N_3811,N_3726,N_3613);
xnor U3812 (N_3812,N_3757,N_3761);
nand U3813 (N_3813,N_3718,N_3719);
or U3814 (N_3814,N_3703,N_3662);
nand U3815 (N_3815,N_3698,N_3780);
and U3816 (N_3816,N_3664,N_3603);
nor U3817 (N_3817,N_3794,N_3673);
nor U3818 (N_3818,N_3723,N_3634);
nor U3819 (N_3819,N_3769,N_3665);
xor U3820 (N_3820,N_3623,N_3767);
xnor U3821 (N_3821,N_3609,N_3785);
nor U3822 (N_3822,N_3735,N_3733);
xnor U3823 (N_3823,N_3690,N_3675);
xnor U3824 (N_3824,N_3770,N_3689);
or U3825 (N_3825,N_3705,N_3630);
and U3826 (N_3826,N_3727,N_3776);
nor U3827 (N_3827,N_3646,N_3712);
xor U3828 (N_3828,N_3787,N_3699);
and U3829 (N_3829,N_3755,N_3729);
and U3830 (N_3830,N_3671,N_3696);
or U3831 (N_3831,N_3752,N_3622);
and U3832 (N_3832,N_3686,N_3643);
and U3833 (N_3833,N_3728,N_3620);
and U3834 (N_3834,N_3722,N_3791);
and U3835 (N_3835,N_3762,N_3679);
and U3836 (N_3836,N_3692,N_3745);
nand U3837 (N_3837,N_3706,N_3754);
or U3838 (N_3838,N_3777,N_3683);
nor U3839 (N_3839,N_3638,N_3693);
nor U3840 (N_3840,N_3753,N_3624);
or U3841 (N_3841,N_3700,N_3647);
nand U3842 (N_3842,N_3797,N_3608);
nand U3843 (N_3843,N_3654,N_3709);
nand U3844 (N_3844,N_3688,N_3682);
nand U3845 (N_3845,N_3775,N_3740);
or U3846 (N_3846,N_3795,N_3666);
xor U3847 (N_3847,N_3655,N_3669);
or U3848 (N_3848,N_3793,N_3681);
and U3849 (N_3849,N_3645,N_3685);
nand U3850 (N_3850,N_3618,N_3650);
or U3851 (N_3851,N_3672,N_3737);
or U3852 (N_3852,N_3644,N_3612);
nor U3853 (N_3853,N_3702,N_3713);
and U3854 (N_3854,N_3657,N_3784);
and U3855 (N_3855,N_3772,N_3635);
or U3856 (N_3856,N_3680,N_3678);
nor U3857 (N_3857,N_3783,N_3602);
nand U3858 (N_3858,N_3736,N_3610);
nor U3859 (N_3859,N_3615,N_3633);
and U3860 (N_3860,N_3748,N_3607);
and U3861 (N_3861,N_3695,N_3668);
or U3862 (N_3862,N_3714,N_3756);
xor U3863 (N_3863,N_3730,N_3773);
xor U3864 (N_3864,N_3798,N_3742);
and U3865 (N_3865,N_3676,N_3614);
or U3866 (N_3866,N_3641,N_3605);
or U3867 (N_3867,N_3631,N_3759);
nand U3868 (N_3868,N_3606,N_3781);
and U3869 (N_3869,N_3619,N_3738);
xnor U3870 (N_3870,N_3704,N_3691);
or U3871 (N_3871,N_3684,N_3660);
xnor U3872 (N_3872,N_3663,N_3782);
xor U3873 (N_3873,N_3653,N_3739);
and U3874 (N_3874,N_3721,N_3639);
or U3875 (N_3875,N_3743,N_3701);
and U3876 (N_3876,N_3648,N_3779);
or U3877 (N_3877,N_3637,N_3658);
nand U3878 (N_3878,N_3731,N_3760);
or U3879 (N_3879,N_3765,N_3627);
xnor U3880 (N_3880,N_3652,N_3659);
and U3881 (N_3881,N_3711,N_3649);
and U3882 (N_3882,N_3778,N_3720);
nand U3883 (N_3883,N_3670,N_3628);
xor U3884 (N_3884,N_3799,N_3629);
and U3885 (N_3885,N_3710,N_3687);
or U3886 (N_3886,N_3786,N_3741);
xor U3887 (N_3887,N_3766,N_3717);
nand U3888 (N_3888,N_3796,N_3677);
or U3889 (N_3889,N_3667,N_3625);
nand U3890 (N_3890,N_3656,N_3600);
xor U3891 (N_3891,N_3707,N_3715);
nor U3892 (N_3892,N_3611,N_3636);
nor U3893 (N_3893,N_3601,N_3642);
xor U3894 (N_3894,N_3744,N_3694);
nor U3895 (N_3895,N_3790,N_3651);
nand U3896 (N_3896,N_3763,N_3725);
nand U3897 (N_3897,N_3751,N_3604);
nand U3898 (N_3898,N_3792,N_3747);
nor U3899 (N_3899,N_3626,N_3674);
or U3900 (N_3900,N_3778,N_3647);
nand U3901 (N_3901,N_3703,N_3701);
nand U3902 (N_3902,N_3754,N_3732);
xor U3903 (N_3903,N_3777,N_3722);
nand U3904 (N_3904,N_3638,N_3760);
xor U3905 (N_3905,N_3683,N_3756);
and U3906 (N_3906,N_3671,N_3629);
nand U3907 (N_3907,N_3771,N_3777);
nor U3908 (N_3908,N_3659,N_3798);
nand U3909 (N_3909,N_3682,N_3711);
and U3910 (N_3910,N_3756,N_3766);
nand U3911 (N_3911,N_3774,N_3629);
and U3912 (N_3912,N_3646,N_3625);
and U3913 (N_3913,N_3752,N_3739);
nor U3914 (N_3914,N_3729,N_3706);
nor U3915 (N_3915,N_3749,N_3628);
and U3916 (N_3916,N_3747,N_3640);
and U3917 (N_3917,N_3607,N_3725);
nand U3918 (N_3918,N_3717,N_3727);
xor U3919 (N_3919,N_3638,N_3609);
and U3920 (N_3920,N_3608,N_3740);
nand U3921 (N_3921,N_3675,N_3770);
and U3922 (N_3922,N_3761,N_3759);
nor U3923 (N_3923,N_3689,N_3680);
or U3924 (N_3924,N_3684,N_3606);
or U3925 (N_3925,N_3689,N_3643);
nand U3926 (N_3926,N_3751,N_3731);
or U3927 (N_3927,N_3781,N_3635);
or U3928 (N_3928,N_3764,N_3689);
and U3929 (N_3929,N_3659,N_3630);
and U3930 (N_3930,N_3782,N_3744);
nand U3931 (N_3931,N_3668,N_3611);
nand U3932 (N_3932,N_3779,N_3701);
nand U3933 (N_3933,N_3632,N_3772);
or U3934 (N_3934,N_3685,N_3668);
xor U3935 (N_3935,N_3751,N_3788);
nand U3936 (N_3936,N_3733,N_3685);
xor U3937 (N_3937,N_3698,N_3647);
xnor U3938 (N_3938,N_3745,N_3762);
and U3939 (N_3939,N_3690,N_3652);
or U3940 (N_3940,N_3767,N_3723);
nand U3941 (N_3941,N_3769,N_3777);
and U3942 (N_3942,N_3743,N_3694);
and U3943 (N_3943,N_3649,N_3639);
nand U3944 (N_3944,N_3726,N_3784);
or U3945 (N_3945,N_3798,N_3605);
and U3946 (N_3946,N_3718,N_3696);
or U3947 (N_3947,N_3733,N_3714);
or U3948 (N_3948,N_3637,N_3701);
nor U3949 (N_3949,N_3791,N_3761);
and U3950 (N_3950,N_3626,N_3730);
and U3951 (N_3951,N_3627,N_3718);
xor U3952 (N_3952,N_3679,N_3790);
xor U3953 (N_3953,N_3673,N_3737);
nand U3954 (N_3954,N_3713,N_3663);
and U3955 (N_3955,N_3796,N_3799);
nand U3956 (N_3956,N_3612,N_3726);
and U3957 (N_3957,N_3740,N_3741);
nor U3958 (N_3958,N_3762,N_3644);
nor U3959 (N_3959,N_3690,N_3707);
or U3960 (N_3960,N_3623,N_3705);
nor U3961 (N_3961,N_3774,N_3624);
xor U3962 (N_3962,N_3639,N_3643);
and U3963 (N_3963,N_3662,N_3686);
nand U3964 (N_3964,N_3653,N_3664);
nand U3965 (N_3965,N_3702,N_3619);
and U3966 (N_3966,N_3681,N_3702);
nand U3967 (N_3967,N_3606,N_3722);
and U3968 (N_3968,N_3773,N_3731);
and U3969 (N_3969,N_3641,N_3615);
or U3970 (N_3970,N_3610,N_3723);
and U3971 (N_3971,N_3727,N_3739);
nor U3972 (N_3972,N_3712,N_3769);
or U3973 (N_3973,N_3658,N_3687);
nand U3974 (N_3974,N_3611,N_3752);
nor U3975 (N_3975,N_3661,N_3762);
or U3976 (N_3976,N_3642,N_3672);
xnor U3977 (N_3977,N_3702,N_3648);
xor U3978 (N_3978,N_3704,N_3786);
nand U3979 (N_3979,N_3709,N_3663);
xnor U3980 (N_3980,N_3694,N_3681);
and U3981 (N_3981,N_3689,N_3776);
or U3982 (N_3982,N_3630,N_3627);
nor U3983 (N_3983,N_3707,N_3621);
nor U3984 (N_3984,N_3627,N_3679);
nand U3985 (N_3985,N_3744,N_3633);
xor U3986 (N_3986,N_3725,N_3632);
nor U3987 (N_3987,N_3791,N_3721);
nor U3988 (N_3988,N_3734,N_3713);
or U3989 (N_3989,N_3685,N_3697);
and U3990 (N_3990,N_3745,N_3666);
xnor U3991 (N_3991,N_3630,N_3767);
or U3992 (N_3992,N_3686,N_3761);
or U3993 (N_3993,N_3658,N_3602);
xnor U3994 (N_3994,N_3749,N_3728);
nor U3995 (N_3995,N_3715,N_3761);
and U3996 (N_3996,N_3647,N_3645);
and U3997 (N_3997,N_3783,N_3741);
xnor U3998 (N_3998,N_3782,N_3625);
nor U3999 (N_3999,N_3664,N_3646);
and U4000 (N_4000,N_3835,N_3989);
or U4001 (N_4001,N_3990,N_3886);
nor U4002 (N_4002,N_3946,N_3913);
nor U4003 (N_4003,N_3822,N_3965);
or U4004 (N_4004,N_3819,N_3849);
nor U4005 (N_4005,N_3867,N_3961);
or U4006 (N_4006,N_3982,N_3958);
and U4007 (N_4007,N_3941,N_3917);
xnor U4008 (N_4008,N_3978,N_3914);
and U4009 (N_4009,N_3829,N_3907);
or U4010 (N_4010,N_3898,N_3859);
and U4011 (N_4011,N_3836,N_3980);
xnor U4012 (N_4012,N_3940,N_3997);
nor U4013 (N_4013,N_3880,N_3972);
xor U4014 (N_4014,N_3984,N_3820);
and U4015 (N_4015,N_3916,N_3888);
xor U4016 (N_4016,N_3962,N_3887);
or U4017 (N_4017,N_3831,N_3930);
and U4018 (N_4018,N_3973,N_3828);
and U4019 (N_4019,N_3954,N_3900);
nor U4020 (N_4020,N_3994,N_3818);
nand U4021 (N_4021,N_3803,N_3811);
xor U4022 (N_4022,N_3904,N_3842);
xor U4023 (N_4023,N_3933,N_3881);
and U4024 (N_4024,N_3923,N_3868);
or U4025 (N_4025,N_3877,N_3826);
or U4026 (N_4026,N_3834,N_3844);
or U4027 (N_4027,N_3922,N_3896);
xnor U4028 (N_4028,N_3847,N_3816);
and U4029 (N_4029,N_3810,N_3901);
nor U4030 (N_4030,N_3969,N_3956);
or U4031 (N_4031,N_3899,N_3850);
xor U4032 (N_4032,N_3999,N_3976);
or U4033 (N_4033,N_3837,N_3808);
and U4034 (N_4034,N_3921,N_3876);
and U4035 (N_4035,N_3996,N_3906);
nor U4036 (N_4036,N_3945,N_3942);
or U4037 (N_4037,N_3971,N_3944);
xnor U4038 (N_4038,N_3823,N_3866);
and U4039 (N_4039,N_3912,N_3928);
xor U4040 (N_4040,N_3910,N_3932);
or U4041 (N_4041,N_3857,N_3918);
nor U4042 (N_4042,N_3987,N_3915);
or U4043 (N_4043,N_3854,N_3891);
and U4044 (N_4044,N_3953,N_3902);
nor U4045 (N_4045,N_3874,N_3963);
or U4046 (N_4046,N_3919,N_3934);
xnor U4047 (N_4047,N_3838,N_3802);
and U4048 (N_4048,N_3861,N_3840);
nor U4049 (N_4049,N_3884,N_3882);
nor U4050 (N_4050,N_3805,N_3925);
nor U4051 (N_4051,N_3949,N_3960);
nand U4052 (N_4052,N_3903,N_3814);
and U4053 (N_4053,N_3872,N_3991);
and U4054 (N_4054,N_3927,N_3948);
xnor U4055 (N_4055,N_3858,N_3892);
nand U4056 (N_4056,N_3873,N_3852);
nor U4057 (N_4057,N_3890,N_3817);
or U4058 (N_4058,N_3863,N_3998);
or U4059 (N_4059,N_3975,N_3968);
or U4060 (N_4060,N_3855,N_3832);
nor U4061 (N_4061,N_3983,N_3885);
nor U4062 (N_4062,N_3813,N_3889);
or U4063 (N_4063,N_3897,N_3804);
nand U4064 (N_4064,N_3937,N_3950);
xor U4065 (N_4065,N_3806,N_3926);
nand U4066 (N_4066,N_3988,N_3830);
or U4067 (N_4067,N_3827,N_3981);
xnor U4068 (N_4068,N_3812,N_3875);
nand U4069 (N_4069,N_3853,N_3894);
xor U4070 (N_4070,N_3839,N_3977);
nor U4071 (N_4071,N_3909,N_3870);
or U4072 (N_4072,N_3986,N_3871);
xor U4073 (N_4073,N_3865,N_3895);
and U4074 (N_4074,N_3851,N_3964);
and U4075 (N_4075,N_3869,N_3959);
nor U4076 (N_4076,N_3905,N_3943);
nor U4077 (N_4077,N_3936,N_3985);
or U4078 (N_4078,N_3979,N_3995);
nand U4079 (N_4079,N_3807,N_3846);
nand U4080 (N_4080,N_3931,N_3966);
or U4081 (N_4081,N_3929,N_3935);
nand U4082 (N_4082,N_3992,N_3800);
xor U4083 (N_4083,N_3821,N_3952);
nand U4084 (N_4084,N_3825,N_3845);
nand U4085 (N_4085,N_3841,N_3967);
xor U4086 (N_4086,N_3974,N_3862);
nand U4087 (N_4087,N_3893,N_3856);
or U4088 (N_4088,N_3833,N_3864);
xnor U4089 (N_4089,N_3951,N_3957);
nand U4090 (N_4090,N_3955,N_3924);
nor U4091 (N_4091,N_3947,N_3920);
xnor U4092 (N_4092,N_3879,N_3809);
or U4093 (N_4093,N_3824,N_3993);
and U4094 (N_4094,N_3860,N_3878);
xor U4095 (N_4095,N_3938,N_3815);
nor U4096 (N_4096,N_3908,N_3848);
nand U4097 (N_4097,N_3911,N_3883);
nor U4098 (N_4098,N_3843,N_3939);
nand U4099 (N_4099,N_3970,N_3801);
or U4100 (N_4100,N_3858,N_3919);
xnor U4101 (N_4101,N_3988,N_3861);
and U4102 (N_4102,N_3908,N_3904);
nor U4103 (N_4103,N_3823,N_3873);
nor U4104 (N_4104,N_3826,N_3839);
and U4105 (N_4105,N_3865,N_3937);
nand U4106 (N_4106,N_3819,N_3920);
xor U4107 (N_4107,N_3840,N_3815);
nor U4108 (N_4108,N_3942,N_3822);
xor U4109 (N_4109,N_3886,N_3938);
or U4110 (N_4110,N_3843,N_3954);
xnor U4111 (N_4111,N_3893,N_3873);
nand U4112 (N_4112,N_3954,N_3923);
nor U4113 (N_4113,N_3922,N_3866);
nor U4114 (N_4114,N_3947,N_3861);
nor U4115 (N_4115,N_3819,N_3860);
nand U4116 (N_4116,N_3884,N_3869);
or U4117 (N_4117,N_3928,N_3873);
and U4118 (N_4118,N_3920,N_3851);
nand U4119 (N_4119,N_3911,N_3820);
nor U4120 (N_4120,N_3887,N_3896);
nor U4121 (N_4121,N_3928,N_3989);
xnor U4122 (N_4122,N_3947,N_3898);
and U4123 (N_4123,N_3988,N_3957);
xnor U4124 (N_4124,N_3959,N_3963);
xor U4125 (N_4125,N_3919,N_3921);
and U4126 (N_4126,N_3818,N_3891);
or U4127 (N_4127,N_3913,N_3921);
xnor U4128 (N_4128,N_3956,N_3921);
and U4129 (N_4129,N_3829,N_3995);
nor U4130 (N_4130,N_3827,N_3851);
or U4131 (N_4131,N_3835,N_3954);
xnor U4132 (N_4132,N_3991,N_3964);
and U4133 (N_4133,N_3875,N_3940);
or U4134 (N_4134,N_3972,N_3887);
nand U4135 (N_4135,N_3957,N_3899);
xnor U4136 (N_4136,N_3961,N_3868);
and U4137 (N_4137,N_3942,N_3991);
or U4138 (N_4138,N_3890,N_3982);
xnor U4139 (N_4139,N_3854,N_3958);
xnor U4140 (N_4140,N_3919,N_3886);
or U4141 (N_4141,N_3981,N_3834);
xor U4142 (N_4142,N_3951,N_3835);
nand U4143 (N_4143,N_3928,N_3927);
and U4144 (N_4144,N_3825,N_3867);
xnor U4145 (N_4145,N_3860,N_3871);
nand U4146 (N_4146,N_3879,N_3986);
or U4147 (N_4147,N_3892,N_3864);
nand U4148 (N_4148,N_3952,N_3938);
xnor U4149 (N_4149,N_3945,N_3892);
and U4150 (N_4150,N_3927,N_3808);
xnor U4151 (N_4151,N_3863,N_3920);
nand U4152 (N_4152,N_3955,N_3929);
nand U4153 (N_4153,N_3853,N_3877);
and U4154 (N_4154,N_3908,N_3879);
nand U4155 (N_4155,N_3973,N_3980);
or U4156 (N_4156,N_3984,N_3890);
nor U4157 (N_4157,N_3992,N_3940);
and U4158 (N_4158,N_3934,N_3986);
xor U4159 (N_4159,N_3807,N_3999);
nor U4160 (N_4160,N_3821,N_3966);
nor U4161 (N_4161,N_3883,N_3884);
nand U4162 (N_4162,N_3960,N_3843);
or U4163 (N_4163,N_3939,N_3869);
and U4164 (N_4164,N_3921,N_3916);
nand U4165 (N_4165,N_3916,N_3907);
nand U4166 (N_4166,N_3935,N_3904);
nor U4167 (N_4167,N_3894,N_3847);
xnor U4168 (N_4168,N_3827,N_3855);
nand U4169 (N_4169,N_3811,N_3879);
xnor U4170 (N_4170,N_3940,N_3835);
nand U4171 (N_4171,N_3980,N_3823);
nand U4172 (N_4172,N_3830,N_3833);
nand U4173 (N_4173,N_3890,N_3886);
xor U4174 (N_4174,N_3867,N_3997);
nor U4175 (N_4175,N_3838,N_3959);
xor U4176 (N_4176,N_3912,N_3976);
and U4177 (N_4177,N_3876,N_3869);
and U4178 (N_4178,N_3947,N_3839);
nand U4179 (N_4179,N_3865,N_3906);
and U4180 (N_4180,N_3960,N_3802);
nand U4181 (N_4181,N_3990,N_3843);
and U4182 (N_4182,N_3995,N_3873);
nand U4183 (N_4183,N_3924,N_3805);
nand U4184 (N_4184,N_3961,N_3848);
and U4185 (N_4185,N_3934,N_3837);
and U4186 (N_4186,N_3850,N_3990);
nor U4187 (N_4187,N_3919,N_3815);
and U4188 (N_4188,N_3929,N_3855);
and U4189 (N_4189,N_3889,N_3837);
or U4190 (N_4190,N_3950,N_3919);
or U4191 (N_4191,N_3916,N_3923);
nor U4192 (N_4192,N_3964,N_3808);
or U4193 (N_4193,N_3988,N_3851);
xor U4194 (N_4194,N_3818,N_3803);
xnor U4195 (N_4195,N_3999,N_3944);
and U4196 (N_4196,N_3820,N_3930);
nand U4197 (N_4197,N_3928,N_3992);
nand U4198 (N_4198,N_3865,N_3806);
nor U4199 (N_4199,N_3820,N_3955);
xor U4200 (N_4200,N_4075,N_4044);
nor U4201 (N_4201,N_4087,N_4155);
xor U4202 (N_4202,N_4016,N_4037);
and U4203 (N_4203,N_4195,N_4191);
nor U4204 (N_4204,N_4109,N_4170);
xnor U4205 (N_4205,N_4073,N_4043);
xor U4206 (N_4206,N_4083,N_4139);
nand U4207 (N_4207,N_4142,N_4179);
nor U4208 (N_4208,N_4159,N_4185);
and U4209 (N_4209,N_4050,N_4114);
and U4210 (N_4210,N_4197,N_4018);
nand U4211 (N_4211,N_4181,N_4060);
nand U4212 (N_4212,N_4117,N_4111);
nor U4213 (N_4213,N_4124,N_4081);
xor U4214 (N_4214,N_4172,N_4144);
or U4215 (N_4215,N_4134,N_4086);
xnor U4216 (N_4216,N_4166,N_4002);
nor U4217 (N_4217,N_4019,N_4072);
xor U4218 (N_4218,N_4032,N_4057);
or U4219 (N_4219,N_4056,N_4175);
nor U4220 (N_4220,N_4198,N_4131);
and U4221 (N_4221,N_4127,N_4165);
xnor U4222 (N_4222,N_4190,N_4076);
or U4223 (N_4223,N_4115,N_4025);
or U4224 (N_4224,N_4151,N_4045);
xnor U4225 (N_4225,N_4186,N_4023);
nand U4226 (N_4226,N_4031,N_4042);
nand U4227 (N_4227,N_4153,N_4145);
or U4228 (N_4228,N_4180,N_4040);
xnor U4229 (N_4229,N_4059,N_4066);
nand U4230 (N_4230,N_4012,N_4123);
xnor U4231 (N_4231,N_4183,N_4022);
and U4232 (N_4232,N_4193,N_4070);
nand U4233 (N_4233,N_4149,N_4026);
and U4234 (N_4234,N_4178,N_4129);
nand U4235 (N_4235,N_4199,N_4116);
xor U4236 (N_4236,N_4108,N_4102);
xnor U4237 (N_4237,N_4015,N_4080);
nor U4238 (N_4238,N_4160,N_4071);
xnor U4239 (N_4239,N_4150,N_4034);
or U4240 (N_4240,N_4000,N_4177);
or U4241 (N_4241,N_4168,N_4138);
and U4242 (N_4242,N_4046,N_4007);
and U4243 (N_4243,N_4152,N_4078);
xnor U4244 (N_4244,N_4122,N_4062);
nor U4245 (N_4245,N_4049,N_4038);
xnor U4246 (N_4246,N_4140,N_4069);
and U4247 (N_4247,N_4157,N_4035);
nor U4248 (N_4248,N_4061,N_4047);
nor U4249 (N_4249,N_4014,N_4005);
nand U4250 (N_4250,N_4112,N_4063);
xnor U4251 (N_4251,N_4068,N_4188);
xnor U4252 (N_4252,N_4029,N_4093);
nor U4253 (N_4253,N_4088,N_4121);
nand U4254 (N_4254,N_4048,N_4132);
or U4255 (N_4255,N_4092,N_4001);
nor U4256 (N_4256,N_4110,N_4135);
xor U4257 (N_4257,N_4085,N_4187);
and U4258 (N_4258,N_4104,N_4182);
and U4259 (N_4259,N_4192,N_4097);
nor U4260 (N_4260,N_4021,N_4171);
nand U4261 (N_4261,N_4008,N_4176);
nor U4262 (N_4262,N_4143,N_4090);
nor U4263 (N_4263,N_4099,N_4010);
xor U4264 (N_4264,N_4125,N_4017);
and U4265 (N_4265,N_4126,N_4128);
or U4266 (N_4266,N_4039,N_4095);
and U4267 (N_4267,N_4130,N_4074);
or U4268 (N_4268,N_4174,N_4079);
nor U4269 (N_4269,N_4058,N_4098);
nor U4270 (N_4270,N_4006,N_4053);
and U4271 (N_4271,N_4133,N_4027);
and U4272 (N_4272,N_4148,N_4082);
nand U4273 (N_4273,N_4094,N_4120);
or U4274 (N_4274,N_4162,N_4100);
and U4275 (N_4275,N_4065,N_4024);
nand U4276 (N_4276,N_4101,N_4137);
nand U4277 (N_4277,N_4004,N_4119);
or U4278 (N_4278,N_4051,N_4009);
and U4279 (N_4279,N_4141,N_4055);
or U4280 (N_4280,N_4028,N_4105);
xnor U4281 (N_4281,N_4052,N_4011);
or U4282 (N_4282,N_4067,N_4030);
nand U4283 (N_4283,N_4020,N_4084);
and U4284 (N_4284,N_4103,N_4096);
or U4285 (N_4285,N_4163,N_4013);
nor U4286 (N_4286,N_4113,N_4003);
or U4287 (N_4287,N_4136,N_4169);
nand U4288 (N_4288,N_4173,N_4033);
nand U4289 (N_4289,N_4091,N_4118);
nor U4290 (N_4290,N_4154,N_4107);
xor U4291 (N_4291,N_4189,N_4106);
nand U4292 (N_4292,N_4196,N_4036);
xnor U4293 (N_4293,N_4184,N_4089);
and U4294 (N_4294,N_4064,N_4077);
or U4295 (N_4295,N_4146,N_4161);
or U4296 (N_4296,N_4164,N_4041);
nand U4297 (N_4297,N_4054,N_4194);
nand U4298 (N_4298,N_4156,N_4167);
nand U4299 (N_4299,N_4158,N_4147);
xor U4300 (N_4300,N_4019,N_4016);
nand U4301 (N_4301,N_4078,N_4107);
nand U4302 (N_4302,N_4006,N_4192);
nand U4303 (N_4303,N_4124,N_4125);
or U4304 (N_4304,N_4110,N_4023);
or U4305 (N_4305,N_4035,N_4117);
nor U4306 (N_4306,N_4081,N_4134);
and U4307 (N_4307,N_4108,N_4157);
or U4308 (N_4308,N_4057,N_4005);
nor U4309 (N_4309,N_4132,N_4126);
and U4310 (N_4310,N_4129,N_4047);
xnor U4311 (N_4311,N_4075,N_4153);
xnor U4312 (N_4312,N_4135,N_4029);
nor U4313 (N_4313,N_4163,N_4130);
xor U4314 (N_4314,N_4154,N_4059);
nand U4315 (N_4315,N_4051,N_4160);
nor U4316 (N_4316,N_4133,N_4197);
nor U4317 (N_4317,N_4132,N_4028);
or U4318 (N_4318,N_4026,N_4151);
nand U4319 (N_4319,N_4126,N_4175);
xnor U4320 (N_4320,N_4125,N_4105);
nor U4321 (N_4321,N_4125,N_4044);
and U4322 (N_4322,N_4122,N_4035);
nand U4323 (N_4323,N_4127,N_4074);
nand U4324 (N_4324,N_4145,N_4121);
nor U4325 (N_4325,N_4095,N_4180);
and U4326 (N_4326,N_4198,N_4173);
and U4327 (N_4327,N_4166,N_4070);
and U4328 (N_4328,N_4118,N_4041);
nand U4329 (N_4329,N_4182,N_4012);
nand U4330 (N_4330,N_4148,N_4059);
xnor U4331 (N_4331,N_4127,N_4068);
nand U4332 (N_4332,N_4134,N_4050);
xor U4333 (N_4333,N_4197,N_4107);
nor U4334 (N_4334,N_4002,N_4188);
or U4335 (N_4335,N_4033,N_4082);
xor U4336 (N_4336,N_4029,N_4138);
xnor U4337 (N_4337,N_4052,N_4091);
nand U4338 (N_4338,N_4144,N_4151);
and U4339 (N_4339,N_4029,N_4126);
or U4340 (N_4340,N_4002,N_4074);
nand U4341 (N_4341,N_4062,N_4144);
and U4342 (N_4342,N_4106,N_4043);
xnor U4343 (N_4343,N_4051,N_4071);
nor U4344 (N_4344,N_4135,N_4069);
or U4345 (N_4345,N_4137,N_4170);
nor U4346 (N_4346,N_4130,N_4063);
nor U4347 (N_4347,N_4081,N_4055);
and U4348 (N_4348,N_4052,N_4078);
xor U4349 (N_4349,N_4044,N_4149);
and U4350 (N_4350,N_4147,N_4003);
xor U4351 (N_4351,N_4011,N_4170);
nand U4352 (N_4352,N_4156,N_4155);
or U4353 (N_4353,N_4145,N_4025);
nor U4354 (N_4354,N_4012,N_4075);
and U4355 (N_4355,N_4075,N_4118);
xnor U4356 (N_4356,N_4043,N_4085);
nand U4357 (N_4357,N_4051,N_4123);
xnor U4358 (N_4358,N_4037,N_4045);
or U4359 (N_4359,N_4046,N_4174);
xor U4360 (N_4360,N_4112,N_4024);
nand U4361 (N_4361,N_4046,N_4011);
nand U4362 (N_4362,N_4097,N_4143);
xor U4363 (N_4363,N_4169,N_4095);
xor U4364 (N_4364,N_4188,N_4100);
xnor U4365 (N_4365,N_4035,N_4118);
or U4366 (N_4366,N_4016,N_4187);
xnor U4367 (N_4367,N_4060,N_4125);
nor U4368 (N_4368,N_4028,N_4169);
and U4369 (N_4369,N_4171,N_4107);
xnor U4370 (N_4370,N_4141,N_4028);
xor U4371 (N_4371,N_4047,N_4163);
nor U4372 (N_4372,N_4107,N_4083);
nand U4373 (N_4373,N_4106,N_4168);
and U4374 (N_4374,N_4009,N_4134);
and U4375 (N_4375,N_4120,N_4118);
nor U4376 (N_4376,N_4075,N_4082);
nand U4377 (N_4377,N_4116,N_4013);
nand U4378 (N_4378,N_4083,N_4079);
nand U4379 (N_4379,N_4060,N_4135);
nor U4380 (N_4380,N_4085,N_4107);
xor U4381 (N_4381,N_4025,N_4071);
or U4382 (N_4382,N_4148,N_4071);
xnor U4383 (N_4383,N_4087,N_4015);
or U4384 (N_4384,N_4062,N_4094);
or U4385 (N_4385,N_4078,N_4117);
nor U4386 (N_4386,N_4132,N_4068);
xor U4387 (N_4387,N_4011,N_4047);
nand U4388 (N_4388,N_4101,N_4163);
and U4389 (N_4389,N_4008,N_4019);
nand U4390 (N_4390,N_4020,N_4045);
and U4391 (N_4391,N_4072,N_4092);
nand U4392 (N_4392,N_4014,N_4140);
nand U4393 (N_4393,N_4057,N_4011);
and U4394 (N_4394,N_4041,N_4183);
and U4395 (N_4395,N_4070,N_4072);
nand U4396 (N_4396,N_4108,N_4059);
xnor U4397 (N_4397,N_4004,N_4110);
nand U4398 (N_4398,N_4072,N_4042);
nand U4399 (N_4399,N_4009,N_4043);
nand U4400 (N_4400,N_4321,N_4350);
xor U4401 (N_4401,N_4353,N_4296);
and U4402 (N_4402,N_4309,N_4303);
nor U4403 (N_4403,N_4203,N_4364);
and U4404 (N_4404,N_4396,N_4289);
nand U4405 (N_4405,N_4392,N_4273);
nor U4406 (N_4406,N_4233,N_4231);
nand U4407 (N_4407,N_4311,N_4307);
nor U4408 (N_4408,N_4376,N_4358);
xnor U4409 (N_4409,N_4221,N_4257);
xnor U4410 (N_4410,N_4371,N_4272);
nor U4411 (N_4411,N_4329,N_4246);
nor U4412 (N_4412,N_4280,N_4290);
xor U4413 (N_4413,N_4327,N_4385);
xnor U4414 (N_4414,N_4305,N_4342);
nand U4415 (N_4415,N_4254,N_4295);
and U4416 (N_4416,N_4359,N_4202);
nand U4417 (N_4417,N_4344,N_4224);
nand U4418 (N_4418,N_4384,N_4217);
xnor U4419 (N_4419,N_4399,N_4235);
and U4420 (N_4420,N_4227,N_4252);
or U4421 (N_4421,N_4300,N_4247);
nor U4422 (N_4422,N_4282,N_4284);
nor U4423 (N_4423,N_4304,N_4220);
xor U4424 (N_4424,N_4346,N_4351);
nand U4425 (N_4425,N_4230,N_4225);
xnor U4426 (N_4426,N_4381,N_4285);
nor U4427 (N_4427,N_4345,N_4356);
and U4428 (N_4428,N_4269,N_4340);
nand U4429 (N_4429,N_4354,N_4395);
xor U4430 (N_4430,N_4315,N_4258);
nor U4431 (N_4431,N_4226,N_4318);
nand U4432 (N_4432,N_4219,N_4347);
or U4433 (N_4433,N_4245,N_4264);
xnor U4434 (N_4434,N_4209,N_4204);
nor U4435 (N_4435,N_4279,N_4301);
xor U4436 (N_4436,N_4242,N_4362);
or U4437 (N_4437,N_4374,N_4387);
xor U4438 (N_4438,N_4383,N_4308);
xor U4439 (N_4439,N_4349,N_4332);
xnor U4440 (N_4440,N_4283,N_4223);
or U4441 (N_4441,N_4368,N_4323);
and U4442 (N_4442,N_4277,N_4286);
xnor U4443 (N_4443,N_4278,N_4299);
nand U4444 (N_4444,N_4302,N_4293);
and U4445 (N_4445,N_4366,N_4357);
and U4446 (N_4446,N_4297,N_4271);
and U4447 (N_4447,N_4201,N_4306);
nand U4448 (N_4448,N_4274,N_4330);
and U4449 (N_4449,N_4207,N_4337);
xnor U4450 (N_4450,N_4328,N_4294);
xor U4451 (N_4451,N_4218,N_4312);
nor U4452 (N_4452,N_4210,N_4326);
or U4453 (N_4453,N_4251,N_4324);
nand U4454 (N_4454,N_4343,N_4390);
nor U4455 (N_4455,N_4243,N_4270);
and U4456 (N_4456,N_4336,N_4338);
xnor U4457 (N_4457,N_4208,N_4240);
nand U4458 (N_4458,N_4335,N_4363);
or U4459 (N_4459,N_4391,N_4263);
and U4460 (N_4460,N_4352,N_4244);
and U4461 (N_4461,N_4222,N_4228);
nand U4462 (N_4462,N_4331,N_4365);
and U4463 (N_4463,N_4388,N_4232);
nor U4464 (N_4464,N_4367,N_4287);
nor U4465 (N_4465,N_4214,N_4375);
or U4466 (N_4466,N_4341,N_4325);
nor U4467 (N_4467,N_4256,N_4268);
or U4468 (N_4468,N_4322,N_4212);
nand U4469 (N_4469,N_4216,N_4259);
xor U4470 (N_4470,N_4265,N_4238);
and U4471 (N_4471,N_4393,N_4253);
nor U4472 (N_4472,N_4211,N_4348);
nand U4473 (N_4473,N_4241,N_4319);
nand U4474 (N_4474,N_4215,N_4267);
xor U4475 (N_4475,N_4260,N_4370);
xnor U4476 (N_4476,N_4361,N_4373);
nor U4477 (N_4477,N_4386,N_4234);
nor U4478 (N_4478,N_4239,N_4229);
or U4479 (N_4479,N_4261,N_4291);
nand U4480 (N_4480,N_4333,N_4248);
xor U4481 (N_4481,N_4334,N_4380);
xor U4482 (N_4482,N_4298,N_4379);
and U4483 (N_4483,N_4317,N_4255);
or U4484 (N_4484,N_4200,N_4310);
xor U4485 (N_4485,N_4313,N_4213);
xnor U4486 (N_4486,N_4394,N_4355);
nor U4487 (N_4487,N_4275,N_4314);
nor U4488 (N_4488,N_4288,N_4369);
and U4489 (N_4489,N_4236,N_4360);
nand U4490 (N_4490,N_4205,N_4398);
and U4491 (N_4491,N_4276,N_4389);
or U4492 (N_4492,N_4372,N_4250);
xnor U4493 (N_4493,N_4377,N_4397);
nand U4494 (N_4494,N_4249,N_4292);
and U4495 (N_4495,N_4262,N_4382);
nand U4496 (N_4496,N_4237,N_4266);
and U4497 (N_4497,N_4281,N_4339);
nand U4498 (N_4498,N_4320,N_4378);
xnor U4499 (N_4499,N_4316,N_4206);
and U4500 (N_4500,N_4270,N_4279);
and U4501 (N_4501,N_4224,N_4204);
nand U4502 (N_4502,N_4372,N_4200);
or U4503 (N_4503,N_4229,N_4281);
nand U4504 (N_4504,N_4278,N_4374);
or U4505 (N_4505,N_4300,N_4318);
nand U4506 (N_4506,N_4333,N_4312);
nor U4507 (N_4507,N_4361,N_4228);
or U4508 (N_4508,N_4281,N_4302);
xnor U4509 (N_4509,N_4208,N_4360);
nor U4510 (N_4510,N_4389,N_4221);
or U4511 (N_4511,N_4374,N_4255);
xor U4512 (N_4512,N_4336,N_4289);
or U4513 (N_4513,N_4228,N_4205);
nand U4514 (N_4514,N_4394,N_4349);
xor U4515 (N_4515,N_4247,N_4349);
xor U4516 (N_4516,N_4223,N_4305);
xor U4517 (N_4517,N_4276,N_4201);
or U4518 (N_4518,N_4298,N_4231);
or U4519 (N_4519,N_4228,N_4285);
nand U4520 (N_4520,N_4218,N_4303);
xnor U4521 (N_4521,N_4398,N_4264);
nor U4522 (N_4522,N_4274,N_4359);
and U4523 (N_4523,N_4289,N_4325);
xnor U4524 (N_4524,N_4248,N_4268);
or U4525 (N_4525,N_4356,N_4338);
nand U4526 (N_4526,N_4218,N_4208);
xnor U4527 (N_4527,N_4233,N_4322);
or U4528 (N_4528,N_4381,N_4340);
xor U4529 (N_4529,N_4314,N_4318);
or U4530 (N_4530,N_4352,N_4307);
nand U4531 (N_4531,N_4237,N_4258);
nor U4532 (N_4532,N_4288,N_4213);
nor U4533 (N_4533,N_4219,N_4398);
nor U4534 (N_4534,N_4245,N_4217);
nand U4535 (N_4535,N_4285,N_4226);
xor U4536 (N_4536,N_4382,N_4294);
nor U4537 (N_4537,N_4383,N_4272);
nand U4538 (N_4538,N_4246,N_4379);
xor U4539 (N_4539,N_4330,N_4363);
or U4540 (N_4540,N_4280,N_4348);
nor U4541 (N_4541,N_4389,N_4351);
or U4542 (N_4542,N_4372,N_4208);
xnor U4543 (N_4543,N_4368,N_4212);
xor U4544 (N_4544,N_4266,N_4210);
nand U4545 (N_4545,N_4235,N_4264);
xnor U4546 (N_4546,N_4314,N_4263);
and U4547 (N_4547,N_4212,N_4214);
and U4548 (N_4548,N_4355,N_4207);
xnor U4549 (N_4549,N_4391,N_4207);
or U4550 (N_4550,N_4254,N_4245);
xnor U4551 (N_4551,N_4396,N_4209);
or U4552 (N_4552,N_4383,N_4370);
nor U4553 (N_4553,N_4243,N_4317);
and U4554 (N_4554,N_4301,N_4317);
nand U4555 (N_4555,N_4283,N_4332);
and U4556 (N_4556,N_4264,N_4336);
and U4557 (N_4557,N_4296,N_4360);
xnor U4558 (N_4558,N_4258,N_4360);
xnor U4559 (N_4559,N_4292,N_4350);
nand U4560 (N_4560,N_4342,N_4321);
xnor U4561 (N_4561,N_4211,N_4270);
or U4562 (N_4562,N_4317,N_4346);
nand U4563 (N_4563,N_4370,N_4214);
or U4564 (N_4564,N_4357,N_4273);
or U4565 (N_4565,N_4204,N_4210);
or U4566 (N_4566,N_4311,N_4309);
and U4567 (N_4567,N_4316,N_4228);
and U4568 (N_4568,N_4341,N_4279);
and U4569 (N_4569,N_4305,N_4303);
nor U4570 (N_4570,N_4221,N_4217);
xnor U4571 (N_4571,N_4383,N_4202);
and U4572 (N_4572,N_4271,N_4255);
or U4573 (N_4573,N_4365,N_4337);
nand U4574 (N_4574,N_4391,N_4348);
nand U4575 (N_4575,N_4348,N_4364);
and U4576 (N_4576,N_4390,N_4335);
nand U4577 (N_4577,N_4393,N_4297);
nand U4578 (N_4578,N_4250,N_4214);
nand U4579 (N_4579,N_4345,N_4371);
and U4580 (N_4580,N_4239,N_4335);
xor U4581 (N_4581,N_4285,N_4380);
and U4582 (N_4582,N_4348,N_4205);
and U4583 (N_4583,N_4280,N_4338);
and U4584 (N_4584,N_4204,N_4222);
nor U4585 (N_4585,N_4323,N_4301);
nand U4586 (N_4586,N_4275,N_4232);
or U4587 (N_4587,N_4350,N_4379);
nor U4588 (N_4588,N_4267,N_4254);
or U4589 (N_4589,N_4250,N_4354);
nor U4590 (N_4590,N_4240,N_4264);
nor U4591 (N_4591,N_4202,N_4352);
nand U4592 (N_4592,N_4333,N_4330);
nand U4593 (N_4593,N_4276,N_4260);
nor U4594 (N_4594,N_4204,N_4250);
nand U4595 (N_4595,N_4254,N_4318);
or U4596 (N_4596,N_4271,N_4260);
nand U4597 (N_4597,N_4315,N_4284);
xnor U4598 (N_4598,N_4244,N_4373);
xnor U4599 (N_4599,N_4297,N_4308);
xnor U4600 (N_4600,N_4430,N_4531);
and U4601 (N_4601,N_4532,N_4591);
or U4602 (N_4602,N_4506,N_4490);
and U4603 (N_4603,N_4465,N_4518);
or U4604 (N_4604,N_4538,N_4508);
nor U4605 (N_4605,N_4553,N_4438);
nor U4606 (N_4606,N_4458,N_4590);
nor U4607 (N_4607,N_4534,N_4405);
nand U4608 (N_4608,N_4510,N_4521);
nor U4609 (N_4609,N_4416,N_4455);
nand U4610 (N_4610,N_4482,N_4486);
nor U4611 (N_4611,N_4504,N_4575);
or U4612 (N_4612,N_4581,N_4428);
or U4613 (N_4613,N_4558,N_4579);
xor U4614 (N_4614,N_4468,N_4561);
or U4615 (N_4615,N_4480,N_4498);
xnor U4616 (N_4616,N_4419,N_4530);
and U4617 (N_4617,N_4592,N_4423);
xor U4618 (N_4618,N_4513,N_4417);
xor U4619 (N_4619,N_4491,N_4516);
nor U4620 (N_4620,N_4559,N_4462);
and U4621 (N_4621,N_4440,N_4477);
and U4622 (N_4622,N_4568,N_4582);
or U4623 (N_4623,N_4500,N_4429);
nor U4624 (N_4624,N_4577,N_4589);
xnor U4625 (N_4625,N_4453,N_4566);
and U4626 (N_4626,N_4596,N_4523);
xor U4627 (N_4627,N_4451,N_4409);
nor U4628 (N_4628,N_4410,N_4584);
nor U4629 (N_4629,N_4552,N_4434);
and U4630 (N_4630,N_4436,N_4535);
and U4631 (N_4631,N_4469,N_4495);
and U4632 (N_4632,N_4570,N_4571);
or U4633 (N_4633,N_4587,N_4402);
nand U4634 (N_4634,N_4488,N_4420);
and U4635 (N_4635,N_4565,N_4404);
xor U4636 (N_4636,N_4586,N_4431);
nand U4637 (N_4637,N_4400,N_4470);
and U4638 (N_4638,N_4569,N_4418);
and U4639 (N_4639,N_4464,N_4427);
and U4640 (N_4640,N_4526,N_4503);
or U4641 (N_4641,N_4524,N_4493);
nand U4642 (N_4642,N_4445,N_4557);
and U4643 (N_4643,N_4460,N_4555);
and U4644 (N_4644,N_4599,N_4414);
nor U4645 (N_4645,N_4507,N_4563);
nor U4646 (N_4646,N_4511,N_4546);
nand U4647 (N_4647,N_4580,N_4594);
and U4648 (N_4648,N_4547,N_4437);
xor U4649 (N_4649,N_4598,N_4496);
nor U4650 (N_4650,N_4467,N_4406);
or U4651 (N_4651,N_4497,N_4567);
nand U4652 (N_4652,N_4595,N_4540);
nor U4653 (N_4653,N_4564,N_4411);
xor U4654 (N_4654,N_4578,N_4501);
nand U4655 (N_4655,N_4583,N_4461);
nor U4656 (N_4656,N_4515,N_4544);
xor U4657 (N_4657,N_4439,N_4441);
nor U4658 (N_4658,N_4519,N_4509);
xnor U4659 (N_4659,N_4444,N_4576);
nand U4660 (N_4660,N_4473,N_4512);
xnor U4661 (N_4661,N_4457,N_4421);
nand U4662 (N_4662,N_4459,N_4499);
or U4663 (N_4663,N_4537,N_4542);
and U4664 (N_4664,N_4505,N_4422);
nor U4665 (N_4665,N_4471,N_4528);
and U4666 (N_4666,N_4489,N_4562);
or U4667 (N_4667,N_4525,N_4549);
xnor U4668 (N_4668,N_4502,N_4425);
or U4669 (N_4669,N_4485,N_4448);
xor U4670 (N_4670,N_4446,N_4415);
nor U4671 (N_4671,N_4533,N_4478);
xnor U4672 (N_4672,N_4452,N_4574);
or U4673 (N_4673,N_4539,N_4442);
and U4674 (N_4674,N_4449,N_4517);
xor U4675 (N_4675,N_4408,N_4551);
nor U4676 (N_4676,N_4407,N_4494);
and U4677 (N_4677,N_4585,N_4597);
nor U4678 (N_4678,N_4433,N_4527);
or U4679 (N_4679,N_4573,N_4548);
nor U4680 (N_4680,N_4483,N_4424);
and U4681 (N_4681,N_4484,N_4536);
nor U4682 (N_4682,N_4514,N_4572);
xnor U4683 (N_4683,N_4426,N_4541);
nand U4684 (N_4684,N_4403,N_4481);
nor U4685 (N_4685,N_4560,N_4435);
or U4686 (N_4686,N_4401,N_4554);
nand U4687 (N_4687,N_4520,N_4556);
xnor U4688 (N_4688,N_4529,N_4413);
nand U4689 (N_4689,N_4450,N_4479);
and U4690 (N_4690,N_4466,N_4593);
xnor U4691 (N_4691,N_4456,N_4487);
or U4692 (N_4692,N_4463,N_4550);
xor U4693 (N_4693,N_4492,N_4588);
nor U4694 (N_4694,N_4472,N_4454);
and U4695 (N_4695,N_4432,N_4476);
and U4696 (N_4696,N_4522,N_4412);
nor U4697 (N_4697,N_4475,N_4474);
or U4698 (N_4698,N_4545,N_4543);
nand U4699 (N_4699,N_4443,N_4447);
nor U4700 (N_4700,N_4526,N_4415);
or U4701 (N_4701,N_4473,N_4466);
xnor U4702 (N_4702,N_4481,N_4429);
nor U4703 (N_4703,N_4469,N_4465);
xnor U4704 (N_4704,N_4543,N_4591);
nor U4705 (N_4705,N_4546,N_4535);
nand U4706 (N_4706,N_4414,N_4550);
and U4707 (N_4707,N_4465,N_4510);
or U4708 (N_4708,N_4523,N_4597);
and U4709 (N_4709,N_4469,N_4402);
nor U4710 (N_4710,N_4538,N_4430);
and U4711 (N_4711,N_4472,N_4432);
or U4712 (N_4712,N_4591,N_4593);
nor U4713 (N_4713,N_4514,N_4483);
and U4714 (N_4714,N_4521,N_4524);
xnor U4715 (N_4715,N_4508,N_4460);
xnor U4716 (N_4716,N_4592,N_4572);
nor U4717 (N_4717,N_4417,N_4589);
and U4718 (N_4718,N_4574,N_4503);
nand U4719 (N_4719,N_4590,N_4475);
nor U4720 (N_4720,N_4428,N_4434);
nand U4721 (N_4721,N_4427,N_4515);
xnor U4722 (N_4722,N_4417,N_4495);
nor U4723 (N_4723,N_4415,N_4485);
or U4724 (N_4724,N_4422,N_4414);
and U4725 (N_4725,N_4445,N_4591);
xor U4726 (N_4726,N_4509,N_4466);
nor U4727 (N_4727,N_4494,N_4401);
nor U4728 (N_4728,N_4537,N_4460);
and U4729 (N_4729,N_4508,N_4487);
nand U4730 (N_4730,N_4551,N_4506);
nand U4731 (N_4731,N_4568,N_4442);
xnor U4732 (N_4732,N_4501,N_4590);
xor U4733 (N_4733,N_4488,N_4527);
xor U4734 (N_4734,N_4487,N_4470);
nand U4735 (N_4735,N_4573,N_4422);
or U4736 (N_4736,N_4508,N_4498);
nor U4737 (N_4737,N_4523,N_4564);
and U4738 (N_4738,N_4514,N_4439);
and U4739 (N_4739,N_4474,N_4409);
nor U4740 (N_4740,N_4496,N_4471);
nor U4741 (N_4741,N_4442,N_4428);
xor U4742 (N_4742,N_4414,N_4551);
nor U4743 (N_4743,N_4594,N_4488);
xor U4744 (N_4744,N_4587,N_4492);
xor U4745 (N_4745,N_4464,N_4588);
xnor U4746 (N_4746,N_4516,N_4573);
xor U4747 (N_4747,N_4475,N_4503);
or U4748 (N_4748,N_4436,N_4498);
nor U4749 (N_4749,N_4442,N_4530);
nor U4750 (N_4750,N_4503,N_4463);
nand U4751 (N_4751,N_4461,N_4513);
nor U4752 (N_4752,N_4436,N_4525);
xnor U4753 (N_4753,N_4457,N_4458);
nor U4754 (N_4754,N_4453,N_4495);
xnor U4755 (N_4755,N_4495,N_4557);
or U4756 (N_4756,N_4554,N_4470);
and U4757 (N_4757,N_4501,N_4427);
xor U4758 (N_4758,N_4598,N_4426);
nor U4759 (N_4759,N_4487,N_4452);
and U4760 (N_4760,N_4524,N_4459);
xnor U4761 (N_4761,N_4583,N_4481);
or U4762 (N_4762,N_4469,N_4443);
xnor U4763 (N_4763,N_4533,N_4497);
or U4764 (N_4764,N_4481,N_4422);
nand U4765 (N_4765,N_4572,N_4460);
nor U4766 (N_4766,N_4513,N_4548);
and U4767 (N_4767,N_4559,N_4522);
or U4768 (N_4768,N_4506,N_4486);
and U4769 (N_4769,N_4410,N_4488);
xor U4770 (N_4770,N_4430,N_4583);
nand U4771 (N_4771,N_4505,N_4496);
nand U4772 (N_4772,N_4520,N_4418);
and U4773 (N_4773,N_4506,N_4453);
nand U4774 (N_4774,N_4526,N_4491);
or U4775 (N_4775,N_4406,N_4489);
xor U4776 (N_4776,N_4554,N_4537);
or U4777 (N_4777,N_4499,N_4445);
nor U4778 (N_4778,N_4542,N_4504);
nand U4779 (N_4779,N_4588,N_4565);
or U4780 (N_4780,N_4424,N_4466);
and U4781 (N_4781,N_4514,N_4524);
nand U4782 (N_4782,N_4560,N_4567);
nor U4783 (N_4783,N_4550,N_4426);
or U4784 (N_4784,N_4527,N_4508);
xor U4785 (N_4785,N_4500,N_4545);
and U4786 (N_4786,N_4401,N_4455);
xor U4787 (N_4787,N_4403,N_4454);
xor U4788 (N_4788,N_4501,N_4597);
xor U4789 (N_4789,N_4493,N_4587);
xnor U4790 (N_4790,N_4472,N_4401);
or U4791 (N_4791,N_4588,N_4490);
nor U4792 (N_4792,N_4575,N_4559);
nor U4793 (N_4793,N_4494,N_4481);
nand U4794 (N_4794,N_4590,N_4563);
nand U4795 (N_4795,N_4570,N_4469);
xor U4796 (N_4796,N_4402,N_4457);
nor U4797 (N_4797,N_4527,N_4571);
xor U4798 (N_4798,N_4441,N_4463);
xnor U4799 (N_4799,N_4494,N_4496);
or U4800 (N_4800,N_4624,N_4687);
xor U4801 (N_4801,N_4762,N_4710);
xor U4802 (N_4802,N_4705,N_4632);
nor U4803 (N_4803,N_4652,N_4623);
and U4804 (N_4804,N_4664,N_4747);
nand U4805 (N_4805,N_4775,N_4699);
xnor U4806 (N_4806,N_4650,N_4691);
or U4807 (N_4807,N_4731,N_4689);
or U4808 (N_4808,N_4784,N_4753);
and U4809 (N_4809,N_4630,N_4782);
nand U4810 (N_4810,N_4777,N_4785);
xnor U4811 (N_4811,N_4609,N_4732);
nor U4812 (N_4812,N_4667,N_4702);
nand U4813 (N_4813,N_4757,N_4636);
nand U4814 (N_4814,N_4659,N_4799);
nand U4815 (N_4815,N_4749,N_4616);
nor U4816 (N_4816,N_4717,N_4612);
nand U4817 (N_4817,N_4605,N_4673);
nand U4818 (N_4818,N_4764,N_4637);
or U4819 (N_4819,N_4703,N_4669);
and U4820 (N_4820,N_4648,N_4627);
nand U4821 (N_4821,N_4773,N_4788);
nor U4822 (N_4822,N_4769,N_4614);
nand U4823 (N_4823,N_4653,N_4608);
and U4824 (N_4824,N_4647,N_4640);
xor U4825 (N_4825,N_4727,N_4660);
or U4826 (N_4826,N_4682,N_4685);
or U4827 (N_4827,N_4744,N_4633);
nand U4828 (N_4828,N_4792,N_4666);
nor U4829 (N_4829,N_4663,N_4750);
or U4830 (N_4830,N_4745,N_4670);
nor U4831 (N_4831,N_4754,N_4665);
xor U4832 (N_4832,N_4628,N_4629);
nand U4833 (N_4833,N_4790,N_4722);
nand U4834 (N_4834,N_4655,N_4704);
xor U4835 (N_4835,N_4671,N_4766);
and U4836 (N_4836,N_4761,N_4774);
nor U4837 (N_4837,N_4720,N_4626);
and U4838 (N_4838,N_4668,N_4778);
nor U4839 (N_4839,N_4672,N_4613);
and U4840 (N_4840,N_4716,N_4742);
xnor U4841 (N_4841,N_4729,N_4676);
or U4842 (N_4842,N_4641,N_4780);
and U4843 (N_4843,N_4617,N_4625);
xnor U4844 (N_4844,N_4736,N_4798);
or U4845 (N_4845,N_4601,N_4765);
xnor U4846 (N_4846,N_4606,N_4679);
and U4847 (N_4847,N_4635,N_4796);
or U4848 (N_4848,N_4724,N_4719);
or U4849 (N_4849,N_4781,N_4795);
or U4850 (N_4850,N_4657,N_4739);
nor U4851 (N_4851,N_4768,N_4758);
xor U4852 (N_4852,N_4674,N_4645);
or U4853 (N_4853,N_4728,N_4725);
xor U4854 (N_4854,N_4708,N_4791);
or U4855 (N_4855,N_4639,N_4734);
nor U4856 (N_4856,N_4735,N_4707);
nand U4857 (N_4857,N_4783,N_4662);
xor U4858 (N_4858,N_4686,N_4638);
xor U4859 (N_4859,N_4693,N_4772);
or U4860 (N_4860,N_4748,N_4763);
or U4861 (N_4861,N_4610,N_4711);
and U4862 (N_4862,N_4654,N_4713);
or U4863 (N_4863,N_4684,N_4730);
and U4864 (N_4864,N_4631,N_4793);
nor U4865 (N_4865,N_4771,N_4794);
and U4866 (N_4866,N_4618,N_4770);
or U4867 (N_4867,N_4603,N_4726);
nand U4868 (N_4868,N_4714,N_4619);
nand U4869 (N_4869,N_4602,N_4642);
xnor U4870 (N_4870,N_4706,N_4677);
xnor U4871 (N_4871,N_4738,N_4643);
or U4872 (N_4872,N_4701,N_4733);
nand U4873 (N_4873,N_4767,N_4737);
xor U4874 (N_4874,N_4644,N_4789);
and U4875 (N_4875,N_4658,N_4651);
and U4876 (N_4876,N_4759,N_4611);
nor U4877 (N_4877,N_4680,N_4600);
and U4878 (N_4878,N_4786,N_4746);
and U4879 (N_4879,N_4697,N_4751);
and U4880 (N_4880,N_4760,N_4607);
or U4881 (N_4881,N_4787,N_4776);
nor U4882 (N_4882,N_4696,N_4698);
nor U4883 (N_4883,N_4752,N_4661);
and U4884 (N_4884,N_4646,N_4743);
xnor U4885 (N_4885,N_4712,N_4718);
and U4886 (N_4886,N_4656,N_4622);
nor U4887 (N_4887,N_4615,N_4675);
and U4888 (N_4888,N_4700,N_4755);
or U4889 (N_4889,N_4649,N_4692);
nor U4890 (N_4890,N_4695,N_4740);
xor U4891 (N_4891,N_4715,N_4723);
or U4892 (N_4892,N_4634,N_4621);
and U4893 (N_4893,N_4620,N_4721);
xor U4894 (N_4894,N_4779,N_4756);
or U4895 (N_4895,N_4681,N_4709);
or U4896 (N_4896,N_4688,N_4741);
xnor U4897 (N_4897,N_4678,N_4694);
and U4898 (N_4898,N_4604,N_4690);
or U4899 (N_4899,N_4797,N_4683);
nor U4900 (N_4900,N_4738,N_4655);
xor U4901 (N_4901,N_4738,N_4795);
and U4902 (N_4902,N_4651,N_4724);
nand U4903 (N_4903,N_4755,N_4612);
xnor U4904 (N_4904,N_4644,N_4641);
and U4905 (N_4905,N_4761,N_4616);
and U4906 (N_4906,N_4771,N_4605);
xor U4907 (N_4907,N_4645,N_4762);
and U4908 (N_4908,N_4671,N_4705);
and U4909 (N_4909,N_4776,N_4732);
or U4910 (N_4910,N_4619,N_4604);
or U4911 (N_4911,N_4606,N_4751);
or U4912 (N_4912,N_4679,N_4783);
and U4913 (N_4913,N_4710,N_4652);
or U4914 (N_4914,N_4774,N_4606);
and U4915 (N_4915,N_4603,N_4725);
and U4916 (N_4916,N_4674,N_4738);
nand U4917 (N_4917,N_4657,N_4794);
nor U4918 (N_4918,N_4684,N_4677);
or U4919 (N_4919,N_4680,N_4746);
nor U4920 (N_4920,N_4602,N_4795);
xor U4921 (N_4921,N_4601,N_4738);
or U4922 (N_4922,N_4777,N_4660);
xnor U4923 (N_4923,N_4798,N_4622);
nor U4924 (N_4924,N_4614,N_4679);
nand U4925 (N_4925,N_4747,N_4786);
xnor U4926 (N_4926,N_4641,N_4666);
nand U4927 (N_4927,N_4636,N_4653);
nand U4928 (N_4928,N_4757,N_4766);
and U4929 (N_4929,N_4732,N_4620);
nand U4930 (N_4930,N_4640,N_4654);
nand U4931 (N_4931,N_4602,N_4722);
or U4932 (N_4932,N_4621,N_4618);
and U4933 (N_4933,N_4642,N_4760);
or U4934 (N_4934,N_4609,N_4793);
and U4935 (N_4935,N_4764,N_4744);
nand U4936 (N_4936,N_4632,N_4788);
xnor U4937 (N_4937,N_4660,N_4618);
xnor U4938 (N_4938,N_4660,N_4737);
nand U4939 (N_4939,N_4772,N_4602);
nor U4940 (N_4940,N_4648,N_4634);
or U4941 (N_4941,N_4788,N_4628);
nor U4942 (N_4942,N_4671,N_4645);
nand U4943 (N_4943,N_4739,N_4748);
nor U4944 (N_4944,N_4760,N_4695);
xnor U4945 (N_4945,N_4692,N_4728);
or U4946 (N_4946,N_4650,N_4731);
and U4947 (N_4947,N_4620,N_4678);
or U4948 (N_4948,N_4762,N_4621);
nand U4949 (N_4949,N_4685,N_4700);
xor U4950 (N_4950,N_4626,N_4605);
nand U4951 (N_4951,N_4693,N_4700);
nand U4952 (N_4952,N_4680,N_4697);
xnor U4953 (N_4953,N_4665,N_4678);
and U4954 (N_4954,N_4797,N_4792);
xnor U4955 (N_4955,N_4755,N_4649);
and U4956 (N_4956,N_4667,N_4781);
or U4957 (N_4957,N_4665,N_4771);
nor U4958 (N_4958,N_4659,N_4605);
or U4959 (N_4959,N_4791,N_4756);
or U4960 (N_4960,N_4680,N_4672);
and U4961 (N_4961,N_4744,N_4703);
nor U4962 (N_4962,N_4605,N_4756);
xor U4963 (N_4963,N_4791,N_4788);
and U4964 (N_4964,N_4700,N_4754);
xor U4965 (N_4965,N_4798,N_4781);
nor U4966 (N_4966,N_4682,N_4667);
nor U4967 (N_4967,N_4685,N_4758);
or U4968 (N_4968,N_4678,N_4780);
nor U4969 (N_4969,N_4688,N_4648);
nand U4970 (N_4970,N_4784,N_4730);
nand U4971 (N_4971,N_4783,N_4664);
nor U4972 (N_4972,N_4767,N_4715);
xnor U4973 (N_4973,N_4758,N_4762);
or U4974 (N_4974,N_4713,N_4724);
or U4975 (N_4975,N_4691,N_4760);
and U4976 (N_4976,N_4691,N_4737);
nand U4977 (N_4977,N_4644,N_4666);
nor U4978 (N_4978,N_4642,N_4603);
or U4979 (N_4979,N_4645,N_4746);
or U4980 (N_4980,N_4631,N_4724);
or U4981 (N_4981,N_4784,N_4645);
and U4982 (N_4982,N_4648,N_4793);
nor U4983 (N_4983,N_4790,N_4601);
nand U4984 (N_4984,N_4707,N_4671);
nand U4985 (N_4985,N_4728,N_4796);
nand U4986 (N_4986,N_4604,N_4727);
nand U4987 (N_4987,N_4699,N_4719);
nand U4988 (N_4988,N_4758,N_4642);
nor U4989 (N_4989,N_4786,N_4718);
or U4990 (N_4990,N_4690,N_4668);
or U4991 (N_4991,N_4731,N_4706);
nor U4992 (N_4992,N_4768,N_4606);
nand U4993 (N_4993,N_4741,N_4718);
and U4994 (N_4994,N_4620,N_4769);
and U4995 (N_4995,N_4749,N_4607);
and U4996 (N_4996,N_4647,N_4657);
nor U4997 (N_4997,N_4616,N_4709);
or U4998 (N_4998,N_4645,N_4747);
xnor U4999 (N_4999,N_4605,N_4672);
xor U5000 (N_5000,N_4874,N_4838);
xnor U5001 (N_5001,N_4972,N_4929);
xor U5002 (N_5002,N_4861,N_4832);
xor U5003 (N_5003,N_4833,N_4999);
or U5004 (N_5004,N_4976,N_4961);
nor U5005 (N_5005,N_4856,N_4969);
nor U5006 (N_5006,N_4947,N_4801);
or U5007 (N_5007,N_4864,N_4964);
and U5008 (N_5008,N_4867,N_4931);
or U5009 (N_5009,N_4873,N_4809);
or U5010 (N_5010,N_4953,N_4994);
nor U5011 (N_5011,N_4876,N_4883);
xor U5012 (N_5012,N_4828,N_4889);
xnor U5013 (N_5013,N_4990,N_4979);
xor U5014 (N_5014,N_4997,N_4862);
or U5015 (N_5015,N_4888,N_4875);
nand U5016 (N_5016,N_4939,N_4967);
or U5017 (N_5017,N_4869,N_4818);
nand U5018 (N_5018,N_4954,N_4943);
or U5019 (N_5019,N_4917,N_4842);
nor U5020 (N_5020,N_4813,N_4891);
or U5021 (N_5021,N_4894,N_4982);
nor U5022 (N_5022,N_4902,N_4918);
and U5023 (N_5023,N_4870,N_4837);
nor U5024 (N_5024,N_4987,N_4877);
nand U5025 (N_5025,N_4806,N_4965);
and U5026 (N_5026,N_4886,N_4957);
and U5027 (N_5027,N_4951,N_4904);
or U5028 (N_5028,N_4985,N_4908);
nand U5029 (N_5029,N_4899,N_4909);
nand U5030 (N_5030,N_4978,N_4826);
xnor U5031 (N_5031,N_4991,N_4932);
xnor U5032 (N_5032,N_4919,N_4924);
nor U5033 (N_5033,N_4984,N_4846);
nand U5034 (N_5034,N_4808,N_4973);
nor U5035 (N_5035,N_4851,N_4863);
xnor U5036 (N_5036,N_4836,N_4956);
and U5037 (N_5037,N_4887,N_4988);
nand U5038 (N_5038,N_4952,N_4921);
nor U5039 (N_5039,N_4983,N_4892);
nand U5040 (N_5040,N_4849,N_4933);
or U5041 (N_5041,N_4900,N_4895);
xnor U5042 (N_5042,N_4854,N_4814);
or U5043 (N_5043,N_4903,N_4940);
and U5044 (N_5044,N_4884,N_4948);
or U5045 (N_5045,N_4996,N_4949);
nor U5046 (N_5046,N_4866,N_4914);
xor U5047 (N_5047,N_4946,N_4871);
xor U5048 (N_5048,N_4859,N_4812);
nor U5049 (N_5049,N_4807,N_4975);
xor U5050 (N_5050,N_4959,N_4845);
xnor U5051 (N_5051,N_4989,N_4811);
nand U5052 (N_5052,N_4936,N_4893);
xnor U5053 (N_5053,N_4852,N_4880);
and U5054 (N_5054,N_4890,N_4906);
or U5055 (N_5055,N_4850,N_4968);
nand U5056 (N_5056,N_4885,N_4821);
and U5057 (N_5057,N_4944,N_4942);
or U5058 (N_5058,N_4920,N_4963);
xor U5059 (N_5059,N_4926,N_4824);
xor U5060 (N_5060,N_4868,N_4977);
nor U5061 (N_5061,N_4927,N_4901);
or U5062 (N_5062,N_4802,N_4839);
nand U5063 (N_5063,N_4841,N_4882);
and U5064 (N_5064,N_4804,N_4855);
nand U5065 (N_5065,N_4911,N_4848);
xnor U5066 (N_5066,N_4815,N_4853);
xor U5067 (N_5067,N_4827,N_4817);
and U5068 (N_5068,N_4981,N_4872);
or U5069 (N_5069,N_4847,N_4881);
nor U5070 (N_5070,N_4960,N_4835);
nand U5071 (N_5071,N_4843,N_4865);
or U5072 (N_5072,N_4974,N_4980);
or U5073 (N_5073,N_4910,N_4857);
or U5074 (N_5074,N_4907,N_4834);
nor U5075 (N_5075,N_4879,N_4831);
xor U5076 (N_5076,N_4878,N_4896);
nor U5077 (N_5077,N_4941,N_4966);
xor U5078 (N_5078,N_4800,N_4822);
nor U5079 (N_5079,N_4816,N_4860);
or U5080 (N_5080,N_4803,N_4934);
xor U5081 (N_5081,N_4819,N_4898);
nand U5082 (N_5082,N_4958,N_4986);
nand U5083 (N_5083,N_4950,N_4962);
or U5084 (N_5084,N_4998,N_4928);
or U5085 (N_5085,N_4971,N_4829);
nor U5086 (N_5086,N_4830,N_4923);
nor U5087 (N_5087,N_4955,N_4992);
nand U5088 (N_5088,N_4905,N_4930);
xor U5089 (N_5089,N_4937,N_4945);
nor U5090 (N_5090,N_4810,N_4916);
nand U5091 (N_5091,N_4844,N_4825);
and U5092 (N_5092,N_4995,N_4840);
or U5093 (N_5093,N_4993,N_4970);
xnor U5094 (N_5094,N_4925,N_4805);
or U5095 (N_5095,N_4858,N_4938);
nand U5096 (N_5096,N_4912,N_4915);
xnor U5097 (N_5097,N_4823,N_4935);
xor U5098 (N_5098,N_4913,N_4922);
or U5099 (N_5099,N_4820,N_4897);
xor U5100 (N_5100,N_4941,N_4885);
xnor U5101 (N_5101,N_4999,N_4837);
and U5102 (N_5102,N_4853,N_4890);
nand U5103 (N_5103,N_4883,N_4857);
or U5104 (N_5104,N_4900,N_4924);
nor U5105 (N_5105,N_4990,N_4883);
nand U5106 (N_5106,N_4840,N_4873);
xor U5107 (N_5107,N_4989,N_4987);
nor U5108 (N_5108,N_4975,N_4880);
or U5109 (N_5109,N_4971,N_4969);
and U5110 (N_5110,N_4831,N_4833);
and U5111 (N_5111,N_4984,N_4998);
xor U5112 (N_5112,N_4956,N_4829);
xnor U5113 (N_5113,N_4824,N_4946);
and U5114 (N_5114,N_4924,N_4813);
or U5115 (N_5115,N_4941,N_4895);
and U5116 (N_5116,N_4826,N_4870);
and U5117 (N_5117,N_4804,N_4833);
or U5118 (N_5118,N_4856,N_4912);
nor U5119 (N_5119,N_4881,N_4886);
xor U5120 (N_5120,N_4861,N_4931);
nor U5121 (N_5121,N_4931,N_4822);
xnor U5122 (N_5122,N_4986,N_4943);
xor U5123 (N_5123,N_4958,N_4835);
nand U5124 (N_5124,N_4982,N_4905);
or U5125 (N_5125,N_4959,N_4806);
nand U5126 (N_5126,N_4893,N_4874);
and U5127 (N_5127,N_4818,N_4832);
or U5128 (N_5128,N_4942,N_4877);
and U5129 (N_5129,N_4931,N_4988);
or U5130 (N_5130,N_4848,N_4818);
xnor U5131 (N_5131,N_4815,N_4894);
nand U5132 (N_5132,N_4834,N_4947);
nor U5133 (N_5133,N_4833,N_4822);
nand U5134 (N_5134,N_4935,N_4808);
and U5135 (N_5135,N_4850,N_4969);
or U5136 (N_5136,N_4902,N_4859);
and U5137 (N_5137,N_4891,N_4898);
nor U5138 (N_5138,N_4883,N_4956);
xor U5139 (N_5139,N_4923,N_4804);
and U5140 (N_5140,N_4820,N_4825);
nand U5141 (N_5141,N_4850,N_4933);
or U5142 (N_5142,N_4813,N_4810);
or U5143 (N_5143,N_4824,N_4808);
xnor U5144 (N_5144,N_4893,N_4869);
nor U5145 (N_5145,N_4899,N_4941);
xor U5146 (N_5146,N_4813,N_4931);
xor U5147 (N_5147,N_4961,N_4831);
nor U5148 (N_5148,N_4936,N_4841);
or U5149 (N_5149,N_4964,N_4934);
or U5150 (N_5150,N_4858,N_4993);
nor U5151 (N_5151,N_4933,N_4895);
nand U5152 (N_5152,N_4931,N_4812);
nor U5153 (N_5153,N_4836,N_4959);
nand U5154 (N_5154,N_4876,N_4837);
nand U5155 (N_5155,N_4905,N_4896);
nor U5156 (N_5156,N_4990,N_4907);
nand U5157 (N_5157,N_4891,N_4841);
nor U5158 (N_5158,N_4905,N_4825);
or U5159 (N_5159,N_4843,N_4879);
xnor U5160 (N_5160,N_4930,N_4848);
or U5161 (N_5161,N_4934,N_4909);
nand U5162 (N_5162,N_4998,N_4983);
and U5163 (N_5163,N_4976,N_4898);
or U5164 (N_5164,N_4957,N_4912);
nor U5165 (N_5165,N_4962,N_4894);
and U5166 (N_5166,N_4987,N_4972);
nand U5167 (N_5167,N_4855,N_4840);
and U5168 (N_5168,N_4888,N_4985);
or U5169 (N_5169,N_4817,N_4897);
nor U5170 (N_5170,N_4979,N_4989);
nand U5171 (N_5171,N_4912,N_4836);
and U5172 (N_5172,N_4951,N_4877);
nor U5173 (N_5173,N_4890,N_4918);
xor U5174 (N_5174,N_4948,N_4834);
xor U5175 (N_5175,N_4962,N_4988);
nor U5176 (N_5176,N_4820,N_4891);
or U5177 (N_5177,N_4846,N_4867);
and U5178 (N_5178,N_4811,N_4919);
nand U5179 (N_5179,N_4914,N_4806);
and U5180 (N_5180,N_4862,N_4920);
or U5181 (N_5181,N_4884,N_4972);
nor U5182 (N_5182,N_4883,N_4870);
nand U5183 (N_5183,N_4909,N_4963);
xor U5184 (N_5184,N_4873,N_4916);
or U5185 (N_5185,N_4852,N_4955);
nand U5186 (N_5186,N_4806,N_4969);
nor U5187 (N_5187,N_4932,N_4938);
and U5188 (N_5188,N_4839,N_4816);
and U5189 (N_5189,N_4954,N_4907);
or U5190 (N_5190,N_4866,N_4956);
nor U5191 (N_5191,N_4906,N_4951);
nor U5192 (N_5192,N_4902,N_4919);
nor U5193 (N_5193,N_4927,N_4911);
and U5194 (N_5194,N_4978,N_4977);
xnor U5195 (N_5195,N_4805,N_4940);
xnor U5196 (N_5196,N_4904,N_4854);
and U5197 (N_5197,N_4804,N_4937);
or U5198 (N_5198,N_4898,N_4956);
xor U5199 (N_5199,N_4903,N_4971);
nand U5200 (N_5200,N_5168,N_5154);
nor U5201 (N_5201,N_5134,N_5025);
and U5202 (N_5202,N_5086,N_5064);
xnor U5203 (N_5203,N_5094,N_5116);
nand U5204 (N_5204,N_5126,N_5118);
nor U5205 (N_5205,N_5138,N_5114);
and U5206 (N_5206,N_5111,N_5136);
or U5207 (N_5207,N_5084,N_5110);
and U5208 (N_5208,N_5083,N_5120);
nor U5209 (N_5209,N_5040,N_5146);
xor U5210 (N_5210,N_5055,N_5190);
xnor U5211 (N_5211,N_5062,N_5013);
nor U5212 (N_5212,N_5035,N_5038);
nand U5213 (N_5213,N_5155,N_5087);
xnor U5214 (N_5214,N_5117,N_5031);
xor U5215 (N_5215,N_5058,N_5182);
xnor U5216 (N_5216,N_5073,N_5039);
xor U5217 (N_5217,N_5063,N_5145);
and U5218 (N_5218,N_5106,N_5172);
nor U5219 (N_5219,N_5027,N_5131);
and U5220 (N_5220,N_5036,N_5034);
nor U5221 (N_5221,N_5121,N_5060);
nor U5222 (N_5222,N_5077,N_5011);
nand U5223 (N_5223,N_5105,N_5159);
or U5224 (N_5224,N_5191,N_5071);
xor U5225 (N_5225,N_5141,N_5122);
xor U5226 (N_5226,N_5001,N_5183);
xor U5227 (N_5227,N_5167,N_5163);
nand U5228 (N_5228,N_5096,N_5028);
nand U5229 (N_5229,N_5198,N_5107);
and U5230 (N_5230,N_5143,N_5133);
nand U5231 (N_5231,N_5142,N_5095);
and U5232 (N_5232,N_5147,N_5012);
nand U5233 (N_5233,N_5165,N_5014);
and U5234 (N_5234,N_5043,N_5150);
xnor U5235 (N_5235,N_5074,N_5021);
or U5236 (N_5236,N_5079,N_5051);
xnor U5237 (N_5237,N_5042,N_5080);
xnor U5238 (N_5238,N_5192,N_5023);
and U5239 (N_5239,N_5137,N_5066);
or U5240 (N_5240,N_5092,N_5196);
nor U5241 (N_5241,N_5022,N_5157);
xor U5242 (N_5242,N_5171,N_5135);
nand U5243 (N_5243,N_5162,N_5024);
nand U5244 (N_5244,N_5148,N_5197);
or U5245 (N_5245,N_5102,N_5056);
and U5246 (N_5246,N_5176,N_5002);
nor U5247 (N_5247,N_5153,N_5139);
nand U5248 (N_5248,N_5166,N_5091);
xnor U5249 (N_5249,N_5177,N_5123);
nor U5250 (N_5250,N_5124,N_5113);
xor U5251 (N_5251,N_5088,N_5008);
xor U5252 (N_5252,N_5119,N_5109);
or U5253 (N_5253,N_5020,N_5044);
nor U5254 (N_5254,N_5175,N_5030);
or U5255 (N_5255,N_5005,N_5188);
nor U5256 (N_5256,N_5103,N_5082);
or U5257 (N_5257,N_5127,N_5161);
xnor U5258 (N_5258,N_5033,N_5004);
xnor U5259 (N_5259,N_5187,N_5151);
nor U5260 (N_5260,N_5076,N_5170);
nor U5261 (N_5261,N_5000,N_5132);
nand U5262 (N_5262,N_5098,N_5019);
nand U5263 (N_5263,N_5037,N_5067);
xor U5264 (N_5264,N_5164,N_5045);
xnor U5265 (N_5265,N_5041,N_5101);
nand U5266 (N_5266,N_5160,N_5029);
or U5267 (N_5267,N_5169,N_5089);
xor U5268 (N_5268,N_5059,N_5069);
or U5269 (N_5269,N_5090,N_5181);
nand U5270 (N_5270,N_5125,N_5174);
nor U5271 (N_5271,N_5003,N_5097);
or U5272 (N_5272,N_5178,N_5015);
nand U5273 (N_5273,N_5068,N_5065);
nor U5274 (N_5274,N_5112,N_5149);
nor U5275 (N_5275,N_5130,N_5057);
and U5276 (N_5276,N_5152,N_5199);
xor U5277 (N_5277,N_5115,N_5017);
and U5278 (N_5278,N_5195,N_5129);
xnor U5279 (N_5279,N_5070,N_5054);
nor U5280 (N_5280,N_5072,N_5052);
nand U5281 (N_5281,N_5047,N_5140);
nand U5282 (N_5282,N_5186,N_5018);
or U5283 (N_5283,N_5093,N_5104);
nor U5284 (N_5284,N_5081,N_5032);
and U5285 (N_5285,N_5050,N_5158);
nand U5286 (N_5286,N_5185,N_5144);
nand U5287 (N_5287,N_5049,N_5108);
and U5288 (N_5288,N_5053,N_5010);
nor U5289 (N_5289,N_5100,N_5128);
nand U5290 (N_5290,N_5179,N_5194);
or U5291 (N_5291,N_5184,N_5046);
nand U5292 (N_5292,N_5156,N_5075);
xor U5293 (N_5293,N_5009,N_5026);
or U5294 (N_5294,N_5180,N_5061);
nand U5295 (N_5295,N_5078,N_5193);
xor U5296 (N_5296,N_5016,N_5048);
and U5297 (N_5297,N_5085,N_5189);
nor U5298 (N_5298,N_5006,N_5007);
and U5299 (N_5299,N_5173,N_5099);
or U5300 (N_5300,N_5064,N_5144);
xor U5301 (N_5301,N_5041,N_5153);
or U5302 (N_5302,N_5164,N_5142);
nor U5303 (N_5303,N_5067,N_5068);
nand U5304 (N_5304,N_5039,N_5194);
xnor U5305 (N_5305,N_5036,N_5153);
xor U5306 (N_5306,N_5095,N_5052);
nor U5307 (N_5307,N_5088,N_5142);
nand U5308 (N_5308,N_5153,N_5144);
nand U5309 (N_5309,N_5120,N_5164);
nor U5310 (N_5310,N_5111,N_5060);
xor U5311 (N_5311,N_5183,N_5037);
nor U5312 (N_5312,N_5129,N_5031);
and U5313 (N_5313,N_5095,N_5008);
or U5314 (N_5314,N_5157,N_5130);
xor U5315 (N_5315,N_5003,N_5028);
xnor U5316 (N_5316,N_5186,N_5148);
or U5317 (N_5317,N_5075,N_5013);
xnor U5318 (N_5318,N_5113,N_5048);
nand U5319 (N_5319,N_5078,N_5068);
xor U5320 (N_5320,N_5058,N_5094);
xnor U5321 (N_5321,N_5083,N_5101);
nand U5322 (N_5322,N_5133,N_5104);
nand U5323 (N_5323,N_5020,N_5074);
nor U5324 (N_5324,N_5063,N_5088);
nand U5325 (N_5325,N_5151,N_5007);
and U5326 (N_5326,N_5182,N_5170);
nor U5327 (N_5327,N_5039,N_5191);
nand U5328 (N_5328,N_5124,N_5042);
nand U5329 (N_5329,N_5164,N_5121);
or U5330 (N_5330,N_5182,N_5142);
and U5331 (N_5331,N_5089,N_5130);
nor U5332 (N_5332,N_5142,N_5075);
or U5333 (N_5333,N_5010,N_5134);
nand U5334 (N_5334,N_5107,N_5138);
nor U5335 (N_5335,N_5167,N_5194);
nor U5336 (N_5336,N_5095,N_5022);
or U5337 (N_5337,N_5061,N_5070);
xnor U5338 (N_5338,N_5160,N_5093);
nor U5339 (N_5339,N_5088,N_5065);
and U5340 (N_5340,N_5108,N_5161);
and U5341 (N_5341,N_5022,N_5050);
nand U5342 (N_5342,N_5122,N_5152);
or U5343 (N_5343,N_5166,N_5036);
or U5344 (N_5344,N_5113,N_5027);
nor U5345 (N_5345,N_5130,N_5073);
nor U5346 (N_5346,N_5013,N_5156);
and U5347 (N_5347,N_5186,N_5146);
and U5348 (N_5348,N_5163,N_5149);
nand U5349 (N_5349,N_5195,N_5198);
and U5350 (N_5350,N_5087,N_5160);
xor U5351 (N_5351,N_5005,N_5061);
xor U5352 (N_5352,N_5032,N_5142);
nand U5353 (N_5353,N_5154,N_5132);
xor U5354 (N_5354,N_5072,N_5159);
and U5355 (N_5355,N_5048,N_5099);
or U5356 (N_5356,N_5016,N_5188);
nand U5357 (N_5357,N_5198,N_5023);
xnor U5358 (N_5358,N_5195,N_5075);
nand U5359 (N_5359,N_5060,N_5157);
xor U5360 (N_5360,N_5032,N_5126);
nand U5361 (N_5361,N_5120,N_5110);
nand U5362 (N_5362,N_5162,N_5090);
and U5363 (N_5363,N_5148,N_5124);
and U5364 (N_5364,N_5145,N_5198);
nor U5365 (N_5365,N_5110,N_5117);
xor U5366 (N_5366,N_5046,N_5174);
and U5367 (N_5367,N_5196,N_5122);
or U5368 (N_5368,N_5148,N_5039);
nand U5369 (N_5369,N_5156,N_5086);
nand U5370 (N_5370,N_5181,N_5178);
or U5371 (N_5371,N_5109,N_5093);
or U5372 (N_5372,N_5179,N_5063);
and U5373 (N_5373,N_5076,N_5032);
nand U5374 (N_5374,N_5149,N_5015);
or U5375 (N_5375,N_5080,N_5151);
or U5376 (N_5376,N_5045,N_5084);
nor U5377 (N_5377,N_5124,N_5051);
and U5378 (N_5378,N_5014,N_5168);
nor U5379 (N_5379,N_5131,N_5133);
or U5380 (N_5380,N_5163,N_5119);
nor U5381 (N_5381,N_5071,N_5087);
nand U5382 (N_5382,N_5091,N_5097);
xor U5383 (N_5383,N_5071,N_5066);
nor U5384 (N_5384,N_5017,N_5145);
or U5385 (N_5385,N_5006,N_5064);
and U5386 (N_5386,N_5086,N_5081);
and U5387 (N_5387,N_5048,N_5093);
xor U5388 (N_5388,N_5110,N_5187);
xor U5389 (N_5389,N_5086,N_5009);
xor U5390 (N_5390,N_5191,N_5077);
nand U5391 (N_5391,N_5145,N_5186);
nand U5392 (N_5392,N_5019,N_5093);
and U5393 (N_5393,N_5096,N_5155);
nand U5394 (N_5394,N_5185,N_5156);
nor U5395 (N_5395,N_5160,N_5076);
nand U5396 (N_5396,N_5086,N_5041);
nand U5397 (N_5397,N_5163,N_5191);
and U5398 (N_5398,N_5087,N_5179);
nand U5399 (N_5399,N_5086,N_5177);
and U5400 (N_5400,N_5355,N_5334);
and U5401 (N_5401,N_5299,N_5211);
nand U5402 (N_5402,N_5223,N_5390);
xnor U5403 (N_5403,N_5388,N_5216);
nand U5404 (N_5404,N_5227,N_5338);
nor U5405 (N_5405,N_5283,N_5336);
and U5406 (N_5406,N_5207,N_5348);
nor U5407 (N_5407,N_5228,N_5221);
xnor U5408 (N_5408,N_5230,N_5340);
and U5409 (N_5409,N_5300,N_5384);
and U5410 (N_5410,N_5289,N_5247);
nand U5411 (N_5411,N_5327,N_5383);
or U5412 (N_5412,N_5273,N_5262);
xor U5413 (N_5413,N_5234,N_5345);
xor U5414 (N_5414,N_5220,N_5368);
or U5415 (N_5415,N_5328,N_5297);
nand U5416 (N_5416,N_5367,N_5218);
and U5417 (N_5417,N_5315,N_5369);
xnor U5418 (N_5418,N_5275,N_5375);
and U5419 (N_5419,N_5378,N_5250);
nand U5420 (N_5420,N_5226,N_5224);
nand U5421 (N_5421,N_5360,N_5358);
or U5422 (N_5422,N_5241,N_5280);
xor U5423 (N_5423,N_5255,N_5361);
xor U5424 (N_5424,N_5201,N_5214);
and U5425 (N_5425,N_5397,N_5265);
xnor U5426 (N_5426,N_5364,N_5212);
or U5427 (N_5427,N_5399,N_5319);
nor U5428 (N_5428,N_5274,N_5222);
and U5429 (N_5429,N_5341,N_5264);
or U5430 (N_5430,N_5237,N_5286);
nand U5431 (N_5431,N_5206,N_5318);
or U5432 (N_5432,N_5308,N_5310);
or U5433 (N_5433,N_5219,N_5233);
or U5434 (N_5434,N_5277,N_5394);
nand U5435 (N_5435,N_5331,N_5245);
or U5436 (N_5436,N_5349,N_5272);
or U5437 (N_5437,N_5393,N_5240);
nor U5438 (N_5438,N_5295,N_5257);
nor U5439 (N_5439,N_5303,N_5267);
or U5440 (N_5440,N_5365,N_5339);
or U5441 (N_5441,N_5266,N_5270);
or U5442 (N_5442,N_5243,N_5296);
or U5443 (N_5443,N_5372,N_5244);
or U5444 (N_5444,N_5380,N_5391);
nand U5445 (N_5445,N_5261,N_5202);
nand U5446 (N_5446,N_5268,N_5343);
nor U5447 (N_5447,N_5386,N_5210);
nor U5448 (N_5448,N_5342,N_5232);
and U5449 (N_5449,N_5322,N_5387);
xnor U5450 (N_5450,N_5304,N_5254);
and U5451 (N_5451,N_5238,N_5205);
xnor U5452 (N_5452,N_5371,N_5284);
or U5453 (N_5453,N_5385,N_5382);
nor U5454 (N_5454,N_5290,N_5288);
nor U5455 (N_5455,N_5305,N_5302);
nor U5456 (N_5456,N_5350,N_5344);
nor U5457 (N_5457,N_5395,N_5398);
or U5458 (N_5458,N_5209,N_5373);
nand U5459 (N_5459,N_5236,N_5271);
xor U5460 (N_5460,N_5251,N_5291);
or U5461 (N_5461,N_5396,N_5329);
and U5462 (N_5462,N_5379,N_5377);
or U5463 (N_5463,N_5313,N_5337);
or U5464 (N_5464,N_5352,N_5311);
and U5465 (N_5465,N_5325,N_5335);
and U5466 (N_5466,N_5203,N_5293);
and U5467 (N_5467,N_5292,N_5256);
nor U5468 (N_5468,N_5242,N_5332);
xnor U5469 (N_5469,N_5259,N_5309);
nand U5470 (N_5470,N_5279,N_5370);
xnor U5471 (N_5471,N_5321,N_5246);
and U5472 (N_5472,N_5363,N_5333);
xnor U5473 (N_5473,N_5351,N_5356);
nor U5474 (N_5474,N_5326,N_5269);
nand U5475 (N_5475,N_5298,N_5294);
nor U5476 (N_5476,N_5376,N_5301);
and U5477 (N_5477,N_5353,N_5225);
nand U5478 (N_5478,N_5231,N_5263);
and U5479 (N_5479,N_5320,N_5215);
xor U5480 (N_5480,N_5204,N_5312);
or U5481 (N_5481,N_5324,N_5278);
nand U5482 (N_5482,N_5374,N_5253);
nand U5483 (N_5483,N_5347,N_5285);
xnor U5484 (N_5484,N_5235,N_5260);
or U5485 (N_5485,N_5249,N_5281);
nand U5486 (N_5486,N_5217,N_5213);
nor U5487 (N_5487,N_5306,N_5323);
xor U5488 (N_5488,N_5307,N_5316);
and U5489 (N_5489,N_5276,N_5252);
or U5490 (N_5490,N_5357,N_5346);
nand U5491 (N_5491,N_5362,N_5200);
xnor U5492 (N_5492,N_5229,N_5330);
xor U5493 (N_5493,N_5317,N_5381);
xnor U5494 (N_5494,N_5359,N_5314);
nand U5495 (N_5495,N_5389,N_5392);
nand U5496 (N_5496,N_5239,N_5208);
nand U5497 (N_5497,N_5282,N_5287);
nand U5498 (N_5498,N_5354,N_5258);
or U5499 (N_5499,N_5366,N_5248);
or U5500 (N_5500,N_5259,N_5314);
xor U5501 (N_5501,N_5220,N_5315);
or U5502 (N_5502,N_5221,N_5274);
or U5503 (N_5503,N_5263,N_5297);
or U5504 (N_5504,N_5274,N_5214);
nor U5505 (N_5505,N_5253,N_5326);
and U5506 (N_5506,N_5397,N_5274);
or U5507 (N_5507,N_5312,N_5339);
nor U5508 (N_5508,N_5346,N_5366);
xor U5509 (N_5509,N_5212,N_5288);
nand U5510 (N_5510,N_5387,N_5397);
xor U5511 (N_5511,N_5258,N_5316);
nand U5512 (N_5512,N_5248,N_5259);
and U5513 (N_5513,N_5344,N_5305);
nand U5514 (N_5514,N_5355,N_5304);
xor U5515 (N_5515,N_5374,N_5252);
xor U5516 (N_5516,N_5292,N_5390);
and U5517 (N_5517,N_5257,N_5343);
xor U5518 (N_5518,N_5298,N_5284);
or U5519 (N_5519,N_5320,N_5291);
xor U5520 (N_5520,N_5286,N_5272);
xnor U5521 (N_5521,N_5287,N_5396);
and U5522 (N_5522,N_5302,N_5351);
xor U5523 (N_5523,N_5316,N_5240);
or U5524 (N_5524,N_5227,N_5260);
or U5525 (N_5525,N_5367,N_5347);
xnor U5526 (N_5526,N_5282,N_5288);
and U5527 (N_5527,N_5304,N_5271);
and U5528 (N_5528,N_5272,N_5201);
nor U5529 (N_5529,N_5338,N_5236);
and U5530 (N_5530,N_5286,N_5263);
xor U5531 (N_5531,N_5364,N_5360);
and U5532 (N_5532,N_5268,N_5301);
and U5533 (N_5533,N_5330,N_5253);
and U5534 (N_5534,N_5291,N_5256);
or U5535 (N_5535,N_5396,N_5235);
and U5536 (N_5536,N_5217,N_5257);
nand U5537 (N_5537,N_5345,N_5230);
nor U5538 (N_5538,N_5372,N_5209);
xor U5539 (N_5539,N_5227,N_5247);
xor U5540 (N_5540,N_5253,N_5204);
nor U5541 (N_5541,N_5224,N_5252);
xnor U5542 (N_5542,N_5387,N_5388);
nand U5543 (N_5543,N_5260,N_5316);
nor U5544 (N_5544,N_5356,N_5366);
nor U5545 (N_5545,N_5260,N_5217);
nand U5546 (N_5546,N_5225,N_5349);
nor U5547 (N_5547,N_5254,N_5313);
and U5548 (N_5548,N_5378,N_5328);
xor U5549 (N_5549,N_5287,N_5255);
and U5550 (N_5550,N_5374,N_5214);
and U5551 (N_5551,N_5265,N_5345);
xor U5552 (N_5552,N_5263,N_5374);
nor U5553 (N_5553,N_5218,N_5241);
and U5554 (N_5554,N_5221,N_5318);
or U5555 (N_5555,N_5336,N_5258);
nand U5556 (N_5556,N_5333,N_5224);
nor U5557 (N_5557,N_5246,N_5273);
nor U5558 (N_5558,N_5366,N_5281);
xnor U5559 (N_5559,N_5386,N_5345);
or U5560 (N_5560,N_5252,N_5280);
or U5561 (N_5561,N_5247,N_5371);
xnor U5562 (N_5562,N_5253,N_5357);
or U5563 (N_5563,N_5342,N_5286);
or U5564 (N_5564,N_5389,N_5295);
nand U5565 (N_5565,N_5325,N_5309);
nand U5566 (N_5566,N_5204,N_5290);
nand U5567 (N_5567,N_5265,N_5219);
nand U5568 (N_5568,N_5214,N_5309);
nor U5569 (N_5569,N_5227,N_5301);
and U5570 (N_5570,N_5221,N_5331);
and U5571 (N_5571,N_5352,N_5332);
or U5572 (N_5572,N_5296,N_5249);
nor U5573 (N_5573,N_5281,N_5370);
nor U5574 (N_5574,N_5260,N_5364);
or U5575 (N_5575,N_5354,N_5212);
nor U5576 (N_5576,N_5230,N_5362);
nand U5577 (N_5577,N_5392,N_5364);
nand U5578 (N_5578,N_5245,N_5335);
or U5579 (N_5579,N_5231,N_5391);
and U5580 (N_5580,N_5348,N_5232);
and U5581 (N_5581,N_5258,N_5226);
or U5582 (N_5582,N_5359,N_5347);
nand U5583 (N_5583,N_5200,N_5286);
nand U5584 (N_5584,N_5319,N_5205);
or U5585 (N_5585,N_5367,N_5290);
and U5586 (N_5586,N_5298,N_5375);
xnor U5587 (N_5587,N_5263,N_5237);
or U5588 (N_5588,N_5289,N_5296);
or U5589 (N_5589,N_5297,N_5361);
or U5590 (N_5590,N_5289,N_5228);
nand U5591 (N_5591,N_5275,N_5274);
nor U5592 (N_5592,N_5310,N_5386);
or U5593 (N_5593,N_5261,N_5259);
nand U5594 (N_5594,N_5205,N_5380);
and U5595 (N_5595,N_5201,N_5305);
and U5596 (N_5596,N_5270,N_5349);
nor U5597 (N_5597,N_5385,N_5286);
or U5598 (N_5598,N_5222,N_5330);
nor U5599 (N_5599,N_5397,N_5221);
nor U5600 (N_5600,N_5537,N_5482);
and U5601 (N_5601,N_5419,N_5509);
or U5602 (N_5602,N_5439,N_5458);
nand U5603 (N_5603,N_5498,N_5599);
nor U5604 (N_5604,N_5483,N_5581);
and U5605 (N_5605,N_5414,N_5400);
xnor U5606 (N_5606,N_5513,N_5531);
nand U5607 (N_5607,N_5427,N_5582);
and U5608 (N_5608,N_5487,N_5592);
nor U5609 (N_5609,N_5579,N_5437);
xnor U5610 (N_5610,N_5584,N_5429);
nor U5611 (N_5611,N_5523,N_5410);
and U5612 (N_5612,N_5535,N_5442);
xor U5613 (N_5613,N_5467,N_5401);
or U5614 (N_5614,N_5463,N_5445);
or U5615 (N_5615,N_5473,N_5415);
and U5616 (N_5616,N_5516,N_5542);
xnor U5617 (N_5617,N_5594,N_5540);
nand U5618 (N_5618,N_5580,N_5559);
nor U5619 (N_5619,N_5459,N_5511);
or U5620 (N_5620,N_5480,N_5461);
nor U5621 (N_5621,N_5472,N_5454);
xnor U5622 (N_5622,N_5424,N_5533);
xnor U5623 (N_5623,N_5402,N_5507);
and U5624 (N_5624,N_5525,N_5541);
xnor U5625 (N_5625,N_5563,N_5405);
nand U5626 (N_5626,N_5478,N_5574);
and U5627 (N_5627,N_5456,N_5460);
and U5628 (N_5628,N_5404,N_5502);
or U5629 (N_5629,N_5481,N_5505);
xor U5630 (N_5630,N_5500,N_5522);
and U5631 (N_5631,N_5504,N_5521);
nor U5632 (N_5632,N_5566,N_5543);
nor U5633 (N_5633,N_5553,N_5565);
xnor U5634 (N_5634,N_5422,N_5518);
and U5635 (N_5635,N_5433,N_5477);
nand U5636 (N_5636,N_5474,N_5564);
and U5637 (N_5637,N_5508,N_5434);
and U5638 (N_5638,N_5471,N_5587);
nor U5639 (N_5639,N_5417,N_5552);
xnor U5640 (N_5640,N_5503,N_5577);
xnor U5641 (N_5641,N_5519,N_5440);
nand U5642 (N_5642,N_5538,N_5554);
or U5643 (N_5643,N_5556,N_5493);
nor U5644 (N_5644,N_5598,N_5451);
and U5645 (N_5645,N_5431,N_5496);
and U5646 (N_5646,N_5506,N_5466);
nand U5647 (N_5647,N_5562,N_5444);
and U5648 (N_5648,N_5557,N_5425);
and U5649 (N_5649,N_5569,N_5452);
nor U5650 (N_5650,N_5426,N_5408);
or U5651 (N_5651,N_5485,N_5476);
xnor U5652 (N_5652,N_5443,N_5585);
and U5653 (N_5653,N_5413,N_5416);
or U5654 (N_5654,N_5561,N_5406);
nor U5655 (N_5655,N_5526,N_5407);
xor U5656 (N_5656,N_5589,N_5462);
nand U5657 (N_5657,N_5573,N_5436);
xnor U5658 (N_5658,N_5515,N_5491);
nand U5659 (N_5659,N_5501,N_5583);
nand U5660 (N_5660,N_5517,N_5484);
or U5661 (N_5661,N_5418,N_5403);
and U5662 (N_5662,N_5586,N_5411);
nand U5663 (N_5663,N_5597,N_5490);
xor U5664 (N_5664,N_5441,N_5412);
xnor U5665 (N_5665,N_5530,N_5423);
and U5666 (N_5666,N_5539,N_5568);
or U5667 (N_5667,N_5438,N_5432);
or U5668 (N_5668,N_5534,N_5449);
nand U5669 (N_5669,N_5495,N_5514);
xnor U5670 (N_5670,N_5492,N_5590);
or U5671 (N_5671,N_5486,N_5464);
nor U5672 (N_5672,N_5475,N_5548);
or U5673 (N_5673,N_5567,N_5595);
xnor U5674 (N_5674,N_5497,N_5421);
nand U5675 (N_5675,N_5450,N_5409);
xnor U5676 (N_5676,N_5524,N_5468);
nor U5677 (N_5677,N_5499,N_5494);
or U5678 (N_5678,N_5510,N_5455);
xor U5679 (N_5679,N_5558,N_5544);
nor U5680 (N_5680,N_5520,N_5546);
or U5681 (N_5681,N_5447,N_5536);
and U5682 (N_5682,N_5550,N_5572);
nand U5683 (N_5683,N_5560,N_5465);
and U5684 (N_5684,N_5512,N_5448);
and U5685 (N_5685,N_5470,N_5588);
or U5686 (N_5686,N_5532,N_5469);
nand U5687 (N_5687,N_5578,N_5575);
and U5688 (N_5688,N_5435,N_5527);
nand U5689 (N_5689,N_5571,N_5570);
nand U5690 (N_5690,N_5591,N_5549);
nor U5691 (N_5691,N_5593,N_5420);
and U5692 (N_5692,N_5488,N_5576);
and U5693 (N_5693,N_5430,N_5446);
nand U5694 (N_5694,N_5551,N_5489);
nand U5695 (N_5695,N_5453,N_5457);
or U5696 (N_5696,N_5528,N_5555);
nand U5697 (N_5697,N_5428,N_5547);
and U5698 (N_5698,N_5545,N_5479);
and U5699 (N_5699,N_5529,N_5596);
nor U5700 (N_5700,N_5504,N_5570);
nor U5701 (N_5701,N_5461,N_5539);
nor U5702 (N_5702,N_5581,N_5529);
nor U5703 (N_5703,N_5597,N_5433);
xnor U5704 (N_5704,N_5595,N_5439);
and U5705 (N_5705,N_5495,N_5522);
and U5706 (N_5706,N_5414,N_5520);
xnor U5707 (N_5707,N_5534,N_5549);
or U5708 (N_5708,N_5528,N_5409);
nand U5709 (N_5709,N_5583,N_5498);
xnor U5710 (N_5710,N_5552,N_5411);
or U5711 (N_5711,N_5538,N_5444);
nor U5712 (N_5712,N_5557,N_5470);
and U5713 (N_5713,N_5494,N_5549);
xnor U5714 (N_5714,N_5570,N_5448);
and U5715 (N_5715,N_5437,N_5564);
nand U5716 (N_5716,N_5507,N_5573);
or U5717 (N_5717,N_5513,N_5586);
nand U5718 (N_5718,N_5585,N_5518);
and U5719 (N_5719,N_5412,N_5578);
or U5720 (N_5720,N_5576,N_5515);
xor U5721 (N_5721,N_5422,N_5544);
nor U5722 (N_5722,N_5585,N_5476);
nor U5723 (N_5723,N_5569,N_5491);
xnor U5724 (N_5724,N_5520,N_5458);
xor U5725 (N_5725,N_5466,N_5597);
or U5726 (N_5726,N_5599,N_5442);
and U5727 (N_5727,N_5421,N_5593);
nand U5728 (N_5728,N_5489,N_5506);
and U5729 (N_5729,N_5513,N_5575);
or U5730 (N_5730,N_5526,N_5490);
nand U5731 (N_5731,N_5587,N_5402);
and U5732 (N_5732,N_5453,N_5452);
xnor U5733 (N_5733,N_5574,N_5425);
nor U5734 (N_5734,N_5542,N_5537);
or U5735 (N_5735,N_5509,N_5490);
nor U5736 (N_5736,N_5566,N_5594);
or U5737 (N_5737,N_5442,N_5559);
or U5738 (N_5738,N_5404,N_5570);
nand U5739 (N_5739,N_5430,N_5480);
and U5740 (N_5740,N_5590,N_5497);
and U5741 (N_5741,N_5428,N_5500);
or U5742 (N_5742,N_5484,N_5455);
nand U5743 (N_5743,N_5544,N_5456);
nand U5744 (N_5744,N_5516,N_5571);
or U5745 (N_5745,N_5547,N_5457);
nor U5746 (N_5746,N_5408,N_5404);
nor U5747 (N_5747,N_5524,N_5599);
xor U5748 (N_5748,N_5501,N_5568);
nand U5749 (N_5749,N_5538,N_5571);
nor U5750 (N_5750,N_5417,N_5407);
or U5751 (N_5751,N_5569,N_5550);
or U5752 (N_5752,N_5583,N_5470);
and U5753 (N_5753,N_5433,N_5439);
and U5754 (N_5754,N_5479,N_5415);
nand U5755 (N_5755,N_5443,N_5491);
nor U5756 (N_5756,N_5422,N_5458);
nand U5757 (N_5757,N_5419,N_5428);
nor U5758 (N_5758,N_5485,N_5498);
and U5759 (N_5759,N_5473,N_5512);
or U5760 (N_5760,N_5503,N_5412);
nor U5761 (N_5761,N_5402,N_5421);
and U5762 (N_5762,N_5507,N_5583);
and U5763 (N_5763,N_5520,N_5423);
nor U5764 (N_5764,N_5497,N_5456);
and U5765 (N_5765,N_5536,N_5487);
nand U5766 (N_5766,N_5590,N_5475);
and U5767 (N_5767,N_5435,N_5502);
nor U5768 (N_5768,N_5425,N_5529);
nand U5769 (N_5769,N_5503,N_5405);
nor U5770 (N_5770,N_5551,N_5546);
or U5771 (N_5771,N_5422,N_5438);
nand U5772 (N_5772,N_5445,N_5407);
or U5773 (N_5773,N_5584,N_5494);
and U5774 (N_5774,N_5556,N_5450);
xnor U5775 (N_5775,N_5449,N_5508);
xor U5776 (N_5776,N_5534,N_5598);
nor U5777 (N_5777,N_5460,N_5574);
or U5778 (N_5778,N_5518,N_5418);
nand U5779 (N_5779,N_5426,N_5436);
and U5780 (N_5780,N_5497,N_5515);
nand U5781 (N_5781,N_5431,N_5500);
nor U5782 (N_5782,N_5437,N_5508);
nand U5783 (N_5783,N_5444,N_5586);
nor U5784 (N_5784,N_5473,N_5545);
and U5785 (N_5785,N_5443,N_5436);
nand U5786 (N_5786,N_5521,N_5591);
nand U5787 (N_5787,N_5580,N_5458);
or U5788 (N_5788,N_5465,N_5548);
or U5789 (N_5789,N_5568,N_5547);
nor U5790 (N_5790,N_5421,N_5507);
and U5791 (N_5791,N_5451,N_5446);
or U5792 (N_5792,N_5518,N_5557);
and U5793 (N_5793,N_5488,N_5455);
and U5794 (N_5794,N_5562,N_5544);
nor U5795 (N_5795,N_5520,N_5518);
xor U5796 (N_5796,N_5587,N_5448);
or U5797 (N_5797,N_5545,N_5470);
and U5798 (N_5798,N_5402,N_5556);
and U5799 (N_5799,N_5514,N_5426);
and U5800 (N_5800,N_5670,N_5646);
or U5801 (N_5801,N_5685,N_5633);
xnor U5802 (N_5802,N_5627,N_5796);
nor U5803 (N_5803,N_5775,N_5612);
nand U5804 (N_5804,N_5614,N_5654);
nor U5805 (N_5805,N_5798,N_5689);
xnor U5806 (N_5806,N_5707,N_5648);
nor U5807 (N_5807,N_5766,N_5755);
and U5808 (N_5808,N_5722,N_5601);
nor U5809 (N_5809,N_5708,N_5740);
nand U5810 (N_5810,N_5721,N_5691);
nand U5811 (N_5811,N_5695,N_5692);
or U5812 (N_5812,N_5743,N_5621);
or U5813 (N_5813,N_5784,N_5678);
or U5814 (N_5814,N_5710,N_5651);
or U5815 (N_5815,N_5632,N_5620);
and U5816 (N_5816,N_5616,N_5647);
xor U5817 (N_5817,N_5644,N_5603);
xnor U5818 (N_5818,N_5688,N_5697);
nand U5819 (N_5819,N_5694,N_5676);
xnor U5820 (N_5820,N_5615,N_5609);
or U5821 (N_5821,N_5600,N_5742);
or U5822 (N_5822,N_5667,N_5605);
nor U5823 (N_5823,N_5720,N_5679);
nor U5824 (N_5824,N_5725,N_5636);
and U5825 (N_5825,N_5764,N_5717);
nand U5826 (N_5826,N_5680,N_5690);
or U5827 (N_5827,N_5778,N_5643);
xnor U5828 (N_5828,N_5604,N_5661);
nor U5829 (N_5829,N_5746,N_5650);
nand U5830 (N_5830,N_5738,N_5669);
or U5831 (N_5831,N_5791,N_5788);
or U5832 (N_5832,N_5728,N_5681);
nand U5833 (N_5833,N_5663,N_5682);
and U5834 (N_5834,N_5671,N_5771);
nor U5835 (N_5835,N_5745,N_5630);
or U5836 (N_5836,N_5705,N_5741);
nor U5837 (N_5837,N_5626,N_5727);
xnor U5838 (N_5838,N_5662,N_5629);
or U5839 (N_5839,N_5739,N_5700);
nor U5840 (N_5840,N_5655,N_5625);
xor U5841 (N_5841,N_5729,N_5698);
nand U5842 (N_5842,N_5653,N_5761);
nand U5843 (N_5843,N_5673,N_5706);
nor U5844 (N_5844,N_5696,N_5617);
xor U5845 (N_5845,N_5723,N_5768);
or U5846 (N_5846,N_5731,N_5760);
or U5847 (N_5847,N_5776,N_5749);
and U5848 (N_5848,N_5641,N_5703);
and U5849 (N_5849,N_5767,N_5783);
nor U5850 (N_5850,N_5790,N_5757);
nand U5851 (N_5851,N_5718,N_5726);
nand U5852 (N_5852,N_5715,N_5638);
nand U5853 (N_5853,N_5716,N_5665);
nor U5854 (N_5854,N_5734,N_5787);
or U5855 (N_5855,N_5779,N_5635);
nor U5856 (N_5856,N_5735,N_5704);
xnor U5857 (N_5857,N_5631,N_5730);
nor U5858 (N_5858,N_5782,N_5637);
nand U5859 (N_5859,N_5709,N_5754);
or U5860 (N_5860,N_5756,N_5795);
nand U5861 (N_5861,N_5758,N_5732);
xnor U5862 (N_5862,N_5701,N_5733);
nand U5863 (N_5863,N_5719,N_5724);
nor U5864 (N_5864,N_5780,N_5677);
nor U5865 (N_5865,N_5652,N_5765);
or U5866 (N_5866,N_5659,N_5753);
nor U5867 (N_5867,N_5797,N_5687);
nand U5868 (N_5868,N_5750,N_5640);
and U5869 (N_5869,N_5675,N_5713);
nor U5870 (N_5870,N_5763,N_5759);
or U5871 (N_5871,N_5613,N_5672);
or U5872 (N_5872,N_5785,N_5607);
xor U5873 (N_5873,N_5789,N_5657);
nand U5874 (N_5874,N_5792,N_5628);
or U5875 (N_5875,N_5751,N_5714);
or U5876 (N_5876,N_5793,N_5747);
nand U5877 (N_5877,N_5712,N_5799);
or U5878 (N_5878,N_5611,N_5736);
nand U5879 (N_5879,N_5664,N_5770);
nor U5880 (N_5880,N_5602,N_5666);
or U5881 (N_5881,N_5606,N_5686);
and U5882 (N_5882,N_5610,N_5699);
and U5883 (N_5883,N_5777,N_5711);
or U5884 (N_5884,N_5668,N_5658);
nand U5885 (N_5885,N_5769,N_5656);
or U5886 (N_5886,N_5619,N_5737);
and U5887 (N_5887,N_5649,N_5752);
and U5888 (N_5888,N_5642,N_5702);
nor U5889 (N_5889,N_5773,N_5684);
nand U5890 (N_5890,N_5639,N_5744);
and U5891 (N_5891,N_5634,N_5660);
and U5892 (N_5892,N_5786,N_5618);
xor U5893 (N_5893,N_5683,N_5762);
or U5894 (N_5894,N_5623,N_5645);
and U5895 (N_5895,N_5624,N_5693);
and U5896 (N_5896,N_5748,N_5781);
nand U5897 (N_5897,N_5774,N_5772);
xnor U5898 (N_5898,N_5794,N_5622);
nor U5899 (N_5899,N_5608,N_5674);
or U5900 (N_5900,N_5646,N_5606);
nor U5901 (N_5901,N_5681,N_5695);
nor U5902 (N_5902,N_5758,N_5777);
nand U5903 (N_5903,N_5761,N_5707);
xnor U5904 (N_5904,N_5787,N_5751);
nand U5905 (N_5905,N_5757,N_5674);
xnor U5906 (N_5906,N_5730,N_5731);
nor U5907 (N_5907,N_5750,N_5739);
xnor U5908 (N_5908,N_5750,N_5796);
and U5909 (N_5909,N_5613,N_5733);
xnor U5910 (N_5910,N_5734,N_5649);
xnor U5911 (N_5911,N_5649,N_5756);
or U5912 (N_5912,N_5716,N_5640);
xor U5913 (N_5913,N_5604,N_5675);
nand U5914 (N_5914,N_5677,N_5628);
nand U5915 (N_5915,N_5704,N_5650);
xnor U5916 (N_5916,N_5687,N_5662);
nor U5917 (N_5917,N_5624,N_5750);
or U5918 (N_5918,N_5718,N_5710);
nor U5919 (N_5919,N_5743,N_5674);
nor U5920 (N_5920,N_5677,N_5764);
or U5921 (N_5921,N_5782,N_5689);
and U5922 (N_5922,N_5790,N_5674);
or U5923 (N_5923,N_5711,N_5716);
xor U5924 (N_5924,N_5725,N_5692);
nor U5925 (N_5925,N_5761,N_5658);
nor U5926 (N_5926,N_5662,N_5757);
or U5927 (N_5927,N_5646,N_5647);
or U5928 (N_5928,N_5642,N_5796);
or U5929 (N_5929,N_5675,N_5622);
nand U5930 (N_5930,N_5727,N_5711);
nor U5931 (N_5931,N_5617,N_5782);
nor U5932 (N_5932,N_5660,N_5720);
and U5933 (N_5933,N_5638,N_5664);
and U5934 (N_5934,N_5784,N_5683);
and U5935 (N_5935,N_5716,N_5731);
or U5936 (N_5936,N_5701,N_5646);
nand U5937 (N_5937,N_5761,N_5690);
nand U5938 (N_5938,N_5614,N_5636);
nand U5939 (N_5939,N_5681,N_5730);
and U5940 (N_5940,N_5734,N_5713);
xnor U5941 (N_5941,N_5651,N_5624);
xnor U5942 (N_5942,N_5642,N_5763);
nor U5943 (N_5943,N_5644,N_5733);
xor U5944 (N_5944,N_5649,N_5746);
and U5945 (N_5945,N_5788,N_5674);
nand U5946 (N_5946,N_5710,N_5643);
or U5947 (N_5947,N_5676,N_5697);
and U5948 (N_5948,N_5682,N_5766);
nand U5949 (N_5949,N_5611,N_5673);
nand U5950 (N_5950,N_5738,N_5732);
and U5951 (N_5951,N_5752,N_5778);
xnor U5952 (N_5952,N_5696,N_5686);
nor U5953 (N_5953,N_5679,N_5602);
xor U5954 (N_5954,N_5695,N_5756);
or U5955 (N_5955,N_5794,N_5650);
and U5956 (N_5956,N_5672,N_5619);
and U5957 (N_5957,N_5676,N_5678);
nand U5958 (N_5958,N_5641,N_5672);
xnor U5959 (N_5959,N_5719,N_5725);
and U5960 (N_5960,N_5665,N_5680);
or U5961 (N_5961,N_5646,N_5691);
and U5962 (N_5962,N_5623,N_5627);
nand U5963 (N_5963,N_5731,N_5771);
xor U5964 (N_5964,N_5743,N_5763);
or U5965 (N_5965,N_5684,N_5677);
or U5966 (N_5966,N_5649,N_5791);
nand U5967 (N_5967,N_5627,N_5603);
xnor U5968 (N_5968,N_5715,N_5797);
or U5969 (N_5969,N_5792,N_5780);
or U5970 (N_5970,N_5758,N_5711);
and U5971 (N_5971,N_5672,N_5674);
and U5972 (N_5972,N_5790,N_5673);
nor U5973 (N_5973,N_5674,N_5711);
xnor U5974 (N_5974,N_5644,N_5729);
nand U5975 (N_5975,N_5613,N_5799);
nand U5976 (N_5976,N_5702,N_5711);
and U5977 (N_5977,N_5767,N_5782);
nand U5978 (N_5978,N_5699,N_5619);
nand U5979 (N_5979,N_5702,N_5649);
xnor U5980 (N_5980,N_5638,N_5615);
nor U5981 (N_5981,N_5641,N_5637);
and U5982 (N_5982,N_5695,N_5677);
nor U5983 (N_5983,N_5605,N_5613);
xor U5984 (N_5984,N_5645,N_5659);
xnor U5985 (N_5985,N_5725,N_5710);
or U5986 (N_5986,N_5715,N_5791);
and U5987 (N_5987,N_5695,N_5721);
nand U5988 (N_5988,N_5628,N_5719);
nor U5989 (N_5989,N_5758,N_5753);
nor U5990 (N_5990,N_5658,N_5622);
or U5991 (N_5991,N_5679,N_5702);
xor U5992 (N_5992,N_5640,N_5789);
or U5993 (N_5993,N_5747,N_5666);
nor U5994 (N_5994,N_5640,N_5609);
and U5995 (N_5995,N_5628,N_5740);
xor U5996 (N_5996,N_5737,N_5629);
nor U5997 (N_5997,N_5681,N_5671);
xor U5998 (N_5998,N_5602,N_5655);
or U5999 (N_5999,N_5797,N_5600);
xnor U6000 (N_6000,N_5879,N_5815);
nor U6001 (N_6001,N_5920,N_5900);
nor U6002 (N_6002,N_5910,N_5896);
nand U6003 (N_6003,N_5915,N_5913);
or U6004 (N_6004,N_5931,N_5943);
xnor U6005 (N_6005,N_5829,N_5934);
nand U6006 (N_6006,N_5824,N_5969);
and U6007 (N_6007,N_5924,N_5919);
xor U6008 (N_6008,N_5828,N_5965);
nor U6009 (N_6009,N_5821,N_5908);
nor U6010 (N_6010,N_5987,N_5857);
nand U6011 (N_6011,N_5819,N_5945);
and U6012 (N_6012,N_5817,N_5820);
xor U6013 (N_6013,N_5818,N_5802);
and U6014 (N_6014,N_5894,N_5854);
and U6015 (N_6015,N_5912,N_5923);
xor U6016 (N_6016,N_5993,N_5907);
nand U6017 (N_6017,N_5809,N_5864);
or U6018 (N_6018,N_5921,N_5833);
nor U6019 (N_6019,N_5891,N_5886);
nor U6020 (N_6020,N_5976,N_5994);
nor U6021 (N_6021,N_5823,N_5835);
or U6022 (N_6022,N_5911,N_5939);
nand U6023 (N_6023,N_5850,N_5859);
xor U6024 (N_6024,N_5866,N_5841);
nor U6025 (N_6025,N_5816,N_5812);
nor U6026 (N_6026,N_5909,N_5893);
and U6027 (N_6027,N_5877,N_5884);
nand U6028 (N_6028,N_5989,N_5863);
nand U6029 (N_6029,N_5941,N_5960);
or U6030 (N_6030,N_5839,N_5843);
nor U6031 (N_6031,N_5916,N_5806);
nand U6032 (N_6032,N_5871,N_5831);
or U6033 (N_6033,N_5810,N_5926);
xnor U6034 (N_6034,N_5855,N_5801);
nor U6035 (N_6035,N_5875,N_5992);
nand U6036 (N_6036,N_5914,N_5813);
or U6037 (N_6037,N_5800,N_5996);
and U6038 (N_6038,N_5856,N_5870);
or U6039 (N_6039,N_5984,N_5868);
nand U6040 (N_6040,N_5962,N_5963);
nand U6041 (N_6041,N_5959,N_5917);
nor U6042 (N_6042,N_5957,N_5973);
xor U6043 (N_6043,N_5890,N_5938);
nor U6044 (N_6044,N_5882,N_5929);
and U6045 (N_6045,N_5844,N_5822);
nand U6046 (N_6046,N_5967,N_5972);
nand U6047 (N_6047,N_5861,N_5954);
or U6048 (N_6048,N_5805,N_5807);
xor U6049 (N_6049,N_5979,N_5880);
or U6050 (N_6050,N_5928,N_5885);
nor U6051 (N_6051,N_5949,N_5860);
nand U6052 (N_6052,N_5922,N_5936);
nor U6053 (N_6053,N_5889,N_5899);
and U6054 (N_6054,N_5991,N_5947);
nor U6055 (N_6055,N_5903,N_5955);
or U6056 (N_6056,N_5874,N_5958);
xnor U6057 (N_6057,N_5933,N_5999);
xor U6058 (N_6058,N_5836,N_5966);
nor U6059 (N_6059,N_5825,N_5940);
nor U6060 (N_6060,N_5988,N_5930);
nand U6061 (N_6061,N_5838,N_5853);
or U6062 (N_6062,N_5847,N_5881);
or U6063 (N_6063,N_5851,N_5951);
and U6064 (N_6064,N_5830,N_5873);
or U6065 (N_6065,N_5837,N_5977);
xor U6066 (N_6066,N_5832,N_5937);
xnor U6067 (N_6067,N_5803,N_5983);
or U6068 (N_6068,N_5932,N_5840);
nor U6069 (N_6069,N_5892,N_5804);
nand U6070 (N_6070,N_5953,N_5952);
and U6071 (N_6071,N_5826,N_5998);
and U6072 (N_6072,N_5950,N_5981);
or U6073 (N_6073,N_5901,N_5872);
and U6074 (N_6074,N_5846,N_5865);
nor U6075 (N_6075,N_5867,N_5985);
nor U6076 (N_6076,N_5869,N_5849);
or U6077 (N_6077,N_5942,N_5927);
nor U6078 (N_6078,N_5878,N_5834);
and U6079 (N_6079,N_5898,N_5975);
nor U6080 (N_6080,N_5961,N_5980);
and U6081 (N_6081,N_5814,N_5948);
nor U6082 (N_6082,N_5827,N_5968);
nor U6083 (N_6083,N_5995,N_5997);
nor U6084 (N_6084,N_5862,N_5883);
nand U6085 (N_6085,N_5935,N_5971);
xor U6086 (N_6086,N_5978,N_5842);
nor U6087 (N_6087,N_5974,N_5970);
xnor U6088 (N_6088,N_5904,N_5990);
xor U6089 (N_6089,N_5986,N_5897);
or U6090 (N_6090,N_5876,N_5811);
nand U6091 (N_6091,N_5956,N_5964);
or U6092 (N_6092,N_5888,N_5845);
nor U6093 (N_6093,N_5895,N_5887);
or U6094 (N_6094,N_5905,N_5848);
nand U6095 (N_6095,N_5852,N_5906);
or U6096 (N_6096,N_5982,N_5808);
nand U6097 (N_6097,N_5946,N_5944);
xnor U6098 (N_6098,N_5858,N_5918);
xor U6099 (N_6099,N_5925,N_5902);
or U6100 (N_6100,N_5998,N_5862);
or U6101 (N_6101,N_5936,N_5998);
and U6102 (N_6102,N_5941,N_5858);
and U6103 (N_6103,N_5947,N_5873);
or U6104 (N_6104,N_5994,N_5977);
or U6105 (N_6105,N_5976,N_5956);
nand U6106 (N_6106,N_5878,N_5846);
xnor U6107 (N_6107,N_5896,N_5902);
and U6108 (N_6108,N_5802,N_5955);
and U6109 (N_6109,N_5802,N_5980);
xnor U6110 (N_6110,N_5822,N_5900);
nor U6111 (N_6111,N_5940,N_5894);
or U6112 (N_6112,N_5992,N_5969);
xor U6113 (N_6113,N_5842,N_5876);
and U6114 (N_6114,N_5907,N_5963);
and U6115 (N_6115,N_5928,N_5858);
nand U6116 (N_6116,N_5861,N_5958);
xnor U6117 (N_6117,N_5842,N_5802);
nor U6118 (N_6118,N_5872,N_5810);
nor U6119 (N_6119,N_5855,N_5995);
and U6120 (N_6120,N_5835,N_5991);
nor U6121 (N_6121,N_5832,N_5903);
nand U6122 (N_6122,N_5975,N_5809);
or U6123 (N_6123,N_5890,N_5919);
xnor U6124 (N_6124,N_5845,N_5873);
or U6125 (N_6125,N_5910,N_5820);
or U6126 (N_6126,N_5823,N_5963);
and U6127 (N_6127,N_5866,N_5890);
nor U6128 (N_6128,N_5883,N_5913);
nand U6129 (N_6129,N_5950,N_5965);
nor U6130 (N_6130,N_5858,N_5816);
xor U6131 (N_6131,N_5976,N_5987);
nor U6132 (N_6132,N_5911,N_5871);
and U6133 (N_6133,N_5841,N_5842);
and U6134 (N_6134,N_5911,N_5968);
xor U6135 (N_6135,N_5900,N_5927);
nor U6136 (N_6136,N_5814,N_5959);
or U6137 (N_6137,N_5835,N_5945);
nand U6138 (N_6138,N_5909,N_5905);
nand U6139 (N_6139,N_5804,N_5886);
nor U6140 (N_6140,N_5803,N_5807);
and U6141 (N_6141,N_5934,N_5926);
nor U6142 (N_6142,N_5836,N_5904);
nand U6143 (N_6143,N_5925,N_5907);
nor U6144 (N_6144,N_5822,N_5953);
xor U6145 (N_6145,N_5899,N_5975);
nand U6146 (N_6146,N_5996,N_5938);
and U6147 (N_6147,N_5944,N_5985);
nand U6148 (N_6148,N_5907,N_5912);
nor U6149 (N_6149,N_5813,N_5833);
nand U6150 (N_6150,N_5834,N_5877);
and U6151 (N_6151,N_5859,N_5892);
nor U6152 (N_6152,N_5938,N_5818);
nand U6153 (N_6153,N_5968,N_5937);
or U6154 (N_6154,N_5988,N_5835);
nor U6155 (N_6155,N_5869,N_5982);
nor U6156 (N_6156,N_5840,N_5947);
and U6157 (N_6157,N_5966,N_5936);
nor U6158 (N_6158,N_5935,N_5821);
nand U6159 (N_6159,N_5803,N_5877);
and U6160 (N_6160,N_5874,N_5867);
or U6161 (N_6161,N_5874,N_5853);
nor U6162 (N_6162,N_5914,N_5963);
nor U6163 (N_6163,N_5965,N_5919);
and U6164 (N_6164,N_5849,N_5827);
nand U6165 (N_6165,N_5950,N_5941);
nand U6166 (N_6166,N_5896,N_5909);
nand U6167 (N_6167,N_5998,N_5863);
or U6168 (N_6168,N_5835,N_5854);
xor U6169 (N_6169,N_5823,N_5970);
and U6170 (N_6170,N_5931,N_5867);
xor U6171 (N_6171,N_5806,N_5890);
xnor U6172 (N_6172,N_5861,N_5806);
or U6173 (N_6173,N_5892,N_5884);
or U6174 (N_6174,N_5909,N_5827);
nor U6175 (N_6175,N_5969,N_5918);
xnor U6176 (N_6176,N_5923,N_5835);
and U6177 (N_6177,N_5952,N_5808);
xor U6178 (N_6178,N_5887,N_5821);
or U6179 (N_6179,N_5884,N_5887);
xor U6180 (N_6180,N_5836,N_5954);
or U6181 (N_6181,N_5804,N_5874);
nor U6182 (N_6182,N_5945,N_5816);
nor U6183 (N_6183,N_5931,N_5847);
and U6184 (N_6184,N_5808,N_5936);
xnor U6185 (N_6185,N_5889,N_5942);
or U6186 (N_6186,N_5808,N_5856);
nand U6187 (N_6187,N_5913,N_5804);
or U6188 (N_6188,N_5982,N_5942);
xnor U6189 (N_6189,N_5978,N_5993);
xor U6190 (N_6190,N_5901,N_5971);
nor U6191 (N_6191,N_5844,N_5885);
and U6192 (N_6192,N_5909,N_5924);
nand U6193 (N_6193,N_5825,N_5879);
xor U6194 (N_6194,N_5904,N_5868);
nand U6195 (N_6195,N_5990,N_5961);
and U6196 (N_6196,N_5833,N_5983);
and U6197 (N_6197,N_5838,N_5888);
nand U6198 (N_6198,N_5979,N_5861);
or U6199 (N_6199,N_5917,N_5900);
xor U6200 (N_6200,N_6160,N_6167);
nand U6201 (N_6201,N_6098,N_6179);
or U6202 (N_6202,N_6030,N_6162);
and U6203 (N_6203,N_6174,N_6099);
or U6204 (N_6204,N_6014,N_6156);
nor U6205 (N_6205,N_6053,N_6199);
nor U6206 (N_6206,N_6127,N_6012);
nand U6207 (N_6207,N_6003,N_6103);
and U6208 (N_6208,N_6059,N_6027);
and U6209 (N_6209,N_6018,N_6117);
nand U6210 (N_6210,N_6061,N_6152);
and U6211 (N_6211,N_6133,N_6008);
and U6212 (N_6212,N_6040,N_6191);
and U6213 (N_6213,N_6146,N_6197);
or U6214 (N_6214,N_6187,N_6196);
or U6215 (N_6215,N_6132,N_6121);
nor U6216 (N_6216,N_6138,N_6148);
xor U6217 (N_6217,N_6114,N_6056);
and U6218 (N_6218,N_6048,N_6120);
and U6219 (N_6219,N_6108,N_6131);
nand U6220 (N_6220,N_6021,N_6052);
nand U6221 (N_6221,N_6169,N_6034);
or U6222 (N_6222,N_6136,N_6011);
xor U6223 (N_6223,N_6047,N_6070);
nor U6224 (N_6224,N_6043,N_6150);
or U6225 (N_6225,N_6178,N_6172);
or U6226 (N_6226,N_6147,N_6073);
nand U6227 (N_6227,N_6057,N_6033);
and U6228 (N_6228,N_6084,N_6194);
and U6229 (N_6229,N_6088,N_6062);
or U6230 (N_6230,N_6089,N_6119);
and U6231 (N_6231,N_6016,N_6063);
or U6232 (N_6232,N_6046,N_6159);
and U6233 (N_6233,N_6188,N_6115);
or U6234 (N_6234,N_6015,N_6094);
nand U6235 (N_6235,N_6154,N_6183);
or U6236 (N_6236,N_6175,N_6109);
nor U6237 (N_6237,N_6066,N_6065);
or U6238 (N_6238,N_6190,N_6182);
xnor U6239 (N_6239,N_6102,N_6122);
xnor U6240 (N_6240,N_6134,N_6010);
nor U6241 (N_6241,N_6141,N_6041);
or U6242 (N_6242,N_6130,N_6069);
or U6243 (N_6243,N_6013,N_6139);
xnor U6244 (N_6244,N_6144,N_6051);
and U6245 (N_6245,N_6189,N_6118);
nor U6246 (N_6246,N_6195,N_6123);
nand U6247 (N_6247,N_6017,N_6142);
nor U6248 (N_6248,N_6129,N_6180);
and U6249 (N_6249,N_6153,N_6166);
or U6250 (N_6250,N_6173,N_6105);
and U6251 (N_6251,N_6028,N_6185);
nor U6252 (N_6252,N_6145,N_6002);
xor U6253 (N_6253,N_6176,N_6091);
nor U6254 (N_6254,N_6093,N_6067);
nand U6255 (N_6255,N_6083,N_6022);
and U6256 (N_6256,N_6023,N_6079);
nor U6257 (N_6257,N_6072,N_6006);
or U6258 (N_6258,N_6076,N_6192);
or U6259 (N_6259,N_6000,N_6074);
nor U6260 (N_6260,N_6039,N_6135);
or U6261 (N_6261,N_6112,N_6140);
nor U6262 (N_6262,N_6177,N_6110);
nand U6263 (N_6263,N_6025,N_6020);
and U6264 (N_6264,N_6068,N_6042);
nand U6265 (N_6265,N_6029,N_6031);
xor U6266 (N_6266,N_6038,N_6184);
and U6267 (N_6267,N_6071,N_6087);
nand U6268 (N_6268,N_6035,N_6186);
xor U6269 (N_6269,N_6157,N_6168);
or U6270 (N_6270,N_6170,N_6124);
or U6271 (N_6271,N_6004,N_6106);
nor U6272 (N_6272,N_6126,N_6009);
nand U6273 (N_6273,N_6163,N_6045);
and U6274 (N_6274,N_6155,N_6007);
and U6275 (N_6275,N_6037,N_6036);
nor U6276 (N_6276,N_6100,N_6097);
nor U6277 (N_6277,N_6113,N_6104);
xor U6278 (N_6278,N_6151,N_6095);
and U6279 (N_6279,N_6143,N_6198);
xnor U6280 (N_6280,N_6181,N_6060);
xor U6281 (N_6281,N_6055,N_6081);
or U6282 (N_6282,N_6077,N_6049);
nor U6283 (N_6283,N_6161,N_6001);
or U6284 (N_6284,N_6086,N_6085);
and U6285 (N_6285,N_6024,N_6050);
or U6286 (N_6286,N_6075,N_6107);
nor U6287 (N_6287,N_6044,N_6054);
or U6288 (N_6288,N_6090,N_6101);
or U6289 (N_6289,N_6082,N_6137);
xor U6290 (N_6290,N_6019,N_6171);
nand U6291 (N_6291,N_6026,N_6096);
nor U6292 (N_6292,N_6064,N_6165);
nor U6293 (N_6293,N_6193,N_6032);
nand U6294 (N_6294,N_6092,N_6111);
nor U6295 (N_6295,N_6125,N_6078);
xor U6296 (N_6296,N_6164,N_6005);
xor U6297 (N_6297,N_6058,N_6116);
or U6298 (N_6298,N_6158,N_6149);
or U6299 (N_6299,N_6128,N_6080);
or U6300 (N_6300,N_6118,N_6019);
or U6301 (N_6301,N_6144,N_6031);
and U6302 (N_6302,N_6047,N_6129);
or U6303 (N_6303,N_6166,N_6119);
or U6304 (N_6304,N_6147,N_6199);
nand U6305 (N_6305,N_6034,N_6089);
and U6306 (N_6306,N_6086,N_6132);
and U6307 (N_6307,N_6045,N_6150);
and U6308 (N_6308,N_6012,N_6040);
nand U6309 (N_6309,N_6121,N_6037);
nor U6310 (N_6310,N_6180,N_6015);
or U6311 (N_6311,N_6176,N_6029);
nor U6312 (N_6312,N_6096,N_6183);
or U6313 (N_6313,N_6135,N_6084);
and U6314 (N_6314,N_6138,N_6046);
nand U6315 (N_6315,N_6156,N_6044);
xor U6316 (N_6316,N_6110,N_6132);
or U6317 (N_6317,N_6121,N_6035);
xnor U6318 (N_6318,N_6053,N_6181);
nor U6319 (N_6319,N_6051,N_6016);
or U6320 (N_6320,N_6083,N_6155);
or U6321 (N_6321,N_6113,N_6077);
xor U6322 (N_6322,N_6146,N_6147);
and U6323 (N_6323,N_6070,N_6062);
or U6324 (N_6324,N_6163,N_6115);
or U6325 (N_6325,N_6056,N_6141);
nor U6326 (N_6326,N_6168,N_6084);
xor U6327 (N_6327,N_6157,N_6146);
and U6328 (N_6328,N_6098,N_6196);
nand U6329 (N_6329,N_6039,N_6003);
xnor U6330 (N_6330,N_6168,N_6102);
nand U6331 (N_6331,N_6118,N_6040);
nand U6332 (N_6332,N_6022,N_6018);
xor U6333 (N_6333,N_6180,N_6062);
and U6334 (N_6334,N_6003,N_6038);
nor U6335 (N_6335,N_6198,N_6055);
nand U6336 (N_6336,N_6065,N_6199);
nand U6337 (N_6337,N_6121,N_6186);
nand U6338 (N_6338,N_6032,N_6111);
nor U6339 (N_6339,N_6161,N_6185);
or U6340 (N_6340,N_6009,N_6139);
nand U6341 (N_6341,N_6011,N_6115);
and U6342 (N_6342,N_6134,N_6152);
or U6343 (N_6343,N_6199,N_6074);
and U6344 (N_6344,N_6021,N_6048);
or U6345 (N_6345,N_6002,N_6015);
or U6346 (N_6346,N_6015,N_6197);
and U6347 (N_6347,N_6027,N_6041);
nor U6348 (N_6348,N_6190,N_6155);
nand U6349 (N_6349,N_6088,N_6161);
or U6350 (N_6350,N_6148,N_6062);
and U6351 (N_6351,N_6089,N_6031);
and U6352 (N_6352,N_6198,N_6085);
or U6353 (N_6353,N_6128,N_6178);
or U6354 (N_6354,N_6065,N_6116);
nor U6355 (N_6355,N_6045,N_6004);
nor U6356 (N_6356,N_6037,N_6138);
xor U6357 (N_6357,N_6155,N_6008);
nand U6358 (N_6358,N_6188,N_6101);
xor U6359 (N_6359,N_6124,N_6096);
or U6360 (N_6360,N_6075,N_6074);
xnor U6361 (N_6361,N_6134,N_6024);
and U6362 (N_6362,N_6047,N_6192);
nor U6363 (N_6363,N_6057,N_6058);
xnor U6364 (N_6364,N_6011,N_6023);
nor U6365 (N_6365,N_6116,N_6063);
or U6366 (N_6366,N_6103,N_6087);
xor U6367 (N_6367,N_6185,N_6175);
nand U6368 (N_6368,N_6041,N_6037);
or U6369 (N_6369,N_6074,N_6116);
nand U6370 (N_6370,N_6123,N_6196);
or U6371 (N_6371,N_6147,N_6001);
or U6372 (N_6372,N_6122,N_6167);
nor U6373 (N_6373,N_6138,N_6146);
and U6374 (N_6374,N_6028,N_6135);
and U6375 (N_6375,N_6093,N_6189);
nand U6376 (N_6376,N_6148,N_6118);
nand U6377 (N_6377,N_6133,N_6159);
nor U6378 (N_6378,N_6078,N_6023);
or U6379 (N_6379,N_6015,N_6006);
nor U6380 (N_6380,N_6040,N_6058);
nor U6381 (N_6381,N_6139,N_6058);
nor U6382 (N_6382,N_6153,N_6081);
nand U6383 (N_6383,N_6080,N_6038);
and U6384 (N_6384,N_6148,N_6105);
or U6385 (N_6385,N_6124,N_6073);
xnor U6386 (N_6386,N_6168,N_6113);
nand U6387 (N_6387,N_6061,N_6009);
or U6388 (N_6388,N_6019,N_6076);
nand U6389 (N_6389,N_6130,N_6171);
xor U6390 (N_6390,N_6126,N_6045);
xnor U6391 (N_6391,N_6180,N_6001);
nor U6392 (N_6392,N_6073,N_6022);
xnor U6393 (N_6393,N_6056,N_6171);
nand U6394 (N_6394,N_6022,N_6157);
xor U6395 (N_6395,N_6037,N_6161);
nand U6396 (N_6396,N_6058,N_6110);
xnor U6397 (N_6397,N_6166,N_6102);
nor U6398 (N_6398,N_6199,N_6110);
nand U6399 (N_6399,N_6124,N_6008);
or U6400 (N_6400,N_6267,N_6340);
and U6401 (N_6401,N_6308,N_6322);
and U6402 (N_6402,N_6235,N_6251);
nand U6403 (N_6403,N_6239,N_6290);
and U6404 (N_6404,N_6215,N_6247);
and U6405 (N_6405,N_6213,N_6310);
xnor U6406 (N_6406,N_6311,N_6266);
or U6407 (N_6407,N_6362,N_6349);
and U6408 (N_6408,N_6216,N_6202);
xor U6409 (N_6409,N_6241,N_6363);
and U6410 (N_6410,N_6350,N_6384);
xnor U6411 (N_6411,N_6209,N_6244);
or U6412 (N_6412,N_6254,N_6307);
or U6413 (N_6413,N_6393,N_6212);
xor U6414 (N_6414,N_6395,N_6364);
or U6415 (N_6415,N_6260,N_6283);
and U6416 (N_6416,N_6242,N_6268);
or U6417 (N_6417,N_6305,N_6234);
nand U6418 (N_6418,N_6361,N_6275);
and U6419 (N_6419,N_6385,N_6342);
nand U6420 (N_6420,N_6288,N_6371);
and U6421 (N_6421,N_6358,N_6348);
or U6422 (N_6422,N_6324,N_6331);
xor U6423 (N_6423,N_6316,N_6299);
and U6424 (N_6424,N_6300,N_6294);
or U6425 (N_6425,N_6214,N_6200);
and U6426 (N_6426,N_6265,N_6336);
nand U6427 (N_6427,N_6238,N_6204);
nand U6428 (N_6428,N_6327,N_6297);
or U6429 (N_6429,N_6313,N_6296);
nand U6430 (N_6430,N_6286,N_6326);
or U6431 (N_6431,N_6383,N_6298);
nor U6432 (N_6432,N_6236,N_6328);
and U6433 (N_6433,N_6323,N_6388);
xor U6434 (N_6434,N_6334,N_6227);
or U6435 (N_6435,N_6245,N_6220);
and U6436 (N_6436,N_6381,N_6271);
and U6437 (N_6437,N_6315,N_6356);
xor U6438 (N_6438,N_6232,N_6255);
nand U6439 (N_6439,N_6201,N_6289);
and U6440 (N_6440,N_6351,N_6221);
or U6441 (N_6441,N_6240,N_6355);
nor U6442 (N_6442,N_6284,N_6366);
nand U6443 (N_6443,N_6357,N_6376);
and U6444 (N_6444,N_6344,N_6317);
and U6445 (N_6445,N_6225,N_6330);
xor U6446 (N_6446,N_6335,N_6332);
nor U6447 (N_6447,N_6229,N_6375);
xnor U6448 (N_6448,N_6231,N_6285);
and U6449 (N_6449,N_6382,N_6329);
and U6450 (N_6450,N_6346,N_6368);
nand U6451 (N_6451,N_6250,N_6274);
nor U6452 (N_6452,N_6304,N_6321);
and U6453 (N_6453,N_6392,N_6374);
nand U6454 (N_6454,N_6397,N_6291);
nand U6455 (N_6455,N_6399,N_6269);
xnor U6456 (N_6456,N_6282,N_6302);
xnor U6457 (N_6457,N_6248,N_6280);
or U6458 (N_6458,N_6339,N_6309);
nand U6459 (N_6459,N_6237,N_6306);
or U6460 (N_6460,N_6352,N_6303);
xnor U6461 (N_6461,N_6387,N_6301);
nor U6462 (N_6462,N_6333,N_6249);
and U6463 (N_6463,N_6367,N_6320);
nand U6464 (N_6464,N_6360,N_6354);
xor U6465 (N_6465,N_6390,N_6369);
nand U6466 (N_6466,N_6264,N_6270);
or U6467 (N_6467,N_6261,N_6341);
xnor U6468 (N_6468,N_6391,N_6314);
xor U6469 (N_6469,N_6377,N_6318);
nand U6470 (N_6470,N_6219,N_6205);
and U6471 (N_6471,N_6218,N_6230);
xor U6472 (N_6472,N_6365,N_6273);
xor U6473 (N_6473,N_6337,N_6208);
or U6474 (N_6474,N_6223,N_6338);
xnor U6475 (N_6475,N_6281,N_6396);
nand U6476 (N_6476,N_6207,N_6378);
xor U6477 (N_6477,N_6312,N_6262);
nor U6478 (N_6478,N_6277,N_6252);
nor U6479 (N_6479,N_6211,N_6319);
and U6480 (N_6480,N_6222,N_6379);
or U6481 (N_6481,N_6292,N_6257);
or U6482 (N_6482,N_6373,N_6372);
nand U6483 (N_6483,N_6278,N_6394);
nand U6484 (N_6484,N_6228,N_6263);
xor U6485 (N_6485,N_6347,N_6243);
nor U6486 (N_6486,N_6293,N_6398);
xnor U6487 (N_6487,N_6203,N_6210);
or U6488 (N_6488,N_6259,N_6325);
or U6489 (N_6489,N_6389,N_6279);
and U6490 (N_6490,N_6224,N_6345);
nand U6491 (N_6491,N_6226,N_6370);
or U6492 (N_6492,N_6206,N_6359);
or U6493 (N_6493,N_6233,N_6217);
or U6494 (N_6494,N_6295,N_6343);
nand U6495 (N_6495,N_6386,N_6287);
and U6496 (N_6496,N_6253,N_6258);
and U6497 (N_6497,N_6276,N_6380);
nand U6498 (N_6498,N_6256,N_6272);
or U6499 (N_6499,N_6353,N_6246);
or U6500 (N_6500,N_6229,N_6265);
xor U6501 (N_6501,N_6384,N_6261);
nor U6502 (N_6502,N_6219,N_6216);
nor U6503 (N_6503,N_6372,N_6363);
xor U6504 (N_6504,N_6287,N_6384);
nand U6505 (N_6505,N_6233,N_6389);
nand U6506 (N_6506,N_6200,N_6276);
and U6507 (N_6507,N_6236,N_6303);
and U6508 (N_6508,N_6369,N_6205);
xor U6509 (N_6509,N_6326,N_6388);
nand U6510 (N_6510,N_6300,N_6359);
or U6511 (N_6511,N_6354,N_6205);
nand U6512 (N_6512,N_6384,N_6274);
or U6513 (N_6513,N_6293,N_6270);
nand U6514 (N_6514,N_6253,N_6251);
or U6515 (N_6515,N_6343,N_6377);
nor U6516 (N_6516,N_6390,N_6242);
and U6517 (N_6517,N_6273,N_6235);
or U6518 (N_6518,N_6308,N_6361);
xor U6519 (N_6519,N_6367,N_6387);
and U6520 (N_6520,N_6334,N_6241);
nor U6521 (N_6521,N_6339,N_6240);
or U6522 (N_6522,N_6301,N_6360);
xnor U6523 (N_6523,N_6336,N_6277);
or U6524 (N_6524,N_6256,N_6295);
or U6525 (N_6525,N_6256,N_6328);
nand U6526 (N_6526,N_6322,N_6217);
xor U6527 (N_6527,N_6362,N_6233);
and U6528 (N_6528,N_6274,N_6284);
or U6529 (N_6529,N_6296,N_6334);
and U6530 (N_6530,N_6345,N_6359);
xor U6531 (N_6531,N_6337,N_6330);
xnor U6532 (N_6532,N_6257,N_6321);
or U6533 (N_6533,N_6256,N_6289);
and U6534 (N_6534,N_6373,N_6379);
nor U6535 (N_6535,N_6256,N_6236);
or U6536 (N_6536,N_6284,N_6334);
nand U6537 (N_6537,N_6378,N_6383);
xor U6538 (N_6538,N_6304,N_6398);
nor U6539 (N_6539,N_6311,N_6209);
nand U6540 (N_6540,N_6201,N_6319);
and U6541 (N_6541,N_6230,N_6245);
xnor U6542 (N_6542,N_6394,N_6365);
nor U6543 (N_6543,N_6271,N_6292);
nand U6544 (N_6544,N_6267,N_6218);
or U6545 (N_6545,N_6285,N_6251);
and U6546 (N_6546,N_6351,N_6207);
xor U6547 (N_6547,N_6300,N_6247);
or U6548 (N_6548,N_6265,N_6242);
xor U6549 (N_6549,N_6293,N_6279);
nand U6550 (N_6550,N_6224,N_6353);
and U6551 (N_6551,N_6257,N_6212);
nor U6552 (N_6552,N_6272,N_6278);
nand U6553 (N_6553,N_6376,N_6323);
xnor U6554 (N_6554,N_6299,N_6335);
and U6555 (N_6555,N_6372,N_6399);
nor U6556 (N_6556,N_6283,N_6220);
and U6557 (N_6557,N_6383,N_6333);
xor U6558 (N_6558,N_6207,N_6297);
xnor U6559 (N_6559,N_6244,N_6390);
nand U6560 (N_6560,N_6293,N_6288);
nor U6561 (N_6561,N_6225,N_6208);
xnor U6562 (N_6562,N_6216,N_6243);
or U6563 (N_6563,N_6329,N_6248);
nand U6564 (N_6564,N_6290,N_6260);
nor U6565 (N_6565,N_6221,N_6217);
xor U6566 (N_6566,N_6226,N_6244);
nand U6567 (N_6567,N_6355,N_6319);
or U6568 (N_6568,N_6280,N_6288);
xnor U6569 (N_6569,N_6288,N_6393);
nand U6570 (N_6570,N_6298,N_6368);
nor U6571 (N_6571,N_6356,N_6384);
and U6572 (N_6572,N_6249,N_6235);
nor U6573 (N_6573,N_6388,N_6250);
xor U6574 (N_6574,N_6371,N_6343);
nand U6575 (N_6575,N_6322,N_6281);
nand U6576 (N_6576,N_6380,N_6232);
nand U6577 (N_6577,N_6205,N_6281);
nor U6578 (N_6578,N_6242,N_6321);
and U6579 (N_6579,N_6295,N_6342);
nor U6580 (N_6580,N_6202,N_6393);
nand U6581 (N_6581,N_6244,N_6212);
nand U6582 (N_6582,N_6216,N_6290);
and U6583 (N_6583,N_6323,N_6318);
nand U6584 (N_6584,N_6333,N_6300);
nor U6585 (N_6585,N_6353,N_6323);
nand U6586 (N_6586,N_6292,N_6212);
nand U6587 (N_6587,N_6318,N_6284);
or U6588 (N_6588,N_6297,N_6382);
nor U6589 (N_6589,N_6213,N_6265);
nor U6590 (N_6590,N_6278,N_6316);
or U6591 (N_6591,N_6357,N_6365);
or U6592 (N_6592,N_6229,N_6217);
or U6593 (N_6593,N_6327,N_6340);
and U6594 (N_6594,N_6269,N_6309);
xor U6595 (N_6595,N_6203,N_6231);
or U6596 (N_6596,N_6276,N_6398);
nand U6597 (N_6597,N_6357,N_6269);
nand U6598 (N_6598,N_6270,N_6316);
and U6599 (N_6599,N_6220,N_6247);
or U6600 (N_6600,N_6562,N_6529);
xnor U6601 (N_6601,N_6545,N_6412);
xor U6602 (N_6602,N_6410,N_6466);
nand U6603 (N_6603,N_6577,N_6530);
and U6604 (N_6604,N_6565,N_6514);
nand U6605 (N_6605,N_6421,N_6558);
and U6606 (N_6606,N_6438,N_6472);
nand U6607 (N_6607,N_6549,N_6454);
and U6608 (N_6608,N_6413,N_6433);
nand U6609 (N_6609,N_6507,N_6424);
or U6610 (N_6610,N_6597,N_6556);
or U6611 (N_6611,N_6574,N_6450);
xor U6612 (N_6612,N_6520,N_6489);
and U6613 (N_6613,N_6578,N_6500);
nand U6614 (N_6614,N_6407,N_6587);
nand U6615 (N_6615,N_6504,N_6596);
or U6616 (N_6616,N_6553,N_6510);
nand U6617 (N_6617,N_6502,N_6579);
nor U6618 (N_6618,N_6537,N_6468);
or U6619 (N_6619,N_6492,N_6534);
nand U6620 (N_6620,N_6586,N_6585);
xor U6621 (N_6621,N_6568,N_6431);
or U6622 (N_6622,N_6488,N_6503);
xnor U6623 (N_6623,N_6598,N_6533);
or U6624 (N_6624,N_6443,N_6516);
and U6625 (N_6625,N_6566,N_6559);
xnor U6626 (N_6626,N_6495,N_6547);
and U6627 (N_6627,N_6569,N_6582);
or U6628 (N_6628,N_6469,N_6449);
nand U6629 (N_6629,N_6402,N_6470);
nand U6630 (N_6630,N_6447,N_6526);
nor U6631 (N_6631,N_6480,N_6575);
and U6632 (N_6632,N_6511,N_6573);
nand U6633 (N_6633,N_6595,N_6452);
or U6634 (N_6634,N_6428,N_6440);
and U6635 (N_6635,N_6425,N_6459);
xor U6636 (N_6636,N_6599,N_6437);
nand U6637 (N_6637,N_6481,N_6567);
nor U6638 (N_6638,N_6409,N_6550);
or U6639 (N_6639,N_6554,N_6561);
nor U6640 (N_6640,N_6584,N_6485);
or U6641 (N_6641,N_6501,N_6535);
and U6642 (N_6642,N_6405,N_6475);
nand U6643 (N_6643,N_6416,N_6461);
nand U6644 (N_6644,N_6460,N_6453);
nand U6645 (N_6645,N_6522,N_6486);
and U6646 (N_6646,N_6420,N_6555);
and U6647 (N_6647,N_6427,N_6414);
or U6648 (N_6648,N_6430,N_6429);
or U6649 (N_6649,N_6457,N_6563);
nor U6650 (N_6650,N_6544,N_6476);
or U6651 (N_6651,N_6487,N_6471);
or U6652 (N_6652,N_6557,N_6478);
nand U6653 (N_6653,N_6525,N_6581);
xor U6654 (N_6654,N_6531,N_6423);
or U6655 (N_6655,N_6551,N_6444);
nand U6656 (N_6656,N_6508,N_6515);
xnor U6657 (N_6657,N_6441,N_6426);
nand U6658 (N_6658,N_6446,N_6406);
xnor U6659 (N_6659,N_6509,N_6528);
or U6660 (N_6660,N_6415,N_6498);
nor U6661 (N_6661,N_6540,N_6473);
or U6662 (N_6662,N_6543,N_6465);
nor U6663 (N_6663,N_6512,N_6493);
and U6664 (N_6664,N_6455,N_6506);
or U6665 (N_6665,N_6588,N_6594);
xnor U6666 (N_6666,N_6411,N_6491);
nor U6667 (N_6667,N_6590,N_6524);
and U6668 (N_6668,N_6571,N_6583);
and U6669 (N_6669,N_6403,N_6464);
nand U6670 (N_6670,N_6467,N_6451);
xnor U6671 (N_6671,N_6456,N_6541);
or U6672 (N_6672,N_6560,N_6499);
and U6673 (N_6673,N_6548,N_6474);
nor U6674 (N_6674,N_6400,N_6497);
nor U6675 (N_6675,N_6436,N_6564);
or U6676 (N_6676,N_6479,N_6458);
nor U6677 (N_6677,N_6589,N_6576);
xnor U6678 (N_6678,N_6432,N_6490);
xor U6679 (N_6679,N_6419,N_6570);
xnor U6680 (N_6680,N_6483,N_6496);
nor U6681 (N_6681,N_6513,N_6445);
nand U6682 (N_6682,N_6401,N_6521);
xor U6683 (N_6683,N_6477,N_6552);
or U6684 (N_6684,N_6408,N_6448);
nand U6685 (N_6685,N_6404,N_6418);
nor U6686 (N_6686,N_6505,N_6494);
and U6687 (N_6687,N_6580,N_6484);
nor U6688 (N_6688,N_6442,N_6539);
and U6689 (N_6689,N_6546,N_6542);
and U6690 (N_6690,N_6482,N_6462);
xnor U6691 (N_6691,N_6536,N_6435);
and U6692 (N_6692,N_6591,N_6517);
nor U6693 (N_6693,N_6439,N_6417);
nand U6694 (N_6694,N_6434,N_6532);
xor U6695 (N_6695,N_6523,N_6572);
or U6696 (N_6696,N_6593,N_6519);
or U6697 (N_6697,N_6538,N_6527);
nand U6698 (N_6698,N_6592,N_6518);
xor U6699 (N_6699,N_6422,N_6463);
and U6700 (N_6700,N_6520,N_6523);
xor U6701 (N_6701,N_6443,N_6497);
nor U6702 (N_6702,N_6472,N_6593);
and U6703 (N_6703,N_6427,N_6588);
and U6704 (N_6704,N_6417,N_6481);
and U6705 (N_6705,N_6422,N_6559);
and U6706 (N_6706,N_6405,N_6420);
and U6707 (N_6707,N_6582,N_6463);
nor U6708 (N_6708,N_6550,N_6574);
or U6709 (N_6709,N_6452,N_6518);
and U6710 (N_6710,N_6447,N_6565);
xnor U6711 (N_6711,N_6480,N_6586);
or U6712 (N_6712,N_6451,N_6525);
nor U6713 (N_6713,N_6455,N_6544);
xor U6714 (N_6714,N_6416,N_6486);
nand U6715 (N_6715,N_6523,N_6415);
nand U6716 (N_6716,N_6442,N_6406);
and U6717 (N_6717,N_6553,N_6568);
or U6718 (N_6718,N_6566,N_6522);
or U6719 (N_6719,N_6487,N_6558);
nor U6720 (N_6720,N_6447,N_6489);
and U6721 (N_6721,N_6522,N_6532);
nand U6722 (N_6722,N_6445,N_6506);
nand U6723 (N_6723,N_6504,N_6525);
nor U6724 (N_6724,N_6598,N_6568);
nor U6725 (N_6725,N_6565,N_6585);
nand U6726 (N_6726,N_6556,N_6547);
or U6727 (N_6727,N_6541,N_6435);
and U6728 (N_6728,N_6431,N_6542);
or U6729 (N_6729,N_6404,N_6454);
and U6730 (N_6730,N_6438,N_6447);
or U6731 (N_6731,N_6449,N_6499);
or U6732 (N_6732,N_6585,N_6406);
nand U6733 (N_6733,N_6531,N_6410);
xor U6734 (N_6734,N_6447,N_6589);
and U6735 (N_6735,N_6515,N_6410);
xnor U6736 (N_6736,N_6518,N_6587);
nor U6737 (N_6737,N_6468,N_6541);
and U6738 (N_6738,N_6468,N_6415);
nor U6739 (N_6739,N_6406,N_6454);
nand U6740 (N_6740,N_6507,N_6557);
nor U6741 (N_6741,N_6450,N_6559);
xor U6742 (N_6742,N_6514,N_6483);
or U6743 (N_6743,N_6435,N_6543);
or U6744 (N_6744,N_6560,N_6496);
xor U6745 (N_6745,N_6499,N_6566);
nand U6746 (N_6746,N_6435,N_6482);
xnor U6747 (N_6747,N_6492,N_6400);
xor U6748 (N_6748,N_6413,N_6478);
or U6749 (N_6749,N_6405,N_6546);
nor U6750 (N_6750,N_6465,N_6471);
nand U6751 (N_6751,N_6491,N_6443);
nand U6752 (N_6752,N_6523,N_6552);
and U6753 (N_6753,N_6449,N_6432);
xor U6754 (N_6754,N_6486,N_6502);
nand U6755 (N_6755,N_6515,N_6531);
or U6756 (N_6756,N_6572,N_6431);
and U6757 (N_6757,N_6533,N_6514);
xnor U6758 (N_6758,N_6470,N_6485);
or U6759 (N_6759,N_6407,N_6495);
xor U6760 (N_6760,N_6530,N_6590);
nor U6761 (N_6761,N_6598,N_6432);
nor U6762 (N_6762,N_6429,N_6403);
and U6763 (N_6763,N_6422,N_6445);
nor U6764 (N_6764,N_6579,N_6550);
nand U6765 (N_6765,N_6599,N_6412);
nand U6766 (N_6766,N_6472,N_6483);
and U6767 (N_6767,N_6477,N_6587);
nand U6768 (N_6768,N_6443,N_6545);
nand U6769 (N_6769,N_6400,N_6475);
nand U6770 (N_6770,N_6516,N_6400);
or U6771 (N_6771,N_6556,N_6518);
nand U6772 (N_6772,N_6445,N_6508);
nor U6773 (N_6773,N_6586,N_6490);
xnor U6774 (N_6774,N_6500,N_6510);
xor U6775 (N_6775,N_6422,N_6400);
nand U6776 (N_6776,N_6466,N_6517);
xor U6777 (N_6777,N_6458,N_6469);
and U6778 (N_6778,N_6450,N_6540);
and U6779 (N_6779,N_6551,N_6534);
xor U6780 (N_6780,N_6494,N_6416);
nand U6781 (N_6781,N_6444,N_6540);
and U6782 (N_6782,N_6599,N_6494);
nor U6783 (N_6783,N_6515,N_6549);
nand U6784 (N_6784,N_6500,N_6481);
and U6785 (N_6785,N_6492,N_6587);
xnor U6786 (N_6786,N_6447,N_6555);
or U6787 (N_6787,N_6431,N_6476);
nor U6788 (N_6788,N_6468,N_6464);
or U6789 (N_6789,N_6582,N_6406);
xor U6790 (N_6790,N_6478,N_6544);
nor U6791 (N_6791,N_6505,N_6574);
nor U6792 (N_6792,N_6530,N_6491);
nand U6793 (N_6793,N_6513,N_6460);
and U6794 (N_6794,N_6528,N_6546);
or U6795 (N_6795,N_6579,N_6465);
nand U6796 (N_6796,N_6428,N_6574);
xor U6797 (N_6797,N_6508,N_6488);
or U6798 (N_6798,N_6485,N_6574);
nand U6799 (N_6799,N_6564,N_6402);
or U6800 (N_6800,N_6628,N_6759);
or U6801 (N_6801,N_6649,N_6720);
and U6802 (N_6802,N_6686,N_6749);
or U6803 (N_6803,N_6639,N_6673);
nand U6804 (N_6804,N_6735,N_6634);
and U6805 (N_6805,N_6638,N_6768);
nand U6806 (N_6806,N_6719,N_6695);
nor U6807 (N_6807,N_6678,N_6682);
and U6808 (N_6808,N_6739,N_6797);
nor U6809 (N_6809,N_6601,N_6758);
nand U6810 (N_6810,N_6710,N_6715);
and U6811 (N_6811,N_6640,N_6778);
or U6812 (N_6812,N_6665,N_6748);
xnor U6813 (N_6813,N_6613,N_6674);
and U6814 (N_6814,N_6734,N_6629);
nor U6815 (N_6815,N_6777,N_6775);
xor U6816 (N_6816,N_6684,N_6648);
and U6817 (N_6817,N_6706,N_6799);
or U6818 (N_6818,N_6736,N_6769);
xor U6819 (N_6819,N_6712,N_6658);
xor U6820 (N_6820,N_6750,N_6789);
xnor U6821 (N_6821,N_6667,N_6729);
nand U6822 (N_6822,N_6724,N_6785);
or U6823 (N_6823,N_6651,N_6701);
and U6824 (N_6824,N_6794,N_6611);
xor U6825 (N_6825,N_6631,N_6681);
nand U6826 (N_6826,N_6662,N_6783);
nor U6827 (N_6827,N_6765,N_6763);
and U6828 (N_6828,N_6721,N_6653);
or U6829 (N_6829,N_6669,N_6738);
or U6830 (N_6830,N_6615,N_6725);
or U6831 (N_6831,N_6766,N_6754);
nand U6832 (N_6832,N_6690,N_6700);
nor U6833 (N_6833,N_6643,N_6760);
and U6834 (N_6834,N_6703,N_6707);
xnor U6835 (N_6835,N_6625,N_6642);
xor U6836 (N_6836,N_6600,N_6745);
or U6837 (N_6837,N_6751,N_6767);
xnor U6838 (N_6838,N_6675,N_6795);
nand U6839 (N_6839,N_6752,N_6697);
and U6840 (N_6840,N_6798,N_6731);
or U6841 (N_6841,N_6683,N_6781);
nand U6842 (N_6842,N_6776,N_6713);
nor U6843 (N_6843,N_6657,N_6774);
and U6844 (N_6844,N_6680,N_6694);
or U6845 (N_6845,N_6660,N_6633);
or U6846 (N_6846,N_6627,N_6644);
nand U6847 (N_6847,N_6793,N_6619);
and U6848 (N_6848,N_6732,N_6626);
and U6849 (N_6849,N_6606,N_6666);
xor U6850 (N_6850,N_6698,N_6641);
nand U6851 (N_6851,N_6708,N_6632);
nand U6852 (N_6852,N_6645,N_6779);
or U6853 (N_6853,N_6647,N_6663);
xor U6854 (N_6854,N_6693,N_6671);
and U6855 (N_6855,N_6790,N_6630);
xnor U6856 (N_6856,N_6605,N_6722);
nand U6857 (N_6857,N_6635,N_6689);
nand U6858 (N_6858,N_6786,N_6782);
nor U6859 (N_6859,N_6677,N_6704);
nor U6860 (N_6860,N_6664,N_6614);
nand U6861 (N_6861,N_6646,N_6691);
or U6862 (N_6862,N_6753,N_6618);
nor U6863 (N_6863,N_6705,N_6650);
nor U6864 (N_6864,N_6668,N_6756);
nand U6865 (N_6865,N_6743,N_6636);
and U6866 (N_6866,N_6727,N_6616);
xor U6867 (N_6867,N_6757,N_6612);
or U6868 (N_6868,N_6796,N_6787);
xor U6869 (N_6869,N_6602,N_6659);
nor U6870 (N_6870,N_6737,N_6624);
or U6871 (N_6871,N_6755,N_6728);
nor U6872 (N_6872,N_6610,N_6733);
xor U6873 (N_6873,N_6717,N_6792);
nand U6874 (N_6874,N_6608,N_6770);
or U6875 (N_6875,N_6771,N_6672);
nand U6876 (N_6876,N_6676,N_6692);
or U6877 (N_6877,N_6711,N_6723);
xnor U6878 (N_6878,N_6740,N_6607);
nor U6879 (N_6879,N_6709,N_6655);
nand U6880 (N_6880,N_6742,N_6716);
nand U6881 (N_6881,N_6702,N_6714);
and U6882 (N_6882,N_6726,N_6747);
or U6883 (N_6883,N_6661,N_6654);
nand U6884 (N_6884,N_6617,N_6620);
and U6885 (N_6885,N_6780,N_6656);
or U6886 (N_6886,N_6784,N_6764);
nor U6887 (N_6887,N_6772,N_6718);
and U6888 (N_6888,N_6685,N_6744);
nor U6889 (N_6889,N_6621,N_6791);
or U6890 (N_6890,N_6670,N_6696);
xor U6891 (N_6891,N_6699,N_6679);
and U6892 (N_6892,N_6741,N_6688);
or U6893 (N_6893,N_6637,N_6761);
nor U6894 (N_6894,N_6730,N_6788);
nand U6895 (N_6895,N_6687,N_6746);
or U6896 (N_6896,N_6773,N_6623);
nand U6897 (N_6897,N_6622,N_6603);
xnor U6898 (N_6898,N_6652,N_6762);
and U6899 (N_6899,N_6604,N_6609);
or U6900 (N_6900,N_6666,N_6770);
nand U6901 (N_6901,N_6654,N_6783);
nand U6902 (N_6902,N_6634,N_6675);
nor U6903 (N_6903,N_6679,N_6644);
xnor U6904 (N_6904,N_6617,N_6797);
or U6905 (N_6905,N_6665,N_6749);
and U6906 (N_6906,N_6782,N_6617);
and U6907 (N_6907,N_6649,N_6776);
or U6908 (N_6908,N_6656,N_6637);
nor U6909 (N_6909,N_6799,N_6629);
and U6910 (N_6910,N_6747,N_6794);
xnor U6911 (N_6911,N_6784,N_6704);
or U6912 (N_6912,N_6750,N_6683);
or U6913 (N_6913,N_6636,N_6768);
nor U6914 (N_6914,N_6721,N_6793);
xnor U6915 (N_6915,N_6619,N_6625);
or U6916 (N_6916,N_6654,N_6704);
and U6917 (N_6917,N_6733,N_6681);
nor U6918 (N_6918,N_6757,N_6689);
nand U6919 (N_6919,N_6650,N_6788);
xor U6920 (N_6920,N_6705,N_6714);
nand U6921 (N_6921,N_6694,N_6792);
and U6922 (N_6922,N_6634,N_6775);
nor U6923 (N_6923,N_6694,N_6726);
or U6924 (N_6924,N_6667,N_6785);
xnor U6925 (N_6925,N_6722,N_6699);
nor U6926 (N_6926,N_6774,N_6658);
or U6927 (N_6927,N_6759,N_6701);
or U6928 (N_6928,N_6694,N_6685);
nor U6929 (N_6929,N_6687,N_6714);
nor U6930 (N_6930,N_6646,N_6600);
or U6931 (N_6931,N_6772,N_6770);
and U6932 (N_6932,N_6637,N_6790);
nor U6933 (N_6933,N_6706,N_6673);
or U6934 (N_6934,N_6704,N_6630);
nand U6935 (N_6935,N_6753,N_6738);
and U6936 (N_6936,N_6727,N_6632);
nand U6937 (N_6937,N_6769,N_6686);
and U6938 (N_6938,N_6755,N_6715);
nor U6939 (N_6939,N_6678,N_6749);
nand U6940 (N_6940,N_6681,N_6652);
xnor U6941 (N_6941,N_6642,N_6646);
nor U6942 (N_6942,N_6647,N_6798);
xor U6943 (N_6943,N_6698,N_6717);
xnor U6944 (N_6944,N_6772,N_6683);
or U6945 (N_6945,N_6731,N_6782);
and U6946 (N_6946,N_6735,N_6729);
xor U6947 (N_6947,N_6696,N_6758);
or U6948 (N_6948,N_6718,N_6640);
or U6949 (N_6949,N_6726,N_6646);
nor U6950 (N_6950,N_6788,N_6756);
xnor U6951 (N_6951,N_6746,N_6626);
nand U6952 (N_6952,N_6796,N_6626);
nor U6953 (N_6953,N_6784,N_6695);
nor U6954 (N_6954,N_6753,N_6607);
or U6955 (N_6955,N_6600,N_6779);
and U6956 (N_6956,N_6757,N_6702);
or U6957 (N_6957,N_6628,N_6652);
xor U6958 (N_6958,N_6644,N_6657);
nor U6959 (N_6959,N_6752,N_6793);
nor U6960 (N_6960,N_6726,N_6703);
nand U6961 (N_6961,N_6710,N_6777);
or U6962 (N_6962,N_6678,N_6675);
nor U6963 (N_6963,N_6673,N_6663);
and U6964 (N_6964,N_6778,N_6656);
xnor U6965 (N_6965,N_6717,N_6790);
nor U6966 (N_6966,N_6751,N_6681);
nand U6967 (N_6967,N_6772,N_6676);
xnor U6968 (N_6968,N_6797,N_6785);
xor U6969 (N_6969,N_6726,N_6769);
xnor U6970 (N_6970,N_6791,N_6737);
xnor U6971 (N_6971,N_6692,N_6725);
and U6972 (N_6972,N_6674,N_6738);
nor U6973 (N_6973,N_6708,N_6710);
xnor U6974 (N_6974,N_6763,N_6691);
nand U6975 (N_6975,N_6787,N_6680);
xor U6976 (N_6976,N_6700,N_6725);
nand U6977 (N_6977,N_6659,N_6791);
and U6978 (N_6978,N_6729,N_6675);
nor U6979 (N_6979,N_6781,N_6642);
xnor U6980 (N_6980,N_6799,N_6633);
xor U6981 (N_6981,N_6757,N_6782);
nand U6982 (N_6982,N_6797,N_6723);
xnor U6983 (N_6983,N_6705,N_6751);
nor U6984 (N_6984,N_6687,N_6691);
nand U6985 (N_6985,N_6673,N_6722);
nor U6986 (N_6986,N_6689,N_6653);
xor U6987 (N_6987,N_6680,N_6682);
or U6988 (N_6988,N_6701,N_6735);
xor U6989 (N_6989,N_6755,N_6717);
or U6990 (N_6990,N_6680,N_6695);
nor U6991 (N_6991,N_6763,N_6644);
and U6992 (N_6992,N_6735,N_6660);
or U6993 (N_6993,N_6733,N_6775);
or U6994 (N_6994,N_6682,N_6748);
nor U6995 (N_6995,N_6778,N_6722);
or U6996 (N_6996,N_6687,N_6661);
and U6997 (N_6997,N_6691,N_6726);
nor U6998 (N_6998,N_6656,N_6737);
or U6999 (N_6999,N_6792,N_6620);
nor U7000 (N_7000,N_6816,N_6850);
nor U7001 (N_7001,N_6933,N_6851);
and U7002 (N_7002,N_6891,N_6838);
nand U7003 (N_7003,N_6990,N_6902);
and U7004 (N_7004,N_6818,N_6839);
xor U7005 (N_7005,N_6925,N_6807);
xnor U7006 (N_7006,N_6871,N_6883);
nand U7007 (N_7007,N_6932,N_6840);
nand U7008 (N_7008,N_6824,N_6834);
and U7009 (N_7009,N_6887,N_6975);
and U7010 (N_7010,N_6884,N_6994);
xor U7011 (N_7011,N_6971,N_6913);
xor U7012 (N_7012,N_6998,N_6835);
nand U7013 (N_7013,N_6890,N_6814);
and U7014 (N_7014,N_6825,N_6879);
nor U7015 (N_7015,N_6908,N_6801);
xor U7016 (N_7016,N_6889,N_6940);
xnor U7017 (N_7017,N_6864,N_6921);
and U7018 (N_7018,N_6941,N_6869);
xor U7019 (N_7019,N_6985,N_6922);
and U7020 (N_7020,N_6979,N_6907);
nor U7021 (N_7021,N_6809,N_6837);
or U7022 (N_7022,N_6924,N_6962);
nand U7023 (N_7023,N_6946,N_6942);
nand U7024 (N_7024,N_6833,N_6819);
or U7025 (N_7025,N_6955,N_6939);
and U7026 (N_7026,N_6906,N_6828);
and U7027 (N_7027,N_6927,N_6862);
or U7028 (N_7028,N_6805,N_6956);
and U7029 (N_7029,N_6877,N_6888);
xnor U7030 (N_7030,N_6856,N_6944);
nand U7031 (N_7031,N_6912,N_6993);
nor U7032 (N_7032,N_6812,N_6846);
or U7033 (N_7033,N_6895,N_6968);
xor U7034 (N_7034,N_6992,N_6964);
xnor U7035 (N_7035,N_6920,N_6988);
nor U7036 (N_7036,N_6986,N_6995);
and U7037 (N_7037,N_6896,N_6826);
or U7038 (N_7038,N_6870,N_6899);
xor U7039 (N_7039,N_6863,N_6917);
nor U7040 (N_7040,N_6965,N_6934);
nand U7041 (N_7041,N_6860,N_6916);
and U7042 (N_7042,N_6849,N_6966);
nand U7043 (N_7043,N_6969,N_6943);
or U7044 (N_7044,N_6919,N_6903);
nor U7045 (N_7045,N_6892,N_6960);
xnor U7046 (N_7046,N_6858,N_6853);
nand U7047 (N_7047,N_6949,N_6886);
or U7048 (N_7048,N_6854,N_6802);
xnor U7049 (N_7049,N_6842,N_6859);
xnor U7050 (N_7050,N_6970,N_6904);
and U7051 (N_7051,N_6928,N_6800);
xnor U7052 (N_7052,N_6874,N_6999);
nor U7053 (N_7053,N_6929,N_6841);
xor U7054 (N_7054,N_6836,N_6882);
or U7055 (N_7055,N_6978,N_6981);
xor U7056 (N_7056,N_6950,N_6931);
or U7057 (N_7057,N_6893,N_6865);
and U7058 (N_7058,N_6963,N_6918);
nor U7059 (N_7059,N_6937,N_6980);
or U7060 (N_7060,N_6900,N_6845);
or U7061 (N_7061,N_6972,N_6953);
nor U7062 (N_7062,N_6905,N_6976);
nand U7063 (N_7063,N_6806,N_6973);
nand U7064 (N_7064,N_6901,N_6831);
xnor U7065 (N_7065,N_6848,N_6868);
nor U7066 (N_7066,N_6914,N_6804);
or U7067 (N_7067,N_6873,N_6910);
nor U7068 (N_7068,N_6857,N_6945);
nand U7069 (N_7069,N_6817,N_6977);
nand U7070 (N_7070,N_6983,N_6987);
or U7071 (N_7071,N_6867,N_6866);
or U7072 (N_7072,N_6815,N_6954);
or U7073 (N_7073,N_6989,N_6951);
and U7074 (N_7074,N_6894,N_6881);
nand U7075 (N_7075,N_6855,N_6820);
xnor U7076 (N_7076,N_6911,N_6961);
nand U7077 (N_7077,N_6843,N_6880);
nand U7078 (N_7078,N_6982,N_6959);
and U7079 (N_7079,N_6847,N_6827);
xnor U7080 (N_7080,N_6810,N_6861);
nand U7081 (N_7081,N_6991,N_6967);
nand U7082 (N_7082,N_6947,N_6876);
nand U7083 (N_7083,N_6821,N_6878);
and U7084 (N_7084,N_6938,N_6829);
nand U7085 (N_7085,N_6952,N_6974);
xor U7086 (N_7086,N_6948,N_6926);
or U7087 (N_7087,N_6997,N_6885);
or U7088 (N_7088,N_6958,N_6935);
and U7089 (N_7089,N_6803,N_6875);
nand U7090 (N_7090,N_6823,N_6909);
nor U7091 (N_7091,N_6844,N_6822);
and U7092 (N_7092,N_6936,N_6830);
nand U7093 (N_7093,N_6915,N_6808);
or U7094 (N_7094,N_6813,N_6957);
or U7095 (N_7095,N_6898,N_6832);
and U7096 (N_7096,N_6897,N_6996);
and U7097 (N_7097,N_6872,N_6930);
nand U7098 (N_7098,N_6984,N_6923);
and U7099 (N_7099,N_6811,N_6852);
and U7100 (N_7100,N_6821,N_6924);
and U7101 (N_7101,N_6883,N_6879);
or U7102 (N_7102,N_6910,N_6884);
nor U7103 (N_7103,N_6922,N_6828);
nand U7104 (N_7104,N_6812,N_6860);
nor U7105 (N_7105,N_6830,N_6952);
nand U7106 (N_7106,N_6932,N_6894);
xor U7107 (N_7107,N_6886,N_6852);
nor U7108 (N_7108,N_6997,N_6846);
xor U7109 (N_7109,N_6801,N_6970);
nor U7110 (N_7110,N_6802,N_6920);
nor U7111 (N_7111,N_6825,N_6919);
xnor U7112 (N_7112,N_6904,N_6906);
and U7113 (N_7113,N_6800,N_6925);
and U7114 (N_7114,N_6872,N_6833);
xnor U7115 (N_7115,N_6956,N_6977);
or U7116 (N_7116,N_6915,N_6899);
and U7117 (N_7117,N_6892,N_6832);
nand U7118 (N_7118,N_6949,N_6928);
xor U7119 (N_7119,N_6980,N_6984);
nor U7120 (N_7120,N_6861,N_6869);
or U7121 (N_7121,N_6891,N_6845);
and U7122 (N_7122,N_6968,N_6943);
and U7123 (N_7123,N_6815,N_6989);
or U7124 (N_7124,N_6977,N_6852);
xor U7125 (N_7125,N_6895,N_6936);
nor U7126 (N_7126,N_6819,N_6867);
and U7127 (N_7127,N_6943,N_6810);
nand U7128 (N_7128,N_6868,N_6896);
and U7129 (N_7129,N_6962,N_6853);
and U7130 (N_7130,N_6955,N_6922);
or U7131 (N_7131,N_6922,N_6813);
xor U7132 (N_7132,N_6959,N_6881);
xnor U7133 (N_7133,N_6877,N_6833);
xor U7134 (N_7134,N_6873,N_6997);
or U7135 (N_7135,N_6953,N_6898);
or U7136 (N_7136,N_6814,N_6948);
nand U7137 (N_7137,N_6952,N_6948);
and U7138 (N_7138,N_6923,N_6901);
xor U7139 (N_7139,N_6853,N_6882);
xnor U7140 (N_7140,N_6869,N_6865);
nor U7141 (N_7141,N_6913,N_6938);
xor U7142 (N_7142,N_6964,N_6949);
or U7143 (N_7143,N_6939,N_6822);
and U7144 (N_7144,N_6990,N_6825);
xor U7145 (N_7145,N_6897,N_6995);
nand U7146 (N_7146,N_6921,N_6805);
nor U7147 (N_7147,N_6914,N_6956);
nand U7148 (N_7148,N_6823,N_6885);
and U7149 (N_7149,N_6981,N_6996);
xor U7150 (N_7150,N_6916,N_6971);
nor U7151 (N_7151,N_6920,N_6889);
and U7152 (N_7152,N_6887,N_6819);
and U7153 (N_7153,N_6943,N_6961);
nand U7154 (N_7154,N_6855,N_6879);
and U7155 (N_7155,N_6947,N_6837);
nor U7156 (N_7156,N_6889,N_6868);
and U7157 (N_7157,N_6821,N_6915);
and U7158 (N_7158,N_6839,N_6985);
or U7159 (N_7159,N_6842,N_6935);
or U7160 (N_7160,N_6857,N_6940);
or U7161 (N_7161,N_6810,N_6996);
xor U7162 (N_7162,N_6835,N_6906);
or U7163 (N_7163,N_6986,N_6907);
or U7164 (N_7164,N_6975,N_6806);
nand U7165 (N_7165,N_6903,N_6830);
and U7166 (N_7166,N_6962,N_6915);
or U7167 (N_7167,N_6806,N_6947);
nor U7168 (N_7168,N_6903,N_6822);
nand U7169 (N_7169,N_6806,N_6846);
xnor U7170 (N_7170,N_6800,N_6843);
xnor U7171 (N_7171,N_6911,N_6892);
or U7172 (N_7172,N_6971,N_6890);
and U7173 (N_7173,N_6924,N_6872);
or U7174 (N_7174,N_6899,N_6815);
and U7175 (N_7175,N_6983,N_6992);
nand U7176 (N_7176,N_6816,N_6971);
nor U7177 (N_7177,N_6894,N_6907);
nor U7178 (N_7178,N_6876,N_6944);
and U7179 (N_7179,N_6804,N_6827);
or U7180 (N_7180,N_6836,N_6927);
or U7181 (N_7181,N_6815,N_6980);
and U7182 (N_7182,N_6824,N_6830);
or U7183 (N_7183,N_6814,N_6952);
nor U7184 (N_7184,N_6815,N_6883);
or U7185 (N_7185,N_6926,N_6876);
and U7186 (N_7186,N_6976,N_6819);
and U7187 (N_7187,N_6881,N_6990);
or U7188 (N_7188,N_6918,N_6938);
nand U7189 (N_7189,N_6925,N_6839);
nand U7190 (N_7190,N_6860,N_6876);
nand U7191 (N_7191,N_6931,N_6844);
nand U7192 (N_7192,N_6892,N_6864);
and U7193 (N_7193,N_6973,N_6921);
nand U7194 (N_7194,N_6816,N_6861);
nor U7195 (N_7195,N_6873,N_6875);
or U7196 (N_7196,N_6964,N_6810);
xor U7197 (N_7197,N_6827,N_6818);
or U7198 (N_7198,N_6944,N_6847);
xor U7199 (N_7199,N_6862,N_6986);
or U7200 (N_7200,N_7003,N_7167);
nand U7201 (N_7201,N_7115,N_7016);
xnor U7202 (N_7202,N_7032,N_7017);
or U7203 (N_7203,N_7096,N_7030);
xnor U7204 (N_7204,N_7057,N_7182);
or U7205 (N_7205,N_7143,N_7036);
and U7206 (N_7206,N_7004,N_7107);
nor U7207 (N_7207,N_7061,N_7008);
nor U7208 (N_7208,N_7007,N_7130);
and U7209 (N_7209,N_7116,N_7195);
nand U7210 (N_7210,N_7178,N_7060);
and U7211 (N_7211,N_7020,N_7153);
nor U7212 (N_7212,N_7009,N_7198);
xnor U7213 (N_7213,N_7071,N_7139);
and U7214 (N_7214,N_7014,N_7174);
nand U7215 (N_7215,N_7084,N_7199);
and U7216 (N_7216,N_7147,N_7100);
nand U7217 (N_7217,N_7154,N_7091);
nor U7218 (N_7218,N_7113,N_7186);
nor U7219 (N_7219,N_7138,N_7000);
or U7220 (N_7220,N_7152,N_7104);
and U7221 (N_7221,N_7140,N_7075);
nor U7222 (N_7222,N_7101,N_7041);
nor U7223 (N_7223,N_7034,N_7159);
xnor U7224 (N_7224,N_7103,N_7142);
and U7225 (N_7225,N_7169,N_7048);
xor U7226 (N_7226,N_7062,N_7114);
or U7227 (N_7227,N_7163,N_7108);
or U7228 (N_7228,N_7181,N_7087);
xor U7229 (N_7229,N_7073,N_7192);
xor U7230 (N_7230,N_7149,N_7145);
xnor U7231 (N_7231,N_7090,N_7128);
nand U7232 (N_7232,N_7109,N_7095);
nor U7233 (N_7233,N_7119,N_7111);
xnor U7234 (N_7234,N_7005,N_7082);
nor U7235 (N_7235,N_7053,N_7049);
xnor U7236 (N_7236,N_7045,N_7044);
nand U7237 (N_7237,N_7197,N_7161);
nand U7238 (N_7238,N_7028,N_7166);
xnor U7239 (N_7239,N_7141,N_7122);
xor U7240 (N_7240,N_7136,N_7183);
or U7241 (N_7241,N_7176,N_7013);
nor U7242 (N_7242,N_7012,N_7173);
xor U7243 (N_7243,N_7031,N_7092);
nor U7244 (N_7244,N_7157,N_7121);
or U7245 (N_7245,N_7064,N_7156);
nand U7246 (N_7246,N_7051,N_7043);
nand U7247 (N_7247,N_7112,N_7085);
xor U7248 (N_7248,N_7164,N_7158);
nand U7249 (N_7249,N_7067,N_7069);
or U7250 (N_7250,N_7162,N_7194);
xnor U7251 (N_7251,N_7189,N_7102);
or U7252 (N_7252,N_7076,N_7187);
nand U7253 (N_7253,N_7065,N_7039);
nor U7254 (N_7254,N_7191,N_7177);
and U7255 (N_7255,N_7037,N_7124);
xnor U7256 (N_7256,N_7099,N_7021);
nor U7257 (N_7257,N_7019,N_7106);
nor U7258 (N_7258,N_7135,N_7160);
xnor U7259 (N_7259,N_7047,N_7088);
nor U7260 (N_7260,N_7083,N_7132);
or U7261 (N_7261,N_7080,N_7172);
and U7262 (N_7262,N_7006,N_7059);
or U7263 (N_7263,N_7137,N_7151);
nand U7264 (N_7264,N_7131,N_7110);
or U7265 (N_7265,N_7105,N_7074);
nor U7266 (N_7266,N_7052,N_7118);
nor U7267 (N_7267,N_7190,N_7068);
or U7268 (N_7268,N_7185,N_7077);
nand U7269 (N_7269,N_7148,N_7144);
nand U7270 (N_7270,N_7025,N_7035);
nor U7271 (N_7271,N_7015,N_7072);
nor U7272 (N_7272,N_7127,N_7120);
and U7273 (N_7273,N_7155,N_7040);
or U7274 (N_7274,N_7126,N_7170);
xnor U7275 (N_7275,N_7196,N_7010);
or U7276 (N_7276,N_7134,N_7002);
nor U7277 (N_7277,N_7018,N_7058);
nand U7278 (N_7278,N_7146,N_7171);
or U7279 (N_7279,N_7024,N_7180);
and U7280 (N_7280,N_7094,N_7078);
and U7281 (N_7281,N_7168,N_7117);
xor U7282 (N_7282,N_7029,N_7054);
or U7283 (N_7283,N_7093,N_7188);
nand U7284 (N_7284,N_7097,N_7086);
or U7285 (N_7285,N_7179,N_7098);
nor U7286 (N_7286,N_7022,N_7023);
and U7287 (N_7287,N_7027,N_7175);
and U7288 (N_7288,N_7001,N_7123);
xnor U7289 (N_7289,N_7066,N_7184);
nand U7290 (N_7290,N_7150,N_7063);
xor U7291 (N_7291,N_7133,N_7046);
and U7292 (N_7292,N_7125,N_7081);
and U7293 (N_7293,N_7042,N_7011);
nand U7294 (N_7294,N_7055,N_7129);
nand U7295 (N_7295,N_7056,N_7050);
xnor U7296 (N_7296,N_7033,N_7079);
nor U7297 (N_7297,N_7089,N_7193);
and U7298 (N_7298,N_7038,N_7165);
nor U7299 (N_7299,N_7070,N_7026);
nor U7300 (N_7300,N_7088,N_7077);
or U7301 (N_7301,N_7154,N_7055);
nand U7302 (N_7302,N_7008,N_7066);
nand U7303 (N_7303,N_7153,N_7059);
or U7304 (N_7304,N_7011,N_7130);
nand U7305 (N_7305,N_7174,N_7034);
nand U7306 (N_7306,N_7032,N_7054);
and U7307 (N_7307,N_7142,N_7040);
nor U7308 (N_7308,N_7154,N_7059);
or U7309 (N_7309,N_7052,N_7093);
xnor U7310 (N_7310,N_7054,N_7140);
or U7311 (N_7311,N_7147,N_7043);
nand U7312 (N_7312,N_7099,N_7095);
nor U7313 (N_7313,N_7001,N_7117);
and U7314 (N_7314,N_7002,N_7070);
xnor U7315 (N_7315,N_7027,N_7120);
xnor U7316 (N_7316,N_7163,N_7014);
nor U7317 (N_7317,N_7167,N_7114);
and U7318 (N_7318,N_7024,N_7171);
nand U7319 (N_7319,N_7146,N_7037);
nor U7320 (N_7320,N_7105,N_7146);
nor U7321 (N_7321,N_7171,N_7121);
nand U7322 (N_7322,N_7123,N_7116);
nand U7323 (N_7323,N_7059,N_7199);
nor U7324 (N_7324,N_7147,N_7159);
xnor U7325 (N_7325,N_7124,N_7054);
or U7326 (N_7326,N_7122,N_7010);
nand U7327 (N_7327,N_7023,N_7139);
xnor U7328 (N_7328,N_7015,N_7001);
and U7329 (N_7329,N_7183,N_7038);
nand U7330 (N_7330,N_7157,N_7068);
xor U7331 (N_7331,N_7066,N_7166);
nor U7332 (N_7332,N_7163,N_7077);
and U7333 (N_7333,N_7094,N_7059);
xnor U7334 (N_7334,N_7167,N_7143);
nor U7335 (N_7335,N_7044,N_7056);
and U7336 (N_7336,N_7047,N_7124);
xnor U7337 (N_7337,N_7006,N_7091);
and U7338 (N_7338,N_7075,N_7013);
nor U7339 (N_7339,N_7192,N_7176);
xnor U7340 (N_7340,N_7023,N_7077);
xnor U7341 (N_7341,N_7014,N_7122);
nor U7342 (N_7342,N_7136,N_7055);
xor U7343 (N_7343,N_7084,N_7153);
or U7344 (N_7344,N_7176,N_7046);
and U7345 (N_7345,N_7055,N_7191);
nand U7346 (N_7346,N_7185,N_7113);
and U7347 (N_7347,N_7060,N_7029);
xnor U7348 (N_7348,N_7017,N_7101);
or U7349 (N_7349,N_7036,N_7170);
xor U7350 (N_7350,N_7030,N_7098);
nor U7351 (N_7351,N_7008,N_7036);
or U7352 (N_7352,N_7091,N_7054);
or U7353 (N_7353,N_7046,N_7051);
and U7354 (N_7354,N_7197,N_7086);
nand U7355 (N_7355,N_7194,N_7005);
nor U7356 (N_7356,N_7038,N_7167);
xor U7357 (N_7357,N_7044,N_7153);
nand U7358 (N_7358,N_7063,N_7192);
or U7359 (N_7359,N_7173,N_7149);
and U7360 (N_7360,N_7197,N_7181);
and U7361 (N_7361,N_7034,N_7006);
or U7362 (N_7362,N_7192,N_7188);
xnor U7363 (N_7363,N_7035,N_7168);
or U7364 (N_7364,N_7136,N_7009);
xor U7365 (N_7365,N_7132,N_7157);
xnor U7366 (N_7366,N_7067,N_7171);
and U7367 (N_7367,N_7007,N_7124);
or U7368 (N_7368,N_7054,N_7058);
nor U7369 (N_7369,N_7199,N_7189);
and U7370 (N_7370,N_7146,N_7175);
nor U7371 (N_7371,N_7068,N_7121);
nand U7372 (N_7372,N_7193,N_7018);
nand U7373 (N_7373,N_7185,N_7118);
or U7374 (N_7374,N_7059,N_7026);
and U7375 (N_7375,N_7035,N_7133);
nor U7376 (N_7376,N_7093,N_7156);
nor U7377 (N_7377,N_7198,N_7055);
and U7378 (N_7378,N_7091,N_7195);
nand U7379 (N_7379,N_7172,N_7104);
and U7380 (N_7380,N_7017,N_7001);
and U7381 (N_7381,N_7129,N_7043);
nor U7382 (N_7382,N_7107,N_7059);
nand U7383 (N_7383,N_7001,N_7069);
or U7384 (N_7384,N_7108,N_7195);
or U7385 (N_7385,N_7178,N_7196);
xor U7386 (N_7386,N_7070,N_7141);
and U7387 (N_7387,N_7032,N_7088);
and U7388 (N_7388,N_7145,N_7182);
or U7389 (N_7389,N_7102,N_7003);
xnor U7390 (N_7390,N_7165,N_7087);
nand U7391 (N_7391,N_7184,N_7021);
and U7392 (N_7392,N_7150,N_7061);
or U7393 (N_7393,N_7164,N_7028);
or U7394 (N_7394,N_7037,N_7084);
xor U7395 (N_7395,N_7174,N_7161);
and U7396 (N_7396,N_7145,N_7043);
nand U7397 (N_7397,N_7031,N_7076);
and U7398 (N_7398,N_7125,N_7123);
nor U7399 (N_7399,N_7189,N_7051);
nand U7400 (N_7400,N_7299,N_7387);
or U7401 (N_7401,N_7379,N_7392);
nor U7402 (N_7402,N_7332,N_7258);
and U7403 (N_7403,N_7345,N_7333);
nand U7404 (N_7404,N_7224,N_7334);
xnor U7405 (N_7405,N_7384,N_7239);
or U7406 (N_7406,N_7352,N_7274);
nand U7407 (N_7407,N_7363,N_7243);
nor U7408 (N_7408,N_7336,N_7322);
and U7409 (N_7409,N_7233,N_7253);
and U7410 (N_7410,N_7223,N_7323);
or U7411 (N_7411,N_7225,N_7365);
nor U7412 (N_7412,N_7217,N_7339);
and U7413 (N_7413,N_7201,N_7205);
xnor U7414 (N_7414,N_7285,N_7316);
or U7415 (N_7415,N_7207,N_7354);
nand U7416 (N_7416,N_7222,N_7342);
or U7417 (N_7417,N_7293,N_7314);
xor U7418 (N_7418,N_7238,N_7399);
and U7419 (N_7419,N_7355,N_7208);
nor U7420 (N_7420,N_7278,N_7369);
nand U7421 (N_7421,N_7247,N_7301);
or U7422 (N_7422,N_7300,N_7226);
and U7423 (N_7423,N_7346,N_7357);
and U7424 (N_7424,N_7388,N_7232);
nand U7425 (N_7425,N_7275,N_7305);
nor U7426 (N_7426,N_7270,N_7240);
and U7427 (N_7427,N_7348,N_7335);
nand U7428 (N_7428,N_7267,N_7328);
and U7429 (N_7429,N_7290,N_7244);
and U7430 (N_7430,N_7234,N_7338);
or U7431 (N_7431,N_7343,N_7206);
nand U7432 (N_7432,N_7287,N_7250);
or U7433 (N_7433,N_7254,N_7341);
xor U7434 (N_7434,N_7337,N_7381);
or U7435 (N_7435,N_7200,N_7321);
or U7436 (N_7436,N_7209,N_7308);
and U7437 (N_7437,N_7212,N_7313);
nand U7438 (N_7438,N_7358,N_7350);
or U7439 (N_7439,N_7307,N_7260);
or U7440 (N_7440,N_7303,N_7276);
and U7441 (N_7441,N_7283,N_7359);
nand U7442 (N_7442,N_7386,N_7261);
nand U7443 (N_7443,N_7340,N_7370);
or U7444 (N_7444,N_7320,N_7311);
nand U7445 (N_7445,N_7203,N_7221);
nand U7446 (N_7446,N_7236,N_7282);
or U7447 (N_7447,N_7309,N_7259);
and U7448 (N_7448,N_7296,N_7216);
nand U7449 (N_7449,N_7326,N_7324);
and U7450 (N_7450,N_7297,N_7389);
nand U7451 (N_7451,N_7237,N_7218);
xnor U7452 (N_7452,N_7376,N_7264);
and U7453 (N_7453,N_7393,N_7268);
xor U7454 (N_7454,N_7391,N_7317);
xor U7455 (N_7455,N_7364,N_7255);
nor U7456 (N_7456,N_7310,N_7347);
nor U7457 (N_7457,N_7271,N_7366);
and U7458 (N_7458,N_7227,N_7331);
or U7459 (N_7459,N_7245,N_7390);
nor U7460 (N_7460,N_7213,N_7349);
and U7461 (N_7461,N_7269,N_7279);
nor U7462 (N_7462,N_7288,N_7263);
xnor U7463 (N_7463,N_7395,N_7362);
nand U7464 (N_7464,N_7302,N_7280);
or U7465 (N_7465,N_7266,N_7292);
xor U7466 (N_7466,N_7249,N_7214);
and U7467 (N_7467,N_7398,N_7229);
nand U7468 (N_7468,N_7215,N_7219);
nor U7469 (N_7469,N_7246,N_7318);
and U7470 (N_7470,N_7375,N_7372);
or U7471 (N_7471,N_7256,N_7294);
nor U7472 (N_7472,N_7380,N_7360);
xnor U7473 (N_7473,N_7277,N_7368);
or U7474 (N_7474,N_7248,N_7231);
and U7475 (N_7475,N_7272,N_7394);
or U7476 (N_7476,N_7327,N_7211);
or U7477 (N_7477,N_7329,N_7353);
nor U7478 (N_7478,N_7251,N_7344);
nand U7479 (N_7479,N_7306,N_7235);
nor U7480 (N_7480,N_7289,N_7374);
or U7481 (N_7481,N_7242,N_7319);
xor U7482 (N_7482,N_7356,N_7312);
and U7483 (N_7483,N_7351,N_7202);
or U7484 (N_7484,N_7220,N_7367);
and U7485 (N_7485,N_7265,N_7396);
xnor U7486 (N_7486,N_7204,N_7252);
nor U7487 (N_7487,N_7284,N_7377);
nor U7488 (N_7488,N_7373,N_7385);
and U7489 (N_7489,N_7286,N_7382);
xor U7490 (N_7490,N_7257,N_7315);
nand U7491 (N_7491,N_7291,N_7330);
xnor U7492 (N_7492,N_7273,N_7304);
nand U7493 (N_7493,N_7298,N_7325);
nand U7494 (N_7494,N_7241,N_7281);
or U7495 (N_7495,N_7361,N_7378);
or U7496 (N_7496,N_7397,N_7383);
nor U7497 (N_7497,N_7210,N_7371);
nor U7498 (N_7498,N_7262,N_7295);
xor U7499 (N_7499,N_7228,N_7230);
or U7500 (N_7500,N_7350,N_7220);
nand U7501 (N_7501,N_7333,N_7337);
nand U7502 (N_7502,N_7288,N_7304);
xor U7503 (N_7503,N_7240,N_7387);
nor U7504 (N_7504,N_7232,N_7306);
nor U7505 (N_7505,N_7363,N_7216);
and U7506 (N_7506,N_7232,N_7272);
nor U7507 (N_7507,N_7273,N_7375);
nand U7508 (N_7508,N_7248,N_7255);
nand U7509 (N_7509,N_7206,N_7314);
nand U7510 (N_7510,N_7334,N_7317);
nand U7511 (N_7511,N_7211,N_7268);
xor U7512 (N_7512,N_7244,N_7275);
and U7513 (N_7513,N_7211,N_7233);
or U7514 (N_7514,N_7364,N_7311);
or U7515 (N_7515,N_7228,N_7236);
nor U7516 (N_7516,N_7295,N_7311);
nor U7517 (N_7517,N_7354,N_7316);
nand U7518 (N_7518,N_7319,N_7387);
nor U7519 (N_7519,N_7312,N_7309);
or U7520 (N_7520,N_7216,N_7327);
xor U7521 (N_7521,N_7208,N_7386);
xnor U7522 (N_7522,N_7354,N_7233);
nor U7523 (N_7523,N_7384,N_7396);
nor U7524 (N_7524,N_7230,N_7369);
nor U7525 (N_7525,N_7312,N_7201);
or U7526 (N_7526,N_7354,N_7281);
or U7527 (N_7527,N_7328,N_7398);
xnor U7528 (N_7528,N_7296,N_7336);
nand U7529 (N_7529,N_7332,N_7233);
xor U7530 (N_7530,N_7274,N_7238);
or U7531 (N_7531,N_7295,N_7308);
or U7532 (N_7532,N_7245,N_7366);
or U7533 (N_7533,N_7302,N_7355);
xor U7534 (N_7534,N_7332,N_7225);
nand U7535 (N_7535,N_7258,N_7351);
nand U7536 (N_7536,N_7328,N_7209);
nand U7537 (N_7537,N_7251,N_7261);
and U7538 (N_7538,N_7351,N_7233);
nand U7539 (N_7539,N_7260,N_7297);
and U7540 (N_7540,N_7321,N_7398);
and U7541 (N_7541,N_7306,N_7211);
or U7542 (N_7542,N_7206,N_7254);
nor U7543 (N_7543,N_7397,N_7365);
nand U7544 (N_7544,N_7221,N_7349);
nor U7545 (N_7545,N_7372,N_7242);
or U7546 (N_7546,N_7315,N_7381);
nand U7547 (N_7547,N_7247,N_7263);
and U7548 (N_7548,N_7213,N_7232);
or U7549 (N_7549,N_7221,N_7222);
nand U7550 (N_7550,N_7292,N_7348);
and U7551 (N_7551,N_7252,N_7372);
xnor U7552 (N_7552,N_7204,N_7335);
nor U7553 (N_7553,N_7214,N_7323);
xnor U7554 (N_7554,N_7360,N_7350);
nand U7555 (N_7555,N_7235,N_7293);
and U7556 (N_7556,N_7299,N_7392);
and U7557 (N_7557,N_7274,N_7215);
nor U7558 (N_7558,N_7241,N_7285);
and U7559 (N_7559,N_7268,N_7272);
nand U7560 (N_7560,N_7339,N_7301);
nand U7561 (N_7561,N_7390,N_7295);
nor U7562 (N_7562,N_7367,N_7340);
xor U7563 (N_7563,N_7343,N_7293);
xnor U7564 (N_7564,N_7256,N_7338);
xor U7565 (N_7565,N_7204,N_7269);
or U7566 (N_7566,N_7293,N_7275);
and U7567 (N_7567,N_7338,N_7345);
nand U7568 (N_7568,N_7203,N_7224);
and U7569 (N_7569,N_7382,N_7388);
and U7570 (N_7570,N_7319,N_7253);
nor U7571 (N_7571,N_7202,N_7291);
or U7572 (N_7572,N_7367,N_7336);
nand U7573 (N_7573,N_7280,N_7252);
nor U7574 (N_7574,N_7368,N_7222);
or U7575 (N_7575,N_7390,N_7297);
xnor U7576 (N_7576,N_7258,N_7286);
xnor U7577 (N_7577,N_7277,N_7259);
nand U7578 (N_7578,N_7363,N_7302);
xnor U7579 (N_7579,N_7322,N_7249);
xnor U7580 (N_7580,N_7250,N_7223);
or U7581 (N_7581,N_7252,N_7245);
or U7582 (N_7582,N_7338,N_7364);
nor U7583 (N_7583,N_7222,N_7301);
nand U7584 (N_7584,N_7337,N_7246);
nor U7585 (N_7585,N_7376,N_7266);
and U7586 (N_7586,N_7247,N_7309);
and U7587 (N_7587,N_7240,N_7222);
nor U7588 (N_7588,N_7248,N_7313);
and U7589 (N_7589,N_7359,N_7365);
nand U7590 (N_7590,N_7366,N_7330);
nand U7591 (N_7591,N_7272,N_7287);
xor U7592 (N_7592,N_7299,N_7271);
xor U7593 (N_7593,N_7231,N_7343);
nor U7594 (N_7594,N_7296,N_7269);
xnor U7595 (N_7595,N_7381,N_7207);
xor U7596 (N_7596,N_7317,N_7321);
nor U7597 (N_7597,N_7354,N_7259);
and U7598 (N_7598,N_7245,N_7398);
and U7599 (N_7599,N_7392,N_7206);
nor U7600 (N_7600,N_7556,N_7485);
xor U7601 (N_7601,N_7580,N_7593);
nor U7602 (N_7602,N_7459,N_7406);
or U7603 (N_7603,N_7407,N_7463);
nand U7604 (N_7604,N_7510,N_7426);
or U7605 (N_7605,N_7520,N_7428);
nor U7606 (N_7606,N_7567,N_7470);
nor U7607 (N_7607,N_7517,N_7415);
and U7608 (N_7608,N_7453,N_7478);
or U7609 (N_7609,N_7558,N_7499);
nor U7610 (N_7610,N_7548,N_7482);
nor U7611 (N_7611,N_7448,N_7435);
nand U7612 (N_7612,N_7443,N_7514);
xor U7613 (N_7613,N_7471,N_7466);
or U7614 (N_7614,N_7421,N_7592);
nand U7615 (N_7615,N_7598,N_7531);
nand U7616 (N_7616,N_7454,N_7481);
or U7617 (N_7617,N_7486,N_7461);
or U7618 (N_7618,N_7551,N_7577);
nand U7619 (N_7619,N_7560,N_7405);
nor U7620 (N_7620,N_7535,N_7524);
nor U7621 (N_7621,N_7494,N_7534);
and U7622 (N_7622,N_7501,N_7492);
nand U7623 (N_7623,N_7559,N_7477);
and U7624 (N_7624,N_7500,N_7587);
nand U7625 (N_7625,N_7589,N_7457);
and U7626 (N_7626,N_7410,N_7484);
and U7627 (N_7627,N_7546,N_7458);
xnor U7628 (N_7628,N_7452,N_7409);
xor U7629 (N_7629,N_7432,N_7555);
nand U7630 (N_7630,N_7442,N_7449);
xor U7631 (N_7631,N_7574,N_7515);
nor U7632 (N_7632,N_7430,N_7521);
and U7633 (N_7633,N_7505,N_7586);
nand U7634 (N_7634,N_7411,N_7456);
nor U7635 (N_7635,N_7544,N_7525);
xor U7636 (N_7636,N_7571,N_7402);
or U7637 (N_7637,N_7552,N_7464);
xor U7638 (N_7638,N_7476,N_7455);
nand U7639 (N_7639,N_7532,N_7594);
xnor U7640 (N_7640,N_7422,N_7403);
xor U7641 (N_7641,N_7557,N_7467);
and U7642 (N_7642,N_7599,N_7547);
nor U7643 (N_7643,N_7572,N_7434);
xor U7644 (N_7644,N_7491,N_7446);
xor U7645 (N_7645,N_7427,N_7563);
or U7646 (N_7646,N_7539,N_7550);
nor U7647 (N_7647,N_7549,N_7523);
nand U7648 (N_7648,N_7496,N_7412);
and U7649 (N_7649,N_7538,N_7495);
nor U7650 (N_7650,N_7445,N_7468);
nand U7651 (N_7651,N_7419,N_7502);
or U7652 (N_7652,N_7536,N_7472);
xnor U7653 (N_7653,N_7488,N_7582);
and U7654 (N_7654,N_7424,N_7516);
or U7655 (N_7655,N_7596,N_7584);
and U7656 (N_7656,N_7507,N_7498);
xor U7657 (N_7657,N_7462,N_7565);
nor U7658 (N_7658,N_7444,N_7489);
nand U7659 (N_7659,N_7438,N_7543);
or U7660 (N_7660,N_7423,N_7597);
xor U7661 (N_7661,N_7487,N_7591);
xor U7662 (N_7662,N_7564,N_7511);
xor U7663 (N_7663,N_7588,N_7480);
nor U7664 (N_7664,N_7418,N_7522);
xor U7665 (N_7665,N_7400,N_7429);
and U7666 (N_7666,N_7475,N_7440);
or U7667 (N_7667,N_7583,N_7401);
or U7668 (N_7668,N_7569,N_7519);
and U7669 (N_7669,N_7595,N_7490);
xor U7670 (N_7670,N_7441,N_7545);
nand U7671 (N_7671,N_7469,N_7528);
or U7672 (N_7672,N_7493,N_7568);
xor U7673 (N_7673,N_7433,N_7497);
xor U7674 (N_7674,N_7526,N_7527);
or U7675 (N_7675,N_7578,N_7576);
xor U7676 (N_7676,N_7554,N_7479);
or U7677 (N_7677,N_7590,N_7529);
nand U7678 (N_7678,N_7509,N_7450);
xor U7679 (N_7679,N_7420,N_7447);
xor U7680 (N_7680,N_7416,N_7518);
xnor U7681 (N_7681,N_7451,N_7575);
or U7682 (N_7682,N_7553,N_7436);
xnor U7683 (N_7683,N_7585,N_7542);
or U7684 (N_7684,N_7537,N_7561);
or U7685 (N_7685,N_7540,N_7425);
nor U7686 (N_7686,N_7408,N_7437);
xnor U7687 (N_7687,N_7566,N_7562);
nor U7688 (N_7688,N_7404,N_7581);
and U7689 (N_7689,N_7508,N_7417);
or U7690 (N_7690,N_7465,N_7503);
and U7691 (N_7691,N_7439,N_7414);
nand U7692 (N_7692,N_7473,N_7504);
or U7693 (N_7693,N_7541,N_7530);
xor U7694 (N_7694,N_7474,N_7460);
or U7695 (N_7695,N_7533,N_7513);
nor U7696 (N_7696,N_7570,N_7579);
or U7697 (N_7697,N_7506,N_7573);
or U7698 (N_7698,N_7512,N_7483);
xnor U7699 (N_7699,N_7413,N_7431);
nor U7700 (N_7700,N_7454,N_7412);
and U7701 (N_7701,N_7554,N_7499);
nand U7702 (N_7702,N_7508,N_7542);
xnor U7703 (N_7703,N_7511,N_7463);
nor U7704 (N_7704,N_7449,N_7577);
xor U7705 (N_7705,N_7415,N_7563);
or U7706 (N_7706,N_7515,N_7590);
nand U7707 (N_7707,N_7538,N_7455);
and U7708 (N_7708,N_7542,N_7423);
xnor U7709 (N_7709,N_7482,N_7498);
and U7710 (N_7710,N_7519,N_7597);
nand U7711 (N_7711,N_7541,N_7536);
nor U7712 (N_7712,N_7593,N_7437);
xor U7713 (N_7713,N_7516,N_7531);
nand U7714 (N_7714,N_7439,N_7527);
or U7715 (N_7715,N_7441,N_7516);
or U7716 (N_7716,N_7568,N_7560);
or U7717 (N_7717,N_7415,N_7521);
and U7718 (N_7718,N_7535,N_7585);
nor U7719 (N_7719,N_7427,N_7574);
and U7720 (N_7720,N_7461,N_7506);
and U7721 (N_7721,N_7552,N_7521);
or U7722 (N_7722,N_7479,N_7518);
xnor U7723 (N_7723,N_7401,N_7409);
nand U7724 (N_7724,N_7428,N_7412);
or U7725 (N_7725,N_7522,N_7553);
nand U7726 (N_7726,N_7448,N_7532);
nor U7727 (N_7727,N_7546,N_7425);
xnor U7728 (N_7728,N_7534,N_7402);
and U7729 (N_7729,N_7553,N_7498);
xnor U7730 (N_7730,N_7475,N_7467);
nand U7731 (N_7731,N_7470,N_7599);
xnor U7732 (N_7732,N_7552,N_7569);
nor U7733 (N_7733,N_7588,N_7481);
nand U7734 (N_7734,N_7592,N_7563);
nand U7735 (N_7735,N_7510,N_7592);
nor U7736 (N_7736,N_7515,N_7542);
nor U7737 (N_7737,N_7530,N_7436);
or U7738 (N_7738,N_7532,N_7433);
nand U7739 (N_7739,N_7517,N_7578);
and U7740 (N_7740,N_7445,N_7441);
or U7741 (N_7741,N_7582,N_7473);
nand U7742 (N_7742,N_7501,N_7573);
xor U7743 (N_7743,N_7418,N_7584);
xnor U7744 (N_7744,N_7565,N_7561);
and U7745 (N_7745,N_7512,N_7566);
xor U7746 (N_7746,N_7512,N_7500);
and U7747 (N_7747,N_7571,N_7531);
and U7748 (N_7748,N_7516,N_7522);
xnor U7749 (N_7749,N_7577,N_7546);
nand U7750 (N_7750,N_7567,N_7401);
nand U7751 (N_7751,N_7580,N_7532);
xor U7752 (N_7752,N_7475,N_7542);
nor U7753 (N_7753,N_7495,N_7519);
nand U7754 (N_7754,N_7407,N_7558);
nor U7755 (N_7755,N_7416,N_7588);
nor U7756 (N_7756,N_7546,N_7543);
and U7757 (N_7757,N_7490,N_7489);
or U7758 (N_7758,N_7539,N_7545);
or U7759 (N_7759,N_7533,N_7432);
nor U7760 (N_7760,N_7522,N_7457);
nor U7761 (N_7761,N_7453,N_7598);
nand U7762 (N_7762,N_7571,N_7543);
xor U7763 (N_7763,N_7436,N_7483);
nand U7764 (N_7764,N_7449,N_7486);
nor U7765 (N_7765,N_7428,N_7593);
xor U7766 (N_7766,N_7446,N_7576);
and U7767 (N_7767,N_7598,N_7406);
and U7768 (N_7768,N_7447,N_7416);
and U7769 (N_7769,N_7426,N_7411);
and U7770 (N_7770,N_7505,N_7408);
nor U7771 (N_7771,N_7460,N_7513);
nand U7772 (N_7772,N_7412,N_7555);
nand U7773 (N_7773,N_7449,N_7402);
xor U7774 (N_7774,N_7550,N_7533);
nor U7775 (N_7775,N_7523,N_7526);
nor U7776 (N_7776,N_7449,N_7475);
nor U7777 (N_7777,N_7555,N_7574);
nor U7778 (N_7778,N_7446,N_7536);
xor U7779 (N_7779,N_7519,N_7521);
xor U7780 (N_7780,N_7543,N_7547);
or U7781 (N_7781,N_7471,N_7586);
or U7782 (N_7782,N_7565,N_7566);
xnor U7783 (N_7783,N_7566,N_7523);
or U7784 (N_7784,N_7540,N_7533);
and U7785 (N_7785,N_7477,N_7466);
nor U7786 (N_7786,N_7432,N_7423);
xor U7787 (N_7787,N_7546,N_7549);
xnor U7788 (N_7788,N_7532,N_7432);
and U7789 (N_7789,N_7411,N_7501);
nand U7790 (N_7790,N_7550,N_7545);
and U7791 (N_7791,N_7426,N_7465);
nand U7792 (N_7792,N_7476,N_7460);
or U7793 (N_7793,N_7544,N_7451);
nor U7794 (N_7794,N_7431,N_7569);
xnor U7795 (N_7795,N_7569,N_7572);
or U7796 (N_7796,N_7510,N_7501);
or U7797 (N_7797,N_7464,N_7410);
or U7798 (N_7798,N_7409,N_7469);
nor U7799 (N_7799,N_7445,N_7448);
or U7800 (N_7800,N_7667,N_7715);
and U7801 (N_7801,N_7713,N_7650);
or U7802 (N_7802,N_7770,N_7787);
or U7803 (N_7803,N_7724,N_7632);
xor U7804 (N_7804,N_7683,N_7736);
and U7805 (N_7805,N_7657,N_7615);
xnor U7806 (N_7806,N_7761,N_7705);
and U7807 (N_7807,N_7790,N_7763);
or U7808 (N_7808,N_7660,N_7684);
or U7809 (N_7809,N_7747,N_7737);
nand U7810 (N_7810,N_7612,N_7640);
xor U7811 (N_7811,N_7651,N_7745);
nor U7812 (N_7812,N_7712,N_7799);
and U7813 (N_7813,N_7695,N_7620);
or U7814 (N_7814,N_7607,N_7744);
and U7815 (N_7815,N_7655,N_7642);
nand U7816 (N_7816,N_7796,N_7746);
nor U7817 (N_7817,N_7685,N_7696);
nor U7818 (N_7818,N_7706,N_7728);
xor U7819 (N_7819,N_7639,N_7654);
or U7820 (N_7820,N_7621,N_7791);
or U7821 (N_7821,N_7643,N_7617);
nor U7822 (N_7822,N_7666,N_7623);
or U7823 (N_7823,N_7785,N_7711);
xnor U7824 (N_7824,N_7740,N_7633);
nand U7825 (N_7825,N_7600,N_7648);
and U7826 (N_7826,N_7663,N_7776);
xnor U7827 (N_7827,N_7738,N_7602);
xor U7828 (N_7828,N_7652,N_7754);
xor U7829 (N_7829,N_7760,N_7645);
and U7830 (N_7830,N_7613,N_7694);
xor U7831 (N_7831,N_7622,N_7778);
nand U7832 (N_7832,N_7759,N_7638);
and U7833 (N_7833,N_7668,N_7699);
or U7834 (N_7834,N_7741,N_7606);
or U7835 (N_7835,N_7735,N_7693);
and U7836 (N_7836,N_7777,N_7714);
and U7837 (N_7837,N_7722,N_7686);
or U7838 (N_7838,N_7672,N_7676);
xor U7839 (N_7839,N_7682,N_7749);
nand U7840 (N_7840,N_7700,N_7618);
nand U7841 (N_7841,N_7750,N_7678);
or U7842 (N_7842,N_7730,N_7635);
and U7843 (N_7843,N_7691,N_7644);
or U7844 (N_7844,N_7614,N_7649);
and U7845 (N_7845,N_7679,N_7721);
and U7846 (N_7846,N_7729,N_7637);
nand U7847 (N_7847,N_7688,N_7731);
nor U7848 (N_7848,N_7793,N_7647);
nor U7849 (N_7849,N_7634,N_7681);
nor U7850 (N_7850,N_7718,N_7771);
and U7851 (N_7851,N_7627,N_7701);
nand U7852 (N_7852,N_7739,N_7662);
and U7853 (N_7853,N_7719,N_7727);
xor U7854 (N_7854,N_7603,N_7631);
nor U7855 (N_7855,N_7766,N_7624);
and U7856 (N_7856,N_7628,N_7795);
nand U7857 (N_7857,N_7726,N_7783);
nand U7858 (N_7858,N_7646,N_7773);
and U7859 (N_7859,N_7601,N_7675);
xnor U7860 (N_7860,N_7674,N_7670);
xor U7861 (N_7861,N_7704,N_7797);
nor U7862 (N_7862,N_7774,N_7756);
or U7863 (N_7863,N_7680,N_7702);
nand U7864 (N_7864,N_7608,N_7762);
nand U7865 (N_7865,N_7788,N_7665);
nor U7866 (N_7866,N_7625,N_7708);
and U7867 (N_7867,N_7610,N_7733);
xor U7868 (N_7868,N_7779,N_7619);
nand U7869 (N_7869,N_7629,N_7758);
nand U7870 (N_7870,N_7786,N_7753);
nand U7871 (N_7871,N_7709,N_7604);
nand U7872 (N_7872,N_7653,N_7723);
nand U7873 (N_7873,N_7673,N_7677);
nor U7874 (N_7874,N_7755,N_7768);
and U7875 (N_7875,N_7717,N_7732);
nand U7876 (N_7876,N_7751,N_7687);
or U7877 (N_7877,N_7765,N_7792);
nand U7878 (N_7878,N_7641,N_7703);
nor U7879 (N_7879,N_7764,N_7757);
xnor U7880 (N_7880,N_7767,N_7697);
nor U7881 (N_7881,N_7781,N_7664);
or U7882 (N_7882,N_7775,N_7626);
and U7883 (N_7883,N_7794,N_7636);
nand U7884 (N_7884,N_7690,N_7784);
nand U7885 (N_7885,N_7720,N_7616);
and U7886 (N_7886,N_7782,N_7798);
nor U7887 (N_7887,N_7710,N_7789);
nand U7888 (N_7888,N_7605,N_7659);
or U7889 (N_7889,N_7752,N_7769);
xor U7890 (N_7890,N_7661,N_7716);
nor U7891 (N_7891,N_7780,N_7725);
nand U7892 (N_7892,N_7772,N_7671);
xnor U7893 (N_7893,N_7689,N_7748);
nand U7894 (N_7894,N_7656,N_7611);
and U7895 (N_7895,N_7630,N_7742);
or U7896 (N_7896,N_7658,N_7609);
nor U7897 (N_7897,N_7669,N_7743);
nor U7898 (N_7898,N_7698,N_7707);
xnor U7899 (N_7899,N_7692,N_7734);
nand U7900 (N_7900,N_7734,N_7694);
or U7901 (N_7901,N_7716,N_7659);
nor U7902 (N_7902,N_7729,N_7681);
nor U7903 (N_7903,N_7619,N_7646);
or U7904 (N_7904,N_7666,N_7723);
xor U7905 (N_7905,N_7626,N_7674);
and U7906 (N_7906,N_7797,N_7652);
nand U7907 (N_7907,N_7676,N_7677);
nor U7908 (N_7908,N_7796,N_7772);
nand U7909 (N_7909,N_7732,N_7602);
and U7910 (N_7910,N_7696,N_7615);
nor U7911 (N_7911,N_7690,N_7671);
xnor U7912 (N_7912,N_7698,N_7726);
nand U7913 (N_7913,N_7796,N_7605);
and U7914 (N_7914,N_7755,N_7600);
xor U7915 (N_7915,N_7635,N_7671);
or U7916 (N_7916,N_7676,N_7710);
and U7917 (N_7917,N_7636,N_7798);
and U7918 (N_7918,N_7682,N_7736);
nand U7919 (N_7919,N_7619,N_7716);
and U7920 (N_7920,N_7755,N_7644);
nor U7921 (N_7921,N_7709,N_7745);
or U7922 (N_7922,N_7695,N_7772);
nand U7923 (N_7923,N_7745,N_7725);
and U7924 (N_7924,N_7665,N_7734);
nand U7925 (N_7925,N_7709,N_7635);
nand U7926 (N_7926,N_7671,N_7707);
nand U7927 (N_7927,N_7604,N_7671);
nand U7928 (N_7928,N_7728,N_7646);
nor U7929 (N_7929,N_7658,N_7690);
and U7930 (N_7930,N_7687,N_7698);
and U7931 (N_7931,N_7635,N_7626);
nor U7932 (N_7932,N_7706,N_7723);
and U7933 (N_7933,N_7703,N_7755);
nor U7934 (N_7934,N_7625,N_7773);
or U7935 (N_7935,N_7612,N_7747);
xnor U7936 (N_7936,N_7707,N_7656);
or U7937 (N_7937,N_7673,N_7744);
xnor U7938 (N_7938,N_7609,N_7694);
and U7939 (N_7939,N_7746,N_7763);
or U7940 (N_7940,N_7722,N_7694);
or U7941 (N_7941,N_7730,N_7603);
nand U7942 (N_7942,N_7632,N_7762);
xnor U7943 (N_7943,N_7773,N_7764);
nand U7944 (N_7944,N_7632,N_7613);
nor U7945 (N_7945,N_7785,N_7641);
and U7946 (N_7946,N_7674,N_7782);
xnor U7947 (N_7947,N_7769,N_7700);
nor U7948 (N_7948,N_7638,N_7622);
or U7949 (N_7949,N_7650,N_7743);
xnor U7950 (N_7950,N_7796,N_7745);
and U7951 (N_7951,N_7713,N_7632);
and U7952 (N_7952,N_7601,N_7621);
nor U7953 (N_7953,N_7730,N_7659);
and U7954 (N_7954,N_7641,N_7799);
and U7955 (N_7955,N_7765,N_7628);
or U7956 (N_7956,N_7674,N_7614);
nand U7957 (N_7957,N_7609,N_7704);
nor U7958 (N_7958,N_7766,N_7788);
and U7959 (N_7959,N_7722,N_7687);
nor U7960 (N_7960,N_7661,N_7730);
or U7961 (N_7961,N_7770,N_7778);
and U7962 (N_7962,N_7674,N_7695);
nor U7963 (N_7963,N_7641,N_7752);
and U7964 (N_7964,N_7667,N_7600);
nand U7965 (N_7965,N_7696,N_7666);
xnor U7966 (N_7966,N_7653,N_7793);
nand U7967 (N_7967,N_7608,N_7740);
and U7968 (N_7968,N_7767,N_7671);
and U7969 (N_7969,N_7737,N_7767);
xor U7970 (N_7970,N_7742,N_7792);
nor U7971 (N_7971,N_7758,N_7761);
nor U7972 (N_7972,N_7799,N_7718);
or U7973 (N_7973,N_7662,N_7660);
or U7974 (N_7974,N_7631,N_7721);
xnor U7975 (N_7975,N_7784,N_7767);
xnor U7976 (N_7976,N_7774,N_7666);
nand U7977 (N_7977,N_7680,N_7697);
and U7978 (N_7978,N_7708,N_7733);
nand U7979 (N_7979,N_7612,N_7764);
nand U7980 (N_7980,N_7683,N_7691);
nand U7981 (N_7981,N_7609,N_7701);
nand U7982 (N_7982,N_7768,N_7778);
or U7983 (N_7983,N_7775,N_7666);
nor U7984 (N_7984,N_7744,N_7790);
nand U7985 (N_7985,N_7672,N_7787);
and U7986 (N_7986,N_7686,N_7690);
xor U7987 (N_7987,N_7642,N_7677);
nand U7988 (N_7988,N_7624,N_7750);
nand U7989 (N_7989,N_7714,N_7677);
or U7990 (N_7990,N_7615,N_7602);
xnor U7991 (N_7991,N_7655,N_7632);
or U7992 (N_7992,N_7736,N_7772);
or U7993 (N_7993,N_7782,N_7742);
nor U7994 (N_7994,N_7792,N_7716);
nor U7995 (N_7995,N_7688,N_7790);
nor U7996 (N_7996,N_7657,N_7692);
and U7997 (N_7997,N_7619,N_7743);
or U7998 (N_7998,N_7654,N_7671);
or U7999 (N_7999,N_7707,N_7735);
or U8000 (N_8000,N_7941,N_7860);
xnor U8001 (N_8001,N_7886,N_7882);
and U8002 (N_8002,N_7819,N_7807);
xnor U8003 (N_8003,N_7858,N_7947);
xnor U8004 (N_8004,N_7929,N_7820);
xor U8005 (N_8005,N_7992,N_7922);
and U8006 (N_8006,N_7969,N_7879);
and U8007 (N_8007,N_7822,N_7887);
or U8008 (N_8008,N_7984,N_7883);
and U8009 (N_8009,N_7974,N_7980);
nor U8010 (N_8010,N_7966,N_7872);
and U8011 (N_8011,N_7948,N_7977);
xnor U8012 (N_8012,N_7938,N_7940);
nor U8013 (N_8013,N_7880,N_7821);
xnor U8014 (N_8014,N_7895,N_7812);
nand U8015 (N_8015,N_7874,N_7877);
nand U8016 (N_8016,N_7825,N_7916);
xnor U8017 (N_8017,N_7806,N_7893);
xor U8018 (N_8018,N_7870,N_7962);
nand U8019 (N_8019,N_7926,N_7815);
and U8020 (N_8020,N_7907,N_7934);
xor U8021 (N_8021,N_7976,N_7991);
or U8022 (N_8022,N_7824,N_7891);
or U8023 (N_8023,N_7987,N_7931);
nand U8024 (N_8024,N_7840,N_7867);
and U8025 (N_8025,N_7901,N_7950);
and U8026 (N_8026,N_7855,N_7856);
nand U8027 (N_8027,N_7919,N_7920);
nand U8028 (N_8028,N_7839,N_7906);
nor U8029 (N_8029,N_7888,N_7833);
nor U8030 (N_8030,N_7951,N_7838);
nor U8031 (N_8031,N_7921,N_7939);
xnor U8032 (N_8032,N_7998,N_7881);
nand U8033 (N_8033,N_7981,N_7865);
nor U8034 (N_8034,N_7862,N_7955);
and U8035 (N_8035,N_7971,N_7935);
nor U8036 (N_8036,N_7896,N_7843);
or U8037 (N_8037,N_7917,N_7875);
or U8038 (N_8038,N_7871,N_7829);
and U8039 (N_8039,N_7808,N_7816);
or U8040 (N_8040,N_7996,N_7942);
and U8041 (N_8041,N_7805,N_7944);
nand U8042 (N_8042,N_7831,N_7912);
nor U8043 (N_8043,N_7803,N_7849);
or U8044 (N_8044,N_7817,N_7986);
nand U8045 (N_8045,N_7811,N_7841);
and U8046 (N_8046,N_7924,N_7842);
and U8047 (N_8047,N_7884,N_7964);
xnor U8048 (N_8048,N_7914,N_7837);
nand U8049 (N_8049,N_7994,N_7897);
or U8050 (N_8050,N_7956,N_7848);
xor U8051 (N_8051,N_7900,N_7918);
xor U8052 (N_8052,N_7846,N_7913);
nor U8053 (N_8053,N_7973,N_7970);
nor U8054 (N_8054,N_7930,N_7979);
or U8055 (N_8055,N_7801,N_7937);
or U8056 (N_8056,N_7993,N_7990);
and U8057 (N_8057,N_7864,N_7898);
and U8058 (N_8058,N_7999,N_7863);
nand U8059 (N_8059,N_7835,N_7949);
xnor U8060 (N_8060,N_7857,N_7945);
and U8061 (N_8061,N_7905,N_7818);
and U8062 (N_8062,N_7975,N_7943);
nor U8063 (N_8063,N_7972,N_7902);
xor U8064 (N_8064,N_7978,N_7952);
and U8065 (N_8065,N_7885,N_7845);
or U8066 (N_8066,N_7911,N_7954);
nand U8067 (N_8067,N_7953,N_7989);
nand U8068 (N_8068,N_7910,N_7927);
xnor U8069 (N_8069,N_7894,N_7869);
or U8070 (N_8070,N_7890,N_7866);
xnor U8071 (N_8071,N_7995,N_7960);
nor U8072 (N_8072,N_7915,N_7823);
or U8073 (N_8073,N_7982,N_7853);
nor U8074 (N_8074,N_7832,N_7827);
nand U8075 (N_8075,N_7958,N_7965);
nand U8076 (N_8076,N_7850,N_7988);
xnor U8077 (N_8077,N_7946,N_7925);
xnor U8078 (N_8078,N_7933,N_7903);
or U8079 (N_8079,N_7834,N_7810);
nand U8080 (N_8080,N_7859,N_7923);
nor U8081 (N_8081,N_7861,N_7828);
and U8082 (N_8082,N_7851,N_7813);
or U8083 (N_8083,N_7959,N_7847);
nor U8084 (N_8084,N_7800,N_7968);
and U8085 (N_8085,N_7909,N_7873);
nor U8086 (N_8086,N_7963,N_7876);
xnor U8087 (N_8087,N_7985,N_7868);
nand U8088 (N_8088,N_7928,N_7814);
and U8089 (N_8089,N_7904,N_7899);
and U8090 (N_8090,N_7908,N_7936);
and U8091 (N_8091,N_7967,N_7957);
xor U8092 (N_8092,N_7997,N_7852);
and U8093 (N_8093,N_7804,N_7844);
and U8094 (N_8094,N_7889,N_7892);
nor U8095 (N_8095,N_7961,N_7878);
and U8096 (N_8096,N_7836,N_7802);
and U8097 (N_8097,N_7826,N_7854);
or U8098 (N_8098,N_7932,N_7830);
or U8099 (N_8099,N_7809,N_7983);
nand U8100 (N_8100,N_7817,N_7868);
or U8101 (N_8101,N_7874,N_7978);
nor U8102 (N_8102,N_7817,N_7886);
nor U8103 (N_8103,N_7917,N_7972);
nor U8104 (N_8104,N_7902,N_7869);
nand U8105 (N_8105,N_7806,N_7978);
xor U8106 (N_8106,N_7995,N_7805);
xnor U8107 (N_8107,N_7932,N_7806);
and U8108 (N_8108,N_7989,N_7956);
nor U8109 (N_8109,N_7889,N_7908);
nor U8110 (N_8110,N_7943,N_7914);
or U8111 (N_8111,N_7990,N_7916);
xnor U8112 (N_8112,N_7878,N_7820);
nor U8113 (N_8113,N_7859,N_7977);
nand U8114 (N_8114,N_7943,N_7925);
nand U8115 (N_8115,N_7804,N_7955);
xnor U8116 (N_8116,N_7879,N_7902);
xor U8117 (N_8117,N_7892,N_7989);
xor U8118 (N_8118,N_7841,N_7951);
xnor U8119 (N_8119,N_7899,N_7816);
and U8120 (N_8120,N_7917,N_7895);
or U8121 (N_8121,N_7910,N_7867);
xnor U8122 (N_8122,N_7914,N_7888);
and U8123 (N_8123,N_7932,N_7802);
or U8124 (N_8124,N_7904,N_7906);
or U8125 (N_8125,N_7852,N_7893);
nand U8126 (N_8126,N_7815,N_7953);
nand U8127 (N_8127,N_7833,N_7903);
or U8128 (N_8128,N_7810,N_7988);
nor U8129 (N_8129,N_7806,N_7958);
or U8130 (N_8130,N_7998,N_7968);
xnor U8131 (N_8131,N_7870,N_7925);
nor U8132 (N_8132,N_7971,N_7869);
nor U8133 (N_8133,N_7919,N_7890);
nor U8134 (N_8134,N_7936,N_7938);
xor U8135 (N_8135,N_7938,N_7854);
or U8136 (N_8136,N_7921,N_7890);
or U8137 (N_8137,N_7934,N_7804);
xnor U8138 (N_8138,N_7879,N_7958);
or U8139 (N_8139,N_7815,N_7898);
and U8140 (N_8140,N_7987,N_7834);
or U8141 (N_8141,N_7984,N_7923);
or U8142 (N_8142,N_7880,N_7990);
nor U8143 (N_8143,N_7834,N_7900);
or U8144 (N_8144,N_7884,N_7920);
nand U8145 (N_8145,N_7940,N_7975);
and U8146 (N_8146,N_7891,N_7854);
nand U8147 (N_8147,N_7830,N_7910);
and U8148 (N_8148,N_7902,N_7918);
nand U8149 (N_8149,N_7875,N_7944);
nand U8150 (N_8150,N_7929,N_7878);
nand U8151 (N_8151,N_7836,N_7937);
or U8152 (N_8152,N_7942,N_7972);
nor U8153 (N_8153,N_7855,N_7987);
nor U8154 (N_8154,N_7957,N_7814);
and U8155 (N_8155,N_7992,N_7812);
xnor U8156 (N_8156,N_7959,N_7882);
xor U8157 (N_8157,N_7848,N_7852);
nor U8158 (N_8158,N_7821,N_7828);
nor U8159 (N_8159,N_7820,N_7856);
nor U8160 (N_8160,N_7945,N_7933);
nor U8161 (N_8161,N_7932,N_7903);
nand U8162 (N_8162,N_7886,N_7875);
nor U8163 (N_8163,N_7979,N_7942);
nor U8164 (N_8164,N_7892,N_7817);
nor U8165 (N_8165,N_7919,N_7854);
and U8166 (N_8166,N_7913,N_7866);
nand U8167 (N_8167,N_7934,N_7926);
or U8168 (N_8168,N_7905,N_7963);
xor U8169 (N_8169,N_7806,N_7827);
nand U8170 (N_8170,N_7881,N_7952);
or U8171 (N_8171,N_7996,N_7901);
or U8172 (N_8172,N_7894,N_7946);
nor U8173 (N_8173,N_7875,N_7874);
or U8174 (N_8174,N_7852,N_7901);
nor U8175 (N_8175,N_7887,N_7880);
nor U8176 (N_8176,N_7843,N_7920);
or U8177 (N_8177,N_7834,N_7968);
or U8178 (N_8178,N_7847,N_7985);
nor U8179 (N_8179,N_7921,N_7859);
or U8180 (N_8180,N_7890,N_7821);
nand U8181 (N_8181,N_7811,N_7870);
nor U8182 (N_8182,N_7832,N_7877);
nor U8183 (N_8183,N_7982,N_7927);
xnor U8184 (N_8184,N_7856,N_7933);
nor U8185 (N_8185,N_7903,N_7945);
nor U8186 (N_8186,N_7947,N_7981);
nor U8187 (N_8187,N_7995,N_7934);
and U8188 (N_8188,N_7855,N_7890);
xor U8189 (N_8189,N_7913,N_7805);
nor U8190 (N_8190,N_7847,N_7991);
xnor U8191 (N_8191,N_7877,N_7976);
and U8192 (N_8192,N_7813,N_7806);
nand U8193 (N_8193,N_7992,N_7956);
nor U8194 (N_8194,N_7955,N_7984);
xor U8195 (N_8195,N_7817,N_7943);
nand U8196 (N_8196,N_7821,N_7839);
xor U8197 (N_8197,N_7886,N_7889);
nor U8198 (N_8198,N_7956,N_7962);
xor U8199 (N_8199,N_7999,N_7870);
nand U8200 (N_8200,N_8001,N_8101);
and U8201 (N_8201,N_8022,N_8144);
nand U8202 (N_8202,N_8116,N_8014);
nand U8203 (N_8203,N_8186,N_8032);
or U8204 (N_8204,N_8130,N_8125);
xor U8205 (N_8205,N_8170,N_8058);
or U8206 (N_8206,N_8162,N_8195);
nor U8207 (N_8207,N_8098,N_8018);
and U8208 (N_8208,N_8167,N_8061);
xor U8209 (N_8209,N_8164,N_8077);
nand U8210 (N_8210,N_8154,N_8078);
or U8211 (N_8211,N_8073,N_8013);
and U8212 (N_8212,N_8026,N_8194);
nor U8213 (N_8213,N_8056,N_8159);
and U8214 (N_8214,N_8168,N_8107);
or U8215 (N_8215,N_8131,N_8051);
and U8216 (N_8216,N_8151,N_8057);
and U8217 (N_8217,N_8156,N_8063);
nand U8218 (N_8218,N_8008,N_8119);
and U8219 (N_8219,N_8011,N_8082);
and U8220 (N_8220,N_8071,N_8102);
or U8221 (N_8221,N_8142,N_8070);
nor U8222 (N_8222,N_8065,N_8182);
and U8223 (N_8223,N_8084,N_8104);
nand U8224 (N_8224,N_8190,N_8046);
xor U8225 (N_8225,N_8122,N_8176);
and U8226 (N_8226,N_8062,N_8157);
nand U8227 (N_8227,N_8035,N_8052);
or U8228 (N_8228,N_8113,N_8054);
and U8229 (N_8229,N_8042,N_8089);
and U8230 (N_8230,N_8141,N_8085);
nand U8231 (N_8231,N_8128,N_8185);
and U8232 (N_8232,N_8147,N_8193);
or U8233 (N_8233,N_8036,N_8175);
and U8234 (N_8234,N_8006,N_8152);
or U8235 (N_8235,N_8103,N_8038);
nor U8236 (N_8236,N_8079,N_8124);
or U8237 (N_8237,N_8149,N_8118);
or U8238 (N_8238,N_8110,N_8148);
or U8239 (N_8239,N_8121,N_8187);
or U8240 (N_8240,N_8112,N_8000);
and U8241 (N_8241,N_8015,N_8016);
nor U8242 (N_8242,N_8199,N_8060);
nand U8243 (N_8243,N_8012,N_8120);
xnor U8244 (N_8244,N_8047,N_8091);
nor U8245 (N_8245,N_8109,N_8129);
nor U8246 (N_8246,N_8024,N_8075);
nand U8247 (N_8247,N_8177,N_8096);
xor U8248 (N_8248,N_8068,N_8086);
and U8249 (N_8249,N_8002,N_8053);
and U8250 (N_8250,N_8090,N_8074);
and U8251 (N_8251,N_8066,N_8135);
nor U8252 (N_8252,N_8025,N_8049);
xnor U8253 (N_8253,N_8150,N_8092);
xnor U8254 (N_8254,N_8072,N_8076);
and U8255 (N_8255,N_8048,N_8067);
xor U8256 (N_8256,N_8108,N_8050);
or U8257 (N_8257,N_8095,N_8171);
or U8258 (N_8258,N_8140,N_8181);
xor U8259 (N_8259,N_8059,N_8126);
nand U8260 (N_8260,N_8111,N_8040);
nor U8261 (N_8261,N_8037,N_8044);
or U8262 (N_8262,N_8097,N_8027);
or U8263 (N_8263,N_8146,N_8033);
and U8264 (N_8264,N_8045,N_8180);
and U8265 (N_8265,N_8155,N_8105);
or U8266 (N_8266,N_8117,N_8139);
and U8267 (N_8267,N_8114,N_8158);
nand U8268 (N_8268,N_8138,N_8153);
xnor U8269 (N_8269,N_8030,N_8019);
nand U8270 (N_8270,N_8088,N_8034);
nand U8271 (N_8271,N_8133,N_8161);
nor U8272 (N_8272,N_8198,N_8134);
or U8273 (N_8273,N_8007,N_8132);
nand U8274 (N_8274,N_8173,N_8174);
xor U8275 (N_8275,N_8127,N_8028);
and U8276 (N_8276,N_8010,N_8169);
and U8277 (N_8277,N_8136,N_8023);
or U8278 (N_8278,N_8069,N_8087);
nor U8279 (N_8279,N_8083,N_8172);
nor U8280 (N_8280,N_8183,N_8029);
and U8281 (N_8281,N_8184,N_8005);
nand U8282 (N_8282,N_8137,N_8145);
nand U8283 (N_8283,N_8123,N_8100);
nand U8284 (N_8284,N_8165,N_8009);
xor U8285 (N_8285,N_8039,N_8094);
and U8286 (N_8286,N_8020,N_8031);
and U8287 (N_8287,N_8166,N_8081);
or U8288 (N_8288,N_8163,N_8115);
or U8289 (N_8289,N_8191,N_8080);
xor U8290 (N_8290,N_8017,N_8178);
or U8291 (N_8291,N_8055,N_8192);
nand U8292 (N_8292,N_8043,N_8003);
xnor U8293 (N_8293,N_8099,N_8106);
xor U8294 (N_8294,N_8197,N_8004);
xor U8295 (N_8295,N_8093,N_8064);
xor U8296 (N_8296,N_8196,N_8189);
and U8297 (N_8297,N_8021,N_8160);
or U8298 (N_8298,N_8179,N_8041);
nor U8299 (N_8299,N_8143,N_8188);
or U8300 (N_8300,N_8169,N_8036);
and U8301 (N_8301,N_8029,N_8108);
xnor U8302 (N_8302,N_8147,N_8196);
or U8303 (N_8303,N_8178,N_8142);
nor U8304 (N_8304,N_8165,N_8196);
or U8305 (N_8305,N_8109,N_8055);
xnor U8306 (N_8306,N_8058,N_8176);
and U8307 (N_8307,N_8011,N_8094);
nor U8308 (N_8308,N_8048,N_8068);
or U8309 (N_8309,N_8056,N_8057);
xnor U8310 (N_8310,N_8190,N_8122);
nor U8311 (N_8311,N_8014,N_8073);
xor U8312 (N_8312,N_8161,N_8162);
xor U8313 (N_8313,N_8157,N_8059);
xor U8314 (N_8314,N_8056,N_8023);
xnor U8315 (N_8315,N_8142,N_8192);
xnor U8316 (N_8316,N_8117,N_8085);
xnor U8317 (N_8317,N_8092,N_8154);
xor U8318 (N_8318,N_8059,N_8031);
and U8319 (N_8319,N_8169,N_8089);
and U8320 (N_8320,N_8101,N_8196);
and U8321 (N_8321,N_8009,N_8167);
and U8322 (N_8322,N_8026,N_8006);
or U8323 (N_8323,N_8192,N_8114);
nand U8324 (N_8324,N_8160,N_8078);
nand U8325 (N_8325,N_8134,N_8145);
or U8326 (N_8326,N_8074,N_8044);
xnor U8327 (N_8327,N_8003,N_8032);
or U8328 (N_8328,N_8135,N_8046);
nor U8329 (N_8329,N_8163,N_8145);
nor U8330 (N_8330,N_8034,N_8102);
or U8331 (N_8331,N_8026,N_8054);
xor U8332 (N_8332,N_8004,N_8173);
and U8333 (N_8333,N_8129,N_8173);
nor U8334 (N_8334,N_8182,N_8048);
xnor U8335 (N_8335,N_8153,N_8123);
and U8336 (N_8336,N_8052,N_8067);
nand U8337 (N_8337,N_8015,N_8079);
nand U8338 (N_8338,N_8181,N_8045);
nor U8339 (N_8339,N_8145,N_8012);
and U8340 (N_8340,N_8064,N_8030);
nand U8341 (N_8341,N_8030,N_8054);
and U8342 (N_8342,N_8151,N_8177);
nand U8343 (N_8343,N_8013,N_8017);
and U8344 (N_8344,N_8025,N_8161);
nor U8345 (N_8345,N_8129,N_8116);
or U8346 (N_8346,N_8150,N_8157);
xor U8347 (N_8347,N_8169,N_8166);
or U8348 (N_8348,N_8114,N_8093);
xor U8349 (N_8349,N_8147,N_8152);
nor U8350 (N_8350,N_8120,N_8171);
nand U8351 (N_8351,N_8069,N_8139);
and U8352 (N_8352,N_8109,N_8074);
nand U8353 (N_8353,N_8087,N_8151);
xor U8354 (N_8354,N_8078,N_8119);
nand U8355 (N_8355,N_8071,N_8049);
or U8356 (N_8356,N_8034,N_8110);
nand U8357 (N_8357,N_8123,N_8199);
or U8358 (N_8358,N_8004,N_8033);
nand U8359 (N_8359,N_8148,N_8039);
and U8360 (N_8360,N_8178,N_8196);
nor U8361 (N_8361,N_8114,N_8102);
nor U8362 (N_8362,N_8033,N_8058);
xnor U8363 (N_8363,N_8144,N_8048);
and U8364 (N_8364,N_8023,N_8043);
or U8365 (N_8365,N_8064,N_8181);
xor U8366 (N_8366,N_8051,N_8022);
xnor U8367 (N_8367,N_8140,N_8027);
or U8368 (N_8368,N_8066,N_8165);
or U8369 (N_8369,N_8056,N_8198);
nor U8370 (N_8370,N_8152,N_8017);
xor U8371 (N_8371,N_8150,N_8099);
nor U8372 (N_8372,N_8168,N_8063);
and U8373 (N_8373,N_8157,N_8128);
nor U8374 (N_8374,N_8064,N_8130);
or U8375 (N_8375,N_8136,N_8164);
xor U8376 (N_8376,N_8081,N_8004);
or U8377 (N_8377,N_8045,N_8039);
and U8378 (N_8378,N_8042,N_8015);
xnor U8379 (N_8379,N_8083,N_8120);
and U8380 (N_8380,N_8007,N_8117);
and U8381 (N_8381,N_8123,N_8092);
nand U8382 (N_8382,N_8056,N_8078);
nand U8383 (N_8383,N_8028,N_8146);
nand U8384 (N_8384,N_8102,N_8156);
xor U8385 (N_8385,N_8037,N_8114);
or U8386 (N_8386,N_8011,N_8066);
xnor U8387 (N_8387,N_8091,N_8117);
or U8388 (N_8388,N_8108,N_8196);
nor U8389 (N_8389,N_8164,N_8027);
nand U8390 (N_8390,N_8041,N_8050);
nor U8391 (N_8391,N_8156,N_8024);
nor U8392 (N_8392,N_8125,N_8071);
and U8393 (N_8393,N_8110,N_8002);
and U8394 (N_8394,N_8045,N_8139);
nand U8395 (N_8395,N_8061,N_8008);
nand U8396 (N_8396,N_8159,N_8021);
xnor U8397 (N_8397,N_8129,N_8018);
and U8398 (N_8398,N_8056,N_8065);
xor U8399 (N_8399,N_8027,N_8105);
and U8400 (N_8400,N_8226,N_8374);
nor U8401 (N_8401,N_8280,N_8368);
nand U8402 (N_8402,N_8291,N_8371);
or U8403 (N_8403,N_8246,N_8210);
and U8404 (N_8404,N_8327,N_8223);
nor U8405 (N_8405,N_8243,N_8359);
xor U8406 (N_8406,N_8204,N_8345);
nand U8407 (N_8407,N_8289,N_8317);
or U8408 (N_8408,N_8228,N_8263);
nor U8409 (N_8409,N_8207,N_8253);
xnor U8410 (N_8410,N_8241,N_8252);
xor U8411 (N_8411,N_8342,N_8383);
xnor U8412 (N_8412,N_8202,N_8300);
xnor U8413 (N_8413,N_8259,N_8255);
nand U8414 (N_8414,N_8301,N_8377);
and U8415 (N_8415,N_8331,N_8386);
nor U8416 (N_8416,N_8363,N_8395);
nand U8417 (N_8417,N_8298,N_8311);
nor U8418 (N_8418,N_8360,N_8339);
xnor U8419 (N_8419,N_8308,N_8251);
and U8420 (N_8420,N_8231,N_8355);
and U8421 (N_8421,N_8281,N_8315);
nor U8422 (N_8422,N_8380,N_8296);
or U8423 (N_8423,N_8379,N_8306);
nand U8424 (N_8424,N_8334,N_8325);
xnor U8425 (N_8425,N_8215,N_8320);
and U8426 (N_8426,N_8240,N_8353);
nor U8427 (N_8427,N_8272,N_8235);
and U8428 (N_8428,N_8277,N_8389);
xnor U8429 (N_8429,N_8351,N_8385);
nor U8430 (N_8430,N_8384,N_8218);
or U8431 (N_8431,N_8271,N_8323);
or U8432 (N_8432,N_8273,N_8214);
and U8433 (N_8433,N_8352,N_8347);
nor U8434 (N_8434,N_8248,N_8358);
or U8435 (N_8435,N_8269,N_8237);
xor U8436 (N_8436,N_8330,N_8369);
or U8437 (N_8437,N_8211,N_8344);
nand U8438 (N_8438,N_8373,N_8364);
nor U8439 (N_8439,N_8205,N_8266);
or U8440 (N_8440,N_8387,N_8203);
nand U8441 (N_8441,N_8340,N_8378);
and U8442 (N_8442,N_8314,N_8382);
nor U8443 (N_8443,N_8397,N_8309);
and U8444 (N_8444,N_8396,N_8305);
or U8445 (N_8445,N_8318,N_8260);
nor U8446 (N_8446,N_8362,N_8232);
and U8447 (N_8447,N_8227,N_8265);
nor U8448 (N_8448,N_8322,N_8221);
xor U8449 (N_8449,N_8268,N_8290);
nor U8450 (N_8450,N_8326,N_8287);
nor U8451 (N_8451,N_8254,N_8264);
and U8452 (N_8452,N_8350,N_8367);
nand U8453 (N_8453,N_8299,N_8388);
nand U8454 (N_8454,N_8256,N_8216);
or U8455 (N_8455,N_8302,N_8249);
nor U8456 (N_8456,N_8201,N_8349);
nor U8457 (N_8457,N_8366,N_8206);
nand U8458 (N_8458,N_8233,N_8275);
and U8459 (N_8459,N_8270,N_8357);
nor U8460 (N_8460,N_8348,N_8324);
and U8461 (N_8461,N_8276,N_8295);
xor U8462 (N_8462,N_8332,N_8220);
and U8463 (N_8463,N_8343,N_8200);
xnor U8464 (N_8464,N_8282,N_8274);
or U8465 (N_8465,N_8224,N_8294);
xor U8466 (N_8466,N_8267,N_8244);
xor U8467 (N_8467,N_8297,N_8284);
or U8468 (N_8468,N_8278,N_8335);
or U8469 (N_8469,N_8213,N_8229);
nor U8470 (N_8470,N_8230,N_8336);
nor U8471 (N_8471,N_8285,N_8245);
nand U8472 (N_8472,N_8341,N_8338);
nor U8473 (N_8473,N_8247,N_8392);
nand U8474 (N_8474,N_8319,N_8370);
nand U8475 (N_8475,N_8390,N_8398);
or U8476 (N_8476,N_8279,N_8292);
or U8477 (N_8477,N_8303,N_8293);
nor U8478 (N_8478,N_8288,N_8329);
and U8479 (N_8479,N_8381,N_8310);
xnor U8480 (N_8480,N_8391,N_8219);
xor U8481 (N_8481,N_8394,N_8261);
or U8482 (N_8482,N_8375,N_8250);
nor U8483 (N_8483,N_8234,N_8209);
nand U8484 (N_8484,N_8312,N_8222);
nor U8485 (N_8485,N_8399,N_8337);
or U8486 (N_8486,N_8307,N_8304);
xor U8487 (N_8487,N_8212,N_8217);
and U8488 (N_8488,N_8262,N_8354);
nand U8489 (N_8489,N_8258,N_8238);
and U8490 (N_8490,N_8321,N_8236);
and U8491 (N_8491,N_8286,N_8356);
xor U8492 (N_8492,N_8225,N_8313);
and U8493 (N_8493,N_8242,N_8239);
nor U8494 (N_8494,N_8328,N_8208);
or U8495 (N_8495,N_8372,N_8283);
nand U8496 (N_8496,N_8376,N_8346);
and U8497 (N_8497,N_8365,N_8361);
xnor U8498 (N_8498,N_8257,N_8333);
nor U8499 (N_8499,N_8316,N_8393);
nand U8500 (N_8500,N_8228,N_8395);
or U8501 (N_8501,N_8318,N_8297);
xnor U8502 (N_8502,N_8363,N_8269);
xor U8503 (N_8503,N_8373,N_8272);
or U8504 (N_8504,N_8243,N_8357);
nor U8505 (N_8505,N_8377,N_8356);
xnor U8506 (N_8506,N_8222,N_8369);
xor U8507 (N_8507,N_8251,N_8256);
nor U8508 (N_8508,N_8271,N_8345);
and U8509 (N_8509,N_8270,N_8217);
nor U8510 (N_8510,N_8277,N_8282);
nand U8511 (N_8511,N_8260,N_8340);
xnor U8512 (N_8512,N_8329,N_8255);
and U8513 (N_8513,N_8225,N_8241);
nand U8514 (N_8514,N_8305,N_8383);
and U8515 (N_8515,N_8214,N_8372);
and U8516 (N_8516,N_8369,N_8378);
xnor U8517 (N_8517,N_8247,N_8330);
nor U8518 (N_8518,N_8387,N_8277);
or U8519 (N_8519,N_8258,N_8257);
and U8520 (N_8520,N_8229,N_8310);
nand U8521 (N_8521,N_8275,N_8355);
xor U8522 (N_8522,N_8380,N_8259);
nor U8523 (N_8523,N_8321,N_8314);
nor U8524 (N_8524,N_8252,N_8306);
nand U8525 (N_8525,N_8259,N_8244);
or U8526 (N_8526,N_8376,N_8291);
or U8527 (N_8527,N_8330,N_8381);
and U8528 (N_8528,N_8317,N_8312);
and U8529 (N_8529,N_8218,N_8255);
nor U8530 (N_8530,N_8222,N_8340);
nand U8531 (N_8531,N_8395,N_8331);
and U8532 (N_8532,N_8264,N_8306);
nand U8533 (N_8533,N_8321,N_8292);
nand U8534 (N_8534,N_8259,N_8257);
and U8535 (N_8535,N_8246,N_8339);
nor U8536 (N_8536,N_8241,N_8313);
nor U8537 (N_8537,N_8372,N_8391);
nand U8538 (N_8538,N_8226,N_8348);
nor U8539 (N_8539,N_8224,N_8350);
nand U8540 (N_8540,N_8302,N_8272);
nand U8541 (N_8541,N_8376,N_8279);
nor U8542 (N_8542,N_8266,N_8339);
nor U8543 (N_8543,N_8385,N_8208);
xnor U8544 (N_8544,N_8239,N_8240);
nor U8545 (N_8545,N_8266,N_8382);
or U8546 (N_8546,N_8269,N_8337);
or U8547 (N_8547,N_8316,N_8295);
and U8548 (N_8548,N_8373,N_8307);
and U8549 (N_8549,N_8253,N_8302);
or U8550 (N_8550,N_8280,N_8341);
nand U8551 (N_8551,N_8306,N_8362);
nor U8552 (N_8552,N_8247,N_8274);
nor U8553 (N_8553,N_8300,N_8309);
nand U8554 (N_8554,N_8342,N_8253);
nand U8555 (N_8555,N_8207,N_8316);
nor U8556 (N_8556,N_8255,N_8369);
nor U8557 (N_8557,N_8356,N_8310);
and U8558 (N_8558,N_8245,N_8372);
xnor U8559 (N_8559,N_8272,N_8300);
nor U8560 (N_8560,N_8375,N_8354);
and U8561 (N_8561,N_8363,N_8381);
xnor U8562 (N_8562,N_8347,N_8311);
nand U8563 (N_8563,N_8321,N_8279);
nand U8564 (N_8564,N_8222,N_8350);
and U8565 (N_8565,N_8335,N_8377);
or U8566 (N_8566,N_8332,N_8280);
nor U8567 (N_8567,N_8345,N_8272);
nor U8568 (N_8568,N_8276,N_8247);
nor U8569 (N_8569,N_8286,N_8219);
nor U8570 (N_8570,N_8297,N_8237);
xor U8571 (N_8571,N_8213,N_8274);
nor U8572 (N_8572,N_8294,N_8295);
and U8573 (N_8573,N_8202,N_8308);
or U8574 (N_8574,N_8207,N_8337);
and U8575 (N_8575,N_8206,N_8222);
and U8576 (N_8576,N_8258,N_8324);
or U8577 (N_8577,N_8371,N_8201);
nand U8578 (N_8578,N_8265,N_8263);
nor U8579 (N_8579,N_8300,N_8203);
and U8580 (N_8580,N_8244,N_8390);
and U8581 (N_8581,N_8330,N_8366);
or U8582 (N_8582,N_8233,N_8289);
and U8583 (N_8583,N_8261,N_8205);
or U8584 (N_8584,N_8280,N_8334);
xor U8585 (N_8585,N_8379,N_8347);
nand U8586 (N_8586,N_8331,N_8369);
xnor U8587 (N_8587,N_8280,N_8360);
and U8588 (N_8588,N_8324,N_8305);
nor U8589 (N_8589,N_8333,N_8230);
or U8590 (N_8590,N_8252,N_8282);
xnor U8591 (N_8591,N_8229,N_8328);
xor U8592 (N_8592,N_8380,N_8280);
and U8593 (N_8593,N_8277,N_8304);
and U8594 (N_8594,N_8291,N_8270);
xnor U8595 (N_8595,N_8323,N_8372);
nor U8596 (N_8596,N_8208,N_8389);
xnor U8597 (N_8597,N_8326,N_8201);
nand U8598 (N_8598,N_8369,N_8337);
or U8599 (N_8599,N_8268,N_8221);
xnor U8600 (N_8600,N_8467,N_8435);
nor U8601 (N_8601,N_8520,N_8584);
nand U8602 (N_8602,N_8599,N_8555);
xnor U8603 (N_8603,N_8511,N_8585);
and U8604 (N_8604,N_8544,N_8439);
or U8605 (N_8605,N_8589,N_8592);
and U8606 (N_8606,N_8494,N_8515);
and U8607 (N_8607,N_8455,N_8593);
nand U8608 (N_8608,N_8441,N_8510);
nand U8609 (N_8609,N_8521,N_8597);
and U8610 (N_8610,N_8537,N_8533);
nand U8611 (N_8611,N_8519,N_8575);
xnor U8612 (N_8612,N_8493,N_8424);
nand U8613 (N_8613,N_8480,N_8432);
and U8614 (N_8614,N_8508,N_8417);
or U8615 (N_8615,N_8440,N_8560);
xnor U8616 (N_8616,N_8498,N_8530);
or U8617 (N_8617,N_8454,N_8596);
and U8618 (N_8618,N_8576,N_8431);
nand U8619 (N_8619,N_8578,N_8484);
xnor U8620 (N_8620,N_8542,N_8425);
or U8621 (N_8621,N_8472,N_8583);
nor U8622 (N_8622,N_8476,N_8556);
and U8623 (N_8623,N_8554,N_8577);
and U8624 (N_8624,N_8500,N_8571);
nor U8625 (N_8625,N_8569,N_8489);
and U8626 (N_8626,N_8504,N_8461);
nor U8627 (N_8627,N_8485,N_8551);
or U8628 (N_8628,N_8595,N_8526);
or U8629 (N_8629,N_8513,N_8409);
nor U8630 (N_8630,N_8470,N_8558);
nor U8631 (N_8631,N_8548,N_8525);
and U8632 (N_8632,N_8502,N_8453);
nor U8633 (N_8633,N_8539,N_8549);
nor U8634 (N_8634,N_8570,N_8414);
or U8635 (N_8635,N_8403,N_8567);
and U8636 (N_8636,N_8437,N_8450);
and U8637 (N_8637,N_8566,N_8535);
or U8638 (N_8638,N_8449,N_8443);
xor U8639 (N_8639,N_8562,N_8402);
nand U8640 (N_8640,N_8457,N_8456);
or U8641 (N_8641,N_8499,N_8479);
and U8642 (N_8642,N_8400,N_8422);
nor U8643 (N_8643,N_8475,N_8557);
nor U8644 (N_8644,N_8572,N_8547);
nand U8645 (N_8645,N_8464,N_8404);
nor U8646 (N_8646,N_8574,N_8447);
nand U8647 (N_8647,N_8546,N_8451);
and U8648 (N_8648,N_8445,N_8471);
and U8649 (N_8649,N_8419,N_8591);
nor U8650 (N_8650,N_8468,N_8401);
xnor U8651 (N_8651,N_8408,N_8509);
nand U8652 (N_8652,N_8411,N_8466);
nor U8653 (N_8653,N_8568,N_8421);
nand U8654 (N_8654,N_8415,N_8407);
and U8655 (N_8655,N_8459,N_8405);
nor U8656 (N_8656,N_8488,N_8523);
and U8657 (N_8657,N_8434,N_8590);
nand U8658 (N_8658,N_8506,N_8522);
or U8659 (N_8659,N_8543,N_8473);
nand U8660 (N_8660,N_8426,N_8478);
nand U8661 (N_8661,N_8512,N_8586);
nand U8662 (N_8662,N_8448,N_8532);
nand U8663 (N_8663,N_8527,N_8507);
nor U8664 (N_8664,N_8433,N_8452);
nor U8665 (N_8665,N_8469,N_8550);
xor U8666 (N_8666,N_8430,N_8413);
xnor U8667 (N_8667,N_8580,N_8517);
xnor U8668 (N_8668,N_8458,N_8496);
or U8669 (N_8669,N_8444,N_8428);
xor U8670 (N_8670,N_8534,N_8477);
or U8671 (N_8671,N_8463,N_8462);
nor U8672 (N_8672,N_8505,N_8514);
nor U8673 (N_8673,N_8406,N_8516);
nor U8674 (N_8674,N_8474,N_8538);
nand U8675 (N_8675,N_8487,N_8518);
or U8676 (N_8676,N_8594,N_8492);
and U8677 (N_8677,N_8573,N_8503);
nor U8678 (N_8678,N_8531,N_8490);
nand U8679 (N_8679,N_8501,N_8418);
nand U8680 (N_8680,N_8540,N_8588);
nand U8681 (N_8681,N_8412,N_8524);
and U8682 (N_8682,N_8528,N_8565);
nor U8683 (N_8683,N_8495,N_8483);
nor U8684 (N_8684,N_8429,N_8581);
or U8685 (N_8685,N_8491,N_8438);
xnor U8686 (N_8686,N_8481,N_8436);
nand U8687 (N_8687,N_8563,N_8442);
xnor U8688 (N_8688,N_8553,N_8598);
nor U8689 (N_8689,N_8587,N_8486);
nor U8690 (N_8690,N_8545,N_8420);
or U8691 (N_8691,N_8536,N_8541);
nand U8692 (N_8692,N_8497,N_8427);
nand U8693 (N_8693,N_8465,N_8423);
nand U8694 (N_8694,N_8561,N_8446);
xnor U8695 (N_8695,N_8416,N_8410);
xor U8696 (N_8696,N_8579,N_8582);
and U8697 (N_8697,N_8564,N_8482);
nand U8698 (N_8698,N_8529,N_8460);
and U8699 (N_8699,N_8552,N_8559);
nor U8700 (N_8700,N_8483,N_8540);
or U8701 (N_8701,N_8510,N_8433);
and U8702 (N_8702,N_8514,N_8487);
xnor U8703 (N_8703,N_8494,N_8548);
nand U8704 (N_8704,N_8468,N_8598);
nor U8705 (N_8705,N_8502,N_8593);
nand U8706 (N_8706,N_8466,N_8468);
and U8707 (N_8707,N_8402,N_8596);
nor U8708 (N_8708,N_8454,N_8432);
xor U8709 (N_8709,N_8408,N_8438);
nand U8710 (N_8710,N_8410,N_8409);
xnor U8711 (N_8711,N_8519,N_8439);
and U8712 (N_8712,N_8555,N_8406);
nand U8713 (N_8713,N_8536,N_8511);
or U8714 (N_8714,N_8522,N_8412);
xor U8715 (N_8715,N_8442,N_8474);
nor U8716 (N_8716,N_8483,N_8484);
or U8717 (N_8717,N_8405,N_8594);
and U8718 (N_8718,N_8523,N_8560);
and U8719 (N_8719,N_8412,N_8509);
nand U8720 (N_8720,N_8436,N_8549);
nor U8721 (N_8721,N_8443,N_8439);
or U8722 (N_8722,N_8544,N_8570);
nor U8723 (N_8723,N_8500,N_8435);
nor U8724 (N_8724,N_8461,N_8456);
nor U8725 (N_8725,N_8566,N_8487);
and U8726 (N_8726,N_8471,N_8564);
or U8727 (N_8727,N_8578,N_8566);
and U8728 (N_8728,N_8491,N_8435);
xor U8729 (N_8729,N_8492,N_8583);
nand U8730 (N_8730,N_8591,N_8560);
and U8731 (N_8731,N_8573,N_8541);
and U8732 (N_8732,N_8574,N_8488);
nand U8733 (N_8733,N_8598,N_8457);
or U8734 (N_8734,N_8558,N_8468);
and U8735 (N_8735,N_8503,N_8540);
or U8736 (N_8736,N_8430,N_8488);
nor U8737 (N_8737,N_8574,N_8443);
xnor U8738 (N_8738,N_8413,N_8401);
nor U8739 (N_8739,N_8511,N_8526);
and U8740 (N_8740,N_8522,N_8469);
or U8741 (N_8741,N_8568,N_8562);
and U8742 (N_8742,N_8529,N_8587);
xor U8743 (N_8743,N_8465,N_8440);
xnor U8744 (N_8744,N_8525,N_8488);
nand U8745 (N_8745,N_8585,N_8594);
nor U8746 (N_8746,N_8590,N_8547);
and U8747 (N_8747,N_8481,N_8599);
nand U8748 (N_8748,N_8437,N_8456);
or U8749 (N_8749,N_8529,N_8425);
xor U8750 (N_8750,N_8484,N_8490);
nand U8751 (N_8751,N_8414,N_8447);
nor U8752 (N_8752,N_8499,N_8458);
or U8753 (N_8753,N_8555,N_8553);
nand U8754 (N_8754,N_8401,N_8432);
and U8755 (N_8755,N_8585,N_8452);
nor U8756 (N_8756,N_8553,N_8426);
nor U8757 (N_8757,N_8439,N_8558);
xor U8758 (N_8758,N_8434,N_8461);
xor U8759 (N_8759,N_8589,N_8508);
nand U8760 (N_8760,N_8559,N_8476);
or U8761 (N_8761,N_8507,N_8474);
nand U8762 (N_8762,N_8449,N_8540);
and U8763 (N_8763,N_8515,N_8572);
or U8764 (N_8764,N_8565,N_8470);
xnor U8765 (N_8765,N_8502,N_8478);
xnor U8766 (N_8766,N_8485,N_8534);
nand U8767 (N_8767,N_8509,N_8517);
xor U8768 (N_8768,N_8539,N_8520);
xor U8769 (N_8769,N_8585,N_8534);
and U8770 (N_8770,N_8456,N_8446);
and U8771 (N_8771,N_8450,N_8550);
and U8772 (N_8772,N_8565,N_8424);
or U8773 (N_8773,N_8449,N_8500);
or U8774 (N_8774,N_8524,N_8556);
nor U8775 (N_8775,N_8551,N_8483);
or U8776 (N_8776,N_8430,N_8417);
xor U8777 (N_8777,N_8545,N_8583);
nand U8778 (N_8778,N_8434,N_8446);
and U8779 (N_8779,N_8499,N_8403);
and U8780 (N_8780,N_8584,N_8424);
nand U8781 (N_8781,N_8444,N_8568);
xnor U8782 (N_8782,N_8434,N_8453);
nor U8783 (N_8783,N_8550,N_8439);
nand U8784 (N_8784,N_8547,N_8583);
or U8785 (N_8785,N_8581,N_8411);
and U8786 (N_8786,N_8493,N_8492);
and U8787 (N_8787,N_8520,N_8435);
nor U8788 (N_8788,N_8489,N_8508);
xor U8789 (N_8789,N_8594,N_8468);
and U8790 (N_8790,N_8589,N_8404);
xor U8791 (N_8791,N_8441,N_8451);
or U8792 (N_8792,N_8488,N_8591);
xor U8793 (N_8793,N_8563,N_8430);
and U8794 (N_8794,N_8531,N_8405);
nand U8795 (N_8795,N_8474,N_8457);
nand U8796 (N_8796,N_8529,N_8504);
xor U8797 (N_8797,N_8411,N_8588);
xor U8798 (N_8798,N_8401,N_8595);
or U8799 (N_8799,N_8410,N_8554);
nor U8800 (N_8800,N_8628,N_8757);
nand U8801 (N_8801,N_8799,N_8752);
nand U8802 (N_8802,N_8655,N_8649);
xnor U8803 (N_8803,N_8723,N_8770);
nand U8804 (N_8804,N_8724,N_8766);
nor U8805 (N_8805,N_8636,N_8678);
nand U8806 (N_8806,N_8755,N_8746);
nor U8807 (N_8807,N_8781,N_8753);
nor U8808 (N_8808,N_8730,N_8660);
or U8809 (N_8809,N_8713,N_8677);
nor U8810 (N_8810,N_8710,N_8676);
or U8811 (N_8811,N_8788,N_8773);
and U8812 (N_8812,N_8643,N_8768);
and U8813 (N_8813,N_8789,N_8620);
or U8814 (N_8814,N_8740,N_8637);
xnor U8815 (N_8815,N_8756,N_8646);
nand U8816 (N_8816,N_8604,N_8701);
nand U8817 (N_8817,N_8691,N_8612);
and U8818 (N_8818,N_8661,N_8619);
and U8819 (N_8819,N_8771,N_8689);
nand U8820 (N_8820,N_8682,N_8671);
nor U8821 (N_8821,N_8745,N_8674);
or U8822 (N_8822,N_8725,N_8670);
and U8823 (N_8823,N_8606,N_8785);
nand U8824 (N_8824,N_8647,N_8605);
xnor U8825 (N_8825,N_8632,N_8721);
xor U8826 (N_8826,N_8717,N_8737);
or U8827 (N_8827,N_8615,N_8623);
xnor U8828 (N_8828,N_8754,N_8614);
or U8829 (N_8829,N_8783,N_8607);
xor U8830 (N_8830,N_8767,N_8727);
xnor U8831 (N_8831,N_8625,N_8711);
or U8832 (N_8832,N_8720,N_8673);
or U8833 (N_8833,N_8797,N_8790);
and U8834 (N_8834,N_8787,N_8715);
nor U8835 (N_8835,N_8616,N_8657);
and U8836 (N_8836,N_8610,N_8683);
nand U8837 (N_8837,N_8778,N_8690);
nand U8838 (N_8838,N_8656,N_8716);
nand U8839 (N_8839,N_8784,N_8618);
and U8840 (N_8840,N_8700,N_8705);
xnor U8841 (N_8841,N_8658,N_8780);
and U8842 (N_8842,N_8654,N_8749);
nand U8843 (N_8843,N_8622,N_8760);
or U8844 (N_8844,N_8776,N_8732);
nand U8845 (N_8845,N_8793,N_8751);
or U8846 (N_8846,N_8762,N_8731);
or U8847 (N_8847,N_8764,N_8617);
or U8848 (N_8848,N_8719,N_8791);
nor U8849 (N_8849,N_8664,N_8796);
or U8850 (N_8850,N_8692,N_8663);
or U8851 (N_8851,N_8712,N_8686);
nor U8852 (N_8852,N_8786,N_8679);
or U8853 (N_8853,N_8621,N_8726);
and U8854 (N_8854,N_8699,N_8665);
nand U8855 (N_8855,N_8667,N_8627);
nand U8856 (N_8856,N_8693,N_8645);
nand U8857 (N_8857,N_8769,N_8792);
or U8858 (N_8858,N_8688,N_8659);
nor U8859 (N_8859,N_8696,N_8662);
nor U8860 (N_8860,N_8794,N_8702);
nand U8861 (N_8861,N_8736,N_8704);
nor U8862 (N_8862,N_8774,N_8666);
or U8863 (N_8863,N_8772,N_8765);
and U8864 (N_8864,N_8633,N_8652);
nand U8865 (N_8865,N_8668,N_8718);
xnor U8866 (N_8866,N_8669,N_8608);
nor U8867 (N_8867,N_8775,N_8758);
and U8868 (N_8868,N_8680,N_8644);
and U8869 (N_8869,N_8624,N_8798);
nor U8870 (N_8870,N_8747,N_8782);
or U8871 (N_8871,N_8739,N_8707);
and U8872 (N_8872,N_8687,N_8703);
nand U8873 (N_8873,N_8629,N_8734);
nor U8874 (N_8874,N_8603,N_8735);
nand U8875 (N_8875,N_8706,N_8613);
nand U8876 (N_8876,N_8635,N_8714);
nand U8877 (N_8877,N_8777,N_8729);
xor U8878 (N_8878,N_8602,N_8759);
and U8879 (N_8879,N_8742,N_8638);
and U8880 (N_8880,N_8795,N_8601);
and U8881 (N_8881,N_8641,N_8651);
or U8882 (N_8882,N_8748,N_8631);
and U8883 (N_8883,N_8698,N_8763);
nand U8884 (N_8884,N_8695,N_8733);
nand U8885 (N_8885,N_8684,N_8709);
and U8886 (N_8886,N_8750,N_8728);
and U8887 (N_8887,N_8653,N_8685);
nand U8888 (N_8888,N_8743,N_8761);
xor U8889 (N_8889,N_8642,N_8639);
and U8890 (N_8890,N_8744,N_8650);
nor U8891 (N_8891,N_8738,N_8675);
or U8892 (N_8892,N_8634,N_8609);
or U8893 (N_8893,N_8741,N_8630);
xnor U8894 (N_8894,N_8648,N_8672);
nand U8895 (N_8895,N_8626,N_8640);
nor U8896 (N_8896,N_8611,N_8681);
and U8897 (N_8897,N_8708,N_8694);
nand U8898 (N_8898,N_8697,N_8600);
or U8899 (N_8899,N_8779,N_8722);
nor U8900 (N_8900,N_8702,N_8745);
xnor U8901 (N_8901,N_8748,N_8679);
nand U8902 (N_8902,N_8676,N_8629);
nand U8903 (N_8903,N_8611,N_8685);
nand U8904 (N_8904,N_8665,N_8646);
and U8905 (N_8905,N_8608,N_8745);
xor U8906 (N_8906,N_8616,N_8753);
nor U8907 (N_8907,N_8652,N_8715);
nor U8908 (N_8908,N_8768,N_8699);
or U8909 (N_8909,N_8775,N_8798);
xnor U8910 (N_8910,N_8608,N_8792);
or U8911 (N_8911,N_8612,N_8683);
and U8912 (N_8912,N_8631,N_8693);
xnor U8913 (N_8913,N_8745,N_8701);
xor U8914 (N_8914,N_8795,N_8787);
or U8915 (N_8915,N_8738,N_8603);
or U8916 (N_8916,N_8650,N_8646);
nor U8917 (N_8917,N_8675,N_8760);
nor U8918 (N_8918,N_8604,N_8626);
nand U8919 (N_8919,N_8703,N_8616);
or U8920 (N_8920,N_8773,N_8689);
or U8921 (N_8921,N_8702,N_8792);
or U8922 (N_8922,N_8687,N_8753);
nand U8923 (N_8923,N_8712,N_8744);
and U8924 (N_8924,N_8665,N_8617);
nand U8925 (N_8925,N_8679,N_8757);
xnor U8926 (N_8926,N_8755,N_8617);
nor U8927 (N_8927,N_8696,N_8618);
xnor U8928 (N_8928,N_8653,N_8762);
or U8929 (N_8929,N_8717,N_8799);
nor U8930 (N_8930,N_8655,N_8779);
or U8931 (N_8931,N_8652,N_8667);
xor U8932 (N_8932,N_8789,N_8616);
nor U8933 (N_8933,N_8793,N_8726);
or U8934 (N_8934,N_8781,N_8682);
nor U8935 (N_8935,N_8786,N_8686);
and U8936 (N_8936,N_8649,N_8605);
nand U8937 (N_8937,N_8712,N_8604);
and U8938 (N_8938,N_8701,N_8733);
nand U8939 (N_8939,N_8743,N_8630);
nand U8940 (N_8940,N_8649,N_8793);
or U8941 (N_8941,N_8792,N_8651);
nor U8942 (N_8942,N_8683,N_8777);
or U8943 (N_8943,N_8739,N_8776);
or U8944 (N_8944,N_8662,N_8622);
or U8945 (N_8945,N_8660,N_8640);
and U8946 (N_8946,N_8763,N_8767);
or U8947 (N_8947,N_8703,N_8635);
or U8948 (N_8948,N_8707,N_8614);
nor U8949 (N_8949,N_8665,N_8623);
xnor U8950 (N_8950,N_8753,N_8644);
xnor U8951 (N_8951,N_8730,N_8695);
or U8952 (N_8952,N_8629,N_8721);
xor U8953 (N_8953,N_8656,N_8774);
nor U8954 (N_8954,N_8680,N_8726);
nand U8955 (N_8955,N_8735,N_8653);
xor U8956 (N_8956,N_8680,N_8651);
nor U8957 (N_8957,N_8762,N_8716);
nor U8958 (N_8958,N_8695,N_8785);
or U8959 (N_8959,N_8681,N_8676);
and U8960 (N_8960,N_8700,N_8797);
nor U8961 (N_8961,N_8733,N_8739);
xor U8962 (N_8962,N_8664,N_8716);
and U8963 (N_8963,N_8667,N_8752);
and U8964 (N_8964,N_8739,N_8758);
or U8965 (N_8965,N_8769,N_8736);
nor U8966 (N_8966,N_8753,N_8743);
or U8967 (N_8967,N_8641,N_8646);
xnor U8968 (N_8968,N_8700,N_8641);
nand U8969 (N_8969,N_8619,N_8718);
nand U8970 (N_8970,N_8764,N_8781);
and U8971 (N_8971,N_8614,N_8787);
or U8972 (N_8972,N_8680,N_8676);
nor U8973 (N_8973,N_8704,N_8721);
and U8974 (N_8974,N_8742,N_8665);
and U8975 (N_8975,N_8680,N_8642);
nand U8976 (N_8976,N_8713,N_8755);
or U8977 (N_8977,N_8706,N_8612);
or U8978 (N_8978,N_8625,N_8632);
or U8979 (N_8979,N_8732,N_8633);
xnor U8980 (N_8980,N_8681,N_8679);
nor U8981 (N_8981,N_8780,N_8678);
or U8982 (N_8982,N_8747,N_8670);
xor U8983 (N_8983,N_8719,N_8610);
or U8984 (N_8984,N_8786,N_8727);
or U8985 (N_8985,N_8739,N_8712);
or U8986 (N_8986,N_8702,N_8632);
nand U8987 (N_8987,N_8686,N_8608);
or U8988 (N_8988,N_8626,N_8723);
nor U8989 (N_8989,N_8782,N_8660);
nand U8990 (N_8990,N_8726,N_8601);
or U8991 (N_8991,N_8602,N_8774);
nand U8992 (N_8992,N_8777,N_8733);
and U8993 (N_8993,N_8666,N_8739);
xor U8994 (N_8994,N_8775,N_8778);
nor U8995 (N_8995,N_8740,N_8639);
nor U8996 (N_8996,N_8692,N_8713);
and U8997 (N_8997,N_8603,N_8628);
or U8998 (N_8998,N_8673,N_8668);
nand U8999 (N_8999,N_8609,N_8635);
and U9000 (N_9000,N_8861,N_8839);
nor U9001 (N_9001,N_8844,N_8826);
and U9002 (N_9002,N_8925,N_8917);
xnor U9003 (N_9003,N_8879,N_8910);
and U9004 (N_9004,N_8843,N_8885);
nor U9005 (N_9005,N_8968,N_8828);
nand U9006 (N_9006,N_8813,N_8810);
and U9007 (N_9007,N_8852,N_8963);
xor U9008 (N_9008,N_8833,N_8881);
and U9009 (N_9009,N_8829,N_8937);
and U9010 (N_9010,N_8857,N_8827);
or U9011 (N_9011,N_8883,N_8987);
xor U9012 (N_9012,N_8996,N_8904);
xor U9013 (N_9013,N_8892,N_8915);
xnor U9014 (N_9014,N_8805,N_8990);
or U9015 (N_9015,N_8891,N_8938);
and U9016 (N_9016,N_8919,N_8967);
nor U9017 (N_9017,N_8821,N_8934);
nor U9018 (N_9018,N_8897,N_8901);
nand U9019 (N_9019,N_8809,N_8842);
and U9020 (N_9020,N_8802,N_8835);
xnor U9021 (N_9021,N_8939,N_8847);
xnor U9022 (N_9022,N_8804,N_8929);
xor U9023 (N_9023,N_8999,N_8877);
xor U9024 (N_9024,N_8927,N_8888);
or U9025 (N_9025,N_8903,N_8880);
xnor U9026 (N_9026,N_8923,N_8900);
or U9027 (N_9027,N_8922,N_8986);
and U9028 (N_9028,N_8928,N_8875);
xor U9029 (N_9029,N_8921,N_8882);
nand U9030 (N_9030,N_8871,N_8906);
or U9031 (N_9031,N_8859,N_8893);
and U9032 (N_9032,N_8898,N_8840);
xor U9033 (N_9033,N_8812,N_8918);
and U9034 (N_9034,N_8824,N_8962);
xor U9035 (N_9035,N_8936,N_8869);
nor U9036 (N_9036,N_8801,N_8907);
and U9037 (N_9037,N_8974,N_8931);
nand U9038 (N_9038,N_8849,N_8819);
and U9039 (N_9039,N_8911,N_8887);
or U9040 (N_9040,N_8855,N_8932);
xor U9041 (N_9041,N_8993,N_8834);
or U9042 (N_9042,N_8912,N_8832);
or U9043 (N_9043,N_8961,N_8863);
nand U9044 (N_9044,N_8853,N_8817);
or U9045 (N_9045,N_8965,N_8814);
and U9046 (N_9046,N_8825,N_8924);
nand U9047 (N_9047,N_8926,N_8933);
xor U9048 (N_9048,N_8960,N_8867);
nand U9049 (N_9049,N_8822,N_8908);
nor U9050 (N_9050,N_8808,N_8920);
nand U9051 (N_9051,N_8896,N_8966);
nor U9052 (N_9052,N_8860,N_8868);
nor U9053 (N_9053,N_8950,N_8872);
or U9054 (N_9054,N_8816,N_8820);
and U9055 (N_9055,N_8970,N_8976);
xor U9056 (N_9056,N_8935,N_8989);
and U9057 (N_9057,N_8981,N_8815);
nor U9058 (N_9058,N_8955,N_8971);
or U9059 (N_9059,N_8941,N_8947);
xnor U9060 (N_9060,N_8975,N_8876);
nor U9061 (N_9061,N_8982,N_8836);
or U9062 (N_9062,N_8983,N_8985);
xor U9063 (N_9063,N_8862,N_8914);
and U9064 (N_9064,N_8980,N_8988);
or U9065 (N_9065,N_8818,N_8838);
and U9066 (N_9066,N_8811,N_8972);
nand U9067 (N_9067,N_8823,N_8856);
xor U9068 (N_9068,N_8991,N_8830);
or U9069 (N_9069,N_8884,N_8978);
or U9070 (N_9070,N_8948,N_8984);
nor U9071 (N_9071,N_8951,N_8916);
nor U9072 (N_9072,N_8895,N_8850);
xnor U9073 (N_9073,N_8865,N_8952);
nor U9074 (N_9074,N_8930,N_8889);
nor U9075 (N_9075,N_8949,N_8913);
or U9076 (N_9076,N_8994,N_8886);
and U9077 (N_9077,N_8992,N_8846);
and U9078 (N_9078,N_8954,N_8958);
nor U9079 (N_9079,N_8969,N_8848);
and U9080 (N_9080,N_8870,N_8806);
xnor U9081 (N_9081,N_8998,N_8902);
xor U9082 (N_9082,N_8864,N_8878);
xnor U9083 (N_9083,N_8803,N_8837);
nor U9084 (N_9084,N_8873,N_8874);
xnor U9085 (N_9085,N_8854,N_8942);
nor U9086 (N_9086,N_8800,N_8909);
and U9087 (N_9087,N_8957,N_8940);
nand U9088 (N_9088,N_8807,N_8905);
nor U9089 (N_9089,N_8851,N_8977);
xnor U9090 (N_9090,N_8866,N_8845);
nor U9091 (N_9091,N_8943,N_8959);
nor U9092 (N_9092,N_8944,N_8841);
and U9093 (N_9093,N_8956,N_8995);
nand U9094 (N_9094,N_8953,N_8858);
xor U9095 (N_9095,N_8997,N_8831);
and U9096 (N_9096,N_8899,N_8894);
or U9097 (N_9097,N_8946,N_8890);
and U9098 (N_9098,N_8964,N_8979);
nor U9099 (N_9099,N_8945,N_8973);
nor U9100 (N_9100,N_8973,N_8880);
nand U9101 (N_9101,N_8915,N_8904);
or U9102 (N_9102,N_8880,N_8935);
nor U9103 (N_9103,N_8992,N_8950);
and U9104 (N_9104,N_8835,N_8940);
nor U9105 (N_9105,N_8887,N_8821);
xor U9106 (N_9106,N_8831,N_8994);
nand U9107 (N_9107,N_8966,N_8852);
nand U9108 (N_9108,N_8930,N_8834);
xnor U9109 (N_9109,N_8971,N_8843);
or U9110 (N_9110,N_8970,N_8804);
nor U9111 (N_9111,N_8864,N_8914);
nand U9112 (N_9112,N_8935,N_8905);
or U9113 (N_9113,N_8823,N_8916);
nand U9114 (N_9114,N_8986,N_8976);
xor U9115 (N_9115,N_8893,N_8895);
and U9116 (N_9116,N_8960,N_8918);
xnor U9117 (N_9117,N_8973,N_8932);
nor U9118 (N_9118,N_8896,N_8937);
nand U9119 (N_9119,N_8824,N_8837);
and U9120 (N_9120,N_8879,N_8828);
nand U9121 (N_9121,N_8829,N_8943);
or U9122 (N_9122,N_8900,N_8964);
or U9123 (N_9123,N_8820,N_8967);
nand U9124 (N_9124,N_8874,N_8911);
or U9125 (N_9125,N_8967,N_8957);
nand U9126 (N_9126,N_8832,N_8959);
xor U9127 (N_9127,N_8899,N_8923);
nand U9128 (N_9128,N_8810,N_8883);
nor U9129 (N_9129,N_8914,N_8804);
nor U9130 (N_9130,N_8824,N_8870);
nor U9131 (N_9131,N_8827,N_8972);
or U9132 (N_9132,N_8819,N_8898);
xnor U9133 (N_9133,N_8906,N_8982);
nor U9134 (N_9134,N_8918,N_8995);
xnor U9135 (N_9135,N_8838,N_8866);
and U9136 (N_9136,N_8817,N_8828);
or U9137 (N_9137,N_8843,N_8921);
nand U9138 (N_9138,N_8877,N_8928);
or U9139 (N_9139,N_8924,N_8885);
nor U9140 (N_9140,N_8938,N_8930);
nand U9141 (N_9141,N_8894,N_8829);
and U9142 (N_9142,N_8910,N_8812);
and U9143 (N_9143,N_8817,N_8998);
or U9144 (N_9144,N_8945,N_8830);
nor U9145 (N_9145,N_8972,N_8809);
nand U9146 (N_9146,N_8817,N_8905);
nand U9147 (N_9147,N_8995,N_8943);
and U9148 (N_9148,N_8873,N_8955);
nor U9149 (N_9149,N_8921,N_8811);
nand U9150 (N_9150,N_8964,N_8883);
xor U9151 (N_9151,N_8923,N_8971);
or U9152 (N_9152,N_8969,N_8883);
xnor U9153 (N_9153,N_8887,N_8860);
nand U9154 (N_9154,N_8886,N_8813);
xnor U9155 (N_9155,N_8837,N_8880);
and U9156 (N_9156,N_8907,N_8920);
nand U9157 (N_9157,N_8891,N_8822);
nand U9158 (N_9158,N_8976,N_8820);
or U9159 (N_9159,N_8939,N_8957);
xor U9160 (N_9160,N_8942,N_8856);
xnor U9161 (N_9161,N_8988,N_8927);
and U9162 (N_9162,N_8974,N_8989);
and U9163 (N_9163,N_8968,N_8985);
nor U9164 (N_9164,N_8933,N_8943);
nor U9165 (N_9165,N_8820,N_8803);
and U9166 (N_9166,N_8909,N_8828);
nand U9167 (N_9167,N_8970,N_8913);
xor U9168 (N_9168,N_8983,N_8972);
and U9169 (N_9169,N_8819,N_8802);
or U9170 (N_9170,N_8805,N_8819);
nand U9171 (N_9171,N_8894,N_8955);
xnor U9172 (N_9172,N_8948,N_8957);
nand U9173 (N_9173,N_8871,N_8966);
and U9174 (N_9174,N_8844,N_8800);
or U9175 (N_9175,N_8929,N_8829);
nand U9176 (N_9176,N_8809,N_8818);
and U9177 (N_9177,N_8913,N_8897);
and U9178 (N_9178,N_8862,N_8919);
xnor U9179 (N_9179,N_8964,N_8922);
nor U9180 (N_9180,N_8820,N_8977);
and U9181 (N_9181,N_8897,N_8814);
and U9182 (N_9182,N_8856,N_8968);
xnor U9183 (N_9183,N_8975,N_8823);
nor U9184 (N_9184,N_8991,N_8847);
or U9185 (N_9185,N_8871,N_8965);
nor U9186 (N_9186,N_8851,N_8879);
or U9187 (N_9187,N_8807,N_8963);
nand U9188 (N_9188,N_8950,N_8890);
nor U9189 (N_9189,N_8925,N_8941);
nor U9190 (N_9190,N_8880,N_8835);
or U9191 (N_9191,N_8920,N_8941);
nor U9192 (N_9192,N_8853,N_8887);
nor U9193 (N_9193,N_8976,N_8988);
and U9194 (N_9194,N_8804,N_8936);
or U9195 (N_9195,N_8867,N_8850);
nor U9196 (N_9196,N_8920,N_8992);
or U9197 (N_9197,N_8837,N_8828);
nand U9198 (N_9198,N_8859,N_8934);
or U9199 (N_9199,N_8989,N_8880);
and U9200 (N_9200,N_9012,N_9147);
and U9201 (N_9201,N_9047,N_9176);
nor U9202 (N_9202,N_9057,N_9075);
and U9203 (N_9203,N_9008,N_9197);
xnor U9204 (N_9204,N_9127,N_9090);
xor U9205 (N_9205,N_9000,N_9113);
nor U9206 (N_9206,N_9096,N_9097);
xor U9207 (N_9207,N_9038,N_9188);
nor U9208 (N_9208,N_9148,N_9083);
or U9209 (N_9209,N_9140,N_9035);
or U9210 (N_9210,N_9126,N_9061);
nor U9211 (N_9211,N_9021,N_9106);
or U9212 (N_9212,N_9016,N_9013);
nand U9213 (N_9213,N_9002,N_9175);
nor U9214 (N_9214,N_9181,N_9018);
nor U9215 (N_9215,N_9064,N_9017);
nor U9216 (N_9216,N_9001,N_9019);
or U9217 (N_9217,N_9104,N_9062);
nor U9218 (N_9218,N_9132,N_9118);
nand U9219 (N_9219,N_9023,N_9063);
nand U9220 (N_9220,N_9009,N_9092);
or U9221 (N_9221,N_9117,N_9114);
nor U9222 (N_9222,N_9130,N_9120);
xnor U9223 (N_9223,N_9121,N_9003);
or U9224 (N_9224,N_9071,N_9004);
nor U9225 (N_9225,N_9025,N_9103);
nor U9226 (N_9226,N_9087,N_9081);
and U9227 (N_9227,N_9095,N_9189);
nand U9228 (N_9228,N_9053,N_9046);
and U9229 (N_9229,N_9073,N_9142);
nor U9230 (N_9230,N_9067,N_9159);
nand U9231 (N_9231,N_9033,N_9182);
xnor U9232 (N_9232,N_9169,N_9005);
nor U9233 (N_9233,N_9141,N_9187);
xnor U9234 (N_9234,N_9193,N_9089);
nand U9235 (N_9235,N_9167,N_9020);
xor U9236 (N_9236,N_9125,N_9022);
or U9237 (N_9237,N_9076,N_9010);
and U9238 (N_9238,N_9131,N_9174);
nor U9239 (N_9239,N_9093,N_9146);
and U9240 (N_9240,N_9162,N_9068);
or U9241 (N_9241,N_9007,N_9024);
and U9242 (N_9242,N_9031,N_9066);
or U9243 (N_9243,N_9065,N_9172);
xor U9244 (N_9244,N_9026,N_9136);
nor U9245 (N_9245,N_9108,N_9084);
nand U9246 (N_9246,N_9135,N_9178);
xor U9247 (N_9247,N_9014,N_9042);
and U9248 (N_9248,N_9006,N_9155);
xor U9249 (N_9249,N_9164,N_9185);
xnor U9250 (N_9250,N_9032,N_9105);
xor U9251 (N_9251,N_9166,N_9144);
nand U9252 (N_9252,N_9139,N_9054);
or U9253 (N_9253,N_9036,N_9128);
nor U9254 (N_9254,N_9098,N_9041);
xnor U9255 (N_9255,N_9133,N_9179);
and U9256 (N_9256,N_9111,N_9099);
or U9257 (N_9257,N_9186,N_9109);
xor U9258 (N_9258,N_9078,N_9088);
xnor U9259 (N_9259,N_9183,N_9143);
nand U9260 (N_9260,N_9170,N_9158);
xor U9261 (N_9261,N_9034,N_9198);
nand U9262 (N_9262,N_9137,N_9122);
nor U9263 (N_9263,N_9059,N_9079);
nand U9264 (N_9264,N_9196,N_9129);
xor U9265 (N_9265,N_9037,N_9191);
and U9266 (N_9266,N_9050,N_9151);
xor U9267 (N_9267,N_9040,N_9094);
nor U9268 (N_9268,N_9165,N_9157);
nor U9269 (N_9269,N_9154,N_9145);
nand U9270 (N_9270,N_9028,N_9058);
or U9271 (N_9271,N_9138,N_9051);
nor U9272 (N_9272,N_9056,N_9101);
or U9273 (N_9273,N_9091,N_9123);
nand U9274 (N_9274,N_9168,N_9150);
nand U9275 (N_9275,N_9015,N_9199);
nand U9276 (N_9276,N_9086,N_9027);
and U9277 (N_9277,N_9048,N_9011);
nand U9278 (N_9278,N_9119,N_9177);
nand U9279 (N_9279,N_9171,N_9072);
xnor U9280 (N_9280,N_9039,N_9161);
and U9281 (N_9281,N_9153,N_9030);
and U9282 (N_9282,N_9152,N_9190);
nor U9283 (N_9283,N_9070,N_9077);
or U9284 (N_9284,N_9156,N_9043);
xor U9285 (N_9285,N_9060,N_9192);
xor U9286 (N_9286,N_9085,N_9180);
nor U9287 (N_9287,N_9195,N_9029);
xnor U9288 (N_9288,N_9102,N_9134);
nor U9289 (N_9289,N_9184,N_9045);
nor U9290 (N_9290,N_9107,N_9124);
or U9291 (N_9291,N_9082,N_9163);
xor U9292 (N_9292,N_9044,N_9160);
and U9293 (N_9293,N_9074,N_9055);
or U9294 (N_9294,N_9049,N_9100);
or U9295 (N_9295,N_9110,N_9194);
or U9296 (N_9296,N_9112,N_9115);
xor U9297 (N_9297,N_9080,N_9149);
nand U9298 (N_9298,N_9052,N_9173);
nand U9299 (N_9299,N_9069,N_9116);
nand U9300 (N_9300,N_9029,N_9081);
or U9301 (N_9301,N_9164,N_9098);
nand U9302 (N_9302,N_9098,N_9043);
xor U9303 (N_9303,N_9180,N_9044);
nand U9304 (N_9304,N_9080,N_9014);
and U9305 (N_9305,N_9015,N_9008);
or U9306 (N_9306,N_9089,N_9080);
or U9307 (N_9307,N_9174,N_9180);
xnor U9308 (N_9308,N_9011,N_9106);
nor U9309 (N_9309,N_9150,N_9106);
nor U9310 (N_9310,N_9154,N_9136);
or U9311 (N_9311,N_9127,N_9117);
xor U9312 (N_9312,N_9185,N_9124);
or U9313 (N_9313,N_9149,N_9183);
nand U9314 (N_9314,N_9192,N_9115);
and U9315 (N_9315,N_9026,N_9071);
xor U9316 (N_9316,N_9103,N_9157);
nor U9317 (N_9317,N_9104,N_9018);
xor U9318 (N_9318,N_9071,N_9183);
or U9319 (N_9319,N_9128,N_9001);
nand U9320 (N_9320,N_9042,N_9142);
xnor U9321 (N_9321,N_9102,N_9145);
nor U9322 (N_9322,N_9078,N_9027);
xnor U9323 (N_9323,N_9166,N_9054);
nand U9324 (N_9324,N_9192,N_9017);
nand U9325 (N_9325,N_9125,N_9082);
or U9326 (N_9326,N_9142,N_9123);
xnor U9327 (N_9327,N_9136,N_9036);
xor U9328 (N_9328,N_9092,N_9172);
xnor U9329 (N_9329,N_9026,N_9062);
nor U9330 (N_9330,N_9142,N_9114);
xor U9331 (N_9331,N_9004,N_9140);
xnor U9332 (N_9332,N_9159,N_9112);
nor U9333 (N_9333,N_9025,N_9036);
nor U9334 (N_9334,N_9055,N_9146);
nand U9335 (N_9335,N_9116,N_9057);
and U9336 (N_9336,N_9138,N_9072);
nor U9337 (N_9337,N_9087,N_9167);
or U9338 (N_9338,N_9198,N_9109);
xnor U9339 (N_9339,N_9187,N_9064);
and U9340 (N_9340,N_9151,N_9063);
and U9341 (N_9341,N_9158,N_9180);
nand U9342 (N_9342,N_9070,N_9125);
nor U9343 (N_9343,N_9139,N_9170);
and U9344 (N_9344,N_9026,N_9012);
or U9345 (N_9345,N_9121,N_9057);
nor U9346 (N_9346,N_9113,N_9129);
or U9347 (N_9347,N_9031,N_9079);
or U9348 (N_9348,N_9162,N_9166);
nand U9349 (N_9349,N_9004,N_9141);
nor U9350 (N_9350,N_9115,N_9182);
and U9351 (N_9351,N_9058,N_9170);
xor U9352 (N_9352,N_9085,N_9069);
and U9353 (N_9353,N_9030,N_9123);
nor U9354 (N_9354,N_9077,N_9076);
nor U9355 (N_9355,N_9059,N_9075);
and U9356 (N_9356,N_9162,N_9026);
or U9357 (N_9357,N_9069,N_9199);
xor U9358 (N_9358,N_9139,N_9166);
or U9359 (N_9359,N_9184,N_9110);
xor U9360 (N_9360,N_9037,N_9095);
xnor U9361 (N_9361,N_9128,N_9145);
xnor U9362 (N_9362,N_9027,N_9025);
and U9363 (N_9363,N_9016,N_9184);
or U9364 (N_9364,N_9025,N_9068);
nor U9365 (N_9365,N_9135,N_9009);
and U9366 (N_9366,N_9105,N_9150);
nor U9367 (N_9367,N_9196,N_9019);
and U9368 (N_9368,N_9019,N_9171);
nand U9369 (N_9369,N_9023,N_9149);
nand U9370 (N_9370,N_9073,N_9039);
and U9371 (N_9371,N_9194,N_9112);
nand U9372 (N_9372,N_9093,N_9153);
or U9373 (N_9373,N_9104,N_9077);
xor U9374 (N_9374,N_9047,N_9186);
and U9375 (N_9375,N_9117,N_9067);
or U9376 (N_9376,N_9046,N_9080);
nand U9377 (N_9377,N_9160,N_9002);
xnor U9378 (N_9378,N_9026,N_9027);
or U9379 (N_9379,N_9064,N_9034);
and U9380 (N_9380,N_9183,N_9102);
xor U9381 (N_9381,N_9172,N_9049);
nor U9382 (N_9382,N_9189,N_9102);
and U9383 (N_9383,N_9191,N_9021);
nand U9384 (N_9384,N_9005,N_9164);
and U9385 (N_9385,N_9119,N_9182);
or U9386 (N_9386,N_9185,N_9019);
or U9387 (N_9387,N_9152,N_9191);
or U9388 (N_9388,N_9051,N_9163);
nand U9389 (N_9389,N_9095,N_9002);
nand U9390 (N_9390,N_9015,N_9129);
and U9391 (N_9391,N_9171,N_9106);
or U9392 (N_9392,N_9042,N_9007);
or U9393 (N_9393,N_9180,N_9189);
nand U9394 (N_9394,N_9190,N_9053);
and U9395 (N_9395,N_9084,N_9096);
nand U9396 (N_9396,N_9191,N_9166);
and U9397 (N_9397,N_9194,N_9012);
xnor U9398 (N_9398,N_9197,N_9077);
nand U9399 (N_9399,N_9183,N_9032);
nor U9400 (N_9400,N_9351,N_9331);
or U9401 (N_9401,N_9296,N_9333);
xnor U9402 (N_9402,N_9369,N_9291);
nor U9403 (N_9403,N_9215,N_9207);
nor U9404 (N_9404,N_9300,N_9284);
nand U9405 (N_9405,N_9288,N_9228);
nor U9406 (N_9406,N_9314,N_9307);
or U9407 (N_9407,N_9224,N_9270);
xnor U9408 (N_9408,N_9366,N_9387);
or U9409 (N_9409,N_9203,N_9276);
or U9410 (N_9410,N_9349,N_9273);
nor U9411 (N_9411,N_9233,N_9289);
xor U9412 (N_9412,N_9287,N_9386);
or U9413 (N_9413,N_9247,N_9274);
nand U9414 (N_9414,N_9363,N_9248);
or U9415 (N_9415,N_9392,N_9383);
and U9416 (N_9416,N_9399,N_9285);
and U9417 (N_9417,N_9246,N_9393);
nand U9418 (N_9418,N_9326,N_9372);
xnor U9419 (N_9419,N_9375,N_9234);
nor U9420 (N_9420,N_9292,N_9384);
and U9421 (N_9421,N_9360,N_9279);
nand U9422 (N_9422,N_9275,N_9376);
nand U9423 (N_9423,N_9257,N_9316);
or U9424 (N_9424,N_9319,N_9282);
nor U9425 (N_9425,N_9385,N_9239);
xor U9426 (N_9426,N_9330,N_9322);
and U9427 (N_9427,N_9343,N_9223);
xor U9428 (N_9428,N_9344,N_9213);
nor U9429 (N_9429,N_9252,N_9315);
nor U9430 (N_9430,N_9327,N_9381);
nand U9431 (N_9431,N_9256,N_9310);
nor U9432 (N_9432,N_9394,N_9377);
nand U9433 (N_9433,N_9235,N_9339);
or U9434 (N_9434,N_9323,N_9345);
xnor U9435 (N_9435,N_9295,N_9373);
nor U9436 (N_9436,N_9308,N_9268);
xor U9437 (N_9437,N_9361,N_9202);
nor U9438 (N_9438,N_9320,N_9301);
nand U9439 (N_9439,N_9293,N_9312);
nand U9440 (N_9440,N_9318,N_9281);
and U9441 (N_9441,N_9368,N_9371);
xor U9442 (N_9442,N_9214,N_9396);
nand U9443 (N_9443,N_9258,N_9302);
nand U9444 (N_9444,N_9259,N_9237);
or U9445 (N_9445,N_9388,N_9283);
nand U9446 (N_9446,N_9346,N_9226);
and U9447 (N_9447,N_9210,N_9378);
xnor U9448 (N_9448,N_9370,N_9303);
or U9449 (N_9449,N_9249,N_9306);
nand U9450 (N_9450,N_9251,N_9321);
nand U9451 (N_9451,N_9267,N_9278);
xnor U9452 (N_9452,N_9242,N_9355);
xnor U9453 (N_9453,N_9263,N_9362);
and U9454 (N_9454,N_9391,N_9240);
or U9455 (N_9455,N_9340,N_9338);
nor U9456 (N_9456,N_9364,N_9334);
xnor U9457 (N_9457,N_9398,N_9221);
and U9458 (N_9458,N_9220,N_9230);
nand U9459 (N_9459,N_9261,N_9272);
nand U9460 (N_9460,N_9217,N_9313);
and U9461 (N_9461,N_9297,N_9200);
and U9462 (N_9462,N_9253,N_9211);
xor U9463 (N_9463,N_9260,N_9222);
or U9464 (N_9464,N_9336,N_9238);
and U9465 (N_9465,N_9328,N_9382);
nor U9466 (N_9466,N_9311,N_9350);
and U9467 (N_9467,N_9205,N_9299);
nand U9468 (N_9468,N_9286,N_9219);
or U9469 (N_9469,N_9266,N_9212);
nor U9470 (N_9470,N_9290,N_9337);
nor U9471 (N_9471,N_9354,N_9342);
nand U9472 (N_9472,N_9305,N_9358);
and U9473 (N_9473,N_9329,N_9269);
or U9474 (N_9474,N_9335,N_9324);
nor U9475 (N_9475,N_9277,N_9243);
and U9476 (N_9476,N_9352,N_9379);
xnor U9477 (N_9477,N_9208,N_9365);
or U9478 (N_9478,N_9332,N_9325);
or U9479 (N_9479,N_9245,N_9390);
and U9480 (N_9480,N_9397,N_9255);
xor U9481 (N_9481,N_9341,N_9304);
nor U9482 (N_9482,N_9317,N_9367);
or U9483 (N_9483,N_9227,N_9264);
xor U9484 (N_9484,N_9348,N_9201);
or U9485 (N_9485,N_9357,N_9298);
xor U9486 (N_9486,N_9236,N_9280);
nor U9487 (N_9487,N_9204,N_9209);
or U9488 (N_9488,N_9395,N_9254);
or U9489 (N_9489,N_9359,N_9374);
nor U9490 (N_9490,N_9206,N_9218);
xnor U9491 (N_9491,N_9244,N_9262);
and U9492 (N_9492,N_9309,N_9216);
or U9493 (N_9493,N_9232,N_9231);
nand U9494 (N_9494,N_9229,N_9225);
and U9495 (N_9495,N_9353,N_9356);
nor U9496 (N_9496,N_9294,N_9250);
and U9497 (N_9497,N_9271,N_9347);
nor U9498 (N_9498,N_9389,N_9380);
and U9499 (N_9499,N_9265,N_9241);
nand U9500 (N_9500,N_9216,N_9219);
nand U9501 (N_9501,N_9275,N_9360);
xor U9502 (N_9502,N_9346,N_9297);
xnor U9503 (N_9503,N_9297,N_9278);
or U9504 (N_9504,N_9355,N_9216);
or U9505 (N_9505,N_9359,N_9398);
and U9506 (N_9506,N_9266,N_9358);
and U9507 (N_9507,N_9201,N_9269);
nor U9508 (N_9508,N_9365,N_9360);
nor U9509 (N_9509,N_9362,N_9215);
and U9510 (N_9510,N_9284,N_9279);
or U9511 (N_9511,N_9298,N_9301);
or U9512 (N_9512,N_9382,N_9219);
or U9513 (N_9513,N_9325,N_9362);
or U9514 (N_9514,N_9217,N_9236);
xor U9515 (N_9515,N_9359,N_9237);
nand U9516 (N_9516,N_9353,N_9235);
nor U9517 (N_9517,N_9391,N_9393);
or U9518 (N_9518,N_9216,N_9276);
nor U9519 (N_9519,N_9257,N_9311);
and U9520 (N_9520,N_9307,N_9221);
or U9521 (N_9521,N_9332,N_9351);
nor U9522 (N_9522,N_9392,N_9212);
or U9523 (N_9523,N_9208,N_9355);
xor U9524 (N_9524,N_9395,N_9250);
or U9525 (N_9525,N_9240,N_9211);
nor U9526 (N_9526,N_9279,N_9254);
nor U9527 (N_9527,N_9306,N_9335);
or U9528 (N_9528,N_9288,N_9392);
nand U9529 (N_9529,N_9206,N_9352);
nor U9530 (N_9530,N_9293,N_9227);
nor U9531 (N_9531,N_9273,N_9219);
or U9532 (N_9532,N_9274,N_9263);
xnor U9533 (N_9533,N_9226,N_9246);
nor U9534 (N_9534,N_9353,N_9233);
or U9535 (N_9535,N_9339,N_9205);
nor U9536 (N_9536,N_9385,N_9254);
xor U9537 (N_9537,N_9207,N_9268);
xor U9538 (N_9538,N_9270,N_9216);
or U9539 (N_9539,N_9357,N_9398);
nand U9540 (N_9540,N_9300,N_9332);
nor U9541 (N_9541,N_9236,N_9351);
and U9542 (N_9542,N_9235,N_9245);
and U9543 (N_9543,N_9277,N_9398);
and U9544 (N_9544,N_9270,N_9258);
nor U9545 (N_9545,N_9255,N_9263);
xor U9546 (N_9546,N_9273,N_9374);
xor U9547 (N_9547,N_9350,N_9356);
nand U9548 (N_9548,N_9295,N_9228);
and U9549 (N_9549,N_9211,N_9304);
nor U9550 (N_9550,N_9362,N_9390);
or U9551 (N_9551,N_9334,N_9232);
and U9552 (N_9552,N_9388,N_9291);
or U9553 (N_9553,N_9318,N_9340);
xor U9554 (N_9554,N_9205,N_9216);
nand U9555 (N_9555,N_9248,N_9282);
xnor U9556 (N_9556,N_9314,N_9209);
nor U9557 (N_9557,N_9318,N_9317);
nand U9558 (N_9558,N_9269,N_9211);
nor U9559 (N_9559,N_9375,N_9374);
and U9560 (N_9560,N_9244,N_9265);
and U9561 (N_9561,N_9267,N_9237);
xor U9562 (N_9562,N_9200,N_9216);
nand U9563 (N_9563,N_9235,N_9376);
and U9564 (N_9564,N_9282,N_9265);
and U9565 (N_9565,N_9269,N_9299);
xor U9566 (N_9566,N_9218,N_9255);
xnor U9567 (N_9567,N_9296,N_9222);
or U9568 (N_9568,N_9224,N_9314);
nand U9569 (N_9569,N_9354,N_9293);
or U9570 (N_9570,N_9321,N_9218);
xnor U9571 (N_9571,N_9215,N_9210);
nand U9572 (N_9572,N_9355,N_9214);
and U9573 (N_9573,N_9305,N_9379);
xnor U9574 (N_9574,N_9239,N_9380);
nand U9575 (N_9575,N_9272,N_9221);
xnor U9576 (N_9576,N_9390,N_9283);
and U9577 (N_9577,N_9201,N_9256);
and U9578 (N_9578,N_9236,N_9215);
nand U9579 (N_9579,N_9262,N_9355);
nand U9580 (N_9580,N_9293,N_9363);
xor U9581 (N_9581,N_9368,N_9389);
xor U9582 (N_9582,N_9309,N_9350);
or U9583 (N_9583,N_9273,N_9361);
nand U9584 (N_9584,N_9291,N_9285);
nand U9585 (N_9585,N_9335,N_9207);
or U9586 (N_9586,N_9219,N_9260);
nand U9587 (N_9587,N_9347,N_9338);
xnor U9588 (N_9588,N_9218,N_9326);
nand U9589 (N_9589,N_9283,N_9287);
nand U9590 (N_9590,N_9220,N_9339);
xor U9591 (N_9591,N_9247,N_9389);
xor U9592 (N_9592,N_9209,N_9255);
nor U9593 (N_9593,N_9266,N_9215);
xor U9594 (N_9594,N_9290,N_9301);
or U9595 (N_9595,N_9245,N_9288);
nor U9596 (N_9596,N_9290,N_9309);
nor U9597 (N_9597,N_9245,N_9241);
and U9598 (N_9598,N_9319,N_9266);
nor U9599 (N_9599,N_9341,N_9390);
xnor U9600 (N_9600,N_9506,N_9528);
xor U9601 (N_9601,N_9466,N_9574);
nand U9602 (N_9602,N_9434,N_9560);
or U9603 (N_9603,N_9465,N_9490);
xnor U9604 (N_9604,N_9496,N_9477);
or U9605 (N_9605,N_9495,N_9464);
xnor U9606 (N_9606,N_9597,N_9497);
nand U9607 (N_9607,N_9551,N_9457);
xnor U9608 (N_9608,N_9577,N_9584);
nor U9609 (N_9609,N_9550,N_9582);
nand U9610 (N_9610,N_9454,N_9587);
nor U9611 (N_9611,N_9504,N_9439);
or U9612 (N_9612,N_9478,N_9491);
nor U9613 (N_9613,N_9509,N_9585);
nor U9614 (N_9614,N_9489,N_9554);
or U9615 (N_9615,N_9519,N_9419);
nand U9616 (N_9616,N_9578,N_9426);
or U9617 (N_9617,N_9467,N_9415);
and U9618 (N_9618,N_9532,N_9484);
nand U9619 (N_9619,N_9514,N_9565);
xor U9620 (N_9620,N_9453,N_9499);
nor U9621 (N_9621,N_9428,N_9460);
nor U9622 (N_9622,N_9546,N_9450);
nand U9623 (N_9623,N_9581,N_9479);
nor U9624 (N_9624,N_9570,N_9451);
or U9625 (N_9625,N_9527,N_9518);
xnor U9626 (N_9626,N_9513,N_9517);
xnor U9627 (N_9627,N_9566,N_9521);
nand U9628 (N_9628,N_9595,N_9523);
nor U9629 (N_9629,N_9563,N_9594);
nand U9630 (N_9630,N_9480,N_9403);
or U9631 (N_9631,N_9575,N_9561);
xnor U9632 (N_9632,N_9425,N_9562);
nand U9633 (N_9633,N_9423,N_9441);
or U9634 (N_9634,N_9544,N_9462);
and U9635 (N_9635,N_9427,N_9534);
xor U9636 (N_9636,N_9573,N_9412);
and U9637 (N_9637,N_9458,N_9492);
nor U9638 (N_9638,N_9418,N_9508);
nor U9639 (N_9639,N_9433,N_9515);
nor U9640 (N_9640,N_9413,N_9404);
nand U9641 (N_9641,N_9409,N_9400);
xor U9642 (N_9642,N_9598,N_9535);
or U9643 (N_9643,N_9537,N_9402);
and U9644 (N_9644,N_9420,N_9549);
nor U9645 (N_9645,N_9408,N_9405);
nor U9646 (N_9646,N_9586,N_9445);
nand U9647 (N_9647,N_9564,N_9531);
nor U9648 (N_9648,N_9447,N_9436);
nand U9649 (N_9649,N_9470,N_9569);
or U9650 (N_9650,N_9473,N_9468);
nand U9651 (N_9651,N_9442,N_9599);
and U9652 (N_9652,N_9559,N_9556);
or U9653 (N_9653,N_9505,N_9572);
xnor U9654 (N_9654,N_9596,N_9503);
or U9655 (N_9655,N_9592,N_9590);
nor U9656 (N_9656,N_9540,N_9580);
and U9657 (N_9657,N_9449,N_9576);
nor U9658 (N_9658,N_9401,N_9414);
xnor U9659 (N_9659,N_9583,N_9482);
nand U9660 (N_9660,N_9437,N_9488);
and U9661 (N_9661,N_9456,N_9486);
xnor U9662 (N_9662,N_9406,N_9526);
nor U9663 (N_9663,N_9525,N_9438);
or U9664 (N_9664,N_9455,N_9552);
xor U9665 (N_9665,N_9485,N_9511);
or U9666 (N_9666,N_9507,N_9440);
nand U9667 (N_9667,N_9568,N_9444);
nor U9668 (N_9668,N_9538,N_9475);
nor U9669 (N_9669,N_9463,N_9543);
and U9670 (N_9670,N_9541,N_9494);
and U9671 (N_9671,N_9446,N_9571);
nor U9672 (N_9672,N_9469,N_9424);
and U9673 (N_9673,N_9500,N_9591);
nor U9674 (N_9674,N_9502,N_9530);
nand U9675 (N_9675,N_9472,N_9533);
and U9676 (N_9676,N_9579,N_9452);
or U9677 (N_9677,N_9567,N_9430);
or U9678 (N_9678,N_9548,N_9501);
and U9679 (N_9679,N_9555,N_9510);
xor U9680 (N_9680,N_9593,N_9476);
and U9681 (N_9681,N_9474,N_9588);
xnor U9682 (N_9682,N_9416,N_9520);
and U9683 (N_9683,N_9539,N_9410);
nand U9684 (N_9684,N_9407,N_9553);
nand U9685 (N_9685,N_9512,N_9547);
xor U9686 (N_9686,N_9536,N_9421);
nand U9687 (N_9687,N_9411,N_9417);
xnor U9688 (N_9688,N_9493,N_9422);
and U9689 (N_9689,N_9448,N_9498);
and U9690 (N_9690,N_9435,N_9429);
xnor U9691 (N_9691,N_9522,N_9443);
or U9692 (N_9692,N_9529,N_9558);
and U9693 (N_9693,N_9589,N_9545);
nor U9694 (N_9694,N_9471,N_9542);
nand U9695 (N_9695,N_9461,N_9483);
nor U9696 (N_9696,N_9516,N_9524);
nand U9697 (N_9697,N_9431,N_9432);
xor U9698 (N_9698,N_9481,N_9487);
nand U9699 (N_9699,N_9459,N_9557);
or U9700 (N_9700,N_9578,N_9405);
nand U9701 (N_9701,N_9508,N_9481);
xor U9702 (N_9702,N_9459,N_9562);
xor U9703 (N_9703,N_9581,N_9448);
or U9704 (N_9704,N_9486,N_9458);
nor U9705 (N_9705,N_9401,N_9500);
and U9706 (N_9706,N_9509,N_9413);
and U9707 (N_9707,N_9481,N_9494);
or U9708 (N_9708,N_9458,N_9569);
or U9709 (N_9709,N_9571,N_9534);
nand U9710 (N_9710,N_9593,N_9454);
nor U9711 (N_9711,N_9581,N_9530);
and U9712 (N_9712,N_9569,N_9479);
or U9713 (N_9713,N_9462,N_9445);
nor U9714 (N_9714,N_9480,N_9499);
nor U9715 (N_9715,N_9432,N_9437);
or U9716 (N_9716,N_9457,N_9556);
or U9717 (N_9717,N_9400,N_9541);
xnor U9718 (N_9718,N_9460,N_9424);
nor U9719 (N_9719,N_9437,N_9491);
xor U9720 (N_9720,N_9543,N_9482);
or U9721 (N_9721,N_9523,N_9514);
xnor U9722 (N_9722,N_9423,N_9486);
nor U9723 (N_9723,N_9411,N_9587);
nor U9724 (N_9724,N_9549,N_9491);
or U9725 (N_9725,N_9571,N_9505);
or U9726 (N_9726,N_9481,N_9480);
or U9727 (N_9727,N_9485,N_9510);
and U9728 (N_9728,N_9565,N_9488);
nor U9729 (N_9729,N_9529,N_9452);
xor U9730 (N_9730,N_9577,N_9559);
nor U9731 (N_9731,N_9448,N_9594);
or U9732 (N_9732,N_9572,N_9450);
xor U9733 (N_9733,N_9447,N_9443);
and U9734 (N_9734,N_9447,N_9566);
nand U9735 (N_9735,N_9539,N_9401);
or U9736 (N_9736,N_9469,N_9474);
xnor U9737 (N_9737,N_9534,N_9518);
or U9738 (N_9738,N_9577,N_9505);
nor U9739 (N_9739,N_9488,N_9590);
xnor U9740 (N_9740,N_9433,N_9440);
or U9741 (N_9741,N_9576,N_9531);
nor U9742 (N_9742,N_9594,N_9403);
or U9743 (N_9743,N_9541,N_9571);
nand U9744 (N_9744,N_9550,N_9522);
nand U9745 (N_9745,N_9520,N_9585);
and U9746 (N_9746,N_9458,N_9418);
xnor U9747 (N_9747,N_9460,N_9588);
nor U9748 (N_9748,N_9441,N_9505);
nand U9749 (N_9749,N_9466,N_9518);
nand U9750 (N_9750,N_9580,N_9556);
and U9751 (N_9751,N_9453,N_9521);
or U9752 (N_9752,N_9575,N_9541);
and U9753 (N_9753,N_9531,N_9533);
nand U9754 (N_9754,N_9563,N_9436);
nand U9755 (N_9755,N_9443,N_9400);
and U9756 (N_9756,N_9549,N_9463);
nand U9757 (N_9757,N_9571,N_9434);
or U9758 (N_9758,N_9446,N_9428);
nor U9759 (N_9759,N_9461,N_9593);
or U9760 (N_9760,N_9592,N_9528);
and U9761 (N_9761,N_9599,N_9585);
and U9762 (N_9762,N_9573,N_9580);
and U9763 (N_9763,N_9422,N_9439);
nor U9764 (N_9764,N_9439,N_9487);
xor U9765 (N_9765,N_9407,N_9527);
or U9766 (N_9766,N_9456,N_9415);
nand U9767 (N_9767,N_9505,N_9464);
xnor U9768 (N_9768,N_9503,N_9547);
nor U9769 (N_9769,N_9596,N_9493);
nor U9770 (N_9770,N_9589,N_9516);
nand U9771 (N_9771,N_9558,N_9433);
nor U9772 (N_9772,N_9454,N_9428);
nor U9773 (N_9773,N_9440,N_9550);
xor U9774 (N_9774,N_9585,N_9582);
xor U9775 (N_9775,N_9597,N_9590);
nor U9776 (N_9776,N_9433,N_9582);
xnor U9777 (N_9777,N_9467,N_9542);
and U9778 (N_9778,N_9400,N_9517);
xor U9779 (N_9779,N_9404,N_9542);
and U9780 (N_9780,N_9517,N_9563);
or U9781 (N_9781,N_9584,N_9457);
or U9782 (N_9782,N_9404,N_9557);
xor U9783 (N_9783,N_9576,N_9452);
xnor U9784 (N_9784,N_9515,N_9539);
nand U9785 (N_9785,N_9591,N_9567);
and U9786 (N_9786,N_9436,N_9432);
and U9787 (N_9787,N_9432,N_9416);
nor U9788 (N_9788,N_9500,N_9471);
xnor U9789 (N_9789,N_9461,N_9436);
nor U9790 (N_9790,N_9483,N_9592);
and U9791 (N_9791,N_9409,N_9411);
nor U9792 (N_9792,N_9415,N_9468);
xnor U9793 (N_9793,N_9499,N_9575);
and U9794 (N_9794,N_9584,N_9595);
nor U9795 (N_9795,N_9520,N_9598);
xor U9796 (N_9796,N_9517,N_9421);
nor U9797 (N_9797,N_9440,N_9598);
xnor U9798 (N_9798,N_9421,N_9424);
xnor U9799 (N_9799,N_9423,N_9431);
nand U9800 (N_9800,N_9660,N_9784);
nor U9801 (N_9801,N_9652,N_9766);
or U9802 (N_9802,N_9779,N_9727);
and U9803 (N_9803,N_9631,N_9719);
and U9804 (N_9804,N_9761,N_9681);
or U9805 (N_9805,N_9742,N_9629);
and U9806 (N_9806,N_9703,N_9769);
nand U9807 (N_9807,N_9695,N_9698);
or U9808 (N_9808,N_9635,N_9633);
and U9809 (N_9809,N_9749,N_9697);
nand U9810 (N_9810,N_9632,N_9620);
nor U9811 (N_9811,N_9684,N_9713);
or U9812 (N_9812,N_9638,N_9777);
and U9813 (N_9813,N_9702,N_9630);
xnor U9814 (N_9814,N_9792,N_9772);
nand U9815 (N_9815,N_9600,N_9643);
and U9816 (N_9816,N_9694,N_9641);
nand U9817 (N_9817,N_9640,N_9752);
xnor U9818 (N_9818,N_9607,N_9731);
or U9819 (N_9819,N_9711,N_9778);
and U9820 (N_9820,N_9667,N_9775);
nand U9821 (N_9821,N_9747,N_9647);
xnor U9822 (N_9822,N_9706,N_9745);
xor U9823 (N_9823,N_9648,N_9767);
or U9824 (N_9824,N_9780,N_9798);
or U9825 (N_9825,N_9774,N_9797);
xnor U9826 (N_9826,N_9786,N_9751);
or U9827 (N_9827,N_9645,N_9606);
nor U9828 (N_9828,N_9665,N_9622);
nor U9829 (N_9829,N_9672,N_9678);
nor U9830 (N_9830,N_9714,N_9626);
nor U9831 (N_9831,N_9758,N_9655);
xor U9832 (N_9832,N_9619,N_9612);
nand U9833 (N_9833,N_9674,N_9671);
nor U9834 (N_9834,N_9646,N_9666);
xnor U9835 (N_9835,N_9710,N_9699);
nor U9836 (N_9836,N_9720,N_9611);
nand U9837 (N_9837,N_9615,N_9617);
xor U9838 (N_9838,N_9738,N_9683);
xor U9839 (N_9839,N_9618,N_9680);
nand U9840 (N_9840,N_9729,N_9799);
nand U9841 (N_9841,N_9604,N_9691);
and U9842 (N_9842,N_9675,N_9716);
or U9843 (N_9843,N_9709,N_9781);
nor U9844 (N_9844,N_9726,N_9602);
nand U9845 (N_9845,N_9785,N_9649);
and U9846 (N_9846,N_9768,N_9794);
xnor U9847 (N_9847,N_9613,N_9658);
nor U9848 (N_9848,N_9624,N_9701);
xor U9849 (N_9849,N_9746,N_9670);
nor U9850 (N_9850,N_9627,N_9730);
nand U9851 (N_9851,N_9636,N_9717);
xor U9852 (N_9852,N_9748,N_9705);
and U9853 (N_9853,N_9605,N_9628);
nor U9854 (N_9854,N_9728,N_9621);
nor U9855 (N_9855,N_9759,N_9688);
xnor U9856 (N_9856,N_9686,N_9651);
or U9857 (N_9857,N_9639,N_9789);
nand U9858 (N_9858,N_9608,N_9659);
and U9859 (N_9859,N_9722,N_9669);
nand U9860 (N_9860,N_9744,N_9668);
nand U9861 (N_9861,N_9679,N_9663);
or U9862 (N_9862,N_9650,N_9791);
and U9863 (N_9863,N_9673,N_9754);
nand U9864 (N_9864,N_9707,N_9614);
and U9865 (N_9865,N_9733,N_9740);
nor U9866 (N_9866,N_9708,N_9753);
nor U9867 (N_9867,N_9682,N_9712);
and U9868 (N_9868,N_9757,N_9725);
or U9869 (N_9869,N_9783,N_9718);
xor U9870 (N_9870,N_9715,N_9601);
and U9871 (N_9871,N_9677,N_9692);
xor U9872 (N_9872,N_9637,N_9644);
nand U9873 (N_9873,N_9625,N_9653);
nand U9874 (N_9874,N_9610,N_9734);
nor U9875 (N_9875,N_9762,N_9603);
or U9876 (N_9876,N_9743,N_9661);
nor U9877 (N_9877,N_9737,N_9634);
and U9878 (N_9878,N_9773,N_9750);
nor U9879 (N_9879,N_9771,N_9690);
or U9880 (N_9880,N_9787,N_9782);
xnor U9881 (N_9881,N_9763,N_9623);
or U9882 (N_9882,N_9696,N_9616);
or U9883 (N_9883,N_9664,N_9765);
or U9884 (N_9884,N_9685,N_9656);
nand U9885 (N_9885,N_9642,N_9724);
or U9886 (N_9886,N_9756,N_9704);
and U9887 (N_9887,N_9732,N_9693);
nand U9888 (N_9888,N_9687,N_9662);
nor U9889 (N_9889,N_9609,N_9723);
xnor U9890 (N_9890,N_9770,N_9736);
nand U9891 (N_9891,N_9676,N_9795);
nor U9892 (N_9892,N_9790,N_9764);
nand U9893 (N_9893,N_9776,N_9760);
xnor U9894 (N_9894,N_9793,N_9741);
xor U9895 (N_9895,N_9654,N_9721);
or U9896 (N_9896,N_9788,N_9739);
and U9897 (N_9897,N_9735,N_9689);
or U9898 (N_9898,N_9700,N_9796);
nand U9899 (N_9899,N_9657,N_9755);
nor U9900 (N_9900,N_9675,N_9796);
nor U9901 (N_9901,N_9734,N_9771);
and U9902 (N_9902,N_9773,N_9660);
and U9903 (N_9903,N_9751,N_9666);
nand U9904 (N_9904,N_9698,N_9671);
and U9905 (N_9905,N_9644,N_9613);
nand U9906 (N_9906,N_9785,N_9654);
or U9907 (N_9907,N_9762,N_9725);
or U9908 (N_9908,N_9640,N_9765);
or U9909 (N_9909,N_9780,N_9617);
nor U9910 (N_9910,N_9761,N_9618);
xor U9911 (N_9911,N_9797,N_9641);
and U9912 (N_9912,N_9760,N_9748);
nor U9913 (N_9913,N_9763,N_9684);
nand U9914 (N_9914,N_9799,N_9656);
nor U9915 (N_9915,N_9760,N_9755);
nand U9916 (N_9916,N_9717,N_9693);
and U9917 (N_9917,N_9652,N_9695);
or U9918 (N_9918,N_9620,N_9754);
and U9919 (N_9919,N_9692,N_9691);
xnor U9920 (N_9920,N_9619,N_9774);
or U9921 (N_9921,N_9652,N_9622);
and U9922 (N_9922,N_9659,N_9640);
and U9923 (N_9923,N_9740,N_9783);
and U9924 (N_9924,N_9777,N_9740);
xnor U9925 (N_9925,N_9736,N_9663);
and U9926 (N_9926,N_9625,N_9678);
and U9927 (N_9927,N_9603,N_9746);
nand U9928 (N_9928,N_9744,N_9612);
nand U9929 (N_9929,N_9747,N_9705);
nor U9930 (N_9930,N_9736,N_9757);
or U9931 (N_9931,N_9781,N_9771);
xor U9932 (N_9932,N_9622,N_9762);
or U9933 (N_9933,N_9744,N_9689);
or U9934 (N_9934,N_9754,N_9657);
nor U9935 (N_9935,N_9759,N_9630);
and U9936 (N_9936,N_9645,N_9722);
and U9937 (N_9937,N_9732,N_9703);
nor U9938 (N_9938,N_9755,N_9692);
nor U9939 (N_9939,N_9635,N_9622);
nand U9940 (N_9940,N_9764,N_9778);
or U9941 (N_9941,N_9660,N_9741);
or U9942 (N_9942,N_9612,N_9673);
nor U9943 (N_9943,N_9655,N_9795);
nand U9944 (N_9944,N_9735,N_9764);
xor U9945 (N_9945,N_9733,N_9779);
nand U9946 (N_9946,N_9693,N_9779);
xnor U9947 (N_9947,N_9693,N_9762);
nand U9948 (N_9948,N_9744,N_9625);
xor U9949 (N_9949,N_9783,N_9702);
and U9950 (N_9950,N_9773,N_9612);
and U9951 (N_9951,N_9665,N_9722);
nor U9952 (N_9952,N_9613,N_9602);
and U9953 (N_9953,N_9616,N_9660);
nor U9954 (N_9954,N_9728,N_9629);
nor U9955 (N_9955,N_9710,N_9698);
nor U9956 (N_9956,N_9784,N_9617);
nor U9957 (N_9957,N_9640,N_9766);
or U9958 (N_9958,N_9765,N_9727);
nand U9959 (N_9959,N_9672,N_9710);
nand U9960 (N_9960,N_9616,N_9667);
or U9961 (N_9961,N_9693,N_9769);
xor U9962 (N_9962,N_9738,N_9702);
nor U9963 (N_9963,N_9659,N_9606);
xor U9964 (N_9964,N_9696,N_9627);
nor U9965 (N_9965,N_9600,N_9646);
and U9966 (N_9966,N_9609,N_9631);
or U9967 (N_9967,N_9642,N_9624);
nor U9968 (N_9968,N_9699,N_9652);
or U9969 (N_9969,N_9620,N_9681);
nand U9970 (N_9970,N_9708,N_9768);
nand U9971 (N_9971,N_9660,N_9790);
nor U9972 (N_9972,N_9787,N_9659);
xor U9973 (N_9973,N_9643,N_9758);
nor U9974 (N_9974,N_9788,N_9737);
nor U9975 (N_9975,N_9725,N_9681);
and U9976 (N_9976,N_9699,N_9633);
and U9977 (N_9977,N_9770,N_9623);
nor U9978 (N_9978,N_9678,N_9792);
or U9979 (N_9979,N_9618,N_9714);
nor U9980 (N_9980,N_9766,N_9731);
nand U9981 (N_9981,N_9602,N_9731);
nand U9982 (N_9982,N_9716,N_9646);
nor U9983 (N_9983,N_9759,N_9741);
or U9984 (N_9984,N_9641,N_9602);
nand U9985 (N_9985,N_9769,N_9640);
nand U9986 (N_9986,N_9652,N_9734);
nand U9987 (N_9987,N_9773,N_9752);
and U9988 (N_9988,N_9718,N_9721);
nand U9989 (N_9989,N_9798,N_9778);
and U9990 (N_9990,N_9626,N_9697);
xor U9991 (N_9991,N_9681,N_9716);
nand U9992 (N_9992,N_9657,N_9714);
xor U9993 (N_9993,N_9770,N_9626);
and U9994 (N_9994,N_9617,N_9689);
nand U9995 (N_9995,N_9790,N_9624);
nor U9996 (N_9996,N_9764,N_9711);
and U9997 (N_9997,N_9754,N_9623);
or U9998 (N_9998,N_9653,N_9600);
and U9999 (N_9999,N_9649,N_9713);
or UO_0 (O_0,N_9986,N_9972);
nand UO_1 (O_1,N_9951,N_9922);
nand UO_2 (O_2,N_9858,N_9995);
or UO_3 (O_3,N_9880,N_9833);
and UO_4 (O_4,N_9904,N_9895);
nor UO_5 (O_5,N_9850,N_9965);
and UO_6 (O_6,N_9890,N_9823);
and UO_7 (O_7,N_9982,N_9848);
nand UO_8 (O_8,N_9847,N_9821);
or UO_9 (O_9,N_9942,N_9867);
and UO_10 (O_10,N_9831,N_9881);
nand UO_11 (O_11,N_9876,N_9872);
and UO_12 (O_12,N_9868,N_9884);
or UO_13 (O_13,N_9996,N_9891);
nor UO_14 (O_14,N_9997,N_9844);
or UO_15 (O_15,N_9914,N_9945);
nand UO_16 (O_16,N_9941,N_9985);
or UO_17 (O_17,N_9934,N_9973);
nor UO_18 (O_18,N_9961,N_9912);
xnor UO_19 (O_19,N_9878,N_9936);
nor UO_20 (O_20,N_9988,N_9970);
nor UO_21 (O_21,N_9959,N_9931);
or UO_22 (O_22,N_9851,N_9882);
nor UO_23 (O_23,N_9975,N_9836);
or UO_24 (O_24,N_9856,N_9919);
nand UO_25 (O_25,N_9849,N_9888);
or UO_26 (O_26,N_9929,N_9913);
or UO_27 (O_27,N_9841,N_9933);
or UO_28 (O_28,N_9852,N_9954);
nor UO_29 (O_29,N_9889,N_9886);
nor UO_30 (O_30,N_9800,N_9971);
or UO_31 (O_31,N_9947,N_9864);
xor UO_32 (O_32,N_9815,N_9979);
nand UO_33 (O_33,N_9828,N_9960);
nor UO_34 (O_34,N_9953,N_9955);
and UO_35 (O_35,N_9826,N_9897);
or UO_36 (O_36,N_9926,N_9801);
xor UO_37 (O_37,N_9989,N_9937);
nand UO_38 (O_38,N_9920,N_9976);
nor UO_39 (O_39,N_9869,N_9908);
nand UO_40 (O_40,N_9827,N_9909);
xnor UO_41 (O_41,N_9903,N_9834);
nor UO_42 (O_42,N_9928,N_9984);
or UO_43 (O_43,N_9949,N_9870);
xnor UO_44 (O_44,N_9803,N_9837);
or UO_45 (O_45,N_9863,N_9812);
nor UO_46 (O_46,N_9952,N_9977);
nand UO_47 (O_47,N_9917,N_9906);
nand UO_48 (O_48,N_9840,N_9894);
and UO_49 (O_49,N_9811,N_9855);
and UO_50 (O_50,N_9885,N_9842);
nor UO_51 (O_51,N_9932,N_9939);
and UO_52 (O_52,N_9809,N_9991);
nor UO_53 (O_53,N_9896,N_9946);
nor UO_54 (O_54,N_9963,N_9879);
or UO_55 (O_55,N_9938,N_9822);
nor UO_56 (O_56,N_9899,N_9861);
or UO_57 (O_57,N_9935,N_9887);
or UO_58 (O_58,N_9910,N_9873);
or UO_59 (O_59,N_9839,N_9865);
and UO_60 (O_60,N_9859,N_9829);
or UO_61 (O_61,N_9854,N_9990);
xor UO_62 (O_62,N_9804,N_9916);
xor UO_63 (O_63,N_9962,N_9810);
and UO_64 (O_64,N_9892,N_9980);
xnor UO_65 (O_65,N_9806,N_9925);
xnor UO_66 (O_66,N_9957,N_9808);
or UO_67 (O_67,N_9900,N_9857);
nand UO_68 (O_68,N_9802,N_9969);
nor UO_69 (O_69,N_9958,N_9893);
xnor UO_70 (O_70,N_9898,N_9944);
nand UO_71 (O_71,N_9966,N_9846);
and UO_72 (O_72,N_9871,N_9940);
and UO_73 (O_73,N_9902,N_9983);
and UO_74 (O_74,N_9883,N_9805);
and UO_75 (O_75,N_9999,N_9807);
nand UO_76 (O_76,N_9838,N_9974);
nor UO_77 (O_77,N_9911,N_9998);
nor UO_78 (O_78,N_9927,N_9824);
or UO_79 (O_79,N_9981,N_9905);
nand UO_80 (O_80,N_9921,N_9950);
or UO_81 (O_81,N_9845,N_9964);
xor UO_82 (O_82,N_9866,N_9825);
nand UO_83 (O_83,N_9819,N_9818);
xor UO_84 (O_84,N_9875,N_9874);
nor UO_85 (O_85,N_9814,N_9813);
xor UO_86 (O_86,N_9968,N_9943);
xnor UO_87 (O_87,N_9967,N_9817);
nor UO_88 (O_88,N_9924,N_9862);
and UO_89 (O_89,N_9832,N_9956);
nor UO_90 (O_90,N_9860,N_9915);
and UO_91 (O_91,N_9978,N_9948);
and UO_92 (O_92,N_9820,N_9830);
xnor UO_93 (O_93,N_9901,N_9994);
xor UO_94 (O_94,N_9907,N_9930);
nor UO_95 (O_95,N_9992,N_9816);
or UO_96 (O_96,N_9987,N_9923);
nand UO_97 (O_97,N_9918,N_9843);
nand UO_98 (O_98,N_9877,N_9835);
or UO_99 (O_99,N_9993,N_9853);
xor UO_100 (O_100,N_9980,N_9919);
nand UO_101 (O_101,N_9922,N_9890);
and UO_102 (O_102,N_9939,N_9905);
nand UO_103 (O_103,N_9864,N_9968);
and UO_104 (O_104,N_9944,N_9918);
nand UO_105 (O_105,N_9883,N_9817);
xnor UO_106 (O_106,N_9991,N_9969);
and UO_107 (O_107,N_9986,N_9933);
or UO_108 (O_108,N_9887,N_9911);
nand UO_109 (O_109,N_9934,N_9949);
nand UO_110 (O_110,N_9868,N_9877);
xor UO_111 (O_111,N_9806,N_9894);
nor UO_112 (O_112,N_9824,N_9991);
or UO_113 (O_113,N_9801,N_9944);
nand UO_114 (O_114,N_9888,N_9870);
nand UO_115 (O_115,N_9806,N_9923);
nor UO_116 (O_116,N_9904,N_9823);
and UO_117 (O_117,N_9862,N_9894);
or UO_118 (O_118,N_9820,N_9958);
nand UO_119 (O_119,N_9976,N_9803);
xor UO_120 (O_120,N_9886,N_9816);
or UO_121 (O_121,N_9990,N_9930);
nor UO_122 (O_122,N_9992,N_9956);
nor UO_123 (O_123,N_9946,N_9894);
and UO_124 (O_124,N_9810,N_9864);
nand UO_125 (O_125,N_9949,N_9901);
nor UO_126 (O_126,N_9965,N_9995);
nand UO_127 (O_127,N_9897,N_9912);
xor UO_128 (O_128,N_9875,N_9993);
nor UO_129 (O_129,N_9820,N_9890);
nor UO_130 (O_130,N_9805,N_9825);
or UO_131 (O_131,N_9988,N_9854);
xnor UO_132 (O_132,N_9988,N_9986);
nand UO_133 (O_133,N_9847,N_9842);
and UO_134 (O_134,N_9944,N_9924);
or UO_135 (O_135,N_9893,N_9978);
and UO_136 (O_136,N_9865,N_9827);
nor UO_137 (O_137,N_9812,N_9993);
or UO_138 (O_138,N_9887,N_9828);
xor UO_139 (O_139,N_9861,N_9806);
nor UO_140 (O_140,N_9898,N_9892);
or UO_141 (O_141,N_9824,N_9925);
nor UO_142 (O_142,N_9948,N_9837);
xnor UO_143 (O_143,N_9840,N_9837);
xor UO_144 (O_144,N_9982,N_9952);
nand UO_145 (O_145,N_9870,N_9978);
xor UO_146 (O_146,N_9840,N_9862);
xnor UO_147 (O_147,N_9892,N_9852);
xnor UO_148 (O_148,N_9905,N_9848);
nor UO_149 (O_149,N_9974,N_9949);
xnor UO_150 (O_150,N_9840,N_9851);
nor UO_151 (O_151,N_9810,N_9865);
and UO_152 (O_152,N_9803,N_9915);
or UO_153 (O_153,N_9820,N_9849);
xnor UO_154 (O_154,N_9857,N_9894);
or UO_155 (O_155,N_9987,N_9876);
nor UO_156 (O_156,N_9851,N_9923);
and UO_157 (O_157,N_9843,N_9874);
xor UO_158 (O_158,N_9945,N_9981);
nand UO_159 (O_159,N_9830,N_9923);
and UO_160 (O_160,N_9836,N_9852);
nor UO_161 (O_161,N_9997,N_9963);
and UO_162 (O_162,N_9901,N_9990);
and UO_163 (O_163,N_9802,N_9809);
and UO_164 (O_164,N_9878,N_9923);
nand UO_165 (O_165,N_9869,N_9841);
nor UO_166 (O_166,N_9843,N_9948);
or UO_167 (O_167,N_9934,N_9887);
and UO_168 (O_168,N_9945,N_9860);
xnor UO_169 (O_169,N_9992,N_9942);
xor UO_170 (O_170,N_9935,N_9825);
nor UO_171 (O_171,N_9906,N_9956);
xor UO_172 (O_172,N_9880,N_9879);
nand UO_173 (O_173,N_9828,N_9968);
or UO_174 (O_174,N_9919,N_9950);
nand UO_175 (O_175,N_9879,N_9907);
and UO_176 (O_176,N_9929,N_9837);
xnor UO_177 (O_177,N_9832,N_9953);
nor UO_178 (O_178,N_9897,N_9988);
and UO_179 (O_179,N_9848,N_9936);
and UO_180 (O_180,N_9923,N_9804);
nand UO_181 (O_181,N_9828,N_9903);
or UO_182 (O_182,N_9891,N_9899);
nand UO_183 (O_183,N_9881,N_9885);
nand UO_184 (O_184,N_9915,N_9912);
nand UO_185 (O_185,N_9908,N_9857);
xnor UO_186 (O_186,N_9875,N_9984);
or UO_187 (O_187,N_9947,N_9962);
and UO_188 (O_188,N_9981,N_9885);
nand UO_189 (O_189,N_9899,N_9818);
nor UO_190 (O_190,N_9858,N_9820);
xnor UO_191 (O_191,N_9934,N_9903);
nor UO_192 (O_192,N_9927,N_9985);
nand UO_193 (O_193,N_9939,N_9894);
or UO_194 (O_194,N_9946,N_9817);
nor UO_195 (O_195,N_9987,N_9919);
and UO_196 (O_196,N_9805,N_9841);
nand UO_197 (O_197,N_9940,N_9838);
nor UO_198 (O_198,N_9996,N_9894);
and UO_199 (O_199,N_9850,N_9825);
and UO_200 (O_200,N_9865,N_9983);
or UO_201 (O_201,N_9954,N_9942);
or UO_202 (O_202,N_9978,N_9969);
nand UO_203 (O_203,N_9904,N_9839);
nand UO_204 (O_204,N_9808,N_9939);
or UO_205 (O_205,N_9923,N_9881);
or UO_206 (O_206,N_9859,N_9927);
and UO_207 (O_207,N_9901,N_9823);
xor UO_208 (O_208,N_9997,N_9980);
xor UO_209 (O_209,N_9811,N_9996);
nand UO_210 (O_210,N_9944,N_9891);
or UO_211 (O_211,N_9941,N_9906);
nor UO_212 (O_212,N_9923,N_9909);
xor UO_213 (O_213,N_9924,N_9840);
and UO_214 (O_214,N_9886,N_9899);
xor UO_215 (O_215,N_9845,N_9804);
xor UO_216 (O_216,N_9823,N_9903);
or UO_217 (O_217,N_9856,N_9868);
or UO_218 (O_218,N_9846,N_9901);
nor UO_219 (O_219,N_9835,N_9842);
or UO_220 (O_220,N_9823,N_9942);
nor UO_221 (O_221,N_9903,N_9951);
nand UO_222 (O_222,N_9874,N_9835);
xnor UO_223 (O_223,N_9886,N_9906);
or UO_224 (O_224,N_9932,N_9924);
xor UO_225 (O_225,N_9932,N_9842);
nand UO_226 (O_226,N_9916,N_9973);
xnor UO_227 (O_227,N_9990,N_9820);
nand UO_228 (O_228,N_9862,N_9910);
nor UO_229 (O_229,N_9904,N_9973);
or UO_230 (O_230,N_9989,N_9804);
nand UO_231 (O_231,N_9961,N_9843);
nor UO_232 (O_232,N_9933,N_9810);
nand UO_233 (O_233,N_9876,N_9871);
xnor UO_234 (O_234,N_9843,N_9844);
xnor UO_235 (O_235,N_9827,N_9953);
nor UO_236 (O_236,N_9896,N_9910);
xor UO_237 (O_237,N_9936,N_9817);
xor UO_238 (O_238,N_9835,N_9922);
nand UO_239 (O_239,N_9829,N_9928);
xnor UO_240 (O_240,N_9897,N_9951);
nand UO_241 (O_241,N_9856,N_9822);
or UO_242 (O_242,N_9991,N_9900);
nor UO_243 (O_243,N_9834,N_9981);
xor UO_244 (O_244,N_9920,N_9887);
and UO_245 (O_245,N_9982,N_9908);
xnor UO_246 (O_246,N_9853,N_9940);
nand UO_247 (O_247,N_9972,N_9943);
nor UO_248 (O_248,N_9861,N_9935);
nand UO_249 (O_249,N_9974,N_9836);
or UO_250 (O_250,N_9809,N_9921);
nor UO_251 (O_251,N_9949,N_9933);
xnor UO_252 (O_252,N_9920,N_9815);
xor UO_253 (O_253,N_9844,N_9852);
or UO_254 (O_254,N_9999,N_9820);
nand UO_255 (O_255,N_9809,N_9944);
xnor UO_256 (O_256,N_9953,N_9914);
and UO_257 (O_257,N_9875,N_9915);
nand UO_258 (O_258,N_9849,N_9950);
nand UO_259 (O_259,N_9886,N_9868);
nand UO_260 (O_260,N_9851,N_9975);
and UO_261 (O_261,N_9954,N_9931);
or UO_262 (O_262,N_9981,N_9959);
and UO_263 (O_263,N_9936,N_9824);
or UO_264 (O_264,N_9804,N_9803);
or UO_265 (O_265,N_9969,N_9946);
nand UO_266 (O_266,N_9899,N_9978);
nand UO_267 (O_267,N_9937,N_9985);
xor UO_268 (O_268,N_9954,N_9949);
xor UO_269 (O_269,N_9828,N_9982);
nand UO_270 (O_270,N_9913,N_9920);
xnor UO_271 (O_271,N_9805,N_9817);
nand UO_272 (O_272,N_9937,N_9982);
xnor UO_273 (O_273,N_9949,N_9918);
nand UO_274 (O_274,N_9900,N_9839);
nor UO_275 (O_275,N_9900,N_9845);
xnor UO_276 (O_276,N_9970,N_9971);
xnor UO_277 (O_277,N_9882,N_9812);
nand UO_278 (O_278,N_9819,N_9967);
nand UO_279 (O_279,N_9937,N_9925);
or UO_280 (O_280,N_9880,N_9860);
nand UO_281 (O_281,N_9924,N_9816);
xnor UO_282 (O_282,N_9919,N_9873);
nor UO_283 (O_283,N_9981,N_9837);
or UO_284 (O_284,N_9810,N_9945);
nand UO_285 (O_285,N_9870,N_9835);
nand UO_286 (O_286,N_9805,N_9998);
or UO_287 (O_287,N_9959,N_9890);
xnor UO_288 (O_288,N_9809,N_9925);
xor UO_289 (O_289,N_9852,N_9802);
or UO_290 (O_290,N_9872,N_9831);
nor UO_291 (O_291,N_9968,N_9811);
and UO_292 (O_292,N_9922,N_9969);
nand UO_293 (O_293,N_9991,N_9989);
or UO_294 (O_294,N_9901,N_9975);
or UO_295 (O_295,N_9983,N_9814);
xor UO_296 (O_296,N_9825,N_9857);
xnor UO_297 (O_297,N_9874,N_9926);
nand UO_298 (O_298,N_9838,N_9896);
and UO_299 (O_299,N_9837,N_9933);
and UO_300 (O_300,N_9922,N_9970);
and UO_301 (O_301,N_9819,N_9948);
and UO_302 (O_302,N_9948,N_9820);
xnor UO_303 (O_303,N_9847,N_9859);
or UO_304 (O_304,N_9996,N_9969);
xor UO_305 (O_305,N_9837,N_9957);
and UO_306 (O_306,N_9894,N_9922);
nor UO_307 (O_307,N_9943,N_9832);
nand UO_308 (O_308,N_9976,N_9829);
xor UO_309 (O_309,N_9908,N_9953);
or UO_310 (O_310,N_9981,N_9983);
xor UO_311 (O_311,N_9909,N_9815);
nor UO_312 (O_312,N_9919,N_9835);
xnor UO_313 (O_313,N_9940,N_9866);
nor UO_314 (O_314,N_9821,N_9889);
or UO_315 (O_315,N_9909,N_9916);
and UO_316 (O_316,N_9818,N_9822);
nand UO_317 (O_317,N_9973,N_9845);
nor UO_318 (O_318,N_9983,N_9929);
and UO_319 (O_319,N_9946,N_9905);
and UO_320 (O_320,N_9818,N_9820);
and UO_321 (O_321,N_9832,N_9843);
nor UO_322 (O_322,N_9887,N_9844);
nor UO_323 (O_323,N_9936,N_9982);
nor UO_324 (O_324,N_9891,N_9897);
nor UO_325 (O_325,N_9917,N_9943);
nor UO_326 (O_326,N_9946,N_9976);
or UO_327 (O_327,N_9829,N_9967);
nand UO_328 (O_328,N_9909,N_9890);
xor UO_329 (O_329,N_9949,N_9863);
and UO_330 (O_330,N_9805,N_9889);
and UO_331 (O_331,N_9915,N_9917);
or UO_332 (O_332,N_9806,N_9825);
nand UO_333 (O_333,N_9942,N_9900);
nand UO_334 (O_334,N_9919,N_9944);
xor UO_335 (O_335,N_9831,N_9919);
nand UO_336 (O_336,N_9903,N_9945);
nor UO_337 (O_337,N_9806,N_9813);
and UO_338 (O_338,N_9943,N_9912);
or UO_339 (O_339,N_9941,N_9964);
xor UO_340 (O_340,N_9990,N_9972);
and UO_341 (O_341,N_9927,N_9867);
xnor UO_342 (O_342,N_9940,N_9951);
and UO_343 (O_343,N_9996,N_9869);
nand UO_344 (O_344,N_9904,N_9933);
nand UO_345 (O_345,N_9873,N_9879);
or UO_346 (O_346,N_9951,N_9965);
nand UO_347 (O_347,N_9837,N_9975);
and UO_348 (O_348,N_9981,N_9889);
and UO_349 (O_349,N_9874,N_9923);
xnor UO_350 (O_350,N_9824,N_9838);
xor UO_351 (O_351,N_9844,N_9841);
or UO_352 (O_352,N_9947,N_9818);
or UO_353 (O_353,N_9859,N_9934);
and UO_354 (O_354,N_9995,N_9903);
or UO_355 (O_355,N_9989,N_9926);
or UO_356 (O_356,N_9932,N_9886);
nand UO_357 (O_357,N_9943,N_9930);
or UO_358 (O_358,N_9997,N_9970);
nor UO_359 (O_359,N_9856,N_9927);
or UO_360 (O_360,N_9888,N_9984);
nand UO_361 (O_361,N_9950,N_9942);
nand UO_362 (O_362,N_9808,N_9940);
nand UO_363 (O_363,N_9852,N_9876);
nor UO_364 (O_364,N_9972,N_9870);
nor UO_365 (O_365,N_9815,N_9989);
nor UO_366 (O_366,N_9944,N_9916);
nor UO_367 (O_367,N_9847,N_9947);
and UO_368 (O_368,N_9818,N_9933);
and UO_369 (O_369,N_9814,N_9922);
or UO_370 (O_370,N_9924,N_9836);
xnor UO_371 (O_371,N_9905,N_9890);
xnor UO_372 (O_372,N_9867,N_9827);
and UO_373 (O_373,N_9879,N_9847);
nand UO_374 (O_374,N_9955,N_9908);
nor UO_375 (O_375,N_9902,N_9982);
xor UO_376 (O_376,N_9814,N_9877);
nor UO_377 (O_377,N_9863,N_9818);
or UO_378 (O_378,N_9835,N_9976);
xnor UO_379 (O_379,N_9912,N_9871);
and UO_380 (O_380,N_9932,N_9806);
or UO_381 (O_381,N_9863,N_9813);
xor UO_382 (O_382,N_9807,N_9994);
xnor UO_383 (O_383,N_9972,N_9919);
xnor UO_384 (O_384,N_9990,N_9916);
or UO_385 (O_385,N_9945,N_9822);
nor UO_386 (O_386,N_9882,N_9972);
nand UO_387 (O_387,N_9969,N_9924);
and UO_388 (O_388,N_9843,N_9908);
nor UO_389 (O_389,N_9972,N_9978);
nor UO_390 (O_390,N_9842,N_9928);
and UO_391 (O_391,N_9961,N_9943);
xnor UO_392 (O_392,N_9951,N_9980);
xnor UO_393 (O_393,N_9802,N_9897);
xnor UO_394 (O_394,N_9871,N_9844);
nand UO_395 (O_395,N_9924,N_9824);
xor UO_396 (O_396,N_9985,N_9947);
nand UO_397 (O_397,N_9913,N_9964);
and UO_398 (O_398,N_9815,N_9958);
or UO_399 (O_399,N_9863,N_9916);
nand UO_400 (O_400,N_9914,N_9878);
xnor UO_401 (O_401,N_9867,N_9941);
xnor UO_402 (O_402,N_9903,N_9912);
and UO_403 (O_403,N_9901,N_9872);
nand UO_404 (O_404,N_9948,N_9905);
and UO_405 (O_405,N_9929,N_9948);
nand UO_406 (O_406,N_9851,N_9903);
or UO_407 (O_407,N_9997,N_9860);
nand UO_408 (O_408,N_9822,N_9866);
nor UO_409 (O_409,N_9844,N_9828);
or UO_410 (O_410,N_9857,N_9980);
nor UO_411 (O_411,N_9862,N_9908);
nand UO_412 (O_412,N_9904,N_9870);
nor UO_413 (O_413,N_9979,N_9824);
and UO_414 (O_414,N_9850,N_9838);
nor UO_415 (O_415,N_9812,N_9804);
nor UO_416 (O_416,N_9812,N_9840);
nand UO_417 (O_417,N_9986,N_9887);
or UO_418 (O_418,N_9976,N_9972);
and UO_419 (O_419,N_9861,N_9968);
nand UO_420 (O_420,N_9866,N_9870);
nand UO_421 (O_421,N_9940,N_9907);
nor UO_422 (O_422,N_9861,N_9858);
nand UO_423 (O_423,N_9966,N_9977);
nor UO_424 (O_424,N_9900,N_9952);
xnor UO_425 (O_425,N_9933,N_9972);
or UO_426 (O_426,N_9938,N_9831);
xor UO_427 (O_427,N_9898,N_9816);
nor UO_428 (O_428,N_9896,N_9879);
nand UO_429 (O_429,N_9908,N_9881);
xnor UO_430 (O_430,N_9945,N_9828);
or UO_431 (O_431,N_9845,N_9918);
and UO_432 (O_432,N_9885,N_9920);
or UO_433 (O_433,N_9874,N_9994);
nor UO_434 (O_434,N_9801,N_9823);
or UO_435 (O_435,N_9858,N_9931);
nor UO_436 (O_436,N_9864,N_9829);
nor UO_437 (O_437,N_9900,N_9926);
xor UO_438 (O_438,N_9976,N_9899);
and UO_439 (O_439,N_9985,N_9973);
nor UO_440 (O_440,N_9822,N_9876);
and UO_441 (O_441,N_9924,N_9875);
xor UO_442 (O_442,N_9970,N_9804);
nor UO_443 (O_443,N_9947,N_9964);
nand UO_444 (O_444,N_9901,N_9835);
nor UO_445 (O_445,N_9944,N_9935);
nor UO_446 (O_446,N_9979,N_9932);
and UO_447 (O_447,N_9899,N_9957);
and UO_448 (O_448,N_9948,N_9970);
or UO_449 (O_449,N_9857,N_9879);
or UO_450 (O_450,N_9929,N_9802);
or UO_451 (O_451,N_9870,N_9818);
xnor UO_452 (O_452,N_9891,N_9970);
nor UO_453 (O_453,N_9846,N_9817);
xor UO_454 (O_454,N_9951,N_9889);
nand UO_455 (O_455,N_9891,N_9832);
nor UO_456 (O_456,N_9915,N_9844);
xor UO_457 (O_457,N_9937,N_9810);
nand UO_458 (O_458,N_9843,N_9995);
or UO_459 (O_459,N_9828,N_9874);
or UO_460 (O_460,N_9872,N_9804);
and UO_461 (O_461,N_9811,N_9984);
or UO_462 (O_462,N_9902,N_9808);
or UO_463 (O_463,N_9813,N_9910);
nand UO_464 (O_464,N_9805,N_9993);
nor UO_465 (O_465,N_9833,N_9912);
xnor UO_466 (O_466,N_9878,N_9862);
and UO_467 (O_467,N_9968,N_9902);
or UO_468 (O_468,N_9930,N_9840);
nand UO_469 (O_469,N_9916,N_9875);
nand UO_470 (O_470,N_9935,N_9966);
and UO_471 (O_471,N_9925,N_9883);
or UO_472 (O_472,N_9883,N_9920);
nand UO_473 (O_473,N_9931,N_9821);
xnor UO_474 (O_474,N_9919,N_9915);
nand UO_475 (O_475,N_9984,N_9800);
and UO_476 (O_476,N_9808,N_9875);
nor UO_477 (O_477,N_9833,N_9847);
nor UO_478 (O_478,N_9896,N_9958);
nand UO_479 (O_479,N_9983,N_9882);
nor UO_480 (O_480,N_9815,N_9929);
nand UO_481 (O_481,N_9891,N_9904);
nor UO_482 (O_482,N_9936,N_9907);
nor UO_483 (O_483,N_9907,N_9915);
nand UO_484 (O_484,N_9960,N_9864);
and UO_485 (O_485,N_9931,N_9872);
and UO_486 (O_486,N_9986,N_9916);
nand UO_487 (O_487,N_9856,N_9849);
and UO_488 (O_488,N_9923,N_9815);
and UO_489 (O_489,N_9962,N_9854);
xnor UO_490 (O_490,N_9938,N_9812);
nand UO_491 (O_491,N_9957,N_9862);
nor UO_492 (O_492,N_9860,N_9979);
xnor UO_493 (O_493,N_9984,N_9815);
and UO_494 (O_494,N_9901,N_9887);
nor UO_495 (O_495,N_9821,N_9917);
xor UO_496 (O_496,N_9921,N_9845);
nand UO_497 (O_497,N_9875,N_9872);
and UO_498 (O_498,N_9846,N_9905);
and UO_499 (O_499,N_9995,N_9854);
xor UO_500 (O_500,N_9976,N_9934);
xor UO_501 (O_501,N_9970,N_9989);
xor UO_502 (O_502,N_9878,N_9992);
xor UO_503 (O_503,N_9838,N_9846);
nor UO_504 (O_504,N_9936,N_9910);
xor UO_505 (O_505,N_9849,N_9984);
xor UO_506 (O_506,N_9842,N_9980);
nor UO_507 (O_507,N_9940,N_9858);
and UO_508 (O_508,N_9887,N_9905);
nand UO_509 (O_509,N_9854,N_9853);
nor UO_510 (O_510,N_9812,N_9813);
nand UO_511 (O_511,N_9941,N_9947);
nor UO_512 (O_512,N_9984,N_9877);
and UO_513 (O_513,N_9873,N_9972);
or UO_514 (O_514,N_9880,N_9942);
nand UO_515 (O_515,N_9800,N_9999);
and UO_516 (O_516,N_9841,N_9803);
nor UO_517 (O_517,N_9848,N_9859);
nand UO_518 (O_518,N_9864,N_9844);
and UO_519 (O_519,N_9960,N_9943);
or UO_520 (O_520,N_9937,N_9960);
and UO_521 (O_521,N_9816,N_9978);
and UO_522 (O_522,N_9982,N_9806);
and UO_523 (O_523,N_9990,N_9970);
nor UO_524 (O_524,N_9863,N_9914);
and UO_525 (O_525,N_9841,N_9953);
nand UO_526 (O_526,N_9831,N_9876);
or UO_527 (O_527,N_9979,N_9846);
nand UO_528 (O_528,N_9887,N_9946);
or UO_529 (O_529,N_9859,N_9956);
nor UO_530 (O_530,N_9970,N_9887);
nand UO_531 (O_531,N_9933,N_9832);
xnor UO_532 (O_532,N_9870,N_9913);
and UO_533 (O_533,N_9828,N_9878);
nor UO_534 (O_534,N_9981,N_9811);
and UO_535 (O_535,N_9941,N_9925);
and UO_536 (O_536,N_9898,N_9965);
and UO_537 (O_537,N_9938,N_9804);
or UO_538 (O_538,N_9924,N_9970);
or UO_539 (O_539,N_9969,N_9907);
xor UO_540 (O_540,N_9995,N_9945);
xor UO_541 (O_541,N_9980,N_9863);
nor UO_542 (O_542,N_9967,N_9909);
xnor UO_543 (O_543,N_9873,N_9841);
and UO_544 (O_544,N_9891,N_9993);
and UO_545 (O_545,N_9812,N_9955);
or UO_546 (O_546,N_9935,N_9874);
nand UO_547 (O_547,N_9977,N_9859);
xnor UO_548 (O_548,N_9893,N_9972);
or UO_549 (O_549,N_9943,N_9936);
or UO_550 (O_550,N_9940,N_9978);
and UO_551 (O_551,N_9871,N_9928);
nand UO_552 (O_552,N_9847,N_9939);
xor UO_553 (O_553,N_9852,N_9951);
and UO_554 (O_554,N_9862,N_9813);
nand UO_555 (O_555,N_9899,N_9988);
nor UO_556 (O_556,N_9995,N_9998);
xor UO_557 (O_557,N_9925,N_9863);
nand UO_558 (O_558,N_9821,N_9960);
or UO_559 (O_559,N_9979,N_9962);
nor UO_560 (O_560,N_9827,N_9997);
nor UO_561 (O_561,N_9844,N_9944);
or UO_562 (O_562,N_9999,N_9981);
or UO_563 (O_563,N_9917,N_9989);
and UO_564 (O_564,N_9829,N_9872);
nor UO_565 (O_565,N_9983,N_9828);
or UO_566 (O_566,N_9863,N_9873);
nand UO_567 (O_567,N_9801,N_9986);
or UO_568 (O_568,N_9954,N_9894);
or UO_569 (O_569,N_9810,N_9997);
nand UO_570 (O_570,N_9901,N_9850);
and UO_571 (O_571,N_9985,N_9809);
nor UO_572 (O_572,N_9890,N_9972);
or UO_573 (O_573,N_9873,N_9998);
xnor UO_574 (O_574,N_9918,N_9980);
or UO_575 (O_575,N_9916,N_9984);
and UO_576 (O_576,N_9971,N_9848);
xor UO_577 (O_577,N_9847,N_9860);
xnor UO_578 (O_578,N_9965,N_9932);
and UO_579 (O_579,N_9969,N_9939);
nor UO_580 (O_580,N_9915,N_9841);
and UO_581 (O_581,N_9871,N_9960);
nand UO_582 (O_582,N_9919,N_9876);
or UO_583 (O_583,N_9990,N_9932);
xnor UO_584 (O_584,N_9960,N_9854);
or UO_585 (O_585,N_9897,N_9978);
nand UO_586 (O_586,N_9828,N_9877);
nor UO_587 (O_587,N_9835,N_9814);
or UO_588 (O_588,N_9802,N_9927);
nor UO_589 (O_589,N_9984,N_9867);
nor UO_590 (O_590,N_9989,N_9983);
nor UO_591 (O_591,N_9991,N_9919);
xnor UO_592 (O_592,N_9977,N_9861);
nand UO_593 (O_593,N_9918,N_9894);
nand UO_594 (O_594,N_9944,N_9881);
and UO_595 (O_595,N_9848,N_9913);
xnor UO_596 (O_596,N_9836,N_9942);
and UO_597 (O_597,N_9824,N_9853);
and UO_598 (O_598,N_9922,N_9968);
or UO_599 (O_599,N_9867,N_9939);
nor UO_600 (O_600,N_9842,N_9843);
xnor UO_601 (O_601,N_9932,N_9801);
or UO_602 (O_602,N_9814,N_9929);
nor UO_603 (O_603,N_9814,N_9833);
nand UO_604 (O_604,N_9893,N_9815);
nor UO_605 (O_605,N_9882,N_9911);
xor UO_606 (O_606,N_9867,N_9920);
xnor UO_607 (O_607,N_9906,N_9899);
nor UO_608 (O_608,N_9895,N_9968);
nand UO_609 (O_609,N_9846,N_9999);
and UO_610 (O_610,N_9906,N_9995);
xor UO_611 (O_611,N_9889,N_9905);
xor UO_612 (O_612,N_9981,N_9822);
nor UO_613 (O_613,N_9859,N_9998);
xnor UO_614 (O_614,N_9985,N_9818);
nor UO_615 (O_615,N_9837,N_9804);
nand UO_616 (O_616,N_9888,N_9963);
xor UO_617 (O_617,N_9903,N_9885);
xor UO_618 (O_618,N_9906,N_9842);
nand UO_619 (O_619,N_9947,N_9971);
and UO_620 (O_620,N_9836,N_9806);
and UO_621 (O_621,N_9926,N_9915);
nand UO_622 (O_622,N_9801,N_9830);
nand UO_623 (O_623,N_9921,N_9977);
nand UO_624 (O_624,N_9947,N_9838);
xor UO_625 (O_625,N_9900,N_9994);
nand UO_626 (O_626,N_9826,N_9861);
nand UO_627 (O_627,N_9990,N_9906);
xnor UO_628 (O_628,N_9821,N_9930);
nor UO_629 (O_629,N_9986,N_9871);
xnor UO_630 (O_630,N_9947,N_9870);
nor UO_631 (O_631,N_9918,N_9975);
xnor UO_632 (O_632,N_9936,N_9977);
xnor UO_633 (O_633,N_9870,N_9908);
xor UO_634 (O_634,N_9976,N_9824);
and UO_635 (O_635,N_9970,N_9938);
and UO_636 (O_636,N_9939,N_9886);
or UO_637 (O_637,N_9825,N_9968);
nand UO_638 (O_638,N_9800,N_9819);
xnor UO_639 (O_639,N_9958,N_9830);
and UO_640 (O_640,N_9915,N_9980);
xor UO_641 (O_641,N_9946,N_9839);
nor UO_642 (O_642,N_9845,N_9887);
nor UO_643 (O_643,N_9941,N_9855);
nand UO_644 (O_644,N_9820,N_9951);
nand UO_645 (O_645,N_9976,N_9916);
xor UO_646 (O_646,N_9816,N_9830);
or UO_647 (O_647,N_9950,N_9878);
nor UO_648 (O_648,N_9924,N_9811);
and UO_649 (O_649,N_9827,N_9887);
nand UO_650 (O_650,N_9967,N_9908);
and UO_651 (O_651,N_9892,N_9940);
nand UO_652 (O_652,N_9891,N_9822);
or UO_653 (O_653,N_9936,N_9962);
nor UO_654 (O_654,N_9804,N_9863);
nor UO_655 (O_655,N_9845,N_9854);
and UO_656 (O_656,N_9937,N_9856);
xnor UO_657 (O_657,N_9948,N_9836);
and UO_658 (O_658,N_9985,N_9856);
or UO_659 (O_659,N_9808,N_9854);
nand UO_660 (O_660,N_9949,N_9966);
nor UO_661 (O_661,N_9832,N_9839);
or UO_662 (O_662,N_9918,N_9900);
or UO_663 (O_663,N_9927,N_9924);
or UO_664 (O_664,N_9855,N_9845);
and UO_665 (O_665,N_9950,N_9822);
nand UO_666 (O_666,N_9836,N_9821);
nor UO_667 (O_667,N_9816,N_9906);
nor UO_668 (O_668,N_9807,N_9802);
nor UO_669 (O_669,N_9804,N_9847);
nor UO_670 (O_670,N_9990,N_9868);
xnor UO_671 (O_671,N_9956,N_9985);
and UO_672 (O_672,N_9999,N_9869);
nand UO_673 (O_673,N_9978,N_9875);
nand UO_674 (O_674,N_9986,N_9946);
and UO_675 (O_675,N_9813,N_9979);
nand UO_676 (O_676,N_9850,N_9903);
xnor UO_677 (O_677,N_9985,N_9853);
nand UO_678 (O_678,N_9862,N_9931);
and UO_679 (O_679,N_9971,N_9902);
xor UO_680 (O_680,N_9876,N_9908);
nor UO_681 (O_681,N_9964,N_9992);
nor UO_682 (O_682,N_9837,N_9985);
nand UO_683 (O_683,N_9887,N_9980);
nor UO_684 (O_684,N_9985,N_9944);
nor UO_685 (O_685,N_9838,N_9839);
nor UO_686 (O_686,N_9985,N_9909);
nand UO_687 (O_687,N_9888,N_9986);
or UO_688 (O_688,N_9926,N_9914);
nand UO_689 (O_689,N_9816,N_9847);
or UO_690 (O_690,N_9823,N_9802);
xnor UO_691 (O_691,N_9928,N_9915);
nor UO_692 (O_692,N_9960,N_9995);
and UO_693 (O_693,N_9942,N_9924);
nor UO_694 (O_694,N_9809,N_9908);
xnor UO_695 (O_695,N_9891,N_9911);
nor UO_696 (O_696,N_9813,N_9823);
or UO_697 (O_697,N_9856,N_9807);
xor UO_698 (O_698,N_9961,N_9888);
xnor UO_699 (O_699,N_9979,N_9974);
nor UO_700 (O_700,N_9973,N_9972);
and UO_701 (O_701,N_9877,N_9851);
xor UO_702 (O_702,N_9948,N_9913);
xor UO_703 (O_703,N_9923,N_9926);
or UO_704 (O_704,N_9975,N_9914);
nand UO_705 (O_705,N_9971,N_9849);
and UO_706 (O_706,N_9899,N_9928);
xnor UO_707 (O_707,N_9819,N_9994);
nand UO_708 (O_708,N_9810,N_9875);
nand UO_709 (O_709,N_9844,N_9897);
nand UO_710 (O_710,N_9941,N_9907);
nand UO_711 (O_711,N_9902,N_9962);
and UO_712 (O_712,N_9968,N_9926);
nand UO_713 (O_713,N_9940,N_9931);
nor UO_714 (O_714,N_9883,N_9957);
nor UO_715 (O_715,N_9905,N_9828);
nand UO_716 (O_716,N_9981,N_9952);
nor UO_717 (O_717,N_9991,N_9905);
xnor UO_718 (O_718,N_9992,N_9860);
nor UO_719 (O_719,N_9925,N_9973);
or UO_720 (O_720,N_9948,N_9846);
xor UO_721 (O_721,N_9910,N_9906);
nor UO_722 (O_722,N_9840,N_9928);
and UO_723 (O_723,N_9993,N_9822);
nand UO_724 (O_724,N_9876,N_9839);
or UO_725 (O_725,N_9935,N_9879);
nand UO_726 (O_726,N_9877,N_9991);
nand UO_727 (O_727,N_9937,N_9936);
or UO_728 (O_728,N_9991,N_9933);
or UO_729 (O_729,N_9906,N_9865);
nor UO_730 (O_730,N_9990,N_9942);
nor UO_731 (O_731,N_9811,N_9898);
xor UO_732 (O_732,N_9915,N_9871);
nand UO_733 (O_733,N_9844,N_9819);
or UO_734 (O_734,N_9957,N_9848);
xnor UO_735 (O_735,N_9908,N_9893);
and UO_736 (O_736,N_9973,N_9833);
or UO_737 (O_737,N_9828,N_9896);
nand UO_738 (O_738,N_9869,N_9995);
or UO_739 (O_739,N_9903,N_9856);
nor UO_740 (O_740,N_9911,N_9888);
nor UO_741 (O_741,N_9822,N_9921);
and UO_742 (O_742,N_9991,N_9847);
nand UO_743 (O_743,N_9921,N_9988);
and UO_744 (O_744,N_9829,N_9815);
or UO_745 (O_745,N_9978,N_9817);
and UO_746 (O_746,N_9939,N_9921);
nand UO_747 (O_747,N_9889,N_9847);
nor UO_748 (O_748,N_9820,N_9800);
and UO_749 (O_749,N_9946,N_9873);
xnor UO_750 (O_750,N_9895,N_9815);
nand UO_751 (O_751,N_9820,N_9955);
nor UO_752 (O_752,N_9921,N_9940);
and UO_753 (O_753,N_9886,N_9961);
or UO_754 (O_754,N_9886,N_9998);
and UO_755 (O_755,N_9906,N_9814);
nor UO_756 (O_756,N_9874,N_9826);
nor UO_757 (O_757,N_9990,N_9845);
nor UO_758 (O_758,N_9970,N_9915);
xnor UO_759 (O_759,N_9809,N_9948);
xnor UO_760 (O_760,N_9865,N_9836);
and UO_761 (O_761,N_9919,N_9968);
or UO_762 (O_762,N_9891,N_9926);
or UO_763 (O_763,N_9957,N_9803);
or UO_764 (O_764,N_9852,N_9959);
nand UO_765 (O_765,N_9883,N_9999);
and UO_766 (O_766,N_9818,N_9825);
or UO_767 (O_767,N_9858,N_9870);
and UO_768 (O_768,N_9834,N_9864);
and UO_769 (O_769,N_9800,N_9993);
or UO_770 (O_770,N_9978,N_9867);
xnor UO_771 (O_771,N_9948,N_9841);
nand UO_772 (O_772,N_9832,N_9949);
or UO_773 (O_773,N_9827,N_9818);
nor UO_774 (O_774,N_9853,N_9857);
or UO_775 (O_775,N_9931,N_9985);
xnor UO_776 (O_776,N_9811,N_9854);
and UO_777 (O_777,N_9952,N_9936);
or UO_778 (O_778,N_9851,N_9960);
xor UO_779 (O_779,N_9833,N_9825);
nor UO_780 (O_780,N_9891,N_9985);
nor UO_781 (O_781,N_9982,N_9904);
nand UO_782 (O_782,N_9896,N_9864);
or UO_783 (O_783,N_9829,N_9993);
xnor UO_784 (O_784,N_9864,N_9825);
nor UO_785 (O_785,N_9803,N_9806);
xor UO_786 (O_786,N_9946,N_9863);
or UO_787 (O_787,N_9902,N_9975);
nor UO_788 (O_788,N_9967,N_9927);
or UO_789 (O_789,N_9815,N_9826);
nor UO_790 (O_790,N_9808,N_9908);
and UO_791 (O_791,N_9838,N_9901);
xnor UO_792 (O_792,N_9992,N_9872);
nor UO_793 (O_793,N_9883,N_9933);
nor UO_794 (O_794,N_9973,N_9862);
xnor UO_795 (O_795,N_9927,N_9825);
or UO_796 (O_796,N_9885,N_9973);
or UO_797 (O_797,N_9969,N_9881);
xor UO_798 (O_798,N_9848,N_9973);
nor UO_799 (O_799,N_9809,N_9812);
or UO_800 (O_800,N_9994,N_9980);
or UO_801 (O_801,N_9913,N_9833);
nand UO_802 (O_802,N_9841,N_9949);
or UO_803 (O_803,N_9867,N_9832);
nor UO_804 (O_804,N_9970,N_9986);
or UO_805 (O_805,N_9859,N_9955);
and UO_806 (O_806,N_9911,N_9978);
or UO_807 (O_807,N_9851,N_9907);
and UO_808 (O_808,N_9887,N_9974);
nor UO_809 (O_809,N_9954,N_9830);
and UO_810 (O_810,N_9859,N_9879);
or UO_811 (O_811,N_9822,N_9995);
xnor UO_812 (O_812,N_9860,N_9834);
or UO_813 (O_813,N_9805,N_9898);
and UO_814 (O_814,N_9954,N_9859);
nor UO_815 (O_815,N_9897,N_9808);
and UO_816 (O_816,N_9933,N_9900);
xor UO_817 (O_817,N_9960,N_9977);
nor UO_818 (O_818,N_9927,N_9971);
nand UO_819 (O_819,N_9839,N_9978);
nor UO_820 (O_820,N_9945,N_9851);
nor UO_821 (O_821,N_9812,N_9866);
xor UO_822 (O_822,N_9827,N_9823);
nor UO_823 (O_823,N_9961,N_9838);
nor UO_824 (O_824,N_9829,N_9883);
nor UO_825 (O_825,N_9957,N_9967);
nor UO_826 (O_826,N_9892,N_9837);
xnor UO_827 (O_827,N_9840,N_9802);
nand UO_828 (O_828,N_9886,N_9917);
and UO_829 (O_829,N_9849,N_9915);
or UO_830 (O_830,N_9986,N_9868);
xor UO_831 (O_831,N_9944,N_9977);
xnor UO_832 (O_832,N_9844,N_9951);
xor UO_833 (O_833,N_9881,N_9892);
or UO_834 (O_834,N_9939,N_9897);
and UO_835 (O_835,N_9984,N_9833);
xnor UO_836 (O_836,N_9946,N_9920);
xnor UO_837 (O_837,N_9902,N_9948);
xor UO_838 (O_838,N_9905,N_9966);
nand UO_839 (O_839,N_9826,N_9838);
nor UO_840 (O_840,N_9853,N_9897);
nand UO_841 (O_841,N_9866,N_9847);
xor UO_842 (O_842,N_9934,N_9857);
nor UO_843 (O_843,N_9926,N_9901);
xor UO_844 (O_844,N_9862,N_9917);
and UO_845 (O_845,N_9901,N_9964);
or UO_846 (O_846,N_9994,N_9847);
nor UO_847 (O_847,N_9970,N_9893);
and UO_848 (O_848,N_9846,N_9919);
nor UO_849 (O_849,N_9852,N_9865);
nor UO_850 (O_850,N_9984,N_9874);
xnor UO_851 (O_851,N_9857,N_9886);
nor UO_852 (O_852,N_9810,N_9999);
and UO_853 (O_853,N_9852,N_9958);
xnor UO_854 (O_854,N_9973,N_9923);
nand UO_855 (O_855,N_9994,N_9905);
nor UO_856 (O_856,N_9987,N_9899);
nor UO_857 (O_857,N_9841,N_9955);
nor UO_858 (O_858,N_9973,N_9950);
or UO_859 (O_859,N_9927,N_9925);
or UO_860 (O_860,N_9968,N_9819);
xnor UO_861 (O_861,N_9992,N_9970);
and UO_862 (O_862,N_9917,N_9904);
or UO_863 (O_863,N_9832,N_9966);
nor UO_864 (O_864,N_9979,N_9823);
nor UO_865 (O_865,N_9808,N_9883);
and UO_866 (O_866,N_9867,N_9861);
nor UO_867 (O_867,N_9863,N_9872);
nand UO_868 (O_868,N_9964,N_9995);
nand UO_869 (O_869,N_9812,N_9990);
or UO_870 (O_870,N_9814,N_9959);
or UO_871 (O_871,N_9922,N_9813);
xor UO_872 (O_872,N_9935,N_9852);
and UO_873 (O_873,N_9917,N_9812);
or UO_874 (O_874,N_9873,N_9973);
xnor UO_875 (O_875,N_9905,N_9803);
nor UO_876 (O_876,N_9802,N_9932);
and UO_877 (O_877,N_9850,N_9908);
xor UO_878 (O_878,N_9910,N_9888);
and UO_879 (O_879,N_9919,N_9969);
and UO_880 (O_880,N_9994,N_9817);
nor UO_881 (O_881,N_9819,N_9896);
xor UO_882 (O_882,N_9816,N_9864);
or UO_883 (O_883,N_9843,N_9927);
nor UO_884 (O_884,N_9840,N_9878);
nand UO_885 (O_885,N_9807,N_9811);
or UO_886 (O_886,N_9965,N_9945);
and UO_887 (O_887,N_9852,N_9919);
and UO_888 (O_888,N_9888,N_9903);
nand UO_889 (O_889,N_9902,N_9814);
nor UO_890 (O_890,N_9997,N_9946);
and UO_891 (O_891,N_9836,N_9831);
nand UO_892 (O_892,N_9802,N_9873);
xnor UO_893 (O_893,N_9972,N_9975);
nor UO_894 (O_894,N_9963,N_9981);
or UO_895 (O_895,N_9956,N_9849);
or UO_896 (O_896,N_9902,N_9820);
or UO_897 (O_897,N_9846,N_9847);
or UO_898 (O_898,N_9929,N_9852);
nor UO_899 (O_899,N_9809,N_9923);
xor UO_900 (O_900,N_9821,N_9818);
nand UO_901 (O_901,N_9940,N_9873);
or UO_902 (O_902,N_9868,N_9945);
nand UO_903 (O_903,N_9936,N_9915);
or UO_904 (O_904,N_9865,N_9903);
and UO_905 (O_905,N_9863,N_9831);
nor UO_906 (O_906,N_9909,N_9893);
xor UO_907 (O_907,N_9891,N_9906);
and UO_908 (O_908,N_9910,N_9989);
or UO_909 (O_909,N_9994,N_9967);
and UO_910 (O_910,N_9960,N_9984);
or UO_911 (O_911,N_9879,N_9815);
nand UO_912 (O_912,N_9987,N_9924);
nand UO_913 (O_913,N_9951,N_9874);
nor UO_914 (O_914,N_9823,N_9980);
nor UO_915 (O_915,N_9991,N_9832);
xor UO_916 (O_916,N_9902,N_9803);
and UO_917 (O_917,N_9879,N_9867);
nor UO_918 (O_918,N_9855,N_9925);
xnor UO_919 (O_919,N_9926,N_9992);
nand UO_920 (O_920,N_9821,N_9893);
nand UO_921 (O_921,N_9963,N_9813);
or UO_922 (O_922,N_9929,N_9975);
nor UO_923 (O_923,N_9804,N_9911);
xnor UO_924 (O_924,N_9971,N_9867);
xor UO_925 (O_925,N_9816,N_9937);
nand UO_926 (O_926,N_9945,N_9838);
or UO_927 (O_927,N_9992,N_9859);
nor UO_928 (O_928,N_9848,N_9815);
xnor UO_929 (O_929,N_9964,N_9910);
and UO_930 (O_930,N_9903,N_9919);
nand UO_931 (O_931,N_9906,N_9852);
nor UO_932 (O_932,N_9814,N_9843);
nor UO_933 (O_933,N_9800,N_9876);
xor UO_934 (O_934,N_9836,N_9982);
or UO_935 (O_935,N_9983,N_9961);
nor UO_936 (O_936,N_9968,N_9880);
and UO_937 (O_937,N_9909,N_9928);
and UO_938 (O_938,N_9863,N_9993);
or UO_939 (O_939,N_9861,N_9813);
nor UO_940 (O_940,N_9824,N_9971);
xor UO_941 (O_941,N_9860,N_9893);
or UO_942 (O_942,N_9901,N_9932);
and UO_943 (O_943,N_9840,N_9847);
xor UO_944 (O_944,N_9833,N_9969);
xnor UO_945 (O_945,N_9812,N_9883);
nand UO_946 (O_946,N_9882,N_9821);
or UO_947 (O_947,N_9959,N_9914);
xnor UO_948 (O_948,N_9847,N_9931);
or UO_949 (O_949,N_9944,N_9964);
or UO_950 (O_950,N_9961,N_9889);
xnor UO_951 (O_951,N_9812,N_9857);
nand UO_952 (O_952,N_9918,N_9831);
and UO_953 (O_953,N_9994,N_9989);
and UO_954 (O_954,N_9934,N_9854);
nand UO_955 (O_955,N_9992,N_9803);
xor UO_956 (O_956,N_9875,N_9813);
nor UO_957 (O_957,N_9928,N_9904);
and UO_958 (O_958,N_9899,N_9936);
nand UO_959 (O_959,N_9909,N_9856);
xor UO_960 (O_960,N_9940,N_9982);
nand UO_961 (O_961,N_9841,N_9914);
or UO_962 (O_962,N_9810,N_9974);
or UO_963 (O_963,N_9999,N_9912);
xnor UO_964 (O_964,N_9932,N_9880);
xor UO_965 (O_965,N_9805,N_9855);
nor UO_966 (O_966,N_9827,N_9931);
and UO_967 (O_967,N_9948,N_9987);
and UO_968 (O_968,N_9838,N_9939);
nand UO_969 (O_969,N_9927,N_9840);
xnor UO_970 (O_970,N_9800,N_9905);
nor UO_971 (O_971,N_9803,N_9930);
or UO_972 (O_972,N_9819,N_9976);
and UO_973 (O_973,N_9823,N_9917);
or UO_974 (O_974,N_9801,N_9838);
xor UO_975 (O_975,N_9886,N_9834);
nand UO_976 (O_976,N_9920,N_9923);
or UO_977 (O_977,N_9918,N_9819);
xor UO_978 (O_978,N_9981,N_9990);
nor UO_979 (O_979,N_9877,N_9921);
or UO_980 (O_980,N_9922,N_9983);
or UO_981 (O_981,N_9818,N_9901);
xor UO_982 (O_982,N_9873,N_9839);
and UO_983 (O_983,N_9804,N_9933);
nand UO_984 (O_984,N_9855,N_9958);
xnor UO_985 (O_985,N_9921,N_9871);
and UO_986 (O_986,N_9810,N_9886);
and UO_987 (O_987,N_9924,N_9976);
xnor UO_988 (O_988,N_9895,N_9803);
xor UO_989 (O_989,N_9851,N_9869);
xnor UO_990 (O_990,N_9805,N_9810);
and UO_991 (O_991,N_9906,N_9991);
nand UO_992 (O_992,N_9965,N_9921);
nor UO_993 (O_993,N_9878,N_9883);
xor UO_994 (O_994,N_9875,N_9972);
nand UO_995 (O_995,N_9851,N_9983);
nor UO_996 (O_996,N_9982,N_9877);
nor UO_997 (O_997,N_9910,N_9881);
or UO_998 (O_998,N_9840,N_9832);
or UO_999 (O_999,N_9995,N_9838);
nand UO_1000 (O_1000,N_9979,N_9999);
xnor UO_1001 (O_1001,N_9932,N_9972);
and UO_1002 (O_1002,N_9989,N_9961);
and UO_1003 (O_1003,N_9868,N_9903);
xnor UO_1004 (O_1004,N_9999,N_9879);
nand UO_1005 (O_1005,N_9840,N_9866);
nor UO_1006 (O_1006,N_9905,N_9986);
or UO_1007 (O_1007,N_9998,N_9907);
nor UO_1008 (O_1008,N_9869,N_9812);
nor UO_1009 (O_1009,N_9873,N_9835);
or UO_1010 (O_1010,N_9815,N_9906);
or UO_1011 (O_1011,N_9863,N_9981);
nand UO_1012 (O_1012,N_9996,N_9845);
or UO_1013 (O_1013,N_9825,N_9959);
nor UO_1014 (O_1014,N_9926,N_9871);
xnor UO_1015 (O_1015,N_9908,N_9878);
nand UO_1016 (O_1016,N_9884,N_9809);
nand UO_1017 (O_1017,N_9972,N_9898);
or UO_1018 (O_1018,N_9869,N_9914);
xnor UO_1019 (O_1019,N_9870,N_9845);
or UO_1020 (O_1020,N_9876,N_9981);
or UO_1021 (O_1021,N_9848,N_9863);
xor UO_1022 (O_1022,N_9942,N_9908);
and UO_1023 (O_1023,N_9896,N_9935);
nor UO_1024 (O_1024,N_9925,N_9974);
nor UO_1025 (O_1025,N_9885,N_9871);
and UO_1026 (O_1026,N_9865,N_9928);
xnor UO_1027 (O_1027,N_9831,N_9942);
or UO_1028 (O_1028,N_9978,N_9833);
and UO_1029 (O_1029,N_9958,N_9823);
or UO_1030 (O_1030,N_9949,N_9927);
nand UO_1031 (O_1031,N_9920,N_9985);
nand UO_1032 (O_1032,N_9942,N_9957);
nand UO_1033 (O_1033,N_9888,N_9973);
nand UO_1034 (O_1034,N_9937,N_9921);
nand UO_1035 (O_1035,N_9992,N_9997);
xor UO_1036 (O_1036,N_9808,N_9987);
or UO_1037 (O_1037,N_9889,N_9988);
nand UO_1038 (O_1038,N_9952,N_9813);
xnor UO_1039 (O_1039,N_9960,N_9904);
xor UO_1040 (O_1040,N_9974,N_9878);
or UO_1041 (O_1041,N_9921,N_9874);
xor UO_1042 (O_1042,N_9962,N_9884);
and UO_1043 (O_1043,N_9960,N_9908);
xnor UO_1044 (O_1044,N_9952,N_9949);
nand UO_1045 (O_1045,N_9845,N_9942);
nor UO_1046 (O_1046,N_9825,N_9987);
or UO_1047 (O_1047,N_9842,N_9899);
xor UO_1048 (O_1048,N_9860,N_9918);
nand UO_1049 (O_1049,N_9844,N_9895);
xnor UO_1050 (O_1050,N_9910,N_9917);
and UO_1051 (O_1051,N_9807,N_9927);
nand UO_1052 (O_1052,N_9800,N_9897);
nor UO_1053 (O_1053,N_9985,N_9811);
xor UO_1054 (O_1054,N_9860,N_9949);
xnor UO_1055 (O_1055,N_9930,N_9926);
xnor UO_1056 (O_1056,N_9885,N_9938);
nor UO_1057 (O_1057,N_9823,N_9960);
and UO_1058 (O_1058,N_9871,N_9829);
nor UO_1059 (O_1059,N_9941,N_9948);
xor UO_1060 (O_1060,N_9981,N_9919);
or UO_1061 (O_1061,N_9956,N_9839);
and UO_1062 (O_1062,N_9914,N_9904);
nand UO_1063 (O_1063,N_9838,N_9821);
nand UO_1064 (O_1064,N_9977,N_9979);
or UO_1065 (O_1065,N_9987,N_9911);
and UO_1066 (O_1066,N_9874,N_9867);
and UO_1067 (O_1067,N_9914,N_9934);
nor UO_1068 (O_1068,N_9873,N_9950);
nand UO_1069 (O_1069,N_9873,N_9915);
or UO_1070 (O_1070,N_9970,N_9828);
and UO_1071 (O_1071,N_9917,N_9855);
and UO_1072 (O_1072,N_9882,N_9879);
and UO_1073 (O_1073,N_9812,N_9800);
and UO_1074 (O_1074,N_9853,N_9907);
xnor UO_1075 (O_1075,N_9942,N_9915);
or UO_1076 (O_1076,N_9906,N_9821);
nor UO_1077 (O_1077,N_9834,N_9946);
and UO_1078 (O_1078,N_9801,N_9800);
nand UO_1079 (O_1079,N_9883,N_9986);
and UO_1080 (O_1080,N_9827,N_9806);
nor UO_1081 (O_1081,N_9822,N_9965);
or UO_1082 (O_1082,N_9875,N_9817);
and UO_1083 (O_1083,N_9853,N_9906);
nor UO_1084 (O_1084,N_9894,N_9800);
and UO_1085 (O_1085,N_9926,N_9916);
or UO_1086 (O_1086,N_9953,N_9822);
nand UO_1087 (O_1087,N_9965,N_9993);
or UO_1088 (O_1088,N_9945,N_9858);
nor UO_1089 (O_1089,N_9884,N_9912);
or UO_1090 (O_1090,N_9815,N_9932);
xnor UO_1091 (O_1091,N_9932,N_9850);
and UO_1092 (O_1092,N_9809,N_9964);
nor UO_1093 (O_1093,N_9954,N_9831);
xor UO_1094 (O_1094,N_9947,N_9901);
nand UO_1095 (O_1095,N_9829,N_9873);
xnor UO_1096 (O_1096,N_9901,N_9906);
nand UO_1097 (O_1097,N_9929,N_9955);
nor UO_1098 (O_1098,N_9976,N_9983);
nor UO_1099 (O_1099,N_9985,N_9938);
xor UO_1100 (O_1100,N_9809,N_9983);
nor UO_1101 (O_1101,N_9990,N_9826);
and UO_1102 (O_1102,N_9878,N_9810);
or UO_1103 (O_1103,N_9995,N_9873);
nor UO_1104 (O_1104,N_9890,N_9989);
or UO_1105 (O_1105,N_9823,N_9981);
and UO_1106 (O_1106,N_9848,N_9904);
or UO_1107 (O_1107,N_9865,N_9967);
xnor UO_1108 (O_1108,N_9997,N_9965);
nand UO_1109 (O_1109,N_9801,N_9970);
nand UO_1110 (O_1110,N_9918,N_9840);
nor UO_1111 (O_1111,N_9943,N_9888);
xnor UO_1112 (O_1112,N_9818,N_9816);
nand UO_1113 (O_1113,N_9962,N_9993);
and UO_1114 (O_1114,N_9823,N_9804);
nor UO_1115 (O_1115,N_9884,N_9831);
nor UO_1116 (O_1116,N_9973,N_9960);
xnor UO_1117 (O_1117,N_9931,N_9973);
nor UO_1118 (O_1118,N_9832,N_9971);
or UO_1119 (O_1119,N_9956,N_9894);
or UO_1120 (O_1120,N_9871,N_9806);
xnor UO_1121 (O_1121,N_9973,N_9990);
or UO_1122 (O_1122,N_9996,N_9909);
or UO_1123 (O_1123,N_9914,N_9882);
and UO_1124 (O_1124,N_9888,N_9978);
nor UO_1125 (O_1125,N_9906,N_9823);
xnor UO_1126 (O_1126,N_9975,N_9835);
or UO_1127 (O_1127,N_9997,N_9932);
nand UO_1128 (O_1128,N_9836,N_9877);
xor UO_1129 (O_1129,N_9931,N_9852);
nor UO_1130 (O_1130,N_9822,N_9804);
nor UO_1131 (O_1131,N_9895,N_9823);
and UO_1132 (O_1132,N_9987,N_9938);
or UO_1133 (O_1133,N_9895,N_9972);
nand UO_1134 (O_1134,N_9926,N_9973);
xnor UO_1135 (O_1135,N_9906,N_9883);
nor UO_1136 (O_1136,N_9916,N_9974);
nand UO_1137 (O_1137,N_9927,N_9857);
or UO_1138 (O_1138,N_9915,N_9916);
xor UO_1139 (O_1139,N_9967,N_9943);
and UO_1140 (O_1140,N_9935,N_9920);
nand UO_1141 (O_1141,N_9888,N_9989);
nor UO_1142 (O_1142,N_9812,N_9826);
xnor UO_1143 (O_1143,N_9977,N_9939);
xor UO_1144 (O_1144,N_9983,N_9886);
nor UO_1145 (O_1145,N_9880,N_9850);
nand UO_1146 (O_1146,N_9973,N_9942);
xnor UO_1147 (O_1147,N_9936,N_9946);
or UO_1148 (O_1148,N_9818,N_9879);
nor UO_1149 (O_1149,N_9873,N_9996);
nor UO_1150 (O_1150,N_9891,N_9950);
xnor UO_1151 (O_1151,N_9880,N_9910);
nand UO_1152 (O_1152,N_9858,N_9943);
nand UO_1153 (O_1153,N_9941,N_9882);
and UO_1154 (O_1154,N_9837,N_9942);
xnor UO_1155 (O_1155,N_9812,N_9814);
or UO_1156 (O_1156,N_9901,N_9847);
xor UO_1157 (O_1157,N_9877,N_9890);
and UO_1158 (O_1158,N_9910,N_9953);
xnor UO_1159 (O_1159,N_9949,N_9872);
nand UO_1160 (O_1160,N_9804,N_9848);
nand UO_1161 (O_1161,N_9827,N_9965);
or UO_1162 (O_1162,N_9872,N_9905);
nor UO_1163 (O_1163,N_9879,N_9995);
nand UO_1164 (O_1164,N_9852,N_9927);
nor UO_1165 (O_1165,N_9880,N_9935);
xor UO_1166 (O_1166,N_9930,N_9928);
and UO_1167 (O_1167,N_9822,N_9849);
nand UO_1168 (O_1168,N_9841,N_9968);
nand UO_1169 (O_1169,N_9895,N_9875);
and UO_1170 (O_1170,N_9944,N_9911);
and UO_1171 (O_1171,N_9909,N_9869);
and UO_1172 (O_1172,N_9897,N_9884);
and UO_1173 (O_1173,N_9992,N_9928);
and UO_1174 (O_1174,N_9842,N_9861);
or UO_1175 (O_1175,N_9966,N_9931);
nand UO_1176 (O_1176,N_9832,N_9898);
nand UO_1177 (O_1177,N_9987,N_9868);
xor UO_1178 (O_1178,N_9982,N_9821);
and UO_1179 (O_1179,N_9971,N_9912);
nor UO_1180 (O_1180,N_9932,N_9822);
or UO_1181 (O_1181,N_9864,N_9893);
and UO_1182 (O_1182,N_9897,N_9983);
nand UO_1183 (O_1183,N_9980,N_9882);
nor UO_1184 (O_1184,N_9891,N_9934);
nor UO_1185 (O_1185,N_9956,N_9857);
nor UO_1186 (O_1186,N_9995,N_9961);
nor UO_1187 (O_1187,N_9914,N_9927);
xnor UO_1188 (O_1188,N_9941,N_9899);
and UO_1189 (O_1189,N_9805,N_9806);
and UO_1190 (O_1190,N_9864,N_9804);
xor UO_1191 (O_1191,N_9994,N_9825);
nand UO_1192 (O_1192,N_9931,N_9995);
and UO_1193 (O_1193,N_9883,N_9831);
xor UO_1194 (O_1194,N_9970,N_9882);
xnor UO_1195 (O_1195,N_9865,N_9969);
nor UO_1196 (O_1196,N_9866,N_9820);
or UO_1197 (O_1197,N_9954,N_9973);
and UO_1198 (O_1198,N_9977,N_9932);
nand UO_1199 (O_1199,N_9818,N_9857);
nor UO_1200 (O_1200,N_9824,N_9802);
nor UO_1201 (O_1201,N_9994,N_9929);
nor UO_1202 (O_1202,N_9941,N_9876);
and UO_1203 (O_1203,N_9897,N_9868);
xnor UO_1204 (O_1204,N_9834,N_9815);
nand UO_1205 (O_1205,N_9972,N_9891);
nor UO_1206 (O_1206,N_9916,N_9971);
and UO_1207 (O_1207,N_9926,N_9983);
and UO_1208 (O_1208,N_9998,N_9860);
nor UO_1209 (O_1209,N_9929,N_9906);
xor UO_1210 (O_1210,N_9821,N_9901);
nor UO_1211 (O_1211,N_9995,N_9889);
xor UO_1212 (O_1212,N_9849,N_9944);
or UO_1213 (O_1213,N_9874,N_9959);
and UO_1214 (O_1214,N_9863,N_9944);
and UO_1215 (O_1215,N_9891,N_9967);
xor UO_1216 (O_1216,N_9995,N_9992);
nor UO_1217 (O_1217,N_9841,N_9811);
nand UO_1218 (O_1218,N_9828,N_9822);
nor UO_1219 (O_1219,N_9851,N_9826);
nor UO_1220 (O_1220,N_9834,N_9810);
nand UO_1221 (O_1221,N_9890,N_9901);
nor UO_1222 (O_1222,N_9868,N_9919);
nand UO_1223 (O_1223,N_9888,N_9924);
or UO_1224 (O_1224,N_9841,N_9850);
or UO_1225 (O_1225,N_9910,N_9942);
nor UO_1226 (O_1226,N_9860,N_9845);
or UO_1227 (O_1227,N_9967,N_9901);
and UO_1228 (O_1228,N_9977,N_9883);
or UO_1229 (O_1229,N_9878,N_9933);
and UO_1230 (O_1230,N_9855,N_9927);
and UO_1231 (O_1231,N_9836,N_9871);
nand UO_1232 (O_1232,N_9943,N_9979);
nand UO_1233 (O_1233,N_9838,N_9960);
and UO_1234 (O_1234,N_9861,N_9917);
xor UO_1235 (O_1235,N_9893,N_9949);
nor UO_1236 (O_1236,N_9805,N_9895);
xor UO_1237 (O_1237,N_9890,N_9929);
and UO_1238 (O_1238,N_9960,N_9875);
nand UO_1239 (O_1239,N_9950,N_9958);
nand UO_1240 (O_1240,N_9888,N_9902);
and UO_1241 (O_1241,N_9805,N_9942);
or UO_1242 (O_1242,N_9866,N_9934);
and UO_1243 (O_1243,N_9843,N_9964);
and UO_1244 (O_1244,N_9960,N_9980);
or UO_1245 (O_1245,N_9987,N_9913);
nand UO_1246 (O_1246,N_9961,N_9940);
and UO_1247 (O_1247,N_9877,N_9929);
and UO_1248 (O_1248,N_9857,N_9831);
or UO_1249 (O_1249,N_9897,N_9874);
xnor UO_1250 (O_1250,N_9804,N_9867);
nand UO_1251 (O_1251,N_9947,N_9804);
xor UO_1252 (O_1252,N_9808,N_9905);
and UO_1253 (O_1253,N_9927,N_9879);
or UO_1254 (O_1254,N_9900,N_9899);
nand UO_1255 (O_1255,N_9857,N_9865);
nand UO_1256 (O_1256,N_9835,N_9837);
nor UO_1257 (O_1257,N_9916,N_9811);
or UO_1258 (O_1258,N_9882,N_9842);
nor UO_1259 (O_1259,N_9891,N_9846);
nand UO_1260 (O_1260,N_9890,N_9983);
nor UO_1261 (O_1261,N_9995,N_9988);
xor UO_1262 (O_1262,N_9909,N_9998);
or UO_1263 (O_1263,N_9809,N_9819);
xnor UO_1264 (O_1264,N_9854,N_9837);
xnor UO_1265 (O_1265,N_9969,N_9852);
xnor UO_1266 (O_1266,N_9807,N_9942);
and UO_1267 (O_1267,N_9826,N_9926);
nand UO_1268 (O_1268,N_9983,N_9893);
xor UO_1269 (O_1269,N_9834,N_9853);
or UO_1270 (O_1270,N_9943,N_9965);
nand UO_1271 (O_1271,N_9857,N_9852);
nand UO_1272 (O_1272,N_9934,N_9959);
xnor UO_1273 (O_1273,N_9809,N_9963);
and UO_1274 (O_1274,N_9842,N_9927);
and UO_1275 (O_1275,N_9859,N_9912);
nand UO_1276 (O_1276,N_9909,N_9855);
or UO_1277 (O_1277,N_9874,N_9916);
nand UO_1278 (O_1278,N_9846,N_9973);
nor UO_1279 (O_1279,N_9969,N_9967);
or UO_1280 (O_1280,N_9957,N_9876);
and UO_1281 (O_1281,N_9992,N_9954);
nor UO_1282 (O_1282,N_9842,N_9915);
nand UO_1283 (O_1283,N_9851,N_9991);
or UO_1284 (O_1284,N_9850,N_9944);
and UO_1285 (O_1285,N_9937,N_9830);
xor UO_1286 (O_1286,N_9999,N_9806);
xor UO_1287 (O_1287,N_9995,N_9831);
xnor UO_1288 (O_1288,N_9966,N_9926);
or UO_1289 (O_1289,N_9854,N_9921);
nor UO_1290 (O_1290,N_9865,N_9918);
nand UO_1291 (O_1291,N_9956,N_9955);
or UO_1292 (O_1292,N_9807,N_9892);
nand UO_1293 (O_1293,N_9916,N_9992);
or UO_1294 (O_1294,N_9936,N_9931);
nand UO_1295 (O_1295,N_9897,N_9823);
nor UO_1296 (O_1296,N_9981,N_9861);
and UO_1297 (O_1297,N_9921,N_9993);
xnor UO_1298 (O_1298,N_9804,N_9843);
nor UO_1299 (O_1299,N_9830,N_9845);
nor UO_1300 (O_1300,N_9976,N_9888);
and UO_1301 (O_1301,N_9920,N_9881);
nor UO_1302 (O_1302,N_9928,N_9832);
and UO_1303 (O_1303,N_9951,N_9890);
and UO_1304 (O_1304,N_9894,N_9914);
or UO_1305 (O_1305,N_9848,N_9847);
xnor UO_1306 (O_1306,N_9879,N_9902);
nand UO_1307 (O_1307,N_9935,N_9804);
nand UO_1308 (O_1308,N_9817,N_9837);
nor UO_1309 (O_1309,N_9909,N_9828);
nor UO_1310 (O_1310,N_9854,N_9862);
or UO_1311 (O_1311,N_9960,N_9905);
nand UO_1312 (O_1312,N_9966,N_9894);
nand UO_1313 (O_1313,N_9831,N_9956);
nand UO_1314 (O_1314,N_9867,N_9830);
xor UO_1315 (O_1315,N_9931,N_9875);
nand UO_1316 (O_1316,N_9900,N_9966);
nor UO_1317 (O_1317,N_9999,N_9917);
nand UO_1318 (O_1318,N_9851,N_9884);
nor UO_1319 (O_1319,N_9994,N_9993);
and UO_1320 (O_1320,N_9925,N_9942);
xor UO_1321 (O_1321,N_9937,N_9976);
or UO_1322 (O_1322,N_9849,N_9969);
nand UO_1323 (O_1323,N_9844,N_9872);
xor UO_1324 (O_1324,N_9889,N_9938);
or UO_1325 (O_1325,N_9846,N_9858);
nor UO_1326 (O_1326,N_9890,N_9816);
xnor UO_1327 (O_1327,N_9928,N_9807);
xor UO_1328 (O_1328,N_9808,N_9819);
nor UO_1329 (O_1329,N_9899,N_9923);
and UO_1330 (O_1330,N_9821,N_9959);
nand UO_1331 (O_1331,N_9842,N_9896);
nand UO_1332 (O_1332,N_9857,N_9985);
and UO_1333 (O_1333,N_9864,N_9821);
nor UO_1334 (O_1334,N_9955,N_9826);
xnor UO_1335 (O_1335,N_9826,N_9899);
nand UO_1336 (O_1336,N_9812,N_9951);
nand UO_1337 (O_1337,N_9939,N_9841);
nor UO_1338 (O_1338,N_9837,N_9802);
and UO_1339 (O_1339,N_9848,N_9801);
xnor UO_1340 (O_1340,N_9985,N_9922);
nor UO_1341 (O_1341,N_9976,N_9970);
xnor UO_1342 (O_1342,N_9919,N_9939);
nand UO_1343 (O_1343,N_9837,N_9959);
xor UO_1344 (O_1344,N_9883,N_9887);
and UO_1345 (O_1345,N_9827,N_9870);
nor UO_1346 (O_1346,N_9902,N_9942);
and UO_1347 (O_1347,N_9901,N_9945);
or UO_1348 (O_1348,N_9818,N_9883);
nand UO_1349 (O_1349,N_9859,N_9809);
nor UO_1350 (O_1350,N_9924,N_9889);
and UO_1351 (O_1351,N_9935,N_9951);
and UO_1352 (O_1352,N_9921,N_9855);
or UO_1353 (O_1353,N_9822,N_9969);
nand UO_1354 (O_1354,N_9817,N_9962);
nand UO_1355 (O_1355,N_9955,N_9952);
or UO_1356 (O_1356,N_9965,N_9917);
xnor UO_1357 (O_1357,N_9800,N_9946);
nor UO_1358 (O_1358,N_9824,N_9902);
xor UO_1359 (O_1359,N_9917,N_9979);
nor UO_1360 (O_1360,N_9957,N_9907);
and UO_1361 (O_1361,N_9839,N_9928);
xnor UO_1362 (O_1362,N_9949,N_9807);
and UO_1363 (O_1363,N_9802,N_9862);
and UO_1364 (O_1364,N_9930,N_9835);
nand UO_1365 (O_1365,N_9988,N_9962);
nor UO_1366 (O_1366,N_9994,N_9869);
or UO_1367 (O_1367,N_9871,N_9899);
or UO_1368 (O_1368,N_9875,N_9886);
or UO_1369 (O_1369,N_9958,N_9857);
or UO_1370 (O_1370,N_9807,N_9933);
nor UO_1371 (O_1371,N_9907,N_9928);
xor UO_1372 (O_1372,N_9975,N_9946);
and UO_1373 (O_1373,N_9854,N_9878);
and UO_1374 (O_1374,N_9992,N_9988);
xor UO_1375 (O_1375,N_9976,N_9886);
nand UO_1376 (O_1376,N_9892,N_9879);
and UO_1377 (O_1377,N_9901,N_9874);
nand UO_1378 (O_1378,N_9928,N_9874);
nand UO_1379 (O_1379,N_9954,N_9884);
nand UO_1380 (O_1380,N_9935,N_9863);
nand UO_1381 (O_1381,N_9856,N_9885);
nand UO_1382 (O_1382,N_9837,N_9935);
nor UO_1383 (O_1383,N_9856,N_9954);
nor UO_1384 (O_1384,N_9897,N_9840);
nor UO_1385 (O_1385,N_9953,N_9803);
nand UO_1386 (O_1386,N_9947,N_9988);
or UO_1387 (O_1387,N_9920,N_9900);
and UO_1388 (O_1388,N_9818,N_9843);
nor UO_1389 (O_1389,N_9810,N_9856);
nor UO_1390 (O_1390,N_9846,N_9880);
and UO_1391 (O_1391,N_9809,N_9990);
xnor UO_1392 (O_1392,N_9969,N_9982);
or UO_1393 (O_1393,N_9894,N_9878);
or UO_1394 (O_1394,N_9948,N_9911);
xor UO_1395 (O_1395,N_9860,N_9964);
and UO_1396 (O_1396,N_9945,N_9958);
xnor UO_1397 (O_1397,N_9906,N_9969);
xnor UO_1398 (O_1398,N_9955,N_9914);
xnor UO_1399 (O_1399,N_9917,N_9804);
xor UO_1400 (O_1400,N_9953,N_9858);
xnor UO_1401 (O_1401,N_9882,N_9808);
or UO_1402 (O_1402,N_9855,N_9900);
and UO_1403 (O_1403,N_9987,N_9962);
nor UO_1404 (O_1404,N_9986,N_9878);
or UO_1405 (O_1405,N_9959,N_9878);
nor UO_1406 (O_1406,N_9917,N_9945);
nand UO_1407 (O_1407,N_9852,N_9987);
xnor UO_1408 (O_1408,N_9818,N_9935);
xor UO_1409 (O_1409,N_9980,N_9901);
xor UO_1410 (O_1410,N_9865,N_9806);
and UO_1411 (O_1411,N_9858,N_9823);
xor UO_1412 (O_1412,N_9907,N_9813);
xor UO_1413 (O_1413,N_9966,N_9828);
xnor UO_1414 (O_1414,N_9901,N_9815);
or UO_1415 (O_1415,N_9966,N_9831);
xnor UO_1416 (O_1416,N_9917,N_9967);
nor UO_1417 (O_1417,N_9961,N_9903);
nand UO_1418 (O_1418,N_9805,N_9816);
nor UO_1419 (O_1419,N_9836,N_9800);
nor UO_1420 (O_1420,N_9977,N_9994);
or UO_1421 (O_1421,N_9993,N_9938);
or UO_1422 (O_1422,N_9800,N_9938);
or UO_1423 (O_1423,N_9881,N_9806);
and UO_1424 (O_1424,N_9923,N_9849);
xnor UO_1425 (O_1425,N_9811,N_9839);
nand UO_1426 (O_1426,N_9923,N_9887);
and UO_1427 (O_1427,N_9965,N_9814);
nand UO_1428 (O_1428,N_9910,N_9919);
and UO_1429 (O_1429,N_9836,N_9936);
nand UO_1430 (O_1430,N_9948,N_9883);
xor UO_1431 (O_1431,N_9883,N_9834);
nand UO_1432 (O_1432,N_9926,N_9917);
and UO_1433 (O_1433,N_9996,N_9889);
nand UO_1434 (O_1434,N_9808,N_9847);
nand UO_1435 (O_1435,N_9854,N_9966);
nand UO_1436 (O_1436,N_9984,N_9967);
and UO_1437 (O_1437,N_9892,N_9840);
xnor UO_1438 (O_1438,N_9849,N_9812);
nor UO_1439 (O_1439,N_9818,N_9960);
or UO_1440 (O_1440,N_9971,N_9992);
xor UO_1441 (O_1441,N_9999,N_9843);
nor UO_1442 (O_1442,N_9839,N_9959);
nor UO_1443 (O_1443,N_9937,N_9959);
or UO_1444 (O_1444,N_9854,N_9915);
and UO_1445 (O_1445,N_9909,N_9959);
xor UO_1446 (O_1446,N_9963,N_9948);
xor UO_1447 (O_1447,N_9835,N_9986);
and UO_1448 (O_1448,N_9844,N_9976);
and UO_1449 (O_1449,N_9941,N_9950);
xor UO_1450 (O_1450,N_9812,N_9827);
nand UO_1451 (O_1451,N_9897,N_9971);
and UO_1452 (O_1452,N_9907,N_9839);
nand UO_1453 (O_1453,N_9809,N_9800);
nand UO_1454 (O_1454,N_9838,N_9830);
nand UO_1455 (O_1455,N_9949,N_9878);
nand UO_1456 (O_1456,N_9923,N_9903);
nor UO_1457 (O_1457,N_9919,N_9990);
nand UO_1458 (O_1458,N_9972,N_9962);
nor UO_1459 (O_1459,N_9964,N_9924);
and UO_1460 (O_1460,N_9956,N_9884);
nor UO_1461 (O_1461,N_9893,N_9920);
nor UO_1462 (O_1462,N_9825,N_9846);
and UO_1463 (O_1463,N_9864,N_9830);
and UO_1464 (O_1464,N_9967,N_9807);
nand UO_1465 (O_1465,N_9848,N_9926);
and UO_1466 (O_1466,N_9970,N_9931);
or UO_1467 (O_1467,N_9936,N_9834);
or UO_1468 (O_1468,N_9853,N_9886);
xnor UO_1469 (O_1469,N_9929,N_9842);
nand UO_1470 (O_1470,N_9849,N_9824);
xnor UO_1471 (O_1471,N_9904,N_9984);
or UO_1472 (O_1472,N_9849,N_9979);
nor UO_1473 (O_1473,N_9969,N_9905);
xnor UO_1474 (O_1474,N_9924,N_9988);
nand UO_1475 (O_1475,N_9856,N_9942);
nand UO_1476 (O_1476,N_9891,N_9847);
or UO_1477 (O_1477,N_9911,N_9964);
xnor UO_1478 (O_1478,N_9920,N_9912);
or UO_1479 (O_1479,N_9883,N_9814);
and UO_1480 (O_1480,N_9849,N_9985);
and UO_1481 (O_1481,N_9846,N_9861);
and UO_1482 (O_1482,N_9876,N_9864);
xnor UO_1483 (O_1483,N_9984,N_9847);
nand UO_1484 (O_1484,N_9996,N_9927);
xor UO_1485 (O_1485,N_9996,N_9897);
nor UO_1486 (O_1486,N_9860,N_9981);
or UO_1487 (O_1487,N_9940,N_9905);
xor UO_1488 (O_1488,N_9974,N_9825);
and UO_1489 (O_1489,N_9887,N_9802);
xor UO_1490 (O_1490,N_9834,N_9889);
xor UO_1491 (O_1491,N_9912,N_9979);
or UO_1492 (O_1492,N_9986,N_9904);
xor UO_1493 (O_1493,N_9862,N_9812);
or UO_1494 (O_1494,N_9876,N_9989);
nand UO_1495 (O_1495,N_9998,N_9975);
nand UO_1496 (O_1496,N_9800,N_9802);
xor UO_1497 (O_1497,N_9964,N_9931);
and UO_1498 (O_1498,N_9852,N_9807);
and UO_1499 (O_1499,N_9917,N_9865);
endmodule