module basic_3000_30000_3500_150_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_668,In_29);
or U1 (N_1,In_1948,In_2843);
nor U2 (N_2,In_2393,In_2112);
nor U3 (N_3,In_1769,In_2854);
and U4 (N_4,In_614,In_147);
and U5 (N_5,In_2792,In_571);
and U6 (N_6,In_1765,In_2050);
nor U7 (N_7,In_2981,In_1436);
and U8 (N_8,In_306,In_1697);
xor U9 (N_9,In_532,In_204);
nor U10 (N_10,In_2790,In_1987);
nand U11 (N_11,In_716,In_2830);
and U12 (N_12,In_2667,In_2708);
nand U13 (N_13,In_1045,In_806);
or U14 (N_14,In_1604,In_2334);
nand U15 (N_15,In_1465,In_2009);
nand U16 (N_16,In_2450,In_1949);
nor U17 (N_17,In_2378,In_63);
xor U18 (N_18,In_2104,In_2952);
xor U19 (N_19,In_2846,In_1125);
nor U20 (N_20,In_616,In_206);
xor U21 (N_21,In_2065,In_1348);
nor U22 (N_22,In_1080,In_1652);
and U23 (N_23,In_2093,In_1800);
nand U24 (N_24,In_1651,In_917);
nand U25 (N_25,In_2411,In_2254);
nand U26 (N_26,In_1562,In_2037);
and U27 (N_27,In_1556,In_2182);
and U28 (N_28,In_213,In_901);
or U29 (N_29,In_2731,In_1739);
nand U30 (N_30,In_454,In_2734);
nor U31 (N_31,In_581,In_2933);
and U32 (N_32,In_2818,In_978);
nand U33 (N_33,In_290,In_2754);
and U34 (N_34,In_441,In_9);
nand U35 (N_35,In_1374,In_2817);
or U36 (N_36,In_1736,In_575);
xnor U37 (N_37,In_958,In_804);
and U38 (N_38,In_1257,In_28);
nand U39 (N_39,In_1893,In_57);
nand U40 (N_40,In_475,In_2303);
and U41 (N_41,In_1001,In_1424);
and U42 (N_42,In_799,In_2383);
xnor U43 (N_43,In_300,In_890);
nor U44 (N_44,In_88,In_1646);
xnor U45 (N_45,In_2006,In_1795);
nor U46 (N_46,In_1416,In_2622);
and U47 (N_47,In_503,In_524);
xnor U48 (N_48,In_31,In_982);
nand U49 (N_49,In_623,In_1818);
or U50 (N_50,In_2728,In_24);
nand U51 (N_51,In_2194,In_1835);
xnor U52 (N_52,In_379,In_2351);
and U53 (N_53,In_2090,In_1268);
and U54 (N_54,In_1808,In_1202);
and U55 (N_55,In_989,In_61);
nand U56 (N_56,In_2841,In_2837);
nand U57 (N_57,In_788,In_2935);
or U58 (N_58,In_1370,In_2523);
xnor U59 (N_59,In_1851,In_2575);
and U60 (N_60,In_2513,In_2724);
nor U61 (N_61,In_710,In_2957);
nand U62 (N_62,In_1919,In_1211);
and U63 (N_63,In_2900,In_2689);
and U64 (N_64,In_460,In_162);
nor U65 (N_65,In_1883,In_2291);
nand U66 (N_66,In_2819,In_651);
or U67 (N_67,In_1005,In_1720);
or U68 (N_68,In_2238,In_2323);
nor U69 (N_69,In_1042,In_1732);
nor U70 (N_70,In_181,In_1786);
xnor U71 (N_71,In_2289,In_1250);
nor U72 (N_72,In_2459,In_2167);
nor U73 (N_73,In_1843,In_2056);
or U74 (N_74,In_2906,In_408);
nand U75 (N_75,In_2729,In_462);
nor U76 (N_76,In_2505,In_231);
or U77 (N_77,In_1264,In_612);
and U78 (N_78,In_698,In_156);
and U79 (N_79,In_1583,In_2700);
or U80 (N_80,In_1429,In_1316);
nor U81 (N_81,In_399,In_553);
and U82 (N_82,In_1058,In_1420);
xor U83 (N_83,In_339,In_2597);
and U84 (N_84,In_450,In_513);
nor U85 (N_85,In_2499,In_2814);
and U86 (N_86,In_1597,In_1622);
and U87 (N_87,In_655,In_1997);
or U88 (N_88,In_1350,In_959);
or U89 (N_89,In_520,In_2704);
and U90 (N_90,In_1209,In_1738);
and U91 (N_91,In_1877,In_447);
nand U92 (N_92,In_964,In_2949);
xnor U93 (N_93,In_1285,In_1031);
xnor U94 (N_94,In_146,In_690);
and U95 (N_95,In_1309,In_2117);
xor U96 (N_96,In_301,In_1618);
and U97 (N_97,In_2885,In_552);
xor U98 (N_98,In_2067,In_2177);
nor U99 (N_99,In_2894,In_485);
and U100 (N_100,In_1200,In_107);
nor U101 (N_101,In_1,In_903);
and U102 (N_102,In_1771,In_2613);
or U103 (N_103,In_120,In_2501);
or U104 (N_104,In_2361,In_1298);
nand U105 (N_105,In_201,In_20);
or U106 (N_106,In_1779,In_2966);
xnor U107 (N_107,In_1283,In_1197);
or U108 (N_108,In_2567,In_1419);
or U109 (N_109,In_508,In_2757);
nor U110 (N_110,In_1728,In_68);
or U111 (N_111,In_1759,In_1294);
nand U112 (N_112,In_1628,In_947);
and U113 (N_113,In_1986,In_1733);
nand U114 (N_114,In_2223,In_1519);
nor U115 (N_115,In_1539,In_675);
or U116 (N_116,In_2799,In_894);
nand U117 (N_117,In_2748,In_1974);
nor U118 (N_118,In_1820,In_1051);
nand U119 (N_119,In_1079,In_2207);
nand U120 (N_120,In_2247,In_1601);
xnor U121 (N_121,In_1484,In_1116);
nand U122 (N_122,In_993,In_2861);
xor U123 (N_123,In_1678,In_233);
nor U124 (N_124,In_256,In_2094);
and U125 (N_125,In_2539,In_1144);
nand U126 (N_126,In_1511,In_1661);
nor U127 (N_127,In_502,In_2467);
nand U128 (N_128,In_1970,In_1853);
nor U129 (N_129,In_2532,In_2119);
nor U130 (N_130,In_913,In_669);
xnor U131 (N_131,In_734,In_1222);
nor U132 (N_132,In_2280,In_1060);
or U133 (N_133,In_679,In_963);
nor U134 (N_134,In_2690,In_1399);
nand U135 (N_135,In_230,In_657);
xor U136 (N_136,In_1857,In_1522);
or U137 (N_137,In_1330,In_1109);
or U138 (N_138,In_999,In_2913);
and U139 (N_139,In_2257,In_595);
nor U140 (N_140,In_44,In_782);
nor U141 (N_141,In_1289,In_830);
xnor U142 (N_142,In_1333,In_192);
and U143 (N_143,In_1703,In_2078);
and U144 (N_144,In_1136,In_331);
nor U145 (N_145,In_1660,In_5);
and U146 (N_146,In_2229,In_1068);
or U147 (N_147,In_582,In_2694);
xor U148 (N_148,In_1582,In_1700);
nor U149 (N_149,In_1115,In_190);
nand U150 (N_150,In_2663,In_2477);
nand U151 (N_151,In_795,In_237);
nor U152 (N_152,In_1143,In_238);
xnor U153 (N_153,In_2587,In_1392);
or U154 (N_154,In_2835,In_550);
and U155 (N_155,In_2773,In_354);
nor U156 (N_156,In_704,In_891);
nand U157 (N_157,In_590,In_2472);
nand U158 (N_158,In_2014,In_1010);
nor U159 (N_159,In_243,In_2606);
nand U160 (N_160,In_1306,In_1237);
and U161 (N_161,In_605,In_717);
nand U162 (N_162,In_1224,In_509);
and U163 (N_163,In_2990,In_194);
xnor U164 (N_164,In_2412,In_857);
or U165 (N_165,In_246,In_459);
xnor U166 (N_166,In_1692,In_1899);
or U167 (N_167,In_618,In_2771);
and U168 (N_168,In_850,In_2822);
xnor U169 (N_169,In_228,In_1464);
and U170 (N_170,In_1938,In_574);
nor U171 (N_171,In_292,In_2240);
or U172 (N_172,In_1805,In_496);
nor U173 (N_173,In_1588,In_1811);
nor U174 (N_174,In_1648,In_570);
and U175 (N_175,In_1677,In_702);
nor U176 (N_176,In_2725,In_2747);
or U177 (N_177,In_832,In_411);
nand U178 (N_178,In_2166,In_1391);
nand U179 (N_179,In_227,In_1276);
or U180 (N_180,In_735,In_1870);
or U181 (N_181,In_984,In_2699);
xor U182 (N_182,In_1225,In_2552);
or U183 (N_183,In_2801,In_483);
xnor U184 (N_184,In_887,In_1434);
nor U185 (N_185,In_2088,In_2428);
nor U186 (N_186,In_2216,In_1152);
and U187 (N_187,In_2661,In_67);
or U188 (N_188,In_664,In_1242);
or U189 (N_189,In_1991,In_2127);
xnor U190 (N_190,In_974,In_1561);
or U191 (N_191,In_1980,In_724);
nor U192 (N_192,In_2027,In_787);
xnor U193 (N_193,In_2013,In_262);
nand U194 (N_194,In_1838,In_2162);
xor U195 (N_195,In_436,In_746);
nor U196 (N_196,In_1679,In_2096);
or U197 (N_197,In_1112,In_2187);
xnor U198 (N_198,In_2512,In_1213);
nand U199 (N_199,In_490,In_130);
and U200 (N_200,In_1964,In_404);
nand U201 (N_201,In_1214,In_1662);
nor U202 (N_202,In_537,In_1063);
or U203 (N_203,In_1028,In_1123);
xnor U204 (N_204,In_2039,In_1270);
nor U205 (N_205,In_1117,In_2034);
nand U206 (N_206,In_1907,In_387);
nor U207 (N_207,In_104,In_2521);
and U208 (N_208,In_1352,In_1183);
or U209 (N_209,In_356,In_722);
nor U210 (N_210,In_1252,In_1550);
and U211 (N_211,In_1840,In_2655);
and U212 (N_212,In_1188,In_11);
nand U213 (N_213,In_713,In_2273);
and U214 (N_214,In_2641,N_170);
nand U215 (N_215,In_775,In_62);
and U216 (N_216,N_93,In_41);
xor U217 (N_217,In_990,In_1989);
nor U218 (N_218,In_1866,In_2940);
xnor U219 (N_219,In_1691,In_1207);
nor U220 (N_220,In_2149,In_910);
or U221 (N_221,In_2770,In_2615);
nand U222 (N_222,In_2926,In_1928);
nand U223 (N_223,In_2305,In_2953);
nor U224 (N_224,N_153,In_1274);
or U225 (N_225,In_398,N_28);
xnor U226 (N_226,In_2018,In_895);
xnor U227 (N_227,In_1580,N_126);
xor U228 (N_228,In_2693,In_885);
or U229 (N_229,In_2294,In_2038);
xor U230 (N_230,In_2409,In_1711);
and U231 (N_231,In_2805,In_2654);
nor U232 (N_232,In_1600,In_922);
or U233 (N_233,In_1410,In_572);
and U234 (N_234,In_60,N_112);
or U235 (N_235,In_1199,In_672);
and U236 (N_236,In_2856,In_270);
or U237 (N_237,In_1421,In_1920);
or U238 (N_238,In_1255,In_2463);
and U239 (N_239,In_1329,N_30);
nand U240 (N_240,In_565,In_91);
nor U241 (N_241,In_1755,In_53);
nand U242 (N_242,In_38,In_1346);
or U243 (N_243,In_400,N_151);
xor U244 (N_244,In_1025,In_128);
nand U245 (N_245,In_1272,In_1781);
xnor U246 (N_246,In_2016,In_1249);
and U247 (N_247,In_841,In_1828);
or U248 (N_248,In_2277,In_1915);
nand U249 (N_249,In_211,In_226);
or U250 (N_250,In_1332,In_2121);
nor U251 (N_251,In_2621,In_2300);
or U252 (N_252,In_1514,In_2171);
and U253 (N_253,In_169,In_2902);
nor U254 (N_254,In_1925,In_1072);
or U255 (N_255,In_2259,In_209);
nor U256 (N_256,In_2605,In_1463);
nor U257 (N_257,In_1577,In_149);
or U258 (N_258,In_884,In_2255);
xor U259 (N_259,In_1960,In_1182);
nor U260 (N_260,In_2466,In_564);
or U261 (N_261,In_1740,In_653);
xnor U262 (N_262,N_13,In_2028);
nand U263 (N_263,In_2371,In_176);
or U264 (N_264,N_46,In_2425);
and U265 (N_265,In_2394,N_50);
nor U266 (N_266,In_1389,In_52);
or U267 (N_267,In_487,N_92);
and U268 (N_268,In_2377,In_2691);
xnor U269 (N_269,In_518,In_1638);
nor U270 (N_270,In_1520,In_2331);
xnor U271 (N_271,In_2282,N_71);
xor U272 (N_272,In_185,In_131);
or U273 (N_273,In_479,In_245);
xnor U274 (N_274,In_630,In_1384);
xor U275 (N_275,In_2418,In_1398);
and U276 (N_276,In_51,In_2446);
and U277 (N_277,In_1775,In_2538);
nor U278 (N_278,In_2563,In_1734);
nand U279 (N_279,In_881,In_1337);
nor U280 (N_280,In_80,In_2872);
nand U281 (N_281,In_939,In_1494);
nor U282 (N_282,N_133,In_2565);
or U283 (N_283,In_2877,In_1532);
or U284 (N_284,In_353,In_1564);
nand U285 (N_285,N_0,In_2271);
or U286 (N_286,In_2553,In_2032);
xor U287 (N_287,In_1304,In_210);
nor U288 (N_288,In_2141,In_1515);
or U289 (N_289,In_456,In_119);
and U290 (N_290,In_2707,In_809);
nor U291 (N_291,In_2934,In_2676);
and U292 (N_292,In_494,In_2228);
or U293 (N_293,In_1833,In_2310);
nand U294 (N_294,In_2140,In_2897);
nor U295 (N_295,In_2297,In_617);
nor U296 (N_296,In_10,In_2498);
and U297 (N_297,In_602,In_2941);
xnor U298 (N_298,In_449,In_419);
xor U299 (N_299,In_541,In_1445);
xnor U300 (N_300,N_122,In_1961);
nand U301 (N_301,In_2326,In_2151);
and U302 (N_302,In_1657,In_2503);
xnor U303 (N_303,In_1815,In_1278);
nand U304 (N_304,In_2212,In_1914);
xor U305 (N_305,In_533,In_1018);
xor U306 (N_306,In_1999,In_1449);
or U307 (N_307,In_1359,In_1855);
nand U308 (N_308,In_1021,In_1507);
nand U309 (N_309,In_1760,In_1926);
and U310 (N_310,In_900,In_1869);
nor U311 (N_311,In_295,In_2234);
or U312 (N_312,In_313,In_2666);
or U313 (N_313,In_2284,In_1203);
nor U314 (N_314,In_2647,N_75);
nor U315 (N_315,N_29,In_2898);
xor U316 (N_316,In_2440,In_1166);
or U317 (N_317,In_2278,In_1984);
nor U318 (N_318,In_49,In_317);
xor U319 (N_319,In_1430,In_2033);
xor U320 (N_320,In_1243,In_1048);
or U321 (N_321,In_1852,N_69);
nand U322 (N_322,In_621,In_2239);
nor U323 (N_323,In_343,In_1531);
nand U324 (N_324,In_1095,In_279);
xnor U325 (N_325,In_1489,In_2601);
or U326 (N_326,In_2514,In_1461);
or U327 (N_327,In_2534,In_696);
nor U328 (N_328,In_1590,In_2739);
xnor U329 (N_329,In_567,In_836);
and U330 (N_330,N_11,In_1649);
or U331 (N_331,In_263,In_133);
nor U332 (N_332,In_154,In_1792);
or U333 (N_333,In_2733,In_2786);
xor U334 (N_334,In_888,In_851);
nor U335 (N_335,In_2252,In_2268);
nand U336 (N_336,In_1694,In_2407);
nand U337 (N_337,In_721,In_16);
nand U338 (N_338,In_1574,N_136);
or U339 (N_339,In_932,In_2313);
nor U340 (N_340,In_1376,In_1747);
nor U341 (N_341,In_1655,In_561);
or U342 (N_342,N_139,In_1575);
nor U343 (N_343,In_941,In_2107);
nor U344 (N_344,In_2764,In_180);
and U345 (N_345,In_2645,In_1922);
xnor U346 (N_346,In_2617,N_27);
nand U347 (N_347,N_156,In_482);
xor U348 (N_348,In_1358,In_1947);
xor U349 (N_349,In_1971,In_2634);
or U350 (N_350,In_828,In_2026);
xor U351 (N_351,In_1128,In_166);
xor U352 (N_352,In_2573,In_17);
nor U353 (N_353,In_535,In_2648);
and U354 (N_354,In_1658,In_1168);
xor U355 (N_355,In_2079,In_2946);
or U356 (N_356,In_1036,In_1096);
nand U357 (N_357,In_2508,In_684);
or U358 (N_358,In_432,In_1219);
nor U359 (N_359,In_2916,In_30);
xor U360 (N_360,In_2871,In_2128);
and U361 (N_361,In_2399,In_2763);
nand U362 (N_362,N_150,In_452);
nand U363 (N_363,In_644,In_1171);
or U364 (N_364,In_1415,In_1715);
xor U365 (N_365,In_2518,In_671);
or U366 (N_366,In_272,In_1296);
and U367 (N_367,In_1266,In_1282);
or U368 (N_368,In_2979,In_2329);
and U369 (N_369,In_1617,In_302);
nor U370 (N_370,In_1342,In_2288);
xnor U371 (N_371,In_2643,In_960);
nor U372 (N_372,In_2286,In_2507);
nand U373 (N_373,In_351,In_1287);
xnor U374 (N_374,In_816,In_1367);
nor U375 (N_375,In_1317,In_2680);
and U376 (N_376,In_168,In_2089);
nor U377 (N_377,In_96,In_937);
nor U378 (N_378,In_367,In_744);
nor U379 (N_379,In_2976,In_2920);
and U380 (N_380,In_1823,In_805);
and U381 (N_381,In_862,In_511);
xor U382 (N_382,In_1262,In_2626);
and U383 (N_383,In_36,In_783);
or U384 (N_384,In_2829,In_1718);
or U385 (N_385,In_624,In_992);
xor U386 (N_386,In_1414,In_852);
nor U387 (N_387,In_596,In_1228);
nand U388 (N_388,In_2137,In_2620);
or U389 (N_389,In_2542,In_556);
nand U390 (N_390,In_373,N_182);
and U391 (N_391,N_44,In_1238);
xnor U392 (N_392,In_1396,In_762);
or U393 (N_393,In_2306,In_2596);
nand U394 (N_394,N_61,In_2029);
and U395 (N_395,In_2465,In_1780);
and U396 (N_396,In_2003,In_2103);
nor U397 (N_397,In_85,In_874);
nor U398 (N_398,In_2812,In_370);
xnor U399 (N_399,In_609,In_2347);
nor U400 (N_400,In_1867,In_1902);
nor U401 (N_401,In_1995,N_98);
and U402 (N_402,In_648,In_1773);
or U403 (N_403,In_200,In_1768);
and U404 (N_404,In_2062,In_1295);
nor U405 (N_405,In_2738,N_254);
nand U406 (N_406,In_656,In_1169);
nor U407 (N_407,In_707,In_455);
xnor U408 (N_408,N_237,In_793);
nand U409 (N_409,In_2069,N_144);
or U410 (N_410,In_1088,In_222);
nand U411 (N_411,In_1246,In_2447);
nor U412 (N_412,In_1900,In_2489);
and U413 (N_413,In_1226,In_678);
xnor U414 (N_414,In_2341,In_2405);
nand U415 (N_415,In_1684,In_840);
and U416 (N_416,In_2281,In_1754);
xor U417 (N_417,In_525,In_948);
or U418 (N_418,In_445,In_2308);
and U419 (N_419,In_551,In_99);
or U420 (N_420,In_1560,N_217);
and U421 (N_421,In_534,In_402);
nand U422 (N_422,In_434,In_174);
nor U423 (N_423,In_985,In_1124);
nor U424 (N_424,In_2684,In_1150);
xor U425 (N_425,In_1336,In_2340);
and U426 (N_426,N_8,In_1674);
or U427 (N_427,In_1952,In_2912);
or U428 (N_428,In_1794,In_2717);
nand U429 (N_429,N_286,In_2010);
and U430 (N_430,In_529,In_504);
xnor U431 (N_431,In_1699,In_2806);
nand U432 (N_432,In_643,N_2);
xor U433 (N_433,In_2571,In_468);
xnor U434 (N_434,N_90,N_317);
or U435 (N_435,In_1253,In_1707);
xnor U436 (N_436,In_1895,In_2719);
xor U437 (N_437,N_380,N_255);
nand U438 (N_438,In_2320,In_1813);
and U439 (N_439,In_1433,In_1871);
nand U440 (N_440,In_1606,N_148);
or U441 (N_441,N_327,In_1456);
nor U442 (N_442,In_594,In_1052);
or U443 (N_443,In_972,In_2035);
xor U444 (N_444,In_1944,In_2087);
nand U445 (N_445,In_420,In_2984);
nor U446 (N_446,In_1032,In_654);
nand U447 (N_447,N_180,In_2893);
nand U448 (N_448,In_1040,In_1026);
xnor U449 (N_449,In_1400,In_2091);
nand U450 (N_450,In_559,In_366);
nor U451 (N_451,In_2434,In_308);
nor U452 (N_452,In_1099,N_287);
and U453 (N_453,In_70,N_253);
xnor U454 (N_454,In_2311,In_1898);
nor U455 (N_455,In_2395,In_2114);
and U456 (N_456,In_1156,N_77);
and U457 (N_457,In_2664,In_1625);
and U458 (N_458,In_1544,N_174);
xor U459 (N_459,In_73,In_255);
and U460 (N_460,In_1536,In_1686);
or U461 (N_461,In_480,In_991);
xnor U462 (N_462,In_2068,In_2210);
nor U463 (N_463,In_1066,In_2298);
and U464 (N_464,In_182,In_383);
xor U465 (N_465,In_825,In_208);
and U466 (N_466,In_2604,In_1323);
nor U467 (N_467,In_920,N_155);
or U468 (N_468,In_592,In_2939);
xor U469 (N_469,In_2675,In_1453);
and U470 (N_470,N_393,In_1365);
and U471 (N_471,In_2526,In_2566);
and U472 (N_472,In_797,In_942);
xnor U473 (N_473,N_239,In_25);
or U474 (N_474,N_184,In_1011);
and U475 (N_475,In_1955,In_416);
and U476 (N_476,In_2670,In_1455);
or U477 (N_477,In_1233,In_986);
or U478 (N_478,In_1340,In_1347);
xor U479 (N_479,In_1092,In_2510);
xnor U480 (N_480,In_134,In_1413);
nand U481 (N_481,In_148,In_2490);
and U482 (N_482,In_1770,In_2958);
nor U483 (N_483,In_386,In_1189);
nor U484 (N_484,N_107,In_2787);
and U485 (N_485,In_814,In_898);
xor U486 (N_486,In_1321,In_2954);
and U487 (N_487,In_310,N_378);
or U488 (N_488,In_172,In_2679);
nor U489 (N_489,In_1292,In_1693);
nand U490 (N_490,In_1741,N_49);
and U491 (N_491,N_12,In_2205);
or U492 (N_492,In_2386,In_115);
or U493 (N_493,In_2293,In_1310);
and U494 (N_494,In_909,In_2568);
and U495 (N_495,In_378,In_2304);
xnor U496 (N_496,In_1435,In_1155);
xor U497 (N_497,In_2783,In_1743);
nor U498 (N_498,In_1471,In_975);
nand U499 (N_499,In_1175,N_312);
or U500 (N_500,In_2889,N_307);
nor U501 (N_501,In_414,In_1132);
nand U502 (N_502,In_2154,N_59);
nand U503 (N_503,In_1483,In_2494);
xnor U504 (N_504,In_2315,In_691);
nor U505 (N_505,In_2839,In_2349);
xor U506 (N_506,In_2686,In_855);
and U507 (N_507,In_1406,In_2460);
nand U508 (N_508,In_2390,N_200);
and U509 (N_509,In_2767,In_297);
nor U510 (N_510,In_2765,In_2778);
nand U511 (N_511,In_2095,In_2430);
or U512 (N_512,N_57,In_2064);
and U513 (N_513,In_254,In_1408);
or U514 (N_514,In_1006,N_280);
nor U515 (N_515,In_1581,In_393);
nor U516 (N_516,In_680,In_2662);
nor U517 (N_517,In_2385,In_784);
and U518 (N_518,In_1524,In_2366);
xnor U519 (N_519,In_725,In_318);
nor U520 (N_520,In_1596,In_2398);
or U521 (N_521,In_2796,In_267);
xor U522 (N_522,In_936,In_2183);
or U523 (N_523,N_278,N_210);
or U524 (N_524,N_302,In_792);
nand U525 (N_525,In_701,N_109);
nand U526 (N_526,In_446,In_2479);
xnor U527 (N_527,In_1927,In_730);
or U528 (N_528,In_2942,In_1427);
and U529 (N_529,In_394,In_1320);
nand U530 (N_530,In_1631,In_1886);
xnor U531 (N_531,In_2345,N_295);
or U532 (N_532,In_2849,In_2302);
or U533 (N_533,In_1559,In_1992);
and U534 (N_534,In_1064,In_2001);
nand U535 (N_535,In_2600,In_1127);
and U536 (N_536,In_1345,In_333);
nor U537 (N_537,In_1746,In_1565);
xor U538 (N_538,In_2682,In_2988);
nand U539 (N_539,In_74,In_2665);
and U540 (N_540,In_2080,In_727);
nor U541 (N_541,In_32,In_1847);
nand U542 (N_542,N_83,In_1549);
and U543 (N_543,In_2043,In_1185);
nor U544 (N_544,In_217,In_113);
and U545 (N_545,In_818,In_2461);
nand U546 (N_546,In_2072,In_2695);
xnor U547 (N_547,In_1994,In_2578);
and U548 (N_548,In_1953,In_699);
xor U549 (N_549,In_639,In_1527);
nand U550 (N_550,In_1313,In_908);
or U551 (N_551,In_1275,In_2749);
or U552 (N_552,In_2236,In_2882);
nor U553 (N_553,In_138,In_1569);
nand U554 (N_554,In_558,In_1821);
nand U555 (N_555,In_674,In_1834);
nand U556 (N_556,In_821,In_1557);
or U557 (N_557,In_2716,N_272);
and U558 (N_558,In_1355,N_3);
and U559 (N_559,In_2881,In_521);
nor U560 (N_560,In_970,N_87);
nand U561 (N_561,In_1432,In_1327);
xnor U562 (N_562,In_2217,In_2929);
nand U563 (N_563,In_2823,In_1261);
and U564 (N_564,In_2246,N_171);
or U565 (N_565,In_1506,In_2838);
nand U566 (N_566,In_1158,In_444);
and U567 (N_567,In_776,In_2594);
nand U568 (N_568,N_232,In_996);
xor U569 (N_569,In_1439,N_348);
nand U570 (N_570,N_241,In_859);
nand U571 (N_571,In_1566,In_2517);
nor U572 (N_572,In_2116,In_2290);
xnor U573 (N_573,In_2515,In_2330);
nand U574 (N_574,N_89,In_2970);
nor U575 (N_575,In_778,In_2215);
and U576 (N_576,In_2415,In_2285);
and U577 (N_577,In_412,In_1497);
xnor U578 (N_578,N_363,In_1258);
or U579 (N_579,N_370,In_348);
xor U580 (N_580,In_1814,In_2737);
xnor U581 (N_581,In_124,In_870);
or U582 (N_582,In_1475,In_2369);
or U583 (N_583,In_811,In_823);
nor U584 (N_584,In_2609,In_1377);
nand U585 (N_585,In_2746,In_2588);
xnor U586 (N_586,In_1145,In_1135);
xor U587 (N_587,In_1178,In_1360);
nor U588 (N_588,N_313,In_2408);
nor U589 (N_589,In_2487,In_488);
nor U590 (N_590,In_2433,In_1512);
or U591 (N_591,In_2049,In_377);
and U592 (N_592,In_2030,In_2230);
and U593 (N_593,In_319,In_2357);
xnor U594 (N_594,In_2832,In_2502);
nand U595 (N_595,In_165,In_141);
or U596 (N_596,In_560,In_236);
nor U597 (N_597,N_336,N_331);
nor U598 (N_598,N_243,In_2959);
or U599 (N_599,In_2258,N_134);
or U600 (N_600,In_106,In_1375);
nor U601 (N_601,In_2795,In_47);
xor U602 (N_602,N_439,In_732);
or U603 (N_603,In_2203,N_301);
and U604 (N_604,In_1533,N_502);
xor U605 (N_605,N_518,In_1990);
and U606 (N_606,In_1120,N_205);
nand U607 (N_607,In_293,In_715);
and U608 (N_608,In_2189,In_2911);
nand U609 (N_609,N_143,In_2652);
xor U610 (N_610,In_137,N_402);
xor U611 (N_611,N_34,In_2370);
nor U612 (N_612,N_593,In_925);
and U613 (N_613,N_296,In_303);
and U614 (N_614,In_240,In_2057);
nor U615 (N_615,In_1845,In_1319);
xnor U616 (N_616,N_245,In_18);
xor U617 (N_617,In_1717,In_578);
xor U618 (N_618,In_631,In_1708);
and U619 (N_619,N_599,In_1081);
and U620 (N_620,In_337,In_1591);
or U621 (N_621,N_192,N_465);
nand U622 (N_622,In_2392,In_1850);
xnor U623 (N_623,In_79,In_2673);
xnor U624 (N_624,In_2156,In_2265);
nand U625 (N_625,N_523,In_2172);
xnor U626 (N_626,In_362,In_1299);
nand U627 (N_627,N_473,In_288);
or U628 (N_628,N_6,In_695);
xnor U629 (N_629,In_824,N_460);
or U630 (N_630,N_215,In_225);
and U631 (N_631,In_1858,In_1671);
xnor U632 (N_632,In_248,In_1634);
or U633 (N_633,In_1958,In_323);
nand U634 (N_634,In_352,In_2888);
nor U635 (N_635,In_845,In_335);
or U636 (N_636,In_988,In_2928);
xnor U637 (N_637,In_305,In_157);
nand U638 (N_638,In_1053,In_2628);
nor U639 (N_639,N_110,N_343);
xor U640 (N_640,In_632,N_309);
nor U641 (N_641,In_2875,In_1945);
nor U642 (N_642,In_132,In_904);
or U643 (N_643,In_1874,In_563);
and U644 (N_644,In_733,In_2163);
nor U645 (N_645,N_248,N_339);
and U646 (N_646,In_2709,In_112);
nand U647 (N_647,N_355,In_2382);
xnor U648 (N_648,In_758,N_267);
nand U649 (N_649,In_628,In_767);
xor U650 (N_650,In_2175,In_2544);
xor U651 (N_651,In_2040,In_2206);
or U652 (N_652,N_454,In_2339);
xnor U653 (N_653,In_507,In_2455);
xor U654 (N_654,In_2309,In_2316);
and U655 (N_655,In_2556,In_1498);
or U656 (N_656,In_2997,In_528);
nor U657 (N_657,In_2480,In_1827);
nor U658 (N_658,In_1776,In_661);
xnor U659 (N_659,In_2362,In_2726);
nor U660 (N_660,N_173,In_198);
or U661 (N_661,In_649,In_1545);
nand U662 (N_662,In_2968,In_693);
nor U663 (N_663,In_2243,N_522);
nor U664 (N_664,In_2161,In_790);
nand U665 (N_665,In_2148,In_943);
nor U666 (N_666,In_2139,In_285);
nand U667 (N_667,In_2702,In_345);
and U668 (N_668,N_26,In_1772);
nor U669 (N_669,In_2516,N_70);
xor U670 (N_670,In_2869,N_346);
nand U671 (N_671,In_2186,In_2404);
and U672 (N_672,In_2973,N_503);
and U673 (N_673,In_2047,In_2632);
nor U674 (N_674,In_650,In_2925);
xnor U675 (N_675,In_478,In_430);
xnor U676 (N_676,In_1187,In_1611);
nand U677 (N_677,In_2756,In_1896);
nand U678 (N_678,In_1876,In_2099);
nor U679 (N_679,N_16,N_224);
nand U680 (N_680,In_1468,In_1452);
or U681 (N_681,In_662,In_600);
or U682 (N_682,In_1428,In_1248);
nor U683 (N_683,In_601,In_58);
nand U684 (N_684,N_203,In_794);
nor U685 (N_685,In_0,In_2994);
xor U686 (N_686,In_1946,In_1656);
nor U687 (N_687,N_256,In_252);
or U688 (N_688,In_1173,N_160);
nor U689 (N_689,N_420,In_2011);
or U690 (N_690,In_774,In_916);
and U691 (N_691,In_2956,In_1405);
nor U692 (N_692,In_486,In_69);
or U693 (N_693,In_2760,In_1302);
and U694 (N_694,In_2160,In_2943);
or U695 (N_695,In_2732,In_2705);
nor U696 (N_696,N_557,N_84);
nand U697 (N_697,In_2519,N_17);
nor U698 (N_698,N_43,In_2586);
or U699 (N_699,N_452,In_7);
nand U700 (N_700,In_328,In_1174);
xnor U701 (N_701,In_2904,In_2389);
xor U702 (N_702,In_1731,In_3);
and U703 (N_703,In_2850,In_1280);
or U704 (N_704,In_812,N_190);
xor U705 (N_705,In_1643,In_1887);
nand U706 (N_706,In_2000,In_1929);
nor U707 (N_707,In_2809,In_294);
and U708 (N_708,In_924,In_1615);
xnor U709 (N_709,In_2722,In_2232);
nand U710 (N_710,In_175,In_2400);
nor U711 (N_711,N_449,N_276);
xor U712 (N_712,N_586,In_833);
or U713 (N_713,In_2938,In_2414);
nor U714 (N_714,In_755,N_515);
nand U715 (N_715,In_2081,In_1181);
nand U716 (N_716,In_76,In_1179);
nor U717 (N_717,In_1891,In_2813);
and U718 (N_718,In_2328,In_896);
or U719 (N_719,In_1666,In_2744);
nor U720 (N_720,In_1950,In_1702);
or U721 (N_721,In_2636,In_1418);
or U722 (N_722,In_1386,In_554);
xnor U723 (N_723,In_877,In_2574);
nand U724 (N_724,In_311,In_1735);
nor U725 (N_725,N_472,In_835);
or U726 (N_726,N_356,N_396);
xnor U727 (N_727,In_530,In_2132);
nand U728 (N_728,In_737,In_2312);
or U729 (N_729,In_1312,N_587);
nand U730 (N_730,In_1133,In_1488);
or U731 (N_731,In_1043,In_2333);
or U732 (N_732,In_583,In_218);
nor U733 (N_733,In_1077,In_1089);
nor U734 (N_734,N_326,In_497);
and U735 (N_735,In_1019,In_2602);
nand U736 (N_736,In_580,In_822);
nand U737 (N_737,In_706,N_589);
nor U738 (N_738,In_1114,In_1437);
or U739 (N_739,In_2170,In_1502);
nor U740 (N_740,In_325,N_425);
nand U741 (N_741,In_714,N_394);
nand U742 (N_742,In_2564,In_2384);
or U743 (N_743,In_2698,N_407);
nand U744 (N_744,In_2066,N_72);
or U745 (N_745,In_361,In_1623);
xor U746 (N_746,N_146,In_2901);
or U747 (N_747,N_416,N_323);
xor U748 (N_748,N_226,In_304);
nor U749 (N_749,N_277,In_858);
xor U750 (N_750,In_815,In_2740);
nor U751 (N_751,In_2335,In_711);
or U752 (N_752,In_1909,In_2219);
nor U753 (N_753,In_2401,In_2750);
nand U754 (N_754,In_2569,In_636);
nor U755 (N_755,In_2811,In_2017);
nor U756 (N_756,In_357,N_399);
or U757 (N_757,In_1407,N_175);
or U758 (N_758,In_2999,N_567);
or U759 (N_759,In_2120,In_2368);
nor U760 (N_760,In_2388,In_265);
and U761 (N_761,In_1492,In_606);
or U762 (N_762,In_1022,N_488);
and U763 (N_763,In_2410,N_5);
and U764 (N_764,In_42,N_311);
and U765 (N_765,N_397,In_873);
and U766 (N_766,In_2214,In_92);
nor U767 (N_767,N_162,In_199);
xor U768 (N_768,In_780,N_213);
nand U769 (N_769,In_2980,In_476);
and U770 (N_770,In_1723,In_2777);
or U771 (N_771,In_2299,In_2457);
and U772 (N_772,N_270,In_2005);
xnor U773 (N_773,In_1212,In_1695);
xor U774 (N_774,In_1138,In_2967);
or U775 (N_775,In_1861,In_2962);
or U776 (N_776,N_536,N_315);
xnor U777 (N_777,In_981,In_1885);
or U778 (N_778,N_533,In_1752);
nand U779 (N_779,In_2774,In_1493);
and U780 (N_780,N_265,In_2751);
nor U781 (N_781,In_1343,In_1777);
xor U782 (N_782,N_358,In_2421);
nor U783 (N_783,In_371,In_647);
or U784 (N_784,N_595,In_1354);
or U785 (N_785,N_53,In_1404);
and U786 (N_786,In_278,In_1148);
and U787 (N_787,N_372,In_1417);
nor U788 (N_788,N_403,N_20);
and U789 (N_789,In_1356,In_1841);
or U790 (N_790,In_2874,In_2085);
nand U791 (N_791,In_1943,In_1269);
xor U792 (N_792,In_2106,In_2653);
nand U793 (N_793,N_426,In_13);
xnor U794 (N_794,N_195,In_2603);
nor U795 (N_795,In_2971,In_2364);
nand U796 (N_796,In_2584,N_39);
or U797 (N_797,In_221,In_1745);
nor U798 (N_798,N_165,In_2052);
nand U799 (N_799,In_1217,In_1951);
nand U800 (N_800,In_143,In_1924);
and U801 (N_801,In_46,In_1251);
nand U802 (N_802,In_2402,In_2190);
and U803 (N_803,In_2184,In_1859);
nor U804 (N_804,In_667,N_654);
xor U805 (N_805,In_196,In_2483);
or U806 (N_806,In_863,In_1161);
xnor U807 (N_807,In_2318,In_448);
nor U808 (N_808,In_105,In_2815);
xnor U809 (N_809,In_2554,In_577);
xnor U810 (N_810,N_216,In_244);
or U811 (N_811,In_1108,N_316);
nor U812 (N_812,N_519,N_252);
xor U813 (N_813,In_403,N_294);
nor U814 (N_814,In_1897,In_1002);
nand U815 (N_815,In_50,In_2782);
nand U816 (N_816,N_624,In_646);
nand U817 (N_817,In_2168,In_101);
nor U818 (N_818,In_2380,In_2245);
and U819 (N_819,In_1977,In_1162);
nor U820 (N_820,In_2803,In_1766);
nor U821 (N_821,In_437,In_417);
nand U822 (N_822,In_1301,In_183);
and U823 (N_823,In_1966,N_258);
xnor U824 (N_824,In_223,In_2674);
nor U825 (N_825,N_214,In_2046);
and U826 (N_826,In_2656,In_2836);
nor U827 (N_827,In_2852,N_441);
nor U828 (N_828,N_476,In_1105);
xnor U829 (N_829,In_78,In_2075);
nand U830 (N_830,In_1177,In_607);
nand U831 (N_831,In_2098,N_692);
xnor U832 (N_832,In_1047,In_260);
xor U833 (N_833,N_73,In_291);
or U834 (N_834,In_1856,In_385);
xor U835 (N_835,In_418,In_712);
nand U836 (N_836,In_1901,In_719);
or U837 (N_837,In_709,In_2269);
and U838 (N_838,In_1176,N_504);
nor U839 (N_839,In_1167,In_1023);
xor U840 (N_840,N_9,N_383);
nand U841 (N_841,In_2868,N_138);
xnor U842 (N_842,N_412,In_1750);
nor U843 (N_843,In_2423,In_1481);
xnor U844 (N_844,N_526,In_1756);
nor U845 (N_845,N_546,In_1232);
and U846 (N_846,N_636,N_194);
and U847 (N_847,In_515,In_1035);
or U848 (N_848,In_309,In_2551);
nor U849 (N_849,In_253,In_179);
nand U850 (N_850,In_2963,In_1864);
nand U851 (N_851,In_177,In_1516);
and U852 (N_852,In_1206,In_1791);
or U853 (N_853,In_2509,In_800);
or U854 (N_854,In_235,In_1937);
and U855 (N_855,In_2059,In_1589);
and U856 (N_856,N_268,In_389);
or U857 (N_857,In_1616,In_1535);
nand U858 (N_858,In_2706,N_597);
or U859 (N_859,In_2023,N_176);
xnor U860 (N_860,In_658,In_2267);
nand U861 (N_861,N_545,In_1504);
or U862 (N_862,In_234,In_586);
nand U863 (N_863,In_2439,In_779);
nor U864 (N_864,N_588,In_2181);
or U865 (N_865,In_440,In_421);
or U866 (N_866,In_769,In_1024);
xnor U867 (N_867,N_484,In_645);
or U868 (N_868,In_878,In_216);
and U869 (N_869,In_380,In_2995);
and U870 (N_870,In_2322,In_2158);
xor U871 (N_871,In_259,In_142);
and U872 (N_872,N_482,In_158);
or U873 (N_873,In_1716,In_1062);
and U874 (N_874,N_583,In_770);
or U875 (N_875,In_1229,In_2555);
nand U876 (N_876,In_1074,In_232);
nor U877 (N_877,In_1705,In_949);
or U878 (N_878,N_753,In_2213);
nor U879 (N_879,In_2895,In_1157);
xnor U880 (N_880,N_418,N_392);
nand U881 (N_881,In_2208,In_2358);
nor U882 (N_882,In_499,N_94);
nor U883 (N_883,In_1111,In_869);
nand U884 (N_884,N_308,N_163);
and U885 (N_885,In_673,In_1254);
xor U886 (N_886,In_1101,In_1540);
or U887 (N_887,In_1146,In_1518);
and U888 (N_888,In_406,N_448);
xor U889 (N_889,N_233,N_303);
and U890 (N_890,In_170,In_2196);
and U891 (N_891,In_772,In_980);
nor U892 (N_892,N_609,In_837);
or U893 (N_893,In_2580,In_2624);
xnor U894 (N_894,In_1015,In_2741);
and U895 (N_895,In_2431,In_1165);
or U896 (N_896,In_1647,In_847);
nand U897 (N_897,In_127,N_565);
nor U898 (N_898,In_1630,In_2504);
or U899 (N_899,N_415,N_371);
xnor U900 (N_900,In_919,In_1744);
nand U901 (N_901,N_758,In_1722);
nor U902 (N_902,N_225,In_66);
xor U903 (N_903,In_2701,In_670);
xnor U904 (N_904,In_2886,In_224);
nor U905 (N_905,In_1521,In_12);
nand U906 (N_906,In_886,In_2437);
and U907 (N_907,In_843,In_2883);
and U908 (N_908,In_2244,In_1119);
nor U909 (N_909,In_689,In_1334);
and U910 (N_910,N_495,N_723);
nand U911 (N_911,In_2692,In_1160);
and U912 (N_912,In_1385,In_2924);
nand U913 (N_913,In_2825,In_2061);
or U914 (N_914,N_283,N_41);
and U915 (N_915,In_2077,In_1142);
and U916 (N_916,N_475,In_1231);
and U917 (N_917,In_911,In_2918);
nand U918 (N_918,N_505,In_1796);
nand U919 (N_919,In_43,In_81);
or U920 (N_920,In_2862,In_2559);
nand U921 (N_921,In_1664,N_191);
nand U922 (N_922,In_160,In_2927);
xnor U923 (N_923,In_203,In_381);
and U924 (N_924,In_2157,In_6);
and U925 (N_925,In_1078,In_1490);
nand U926 (N_926,In_114,In_929);
or U927 (N_927,In_1640,In_2985);
nor U928 (N_928,In_2546,In_2915);
and U929 (N_929,N_741,In_2058);
and U930 (N_930,N_657,N_429);
or U931 (N_931,In_2019,N_664);
nand U932 (N_932,N_559,In_555);
nand U933 (N_933,In_1667,In_546);
or U934 (N_934,N_788,In_968);
nand U935 (N_935,In_637,In_791);
or U936 (N_936,In_1608,In_2484);
nand U937 (N_937,In_2880,In_697);
nor U938 (N_938,In_703,N_757);
and U939 (N_939,N_754,In_1087);
nor U940 (N_940,N_596,In_1957);
nor U941 (N_941,In_463,In_1372);
xnor U942 (N_942,In_2758,N_591);
xnor U943 (N_943,In_1639,In_2060);
and U944 (N_944,In_191,N_113);
and U945 (N_945,In_118,In_1879);
nand U946 (N_946,In_1379,In_1084);
nand U947 (N_947,In_1538,In_2287);
xor U948 (N_948,In_2537,N_765);
nand U949 (N_949,In_2896,In_336);
nand U950 (N_950,In_1878,N_566);
nand U951 (N_951,In_368,N_364);
and U952 (N_952,N_486,N_498);
nand U953 (N_953,In_1670,N_65);
nor U954 (N_954,In_1830,In_953);
or U955 (N_955,N_674,In_1094);
xor U956 (N_956,In_542,In_1785);
and U957 (N_957,N_290,In_1369);
or U958 (N_958,N_608,In_453);
nand U959 (N_959,In_608,In_547);
nor U960 (N_960,In_2356,In_2365);
xor U961 (N_961,N_725,N_667);
and U962 (N_962,N_451,In_1000);
and U963 (N_963,In_2449,N_496);
or U964 (N_964,N_679,In_2042);
and U965 (N_965,In_1037,N_761);
nor U966 (N_966,N_406,In_761);
and U967 (N_967,In_59,N_739);
nor U968 (N_968,In_1091,In_2420);
or U969 (N_969,N_594,In_1890);
or U970 (N_970,In_549,In_2721);
and U971 (N_971,In_1846,In_1234);
nor U972 (N_972,In_2864,In_1496);
xor U973 (N_973,In_405,N_456);
and U974 (N_974,N_786,In_1799);
nand U975 (N_975,N_575,In_2590);
or U976 (N_976,N_769,In_2204);
xnor U977 (N_977,In_1454,In_522);
nand U978 (N_978,N_345,In_1614);
xnor U979 (N_979,In_2242,In_1473);
nor U980 (N_980,In_1576,N_510);
or U981 (N_981,In_2086,In_2176);
and U982 (N_982,In_2391,In_591);
and U983 (N_983,In_396,In_1923);
or U984 (N_984,In_205,In_83);
nor U985 (N_985,N_539,In_2413);
xnor U986 (N_986,In_1908,N_708);
nor U987 (N_987,In_1191,In_1778);
nor U988 (N_988,N_639,In_27);
or U989 (N_989,N_104,In_718);
xnor U990 (N_990,In_2611,N_152);
or U991 (N_991,N_333,In_620);
or U992 (N_992,N_748,In_2978);
and U993 (N_993,In_2164,In_1829);
and U994 (N_994,In_545,In_1034);
nor U995 (N_995,In_2581,In_531);
nand U996 (N_996,N_230,In_864);
or U997 (N_997,N_742,In_2360);
nand U998 (N_998,In_2947,In_629);
nor U999 (N_999,In_2720,In_2528);
nand U1000 (N_1000,In_2462,In_282);
nand U1001 (N_1001,In_1650,In_56);
nor U1002 (N_1002,In_965,In_1474);
or U1003 (N_1003,In_481,N_641);
or U1004 (N_1004,In_2443,N_709);
and U1005 (N_1005,N_159,In_135);
nor U1006 (N_1006,In_1141,N_652);
and U1007 (N_1007,N_977,In_1934);
and U1008 (N_1008,In_1286,In_2197);
or U1009 (N_1009,In_2535,In_153);
nand U1010 (N_1010,N_459,N_665);
and U1011 (N_1011,In_754,In_1082);
nand U1012 (N_1012,In_2921,In_2743);
nand U1013 (N_1013,N_55,In_341);
nand U1014 (N_1014,In_2951,In_422);
or U1015 (N_1015,In_1086,N_168);
or U1016 (N_1016,N_227,N_145);
nor U1017 (N_1017,In_1965,In_2923);
nand U1018 (N_1018,In_327,N_902);
nor U1019 (N_1019,In_458,In_682);
nand U1020 (N_1020,N_939,In_470);
or U1021 (N_1021,In_677,In_603);
xnor U1022 (N_1022,N_330,In_2788);
or U1023 (N_1023,N_250,In_1761);
nand U1024 (N_1024,N_980,In_1641);
nand U1025 (N_1025,In_2623,In_1578);
xnor U1026 (N_1026,In_1075,N_873);
and U1027 (N_1027,N_354,N_86);
xor U1028 (N_1028,In_705,N_96);
xnor U1029 (N_1029,N_390,N_530);
nand U1030 (N_1030,In_2180,In_2677);
nor U1031 (N_1031,In_1411,N_578);
and U1032 (N_1032,N_911,In_1911);
or U1033 (N_1033,In_1470,N_728);
nor U1034 (N_1034,N_204,In_2469);
or U1035 (N_1035,In_633,In_1548);
and U1036 (N_1036,N_359,N_273);
xnor U1037 (N_1037,N_992,N_756);
nand U1038 (N_1038,In_687,In_921);
and U1039 (N_1039,In_280,In_409);
and U1040 (N_1040,In_2126,In_2644);
or U1041 (N_1041,N_627,In_1227);
nor U1042 (N_1042,N_740,In_1573);
and U1043 (N_1043,In_2847,In_2438);
nand U1044 (N_1044,In_1605,In_103);
or U1045 (N_1045,In_2669,N_979);
xor U1046 (N_1046,In_2179,In_2865);
or U1047 (N_1047,N_36,In_1534);
nand U1048 (N_1048,In_2688,N_764);
nand U1049 (N_1049,In_1491,In_340);
or U1050 (N_1050,In_1046,In_1325);
or U1051 (N_1051,In_1567,In_829);
nor U1052 (N_1052,In_35,N_831);
or U1053 (N_1053,N_481,N_777);
xnor U1054 (N_1054,N_821,N_961);
or U1055 (N_1055,In_2614,In_1054);
xnor U1056 (N_1056,N_231,In_2685);
xor U1057 (N_1057,N_937,N_837);
nand U1058 (N_1058,In_934,In_875);
nand U1059 (N_1059,In_808,N_576);
or U1060 (N_1060,In_2274,N_931);
xor U1061 (N_1061,N_663,In_2165);
nor U1062 (N_1062,In_264,N_767);
nor U1063 (N_1063,In_1008,N_860);
xor U1064 (N_1064,N_548,In_2276);
and U1065 (N_1065,In_1403,In_2557);
nor U1066 (N_1066,In_2996,In_831);
nor U1067 (N_1067,In_1033,In_2343);
or U1068 (N_1068,In_374,In_251);
or U1069 (N_1069,N_929,N_221);
or U1070 (N_1070,N_18,In_2853);
or U1071 (N_1071,In_1685,In_392);
xnor U1072 (N_1072,In_1245,N_443);
xor U1073 (N_1073,In_122,In_2506);
and U1074 (N_1074,In_2816,In_1371);
and U1075 (N_1075,N_10,In_1988);
nand U1076 (N_1076,In_729,In_2406);
nand U1077 (N_1077,In_1056,In_1293);
and U1078 (N_1078,N_125,In_1585);
nand U1079 (N_1079,N_52,In_2004);
nand U1080 (N_1080,N_417,In_358);
and U1081 (N_1081,In_2560,In_2270);
and U1082 (N_1082,In_126,In_315);
nor U1083 (N_1083,In_2441,In_1730);
nor U1084 (N_1084,N_582,N_497);
or U1085 (N_1085,N_492,N_711);
and U1086 (N_1086,N_714,In_1014);
nor U1087 (N_1087,N_228,In_2633);
nor U1088 (N_1088,In_202,In_2547);
or U1089 (N_1089,N_672,N_590);
xor U1090 (N_1090,N_438,N_491);
nand U1091 (N_1091,In_1542,N_971);
nor U1092 (N_1092,In_151,N_432);
nand U1093 (N_1093,In_2202,In_2768);
nand U1094 (N_1094,N_564,In_1817);
nand U1095 (N_1095,N_169,In_429);
and U1096 (N_1096,In_973,In_125);
and U1097 (N_1097,In_2307,N_376);
xnor U1098 (N_1098,In_2138,In_397);
or U1099 (N_1099,In_2076,In_685);
xnor U1100 (N_1100,In_1873,In_1563);
or U1101 (N_1101,In_2903,N_478);
nor U1102 (N_1102,In_2536,N_770);
nand U1103 (N_1103,In_1787,N_611);
xnor U1104 (N_1104,In_1071,In_2264);
and U1105 (N_1105,N_569,In_1027);
xor U1106 (N_1106,N_968,In_241);
or U1107 (N_1107,In_1704,In_2540);
or U1108 (N_1108,In_1402,In_2152);
and U1109 (N_1109,N_457,N_919);
nor U1110 (N_1110,N_54,N_585);
nand U1111 (N_1111,In_2458,In_2932);
nor U1112 (N_1112,N_352,In_94);
or U1113 (N_1113,In_1526,In_1967);
and U1114 (N_1114,N_264,In_140);
and U1115 (N_1115,In_207,In_2261);
or U1116 (N_1116,In_987,In_1767);
nor U1117 (N_1117,N_389,N_970);
nor U1118 (N_1118,In_2736,N_284);
xor U1119 (N_1119,N_64,N_866);
and U1120 (N_1120,In_2464,In_1547);
nor U1121 (N_1121,N_422,N_858);
xnor U1122 (N_1122,In_2683,In_876);
nor U1123 (N_1123,In_867,N_688);
nand U1124 (N_1124,In_2454,In_1624);
nor U1125 (N_1125,In_312,N_219);
xnor U1126 (N_1126,In_2475,In_1892);
nor U1127 (N_1127,N_694,In_1236);
nand U1128 (N_1128,In_197,In_536);
or U1129 (N_1129,N_798,N_462);
or U1130 (N_1130,N_800,In_443);
or U1131 (N_1131,N_130,In_1842);
or U1132 (N_1132,In_1635,In_1366);
nor U1133 (N_1133,In_1822,In_2914);
or U1134 (N_1134,In_1653,N_446);
nor U1135 (N_1135,N_997,N_419);
xor U1136 (N_1136,N_735,In_2531);
nor U1137 (N_1137,In_2231,N_737);
or U1138 (N_1138,In_743,In_1553);
and U1139 (N_1139,N_781,N_235);
or U1140 (N_1140,N_846,In_1457);
or U1141 (N_1141,In_1218,In_344);
nor U1142 (N_1142,N_644,In_2376);
or U1143 (N_1143,In_1985,In_1762);
or U1144 (N_1144,In_1353,In_2710);
nor U1145 (N_1145,In_2562,In_1706);
nand U1146 (N_1146,In_363,In_760);
nand U1147 (N_1147,In_1300,In_1104);
nor U1148 (N_1148,In_1939,In_195);
nand U1149 (N_1149,N_386,In_1669);
nand U1150 (N_1150,In_1281,In_93);
and U1151 (N_1151,In_2766,In_2630);
nor U1152 (N_1152,In_1205,N_341);
nand U1153 (N_1153,N_67,In_2908);
xnor U1154 (N_1154,In_1505,N_775);
xor U1155 (N_1155,In_2983,In_1485);
and U1156 (N_1156,N_463,In_527);
nor U1157 (N_1157,In_1164,N_782);
nand U1158 (N_1158,In_738,N_605);
nor U1159 (N_1159,In_2073,In_1680);
or U1160 (N_1160,In_2627,In_1826);
or U1161 (N_1161,In_2798,N_868);
and U1162 (N_1162,N_750,In_2387);
xor U1163 (N_1163,In_2342,N_543);
xnor U1164 (N_1164,In_889,In_2859);
and U1165 (N_1165,In_2500,In_2910);
xnor U1166 (N_1166,N_793,N_357);
or U1167 (N_1167,In_1495,In_638);
or U1168 (N_1168,In_2826,In_2616);
nand U1169 (N_1169,N_541,N_579);
or U1170 (N_1170,In_1714,In_983);
xnor U1171 (N_1171,In_1725,In_627);
or U1172 (N_1172,In_2845,In_2975);
or U1173 (N_1173,N_648,N_236);
nand U1174 (N_1174,N_996,N_848);
and U1175 (N_1175,N_832,In_2355);
and U1176 (N_1176,In_1263,N_762);
or U1177 (N_1177,N_527,In_853);
nand U1178 (N_1178,N_435,In_994);
and U1179 (N_1179,In_1442,In_1009);
xnor U1180 (N_1180,N_774,N_822);
nand U1181 (N_1181,In_2263,In_1998);
nand U1182 (N_1182,N_710,In_619);
nand U1183 (N_1183,N_823,In_1831);
or U1184 (N_1184,In_2598,In_2485);
xor U1185 (N_1185,In_121,In_892);
nor U1186 (N_1186,In_1004,In_940);
xor U1187 (N_1187,In_1721,N_332);
and U1188 (N_1188,In_865,N_362);
or U1189 (N_1189,In_1130,N_82);
and U1190 (N_1190,In_1423,N_499);
nand U1191 (N_1191,In_979,N_38);
nand U1192 (N_1192,N_658,In_2779);
xor U1193 (N_1193,N_960,In_2965);
xnor U1194 (N_1194,N_633,In_2930);
or U1195 (N_1195,N_37,In_2642);
nand U1196 (N_1196,In_2292,N_870);
xor U1197 (N_1197,N_819,N_186);
nand U1198 (N_1198,N_938,In_1913);
nand U1199 (N_1199,N_340,In_2481);
nor U1200 (N_1200,In_777,N_801);
or U1201 (N_1201,N_1043,In_681);
and U1202 (N_1202,In_277,N_269);
and U1203 (N_1203,In_1140,In_2185);
xor U1204 (N_1204,In_1832,In_320);
xor U1205 (N_1205,In_1388,In_1764);
xnor U1206 (N_1206,N_1111,N_720);
and U1207 (N_1207,In_756,In_286);
xor U1208 (N_1208,N_1118,N_900);
and U1209 (N_1209,N_494,N_201);
or U1210 (N_1210,N_1172,N_1082);
nand U1211 (N_1211,In_1607,In_764);
or U1212 (N_1212,N_952,N_1029);
nand U1213 (N_1213,In_2226,N_328);
nor U1214 (N_1214,In_1801,N_206);
xnor U1215 (N_1215,N_1140,N_1145);
or U1216 (N_1216,In_296,N_879);
or U1217 (N_1217,In_2262,N_512);
and U1218 (N_1218,In_15,In_1230);
or U1219 (N_1219,N_1103,In_321);
or U1220 (N_1220,N_988,N_129);
or U1221 (N_1221,In_1012,In_1788);
and U1222 (N_1222,N_779,In_2857);
or U1223 (N_1223,N_489,In_817);
nand U1224 (N_1224,N_66,N_1105);
xor U1225 (N_1225,In_1106,In_739);
xnor U1226 (N_1226,In_1482,N_893);
nand U1227 (N_1227,N_101,In_930);
nand U1228 (N_1228,In_1918,N_778);
xor U1229 (N_1229,In_1198,In_384);
xnor U1230 (N_1230,N_1025,N_121);
and U1231 (N_1231,N_365,N_1121);
and U1232 (N_1232,In_2646,N_953);
nor U1233 (N_1233,In_2445,In_86);
xor U1234 (N_1234,N_885,In_2337);
and U1235 (N_1235,In_1975,In_946);
and U1236 (N_1236,In_2295,In_1196);
xnor U1237 (N_1237,In_1931,In_538);
and U1238 (N_1238,In_962,In_427);
nand U1239 (N_1239,N_1045,In_753);
xor U1240 (N_1240,In_1555,N_178);
or U1241 (N_1241,In_1322,N_898);
and U1242 (N_1242,In_1619,In_95);
nor U1243 (N_1243,N_202,N_1027);
nor U1244 (N_1244,N_1134,N_1143);
nand U1245 (N_1245,N_166,In_1546);
xnor U1246 (N_1246,In_2687,N_414);
nand U1247 (N_1247,N_1196,N_623);
nor U1248 (N_1248,In_2143,In_435);
nand U1249 (N_1249,N_935,In_1936);
or U1250 (N_1250,In_660,In_2618);
and U1251 (N_1251,In_1380,In_781);
nand U1252 (N_1252,In_1103,N_1166);
and U1253 (N_1253,In_1941,N_382);
or U1254 (N_1254,In_187,In_1331);
and U1255 (N_1255,In_1810,N_329);
nand U1256 (N_1256,In_451,In_1816);
and U1257 (N_1257,N_521,N_867);
or U1258 (N_1258,N_1095,In_2036);
or U1259 (N_1259,N_915,In_390);
nand U1260 (N_1260,In_2761,N_682);
nand U1261 (N_1261,In_2950,N_572);
nand U1262 (N_1262,In_2199,N_745);
nor U1263 (N_1263,In_2681,In_902);
nor U1264 (N_1264,In_1466,In_879);
or U1265 (N_1265,N_1119,N_379);
and U1266 (N_1266,In_2136,In_423);
nand U1267 (N_1267,N_826,N_285);
nor U1268 (N_1268,In_2150,N_717);
and U1269 (N_1269,In_1682,N_606);
nor U1270 (N_1270,N_991,In_2256);
nor U1271 (N_1271,In_2224,N_483);
or U1272 (N_1272,N_936,In_2473);
or U1273 (N_1273,N_1019,N_716);
or U1274 (N_1274,In_665,In_1351);
nor U1275 (N_1275,In_1973,In_2735);
nand U1276 (N_1276,In_1364,In_1737);
nor U1277 (N_1277,N_794,In_274);
nand U1278 (N_1278,N_183,In_123);
xnor U1279 (N_1279,In_882,N_1167);
and U1280 (N_1280,In_1713,In_2635);
and U1281 (N_1281,In_1552,N_1141);
xor U1282 (N_1282,In_1193,In_849);
and U1283 (N_1283,In_1260,In_1673);
nand U1284 (N_1284,N_68,N_240);
xor U1285 (N_1285,In_1110,In_330);
or U1286 (N_1286,In_2444,N_1127);
xnor U1287 (N_1287,In_1676,N_511);
and U1288 (N_1288,In_839,In_1443);
nor U1289 (N_1289,N_193,In_1387);
nand U1290 (N_1290,In_1668,N_1157);
nor U1291 (N_1291,N_103,In_2118);
xor U1292 (N_1292,N_538,In_1665);
or U1293 (N_1293,In_2781,N_172);
and U1294 (N_1294,In_322,In_700);
nor U1295 (N_1295,In_433,N_683);
or U1296 (N_1296,In_1339,N_966);
xor U1297 (N_1297,N_199,N_637);
xor U1298 (N_1298,In_1837,In_2321);
nand U1299 (N_1299,N_442,In_2249);
nand U1300 (N_1300,In_1942,N_188);
and U1301 (N_1301,N_1093,N_618);
nor U1302 (N_1302,N_116,In_2599);
nor U1303 (N_1303,N_324,In_484);
or U1304 (N_1304,In_2109,In_159);
or U1305 (N_1305,In_1315,In_2549);
nor U1306 (N_1306,N_189,N_974);
and U1307 (N_1307,N_470,In_48);
and U1308 (N_1308,N_1039,In_1978);
nor U1309 (N_1309,N_622,N_616);
nor U1310 (N_1310,N_790,In_2759);
nand U1311 (N_1311,N_673,N_827);
and U1312 (N_1312,N_924,In_1592);
nand U1313 (N_1313,N_244,In_34);
xnor U1314 (N_1314,N_1073,In_1122);
or U1315 (N_1315,N_297,N_705);
or U1316 (N_1316,In_2802,In_2800);
and U1317 (N_1317,N_1046,N_555);
or U1318 (N_1318,In_548,In_1802);
xor U1319 (N_1319,In_145,In_1395);
and U1320 (N_1320,In_1710,In_1070);
and U1321 (N_1321,N_695,In_1137);
or U1322 (N_1322,In_1803,In_2936);
or U1323 (N_1323,In_2909,In_1525);
nand U1324 (N_1324,N_835,In_1361);
nand U1325 (N_1325,N_933,In_1626);
nor U1326 (N_1326,N_573,In_519);
nor U1327 (N_1327,N_836,In_102);
xnor U1328 (N_1328,N_686,In_2488);
nor U1329 (N_1329,In_33,N_398);
nor U1330 (N_1330,In_1793,N_562);
xor U1331 (N_1331,In_842,In_512);
and U1332 (N_1332,In_1881,N_626);
nand U1333 (N_1333,In_220,In_2776);
nor U1334 (N_1334,N_896,In_287);
xnor U1335 (N_1335,In_109,In_846);
and U1336 (N_1336,In_967,In_65);
nand U1337 (N_1337,In_1307,N_901);
nor U1338 (N_1338,N_891,In_1472);
xnor U1339 (N_1339,In_2595,In_22);
nand U1340 (N_1340,N_25,In_933);
nand U1341 (N_1341,In_1134,N_1057);
and U1342 (N_1342,In_111,N_440);
or U1343 (N_1343,In_1610,In_1100);
or U1344 (N_1344,In_276,In_2511);
nor U1345 (N_1345,N_1006,N_759);
nor U1346 (N_1346,In_338,In_2867);
xor U1347 (N_1347,In_314,In_2324);
nor U1348 (N_1348,N_1115,N_773);
and U1349 (N_1349,N_334,N_998);
nor U1350 (N_1350,In_37,N_436);
xnor U1351 (N_1351,In_275,In_1394);
and U1352 (N_1352,In_1798,N_632);
and U1353 (N_1353,N_387,In_1221);
nor U1354 (N_1354,In_2977,N_1124);
and U1355 (N_1355,N_517,In_1477);
nand U1356 (N_1356,N_1178,N_925);
or U1357 (N_1357,N_963,N_926);
and U1358 (N_1358,N_338,In_2577);
xnor U1359 (N_1359,In_1824,In_1503);
and U1360 (N_1360,N_24,N_732);
and U1361 (N_1361,N_646,N_1);
nand U1362 (N_1362,In_1059,N_124);
and U1363 (N_1363,In_413,N_506);
and U1364 (N_1364,N_281,N_854);
nand U1365 (N_1365,N_1065,In_334);
and U1366 (N_1366,N_649,In_652);
or U1367 (N_1367,N_1130,In_1338);
and U1368 (N_1368,N_60,In_1216);
xor U1369 (N_1369,N_535,In_1190);
or U1370 (N_1370,N_74,N_137);
nand U1371 (N_1371,In_54,In_347);
and U1372 (N_1372,In_1151,N_4);
or U1373 (N_1373,In_2041,N_807);
xnor U1374 (N_1374,N_377,In_2211);
or U1375 (N_1375,N_513,N_856);
xnor U1376 (N_1376,In_752,In_1709);
and U1377 (N_1377,N_825,N_142);
and U1378 (N_1378,N_859,N_185);
or U1379 (N_1379,In_826,In_2191);
and U1380 (N_1380,N_405,N_1033);
nor U1381 (N_1381,N_1086,In_2296);
nor U1382 (N_1382,In_2350,N_537);
or U1383 (N_1383,N_1078,In_736);
nand U1384 (N_1384,In_1444,In_2142);
xor U1385 (N_1385,In_945,N_733);
or U1386 (N_1386,N_525,In_956);
or U1387 (N_1387,In_2092,In_584);
nor U1388 (N_1388,In_813,N_941);
xor U1389 (N_1389,N_1176,N_1170);
or U1390 (N_1390,In_740,In_2451);
or U1391 (N_1391,N_266,In_1121);
xnor U1392 (N_1392,In_2608,In_2250);
xor U1393 (N_1393,In_905,N_628);
xor U1394 (N_1394,N_508,N_635);
nand U1395 (N_1395,In_1149,N_274);
nor U1396 (N_1396,In_598,N_275);
and U1397 (N_1397,In_1594,In_1460);
or U1398 (N_1398,N_1191,In_1273);
nand U1399 (N_1399,N_954,N_123);
and U1400 (N_1400,N_1250,N_1323);
or U1401 (N_1401,N_956,In_2022);
or U1402 (N_1402,N_455,In_2222);
or U1403 (N_1403,In_1440,In_2520);
or U1404 (N_1404,In_2561,N_1102);
or U1405 (N_1405,In_663,In_1880);
or U1406 (N_1406,In_2346,N_882);
and U1407 (N_1407,In_1724,In_589);
or U1408 (N_1408,In_2495,N_246);
nand U1409 (N_1409,N_1268,N_1353);
or U1410 (N_1410,In_810,In_604);
xor U1411 (N_1411,In_1644,N_554);
xnor U1412 (N_1412,N_1021,In_1848);
nor U1413 (N_1413,N_1260,N_895);
and U1414 (N_1414,In_45,In_2491);
or U1415 (N_1415,In_2892,N_842);
and U1416 (N_1416,N_983,N_47);
xor U1417 (N_1417,N_617,N_944);
nand U1418 (N_1418,In_1509,In_1256);
nor U1419 (N_1419,N_1224,N_1194);
and U1420 (N_1420,N_7,N_802);
and U1421 (N_1421,In_1930,N_271);
or U1422 (N_1422,N_106,In_2651);
or U1423 (N_1423,In_2153,N_964);
or U1424 (N_1424,In_951,In_1554);
nor U1425 (N_1425,N_411,In_2660);
and U1426 (N_1426,In_2998,In_844);
xnor U1427 (N_1427,In_214,In_1882);
or U1428 (N_1428,In_461,In_765);
and U1429 (N_1429,In_442,N_1060);
nor U1430 (N_1430,N_985,N_1308);
nand U1431 (N_1431,In_1872,In_425);
nor U1432 (N_1432,N_930,In_1170);
or U1433 (N_1433,In_1996,In_1097);
nor U1434 (N_1434,N_861,N_678);
nand U1435 (N_1435,In_2797,In_329);
nor U1436 (N_1436,In_2373,In_1844);
nor U1437 (N_1437,In_1223,In_1102);
nor U1438 (N_1438,N_1158,In_100);
and U1439 (N_1439,In_2821,N_619);
or U1440 (N_1440,N_1381,N_771);
nand U1441 (N_1441,In_2070,N_829);
and U1442 (N_1442,N_561,N_127);
nor U1443 (N_1443,In_2873,In_510);
and U1444 (N_1444,N_1305,In_977);
xnor U1445 (N_1445,In_2492,N_80);
nor U1446 (N_1446,N_817,N_1362);
nor U1447 (N_1447,In_1459,In_2831);
nand U1448 (N_1448,N_1116,In_997);
or U1449 (N_1449,In_1912,N_1149);
or U1450 (N_1450,N_847,In_1016);
or U1451 (N_1451,In_688,In_1041);
or U1452 (N_1452,In_757,In_771);
xor U1453 (N_1453,In_1812,In_242);
nor U1454 (N_1454,In_899,N_1350);
nor U1455 (N_1455,N_1251,In_428);
nand U1456 (N_1456,In_2422,N_1302);
nor U1457 (N_1457,In_2629,In_2325);
and U1458 (N_1458,N_1165,In_72);
and U1459 (N_1459,In_161,N_1316);
or U1460 (N_1460,N_408,In_438);
and U1461 (N_1461,N_118,N_157);
xor U1462 (N_1462,N_31,In_150);
xnor U1463 (N_1463,N_375,In_2785);
xor U1464 (N_1464,N_1375,In_2550);
nand U1465 (N_1465,In_219,In_457);
nor U1466 (N_1466,In_1729,In_1426);
and U1467 (N_1467,N_1233,N_922);
or U1468 (N_1468,In_23,In_893);
nand U1469 (N_1469,N_877,In_324);
nand U1470 (N_1470,N_987,N_1030);
or U1471 (N_1471,In_144,In_2478);
nand U1472 (N_1472,N_1334,N_1063);
nor U1473 (N_1473,In_2396,In_284);
nor U1474 (N_1474,In_382,In_1113);
xor U1475 (N_1475,N_1012,N_897);
or U1476 (N_1476,In_1131,In_773);
or U1477 (N_1477,N_350,N_1364);
nor U1478 (N_1478,N_581,N_1219);
nand U1479 (N_1479,N_1179,In_1486);
and U1480 (N_1480,In_728,In_2713);
or U1481 (N_1481,N_604,In_2543);
xnor U1482 (N_1482,In_543,In_2083);
or U1483 (N_1483,N_949,N_1055);
or U1484 (N_1484,N_841,N_187);
nor U1485 (N_1485,N_876,N_690);
xnor U1486 (N_1486,In_1586,N_428);
xor U1487 (N_1487,N_212,In_1487);
nand U1488 (N_1488,In_1154,In_117);
nor U1489 (N_1489,In_495,N_812);
or U1490 (N_1490,N_1247,In_2048);
nor U1491 (N_1491,In_2607,N_288);
or U1492 (N_1492,In_2097,In_969);
and U1493 (N_1493,N_947,In_803);
xnor U1494 (N_1494,In_2828,N_395);
nor U1495 (N_1495,In_71,In_2367);
nand U1496 (N_1496,In_2031,In_866);
and U1497 (N_1497,In_1875,N_724);
xnor U1498 (N_1498,N_845,In_860);
and U1499 (N_1499,N_811,In_2541);
xnor U1500 (N_1500,In_2209,N_689);
and U1501 (N_1501,N_1397,N_63);
nand U1502 (N_1502,N_1022,In_2002);
xnor U1503 (N_1503,N_1257,N_23);
and U1504 (N_1504,In_2024,N_335);
or U1505 (N_1505,N_1262,N_763);
or U1506 (N_1506,N_816,N_1164);
nor U1507 (N_1507,N_1238,In_2982);
nor U1508 (N_1508,In_215,In_1357);
nand U1509 (N_1509,N_712,N_477);
or U1510 (N_1510,In_2657,In_247);
nand U1511 (N_1511,In_1382,N_1284);
or U1512 (N_1512,N_905,N_208);
or U1513 (N_1513,N_1383,N_1005);
xor U1514 (N_1514,In_1884,N_1286);
and U1515 (N_1515,N_729,In_1976);
nor U1516 (N_1516,In_819,In_1003);
nand U1517 (N_1517,In_915,N_889);
and U1518 (N_1518,In_950,In_1916);
xor U1519 (N_1519,In_1239,N_918);
xnor U1520 (N_1520,In_2986,In_2917);
or U1521 (N_1521,In_1797,In_426);
and U1522 (N_1522,In_97,In_766);
and U1523 (N_1523,In_2650,N_549);
xor U1524 (N_1524,In_557,In_2173);
nor U1525 (N_1525,N_1227,In_407);
or U1526 (N_1526,In_2053,N_1040);
or U1527 (N_1527,N_91,In_2522);
nand U1528 (N_1528,In_2987,In_1159);
nand U1529 (N_1529,N_1177,N_890);
nor U1530 (N_1530,N_1009,N_1207);
and U1531 (N_1531,In_2332,N_917);
xor U1532 (N_1532,In_2671,In_2583);
or U1533 (N_1533,In_666,In_2470);
and U1534 (N_1534,N_1390,N_1263);
nand U1535 (N_1535,N_1342,In_98);
and U1536 (N_1536,N_1135,N_1120);
nand U1537 (N_1537,N_1023,In_1383);
nor U1538 (N_1538,In_708,In_2159);
or U1539 (N_1539,In_2715,In_2063);
or U1540 (N_1540,N_1256,In_2718);
nand U1541 (N_1541,In_1067,N_1265);
nand U1542 (N_1542,N_1097,N_466);
nor U1543 (N_1543,N_367,N_1083);
nor U1544 (N_1544,N_584,In_64);
nor U1545 (N_1545,N_601,N_813);
and U1546 (N_1546,N_928,In_1451);
xnor U1547 (N_1547,N_570,N_300);
or U1548 (N_1548,In_2672,N_1229);
or U1549 (N_1549,In_2225,N_1035);
nand U1550 (N_1550,N_1337,N_659);
nor U1551 (N_1551,In_110,In_995);
or U1552 (N_1552,In_1627,In_1220);
nand U1553 (N_1553,In_1425,N_730);
xnor U1554 (N_1554,N_907,N_914);
nand U1555 (N_1555,In_467,N_314);
or U1556 (N_1556,N_360,In_1007);
or U1557 (N_1557,N_863,In_2317);
or U1558 (N_1558,N_529,N_464);
and U1559 (N_1559,N_843,In_269);
nand U1560 (N_1560,N_540,In_2784);
nand U1561 (N_1561,N_1010,N_282);
nor U1562 (N_1562,In_1210,N_1066);
or U1563 (N_1563,N_404,N_887);
or U1564 (N_1564,N_1321,In_55);
or U1565 (N_1565,In_1904,N_1281);
nand U1566 (N_1566,In_2279,N_1211);
or U1567 (N_1567,In_745,N_1355);
xor U1568 (N_1568,In_1698,In_1235);
xor U1569 (N_1569,In_2668,In_1854);
and U1570 (N_1570,In_2638,In_923);
and U1571 (N_1571,In_801,In_1259);
nand U1572 (N_1572,In_2471,N_799);
or U1573 (N_1573,N_262,N_1289);
nor U1574 (N_1574,In_2960,In_2658);
and U1575 (N_1575,N_1369,In_2969);
nor U1576 (N_1576,In_593,N_361);
or U1577 (N_1577,N_1349,In_613);
nor U1578 (N_1578,In_2548,N_1266);
or U1579 (N_1579,In_848,In_2755);
nand U1580 (N_1580,N_1159,N_1190);
or U1581 (N_1581,N_1218,N_853);
and U1582 (N_1582,In_694,In_1362);
or U1583 (N_1583,N_320,In_931);
nand U1584 (N_1584,N_1340,In_1609);
nand U1585 (N_1585,N_1131,N_14);
and U1586 (N_1586,N_888,N_1259);
nor U1587 (N_1587,In_938,In_2659);
nor U1588 (N_1588,N_981,N_1231);
nand U1589 (N_1589,In_2021,N_1212);
or U1590 (N_1590,N_229,In_2591);
xor U1591 (N_1591,N_869,In_1284);
xnor U1592 (N_1592,N_815,In_2905);
nor U1593 (N_1593,In_2992,In_155);
or U1594 (N_1594,N_932,N_792);
nand U1595 (N_1595,In_2775,In_1969);
and U1596 (N_1596,In_2218,N_1371);
and U1597 (N_1597,N_631,N_1189);
nor U1598 (N_1598,In_307,In_1806);
nor U1599 (N_1599,In_268,In_1917);
xnor U1600 (N_1600,N_1449,In_1688);
nand U1601 (N_1601,N_1173,In_514);
nand U1602 (N_1602,In_152,In_1568);
nand U1603 (N_1603,N_1530,In_642);
nand U1604 (N_1604,In_129,N_131);
and U1605 (N_1605,N_1455,In_1940);
nor U1606 (N_1606,N_1228,In_1478);
nand U1607 (N_1607,N_500,In_1981);
xor U1608 (N_1608,N_1499,In_2145);
nand U1609 (N_1609,N_1114,N_76);
and U1610 (N_1610,In_89,In_401);
and U1611 (N_1611,N_577,N_1405);
or U1612 (N_1612,In_796,N_1155);
nor U1613 (N_1613,N_834,In_2570);
nor U1614 (N_1614,In_87,N_1110);
and U1615 (N_1615,In_1727,In_1083);
and U1616 (N_1616,In_1689,N_603);
xor U1617 (N_1617,In_2855,N_1104);
xnor U1618 (N_1618,In_184,N_1283);
and U1619 (N_1619,In_2876,In_350);
nor U1620 (N_1620,In_517,In_2327);
nor U1621 (N_1621,In_1863,In_1579);
nor U1622 (N_1622,N_342,N_680);
nand U1623 (N_1623,N_849,N_1053);
nor U1624 (N_1624,In_566,N_910);
or U1625 (N_1625,In_763,N_1223);
nand U1626 (N_1626,N_785,In_2435);
nor U1627 (N_1627,In_838,In_854);
nor U1628 (N_1628,N_1548,N_698);
and U1629 (N_1629,N_693,N_894);
or U1630 (N_1630,N_1090,N_1388);
nor U1631 (N_1631,In_2111,N_1365);
nor U1632 (N_1632,In_2344,N_423);
and U1633 (N_1633,N_1456,In_2851);
nor U1634 (N_1634,N_828,N_35);
nand U1635 (N_1635,N_1574,N_1447);
xor U1636 (N_1636,In_1571,N_1142);
nand U1637 (N_1637,N_615,N_1048);
and U1638 (N_1638,N_1199,In_1401);
and U1639 (N_1639,In_523,N_1422);
nor U1640 (N_1640,N_289,N_1129);
xor U1641 (N_1641,N_291,N_746);
or U1642 (N_1642,N_805,In_1501);
xnor U1643 (N_1643,N_662,N_824);
nor U1644 (N_1644,N_318,N_1113);
nor U1645 (N_1645,In_1381,N_943);
nand U1646 (N_1646,N_1493,N_1293);
and U1647 (N_1647,N_1593,N_986);
or U1648 (N_1648,N_976,In_1194);
xor U1649 (N_1649,N_1592,In_2237);
xor U1650 (N_1650,In_1065,N_1413);
nand U1651 (N_1651,N_1325,In_2870);
or U1652 (N_1652,N_223,N_1324);
nand U1653 (N_1653,N_744,N_1377);
nand U1654 (N_1654,N_1357,N_776);
nand U1655 (N_1655,In_2131,N_1287);
or U1656 (N_1656,N_1382,In_1118);
nand U1657 (N_1657,N_1453,N_681);
or U1658 (N_1658,N_167,N_1184);
and U1659 (N_1659,N_198,In_415);
and U1660 (N_1660,N_111,N_948);
nor U1661 (N_1661,N_1152,N_1004);
or U1662 (N_1662,In_1905,In_2833);
nor U1663 (N_1663,N_468,N_1421);
xnor U1664 (N_1664,In_2919,N_1431);
xor U1665 (N_1665,N_1581,In_2429);
nand U1666 (N_1666,N_1156,N_1392);
or U1667 (N_1667,N_940,N_1559);
nor U1668 (N_1668,N_1434,N_653);
nand U1669 (N_1669,N_19,In_1020);
and U1670 (N_1670,In_1603,N_687);
nor U1671 (N_1671,N_1486,N_958);
xor U1672 (N_1672,N_1269,N_1557);
or U1673 (N_1673,In_489,N_1037);
nand U1674 (N_1674,N_373,N_1523);
nor U1675 (N_1675,N_1556,In_2860);
nor U1676 (N_1676,N_625,In_2840);
or U1677 (N_1677,N_1500,N_713);
xnor U1678 (N_1678,In_2752,N_1571);
xor U1679 (N_1679,N_1358,N_1106);
nor U1680 (N_1680,In_2789,N_1311);
and U1681 (N_1681,N_1002,N_804);
or U1682 (N_1682,N_108,N_607);
nand U1683 (N_1683,N_994,In_751);
nand U1684 (N_1684,N_1125,In_2844);
nor U1685 (N_1685,In_588,In_1344);
nor U1686 (N_1686,In_2476,N_1524);
nand U1687 (N_1687,N_1558,N_990);
or U1688 (N_1688,N_507,N_222);
or U1689 (N_1689,N_1506,In_2354);
nand U1690 (N_1690,In_1393,N_978);
and U1691 (N_1691,N_353,In_281);
and U1692 (N_1692,N_1570,N_1249);
nand U1693 (N_1693,In_2762,N_1069);
xnor U1694 (N_1694,In_14,N_1261);
xor U1695 (N_1695,N_1169,In_1701);
nor U1696 (N_1696,N_1061,In_2678);
and U1697 (N_1697,In_731,N_1374);
and U1698 (N_1698,In_2155,N_916);
xor U1699 (N_1699,In_2416,In_139);
nand U1700 (N_1700,N_102,N_1050);
xnor U1701 (N_1701,In_1963,N_1071);
nor U1702 (N_1702,In_2319,N_1451);
xor U1703 (N_1703,N_99,N_727);
and U1704 (N_1704,In_2780,In_2008);
nand U1705 (N_1705,N_1575,In_1954);
and U1706 (N_1706,In_1612,In_1889);
xnor U1707 (N_1707,In_1663,N_1322);
nand U1708 (N_1708,N_1384,In_2372);
nand U1709 (N_1709,N_1237,In_610);
or U1710 (N_1710,In_2379,In_1696);
nor U1711 (N_1711,N_1503,N_731);
or U1712 (N_1712,N_374,In_1328);
or U1713 (N_1713,In_1774,In_827);
nand U1714 (N_1714,In_914,N_1254);
nand U1715 (N_1715,In_359,In_2696);
nor U1716 (N_1716,N_1085,N_1497);
xor U1717 (N_1717,N_1264,N_1175);
or U1718 (N_1718,N_1052,N_128);
or U1719 (N_1719,N_325,N_1563);
or U1720 (N_1720,In_2220,N_1551);
or U1721 (N_1721,N_1533,In_2592);
or U1722 (N_1722,N_1015,N_904);
nor U1723 (N_1723,N_1016,N_15);
nor U1724 (N_1724,In_1126,In_2025);
and U1725 (N_1725,N_1341,N_1122);
xor U1726 (N_1726,N_1536,In_2336);
nor U1727 (N_1727,N_1013,N_1274);
nor U1728 (N_1728,In_585,In_1422);
and U1729 (N_1729,In_1201,N_1344);
xnor U1730 (N_1730,N_1018,In_493);
or U1731 (N_1731,N_1361,In_2123);
or U1732 (N_1732,N_1534,N_972);
xnor U1733 (N_1733,N_514,N_279);
xor U1734 (N_1734,N_1202,N_1042);
nand U1735 (N_1735,N_1525,N_934);
xor U1736 (N_1736,N_1154,N_1351);
nor U1737 (N_1737,N_975,N_322);
xnor U1738 (N_1738,N_85,N_1560);
nand U1739 (N_1739,N_1276,In_471);
or U1740 (N_1740,N_453,In_2730);
nand U1741 (N_1741,N_772,N_1590);
xor U1742 (N_1742,N_1531,N_22);
nor U1743 (N_1743,In_2314,N_1394);
xnor U1744 (N_1744,In_1894,In_2272);
and U1745 (N_1745,In_1860,In_1341);
or U1746 (N_1746,N_1441,N_1094);
nand U1747 (N_1747,N_1288,N_1128);
and U1748 (N_1748,In_1587,N_957);
nor U1749 (N_1749,In_2144,In_1959);
nand U1750 (N_1750,In_579,N_132);
nand U1751 (N_1751,N_1317,N_1468);
or U1752 (N_1752,In_2530,In_410);
and U1753 (N_1753,N_851,N_1304);
or U1754 (N_1754,In_261,N_736);
or U1755 (N_1755,In_2891,N_1187);
nor U1756 (N_1756,In_1599,N_450);
nand U1757 (N_1757,In_2579,In_395);
nor U1758 (N_1758,N_1295,N_1579);
and U1759 (N_1759,In_2834,In_2174);
xor U1760 (N_1760,N_1402,In_1480);
nor U1761 (N_1761,In_316,In_365);
nand U1762 (N_1762,N_1398,N_1391);
and U1763 (N_1763,N_263,In_1849);
nand U1764 (N_1764,In_1790,N_946);
or U1765 (N_1765,N_56,N_722);
nand U1766 (N_1766,N_1414,N_1299);
or U1767 (N_1767,N_1395,N_1424);
or U1768 (N_1768,N_209,In_4);
xor U1769 (N_1769,In_1675,N_1292);
xnor U1770 (N_1770,In_2585,N_1074);
or U1771 (N_1771,N_1282,In_2426);
or U1772 (N_1772,N_580,N_78);
xor U1773 (N_1773,In_492,N_1038);
xor U1774 (N_1774,N_1181,In_289);
and U1775 (N_1775,N_1367,In_2192);
or U1776 (N_1776,In_116,In_1271);
nand U1777 (N_1777,N_598,N_668);
xnor U1778 (N_1778,In_2820,N_1472);
nor U1779 (N_1779,In_861,In_634);
nor U1780 (N_1780,N_528,In_2866);
nor U1781 (N_1781,N_1478,In_750);
or U1782 (N_1782,N_1075,In_1654);
nor U1783 (N_1783,N_1026,N_400);
nor U1784 (N_1784,N_784,N_1535);
nor U1785 (N_1785,N_293,In_587);
and U1786 (N_1786,N_1517,In_2899);
xnor U1787 (N_1787,N_1279,In_2931);
nor U1788 (N_1788,N_1151,In_611);
and U1789 (N_1789,In_2374,N_1185);
and U1790 (N_1790,N_1385,N_1285);
nand U1791 (N_1791,N_1335,N_620);
and U1792 (N_1792,N_969,N_806);
and U1793 (N_1793,N_1183,In_562);
and U1794 (N_1794,N_421,In_1448);
xnor U1795 (N_1795,In_1510,N_638);
and U1796 (N_1796,In_683,N_385);
xor U1797 (N_1797,N_1538,N_1214);
nor U1798 (N_1798,In_372,In_2619);
nand U1799 (N_1799,In_966,In_2074);
nor U1800 (N_1800,N_1748,N_349);
or U1801 (N_1801,N_1051,N_1352);
and U1802 (N_1802,In_2201,N_965);
and U1803 (N_1803,N_1795,In_1172);
and U1804 (N_1804,N_1703,N_1644);
nand U1805 (N_1805,In_1500,In_2403);
nand U1806 (N_1806,N_1688,N_1528);
nor U1807 (N_1807,N_1651,N_1062);
and U1808 (N_1808,N_1514,N_1480);
nand U1809 (N_1809,N_260,N_1628);
nand U1810 (N_1810,In_834,N_1147);
or U1811 (N_1811,N_1632,N_58);
or U1812 (N_1812,In_625,N_1790);
xnor U1813 (N_1813,In_1017,In_332);
or U1814 (N_1814,N_1077,N_531);
nor U1815 (N_1815,In_2640,In_506);
xnor U1816 (N_1816,In_2105,In_229);
nand U1817 (N_1817,N_424,N_1297);
and U1818 (N_1818,N_1682,In_720);
or U1819 (N_1819,In_1290,N_1762);
nor U1820 (N_1820,N_691,N_989);
nand U1821 (N_1821,In_2808,In_928);
xor U1822 (N_1822,N_1403,N_1665);
nor U1823 (N_1823,N_1521,In_723);
or U1824 (N_1824,N_1047,In_2772);
or U1825 (N_1825,In_516,In_1208);
xor U1826 (N_1826,N_485,N_906);
or U1827 (N_1827,In_1633,In_1659);
or U1828 (N_1828,In_360,N_1419);
and U1829 (N_1829,In_807,N_1720);
xor U1830 (N_1830,N_1734,N_660);
nor U1831 (N_1831,N_149,N_1784);
nand U1832 (N_1832,N_1522,N_671);
and U1833 (N_1833,N_1621,N_1485);
or U1834 (N_1834,N_1791,N_1188);
nand U1835 (N_1835,N_1273,In_2115);
nor U1836 (N_1836,In_2533,N_1137);
nor U1837 (N_1837,N_40,N_629);
and U1838 (N_1838,N_1476,N_1691);
xor U1839 (N_1839,N_1603,N_220);
xnor U1840 (N_1840,In_1279,In_2178);
or U1841 (N_1841,In_2436,N_1796);
nor U1842 (N_1842,N_1512,In_2146);
and U1843 (N_1843,N_388,N_558);
nand U1844 (N_1844,In_1195,N_249);
xor U1845 (N_1845,N_1519,In_786);
xor U1846 (N_1846,N_1680,In_1476);
and U1847 (N_1847,N_1408,N_1730);
or U1848 (N_1848,In_2442,N_1221);
nand U1849 (N_1849,N_154,N_640);
xnor U1850 (N_1850,N_1539,N_700);
nor U1851 (N_1851,In_439,In_108);
and U1852 (N_1852,N_726,N_1123);
nor U1853 (N_1853,N_871,N_1561);
nand U1854 (N_1854,In_505,N_1275);
and U1855 (N_1855,In_676,N_927);
or U1856 (N_1856,N_1049,N_431);
nor U1857 (N_1857,N_1649,N_751);
xor U1858 (N_1858,In_1186,N_1595);
nand U1859 (N_1859,N_1003,N_647);
nand U1860 (N_1860,In_474,In_1748);
nand U1861 (N_1861,N_1689,N_1008);
nand U1862 (N_1862,In_250,In_364);
nor U1863 (N_1863,N_1442,N_1686);
or U1864 (N_1864,N_1309,In_741);
or U1865 (N_1865,N_257,N_1461);
or U1866 (N_1866,In_871,N_1108);
nand U1867 (N_1867,N_1240,In_39);
xnor U1868 (N_1868,N_1704,N_1741);
nor U1869 (N_1869,N_1126,N_1604);
nand U1870 (N_1870,In_1247,In_2524);
or U1871 (N_1871,In_1956,N_1630);
xor U1872 (N_1872,In_2113,N_1638);
nand U1873 (N_1873,N_1589,In_1621);
or U1874 (N_1874,In_2260,In_163);
and U1875 (N_1875,N_1246,N_337);
and U1876 (N_1876,In_1513,N_1726);
and U1877 (N_1877,In_1458,N_161);
nand U1878 (N_1878,N_1024,In_2711);
or U1879 (N_1879,In_2753,N_1709);
nand U1880 (N_1880,In_2456,In_907);
or U1881 (N_1881,In_573,In_1636);
nand U1882 (N_1882,N_699,In_1265);
or U1883 (N_1883,N_1700,N_1225);
nor U1884 (N_1884,In_1789,In_2110);
and U1885 (N_1885,N_613,In_2631);
nand U1886 (N_1886,In_1637,N_1412);
xor U1887 (N_1887,N_621,N_1618);
or U1888 (N_1888,N_945,N_1243);
and U1889 (N_1889,N_1457,N_1507);
nor U1890 (N_1890,N_1401,N_1540);
nand U1891 (N_1891,N_886,In_1107);
nor U1892 (N_1892,N_1180,In_1968);
nor U1893 (N_1893,N_1462,N_1301);
nand U1894 (N_1894,In_659,N_1087);
or U1895 (N_1895,N_875,N_1291);
nand U1896 (N_1896,N_1564,In_2810);
nand U1897 (N_1897,N_1775,N_1607);
or U1898 (N_1898,N_1000,In_2100);
nor U1899 (N_1899,N_158,N_766);
nor U1900 (N_1900,In_2993,In_2133);
nand U1901 (N_1901,In_1057,N_1399);
or U1902 (N_1902,N_1089,N_1319);
or U1903 (N_1903,In_1906,N_97);
xor U1904 (N_1904,In_2135,In_2745);
or U1905 (N_1905,N_1711,N_1779);
and U1906 (N_1906,In_77,N_704);
and U1907 (N_1907,N_1277,N_1463);
and U1908 (N_1908,N_479,N_1420);
nand U1909 (N_1909,N_467,N_1109);
and U1910 (N_1910,In_1441,N_1477);
nand U1911 (N_1911,N_1569,In_1318);
and U1912 (N_1912,N_1650,N_1764);
nand U1913 (N_1913,N_117,In_1782);
or U1914 (N_1914,N_1668,N_1495);
nand U1915 (N_1915,In_193,N_1360);
and U1916 (N_1916,N_1745,In_1753);
nor U1917 (N_1917,In_136,N_878);
nor U1918 (N_1918,N_1107,N_1380);
or U1919 (N_1919,N_1161,N_1490);
nand U1920 (N_1920,N_1436,N_1146);
nand U1921 (N_1921,N_1629,N_1655);
xor U1922 (N_1922,In_742,N_1092);
and U1923 (N_1923,N_181,In_957);
and U1924 (N_1924,N_1754,N_1729);
xor U1925 (N_1925,N_1798,N_666);
nor U1926 (N_1926,N_480,N_1492);
nand U1927 (N_1927,In_1593,In_1397);
nor U1928 (N_1928,In_918,N_1437);
or U1929 (N_1929,N_592,N_1488);
and U1930 (N_1930,N_1200,N_1718);
nor U1931 (N_1931,N_1487,In_1184);
and U1932 (N_1932,In_2253,In_880);
nor U1933 (N_1933,N_670,N_1641);
and U1934 (N_1934,N_197,N_1685);
xor U1935 (N_1935,N_1646,In_2452);
and U1936 (N_1936,N_427,N_610);
and U1937 (N_1937,N_1605,N_1732);
nand U1938 (N_1938,In_1683,In_2241);
or U1939 (N_1939,In_1613,N_840);
and U1940 (N_1940,N_542,In_883);
xnor U1941 (N_1941,N_304,N_1706);
nand U1942 (N_1942,In_1742,N_908);
nor U1943 (N_1943,N_1527,N_105);
xor U1944 (N_1944,N_1622,In_491);
or U1945 (N_1945,N_743,In_2227);
or U1946 (N_1946,In_2102,N_1076);
nor U1947 (N_1947,N_950,N_1148);
nor U1948 (N_1948,N_1642,In_748);
nand U1949 (N_1949,In_906,In_2071);
nand U1950 (N_1950,In_1632,N_1572);
and U1951 (N_1951,In_2427,In_2497);
nor U1952 (N_1952,N_1096,N_1160);
nand U1953 (N_1953,N_164,N_1654);
xnor U1954 (N_1954,In_1469,In_1763);
nor U1955 (N_1955,N_675,In_1933);
and U1956 (N_1956,N_384,N_1725);
nand U1957 (N_1957,N_1498,N_1769);
or U1958 (N_1958,In_1192,In_1751);
and U1959 (N_1959,N_1484,N_1634);
xnor U1960 (N_1960,In_2486,In_1479);
nor U1961 (N_1961,N_1144,In_249);
xor U1962 (N_1962,In_375,In_271);
and U1963 (N_1963,N_1370,In_2474);
nor U1964 (N_1964,N_1696,N_1427);
xnor U1965 (N_1965,N_1619,N_1636);
xor U1966 (N_1966,In_2012,N_1195);
or U1967 (N_1967,N_1064,In_1629);
nand U1968 (N_1968,In_1551,In_2101);
nand U1969 (N_1969,N_1584,N_544);
xor U1970 (N_1970,In_188,In_1390);
or U1971 (N_1971,N_1562,N_818);
nor U1972 (N_1972,N_1252,N_857);
nor U1973 (N_1973,N_1739,N_881);
xnor U1974 (N_1974,In_1537,In_961);
xor U1975 (N_1975,N_447,N_780);
or U1976 (N_1976,N_1466,In_472);
nand U1977 (N_1977,N_1652,In_568);
nand U1978 (N_1978,In_2955,N_368);
nor U1979 (N_1979,In_1431,N_1664);
nand U1980 (N_1980,In_1825,In_2972);
or U1981 (N_1981,In_2496,N_305);
and U1982 (N_1982,In_84,N_501);
nor U1983 (N_1983,N_1648,N_685);
xor U1984 (N_1984,N_247,In_802);
nand U1985 (N_1985,In_2375,N_1698);
nor U1986 (N_1986,N_921,In_2944);
nand U1987 (N_1987,N_999,N_1673);
xor U1988 (N_1988,N_755,N_401);
nand U1989 (N_1989,N_509,In_1409);
xor U1990 (N_1990,In_2807,N_1608);
and U1991 (N_1991,N_1489,N_1201);
nor U1992 (N_1992,N_48,In_2848);
xor U1993 (N_1993,N_1438,N_1387);
nand U1994 (N_1994,N_995,In_2572);
nor U1995 (N_1995,In_498,N_1331);
and U1996 (N_1996,In_2714,In_2082);
or U1997 (N_1997,N_1667,In_2235);
nor U1998 (N_1998,N_810,N_1139);
and U1999 (N_1999,N_1598,In_1085);
nor U2000 (N_2000,N_1417,N_1797);
nand U2001 (N_2001,N_1662,N_833);
nand U2002 (N_2002,In_1993,N_119);
and U2003 (N_2003,N_1481,N_493);
or U2004 (N_2004,In_1049,N_789);
and U2005 (N_2005,In_1712,N_1701);
nand U2006 (N_2006,N_1600,N_410);
nor U2007 (N_2007,N_1032,N_1836);
xor U2008 (N_2008,N_1479,N_1885);
or U2009 (N_2009,N_1974,N_1450);
and U2010 (N_2010,N_1210,N_1772);
nor U2011 (N_2011,N_1354,In_1719);
and U2012 (N_2012,N_1515,N_1034);
nand U2013 (N_2013,N_1884,N_1969);
xor U2014 (N_2014,In_1972,N_1966);
or U2015 (N_2015,N_1721,N_862);
xor U2016 (N_2016,N_211,N_1867);
nor U2017 (N_2017,N_1902,N_1921);
and U2018 (N_2018,N_1657,N_1848);
nor U2019 (N_2019,N_1235,N_1555);
xnor U2020 (N_2020,In_1868,N_1971);
or U2021 (N_2021,N_1272,N_684);
xor U2022 (N_2022,In_2129,In_2712);
or U2023 (N_2023,In_1681,N_1714);
or U2024 (N_2024,In_283,N_1471);
nor U2025 (N_2025,In_2424,N_487);
xor U2026 (N_2026,N_1072,N_1386);
nor U2027 (N_2027,N_1957,In_2130);
nand U2028 (N_2028,N_1773,N_1193);
and U2029 (N_2029,N_697,N_1900);
xor U2030 (N_2030,N_1348,N_1928);
nor U2031 (N_2031,N_1491,N_563);
nand U2032 (N_2032,N_1894,N_1861);
and U2033 (N_2033,N_1687,N_1851);
or U2034 (N_2034,N_1941,In_257);
nand U2035 (N_2035,In_1044,N_1812);
or U2036 (N_2036,N_1810,N_1880);
and U2037 (N_2037,In_1508,N_703);
nand U2038 (N_2038,N_1683,N_574);
nor U2039 (N_2039,N_1502,N_1647);
nand U2040 (N_2040,N_1929,In_1529);
xnor U2041 (N_2041,In_2221,In_897);
nor U2042 (N_2042,N_1241,In_952);
and U2043 (N_2043,In_2842,In_26);
xor U2044 (N_2044,In_1572,N_1433);
or U2045 (N_2045,N_1707,N_1098);
and U2046 (N_2046,N_135,N_1984);
xor U2047 (N_2047,In_1314,N_1728);
or U2048 (N_2048,N_830,N_1825);
nand U2049 (N_2049,In_820,In_1450);
xor U2050 (N_2050,In_2582,N_1338);
xor U2051 (N_2051,N_1895,N_1933);
nor U2052 (N_2052,N_1767,N_1326);
xnor U2053 (N_2053,N_433,N_669);
and U2054 (N_2054,In_1888,In_1595);
and U2055 (N_2055,In_2793,N_1831);
xor U2056 (N_2056,N_1837,In_1055);
or U2057 (N_2057,In_2045,N_461);
and U2058 (N_2058,N_612,N_1890);
nand U2059 (N_2059,N_1547,In_1240);
xnor U2060 (N_2060,N_1056,N_445);
xnor U2061 (N_2061,N_715,N_1153);
xnor U2062 (N_2062,In_1558,In_1215);
or U2063 (N_2063,N_1426,In_239);
nor U2064 (N_2064,In_1982,N_1850);
nor U2065 (N_2065,N_551,N_1839);
nor U2066 (N_2066,In_641,N_1955);
nor U2067 (N_2067,In_2742,N_1715);
xor U2068 (N_2068,In_75,N_1084);
nor U2069 (N_2069,N_1011,N_1186);
and U2070 (N_2070,In_1807,N_1920);
and U2071 (N_2071,N_1835,In_21);
xnor U2072 (N_2072,In_369,In_376);
nor U2073 (N_2073,N_1991,N_1758);
and U2074 (N_2074,N_1994,N_1303);
or U2075 (N_2075,N_1959,N_1684);
nand U2076 (N_2076,N_1626,N_1870);
nor U2077 (N_2077,N_1345,In_1076);
or U2078 (N_2078,N_1856,N_1582);
xor U2079 (N_2079,In_2108,N_1913);
xor U2080 (N_2080,N_1793,N_1222);
nor U2081 (N_2081,N_33,N_1203);
nand U2082 (N_2082,N_571,N_1803);
nand U2083 (N_2083,In_1570,N_1520);
or U2084 (N_2084,N_1849,In_1517);
and U2085 (N_2085,N_1864,N_1432);
or U2086 (N_2086,N_880,N_1236);
or U2087 (N_2087,N_1866,In_1069);
and U2088 (N_2088,In_1412,N_1824);
and U2089 (N_2089,In_326,N_1838);
nor U2090 (N_2090,N_1693,N_1973);
and U2091 (N_2091,N_1300,In_622);
xnor U2092 (N_2092,N_430,In_178);
nor U2093 (N_2093,N_1213,N_1749);
or U2094 (N_2094,In_298,N_1736);
xor U2095 (N_2095,In_544,N_306);
nand U2096 (N_2096,In_1910,N_1313);
xor U2097 (N_2097,N_1329,N_1396);
nor U2098 (N_2098,In_1804,N_1914);
nor U2099 (N_2099,N_1862,N_292);
nor U2100 (N_2100,N_1409,N_1901);
and U2101 (N_2101,N_79,N_1742);
nor U2102 (N_2102,N_1809,N_1818);
and U2103 (N_2103,N_391,N_1079);
nor U2104 (N_2104,N_738,N_1513);
or U2105 (N_2105,N_1777,N_140);
nor U2106 (N_2106,N_1518,N_32);
and U2107 (N_2107,N_1830,N_1602);
nand U2108 (N_2108,N_1459,N_1653);
and U2109 (N_2109,N_1162,N_1865);
and U2110 (N_2110,N_1546,In_1204);
or U2111 (N_2111,N_768,N_1670);
and U2112 (N_2112,N_409,In_2794);
nand U2113 (N_2113,In_998,In_2922);
xnor U2114 (N_2114,N_1150,In_2124);
nor U2115 (N_2115,N_1931,In_1903);
nand U2116 (N_2116,In_1093,N_1336);
or U2117 (N_2117,N_520,N_718);
nand U2118 (N_2118,N_645,N_1926);
or U2119 (N_2119,In_1584,N_568);
xor U2120 (N_2120,N_1627,N_1786);
nor U2121 (N_2121,In_2397,N_21);
and U2122 (N_2122,In_173,In_2301);
nor U2123 (N_2123,In_1305,N_1844);
xor U2124 (N_2124,In_1378,In_1163);
xor U2125 (N_2125,N_1452,N_556);
nand U2126 (N_2126,N_1932,N_1494);
nor U2127 (N_2127,In_2188,N_1774);
nand U2128 (N_2128,N_1132,In_1784);
or U2129 (N_2129,N_251,In_2147);
xnor U2130 (N_2130,N_1368,N_1429);
nor U2131 (N_2131,N_1568,N_469);
nor U2132 (N_2132,N_1869,N_1215);
or U2133 (N_2133,N_238,In_2937);
or U2134 (N_2134,N_1333,N_1234);
or U2135 (N_2135,N_1343,N_892);
and U2136 (N_2136,N_1802,In_1147);
nor U2137 (N_2137,N_1904,N_1620);
or U2138 (N_2138,N_100,N_1820);
or U2139 (N_2139,In_2482,N_458);
xnor U2140 (N_2140,In_927,N_814);
xnor U2141 (N_2141,N_1690,N_1635);
nand U2142 (N_2142,N_1800,In_539);
nand U2143 (N_2143,In_1447,In_1758);
and U2144 (N_2144,In_615,N_259);
and U2145 (N_2145,In_2020,In_1839);
nor U2146 (N_2146,In_2589,N_1112);
nand U2147 (N_2147,N_1389,N_1887);
nand U2148 (N_2148,N_1804,N_516);
or U2149 (N_2149,N_1746,In_1098);
nor U2150 (N_2150,N_1782,N_1217);
nor U2151 (N_2151,N_1886,In_1932);
or U2152 (N_2152,In_2044,N_1723);
or U2153 (N_2153,N_1659,In_686);
nor U2154 (N_2154,N_1958,In_349);
or U2155 (N_2155,N_1585,In_1983);
or U2156 (N_2156,In_2084,In_2907);
or U2157 (N_2157,N_655,N_1713);
nand U2158 (N_2158,N_1731,N_808);
xor U2159 (N_2159,In_2727,N_1854);
nor U2160 (N_2160,N_1983,In_2122);
or U2161 (N_2161,N_88,In_1324);
nor U2162 (N_2162,N_1776,N_1624);
nand U2163 (N_2163,N_1934,N_1242);
or U2164 (N_2164,N_1799,N_1230);
and U2165 (N_2165,N_1347,N_321);
and U2166 (N_2166,N_474,N_1460);
or U2167 (N_2167,N_1001,N_1359);
xor U2168 (N_2168,In_424,In_747);
nand U2169 (N_2169,In_2884,N_114);
nor U2170 (N_2170,N_1672,In_2200);
xor U2171 (N_2171,In_1962,N_760);
nand U2172 (N_2172,N_1255,In_1373);
and U2173 (N_2173,N_1738,N_1430);
nand U2174 (N_2174,N_1724,N_1781);
nor U2175 (N_2175,N_1469,N_1761);
nor U2176 (N_2176,N_1044,In_2723);
nor U2177 (N_2177,N_1036,N_602);
xor U2178 (N_2178,N_1633,N_1843);
xnor U2179 (N_2179,N_1314,N_299);
nor U2180 (N_2180,N_1258,In_1921);
nor U2181 (N_2181,N_1379,N_982);
nand U2182 (N_2182,N_1404,N_1192);
nand U2183 (N_2183,N_1537,In_1935);
nand U2184 (N_2184,N_650,In_2359);
nand U2185 (N_2185,N_1091,In_1865);
nor U2186 (N_2186,N_1615,N_1699);
or U2187 (N_2187,In_2887,In_1446);
nand U2188 (N_2188,In_1308,In_258);
or U2189 (N_2189,N_1307,N_797);
nand U2190 (N_2190,N_1406,N_1980);
xnor U2191 (N_2191,N_1925,In_1620);
or U2192 (N_2192,N_1599,N_1733);
or U2193 (N_2193,N_1041,N_1937);
and U2194 (N_2194,In_599,N_614);
nor U2195 (N_2195,In_1499,N_1719);
nor U2196 (N_2196,N_1968,N_1744);
xor U2197 (N_2197,In_1335,N_839);
nand U2198 (N_2198,N_1770,N_1439);
nand U2199 (N_2199,N_560,N_1623);
or U2200 (N_2200,N_1198,In_1809);
nor U2201 (N_2201,N_2026,N_1610);
nor U2202 (N_2202,N_2154,N_1765);
xor U2203 (N_2203,N_1743,N_1875);
nand U2204 (N_2204,N_2123,In_1528);
xnor U2205 (N_2205,N_721,N_2183);
nand U2206 (N_2206,N_2197,N_2182);
xor U2207 (N_2207,N_1373,N_1611);
or U2208 (N_2208,N_1917,N_642);
xnor U2209 (N_2209,N_1578,N_2180);
and U2210 (N_2210,N_2133,N_242);
nand U2211 (N_2211,N_1945,N_1312);
and U2212 (N_2212,N_2087,N_1660);
nor U2213 (N_2213,N_1197,N_2041);
nor U2214 (N_2214,N_1510,N_803);
nor U2215 (N_2215,In_501,N_1989);
nor U2216 (N_2216,In_2353,In_1303);
or U2217 (N_2217,N_1081,In_2251);
or U2218 (N_2218,N_1919,N_973);
xor U2219 (N_2219,N_1444,N_1874);
or U2220 (N_2220,N_1947,N_1617);
or U2221 (N_2221,N_1567,N_1020);
and U2222 (N_2222,N_1747,N_2080);
xor U2223 (N_2223,N_1614,N_1924);
nor U2224 (N_2224,N_2103,N_1529);
nor U2225 (N_2225,N_2090,N_1315);
and U2226 (N_2226,N_1740,N_2010);
nor U2227 (N_2227,N_1995,N_1915);
nand U2228 (N_2228,N_2131,In_692);
nand U2229 (N_2229,N_2153,N_1695);
nor U2230 (N_2230,N_967,N_1816);
or U2231 (N_2231,N_1908,N_2078);
nand U2232 (N_2232,N_2024,N_1163);
and U2233 (N_2233,N_1117,N_2007);
nand U2234 (N_2234,In_1311,N_1088);
nor U2235 (N_2235,N_1882,In_171);
xnor U2236 (N_2236,N_2091,N_702);
and U2237 (N_2237,N_2185,N_1952);
nand U2238 (N_2238,N_1467,N_2119);
nor U2239 (N_2239,N_1458,In_2863);
nand U2240 (N_2240,N_1819,In_1038);
or U2241 (N_2241,N_1411,N_913);
xnor U2242 (N_2242,N_2139,N_2069);
or U2243 (N_2243,N_1857,N_2115);
nand U2244 (N_2244,In_431,In_1462);
or U2245 (N_2245,N_1366,N_2037);
or U2246 (N_2246,N_1661,N_1298);
xor U2247 (N_2247,N_2013,N_2042);
xor U2248 (N_2248,N_2167,N_1905);
or U2249 (N_2249,N_2142,In_1153);
or U2250 (N_2250,N_532,In_2625);
and U2251 (N_2251,N_1671,N_2129);
nand U2252 (N_2252,N_2111,N_2021);
nand U2253 (N_2253,N_552,N_1612);
nand U2254 (N_2254,N_2112,In_2824);
nand U2255 (N_2255,N_1964,N_796);
and U2256 (N_2256,In_2233,N_2181);
and U2257 (N_2257,N_2040,N_1944);
and U2258 (N_2258,N_2020,N_147);
xor U2259 (N_2259,N_2156,N_1133);
or U2260 (N_2260,N_2166,In_2804);
nor U2261 (N_2261,N_2178,N_984);
xnor U2262 (N_2262,In_1297,N_912);
and U2263 (N_2263,N_1988,N_2082);
and U2264 (N_2264,In_346,In_1288);
or U2265 (N_2265,N_2088,N_2061);
and U2266 (N_2266,In_1862,N_838);
or U2267 (N_2267,In_2283,N_2155);
nor U2268 (N_2268,N_677,N_872);
and U2269 (N_2269,N_2172,N_1565);
and U2270 (N_2270,N_413,N_1768);
or U2271 (N_2271,In_2525,N_1978);
nand U2272 (N_2272,N_1829,N_2023);
nand U2273 (N_2273,In_640,N_381);
nor U2274 (N_2274,N_1425,N_1794);
or U2275 (N_2275,N_1332,In_1543);
nand U2276 (N_2276,N_1454,N_1666);
nand U2277 (N_2277,N_1834,N_1805);
xnor U2278 (N_2278,N_1253,In_164);
nor U2279 (N_2279,N_1697,N_1054);
xor U2280 (N_2280,N_2086,In_2275);
nor U2281 (N_2281,N_1923,In_954);
nand U2282 (N_2282,N_1760,N_2191);
xnor U2283 (N_2283,In_944,N_2177);
or U2284 (N_2284,N_2146,In_2527);
or U2285 (N_2285,N_1448,N_1956);
and U2286 (N_2286,In_189,In_2637);
and U2287 (N_2287,In_540,N_1676);
nand U2288 (N_2288,N_1936,N_2004);
and U2289 (N_2289,N_2108,N_1705);
xor U2290 (N_2290,N_434,In_2610);
and U2291 (N_2291,N_1759,In_759);
nand U2292 (N_2292,In_1277,N_955);
nor U2293 (N_2293,N_1868,N_2187);
xnor U2294 (N_2294,N_1596,N_2147);
nor U2295 (N_2295,N_51,In_2961);
nand U2296 (N_2296,N_2150,N_656);
nand U2297 (N_2297,N_643,N_2074);
xor U2298 (N_2298,N_1356,N_2015);
or U2299 (N_2299,N_1833,N_676);
xor U2300 (N_2300,N_2107,In_2015);
or U2301 (N_2301,N_2072,N_2051);
and U2302 (N_2302,In_785,In_1241);
xor U2303 (N_2303,N_850,N_1588);
xnor U2304 (N_2304,N_923,N_2161);
and U2305 (N_2305,In_2134,N_1613);
xor U2306 (N_2306,N_1827,In_465);
and U2307 (N_2307,N_1828,N_2059);
or U2308 (N_2308,In_1757,N_1708);
and U2309 (N_2309,N_2100,In_597);
nand U2310 (N_2310,N_1970,N_2118);
nor U2311 (N_2311,In_2338,N_1516);
nand U2312 (N_2312,N_1859,N_1883);
or U2313 (N_2313,N_2076,N_1267);
or U2314 (N_2314,In_82,N_1544);
nor U2315 (N_2315,N_2134,In_299);
nor U2316 (N_2316,N_2136,N_1640);
nor U2317 (N_2317,N_2175,In_1363);
xnor U2318 (N_2318,In_1073,N_2011);
nand U2319 (N_2319,In_971,N_2012);
nand U2320 (N_2320,N_1860,N_1903);
nand U2321 (N_2321,N_2044,N_1811);
nor U2322 (N_2322,N_1855,N_177);
nand U2323 (N_2323,N_1553,N_1586);
or U2324 (N_2324,N_1591,N_1716);
and U2325 (N_2325,N_1339,N_81);
nor U2326 (N_2326,In_500,N_1609);
nand U2327 (N_2327,In_868,N_1511);
xnor U2328 (N_2328,N_1787,N_1982);
nor U2329 (N_2329,N_1681,N_1939);
nand U2330 (N_2330,N_62,N_1138);
nor U2331 (N_2331,N_1080,In_2432);
nand U2332 (N_2332,In_2348,In_466);
nand U2333 (N_2333,N_1245,N_2179);
and U2334 (N_2334,N_471,N_864);
nor U2335 (N_2335,N_1889,N_2117);
or U2336 (N_2336,N_1840,In_8);
and U2337 (N_2337,In_2545,N_2027);
nand U2338 (N_2338,N_2097,In_1687);
nand U2339 (N_2339,N_1226,N_1296);
nor U2340 (N_2340,N_1942,In_2974);
xor U2341 (N_2341,N_651,N_1702);
and U2342 (N_2342,N_1239,N_1435);
and U2343 (N_2343,N_1378,In_391);
xor U2344 (N_2344,N_2034,N_1692);
or U2345 (N_2345,In_976,N_2164);
nor U2346 (N_2346,N_2073,N_1806);
xor U2347 (N_2347,N_1948,In_2169);
or U2348 (N_2348,N_2031,N_2033);
and U2349 (N_2349,N_1663,N_1543);
or U2350 (N_2350,N_1376,In_1139);
xor U2351 (N_2351,N_1898,N_1938);
or U2352 (N_2352,N_1722,N_1877);
nand U2353 (N_2353,In_273,N_2127);
nand U2354 (N_2354,N_2075,N_1815);
nand U2355 (N_2355,N_1710,N_1845);
nor U2356 (N_2356,In_1050,N_2009);
or U2357 (N_2357,N_1976,N_707);
nor U2358 (N_2358,N_1678,In_2125);
nor U2359 (N_2359,N_1753,In_1783);
or U2360 (N_2360,N_2138,In_2381);
nor U2361 (N_2361,N_2125,N_1935);
nor U2362 (N_2362,N_1168,N_1278);
nand U2363 (N_2363,N_2054,In_1819);
xnor U2364 (N_2364,N_1271,N_1841);
or U2365 (N_2365,N_855,N_437);
xnor U2366 (N_2366,In_1090,N_1766);
and U2367 (N_2367,N_1813,N_2092);
xnor U2368 (N_2368,N_783,N_1778);
nand U2369 (N_2369,N_820,N_2128);
nor U2370 (N_2370,N_344,N_2083);
nor U2371 (N_2371,N_45,N_1290);
and U2372 (N_2372,In_1749,In_2352);
nand U2373 (N_2373,N_1545,N_2018);
and U2374 (N_2374,N_2110,N_1785);
and U2375 (N_2375,N_2122,In_1690);
or U2376 (N_2376,N_1990,N_1136);
nand U2377 (N_2377,In_2419,In_2576);
nor U2378 (N_2378,N_347,N_1549);
and U2379 (N_2379,N_1999,N_1677);
nor U2380 (N_2380,N_1174,N_1440);
and U2381 (N_2381,N_1318,N_2089);
nand U2382 (N_2382,N_1576,N_1953);
and U2383 (N_2383,N_1418,In_576);
xor U2384 (N_2384,N_2014,N_1346);
nor U2385 (N_2385,N_369,N_2099);
xnor U2386 (N_2386,N_2163,N_1909);
nor U2387 (N_2387,N_1101,N_1400);
nand U2388 (N_2388,In_2054,In_1368);
and U2389 (N_2389,N_1998,N_1912);
or U2390 (N_2390,N_1475,N_899);
nand U2391 (N_2391,N_1014,N_1888);
and U2392 (N_2392,N_962,N_1846);
and U2393 (N_2393,N_2198,N_1204);
and U2394 (N_2394,N_1858,N_2169);
nand U2395 (N_2395,N_2116,In_1726);
nand U2396 (N_2396,N_95,N_2049);
nand U2397 (N_2397,N_1616,N_2158);
nor U2398 (N_2398,In_935,N_2000);
or U2399 (N_2399,N_1756,N_1443);
and U2400 (N_2400,N_2106,N_2371);
xor U2401 (N_2401,N_2077,N_2019);
xor U2402 (N_2402,N_2312,N_1587);
or U2403 (N_2403,N_1017,N_2200);
or U2404 (N_2404,N_2144,N_2306);
xor U2405 (N_2405,N_1789,In_2248);
or U2406 (N_2406,N_2228,N_1577);
xnor U2407 (N_2407,N_1896,N_2269);
or U2408 (N_2408,N_884,In_2593);
or U2409 (N_2409,N_2293,N_630);
nor U2410 (N_2410,N_2350,N_600);
xnor U2411 (N_2411,N_1972,N_787);
nand U2412 (N_2412,N_1504,In_464);
xnor U2413 (N_2413,N_1712,N_883);
xnor U2414 (N_2414,N_874,N_2272);
nand U2415 (N_2415,N_2124,In_1467);
nand U2416 (N_2416,N_2190,N_2067);
nand U2417 (N_2417,N_2359,N_2234);
or U2418 (N_2418,N_2196,N_550);
nor U2419 (N_2419,N_2376,N_2380);
xnor U2420 (N_2420,N_1893,N_734);
xnor U2421 (N_2421,N_1892,N_2113);
xnor U2422 (N_2422,N_2102,N_2384);
xor U2423 (N_2423,In_90,N_2159);
nor U2424 (N_2424,N_1946,N_1675);
xnor U2425 (N_2425,N_1445,N_1028);
xnor U2426 (N_2426,N_1658,N_1645);
and U2427 (N_2427,N_1244,N_1393);
and U2428 (N_2428,In_872,N_1232);
nand U2429 (N_2429,N_1910,N_2109);
and U2430 (N_2430,N_2296,N_2145);
nor U2431 (N_2431,N_1879,N_2316);
nand U2432 (N_2432,N_2220,N_2278);
and U2433 (N_2433,N_791,N_2060);
nor U2434 (N_2434,N_1873,N_2275);
and U2435 (N_2435,In_40,N_2056);
or U2436 (N_2436,N_2327,N_2259);
nand U2437 (N_2437,N_2357,In_856);
nor U2438 (N_2438,N_2243,N_2311);
or U2439 (N_2439,N_196,N_1807);
nand U2440 (N_2440,N_1505,N_1583);
xnor U2441 (N_2441,In_1013,N_2137);
and U2442 (N_2442,N_2210,N_2365);
nor U2443 (N_2443,N_2320,N_2317);
nor U2444 (N_2444,N_1496,N_1906);
and U2445 (N_2445,N_1248,N_2120);
and U2446 (N_2446,N_1987,In_749);
nand U2447 (N_2447,N_2141,N_2235);
or U2448 (N_2448,N_1878,In_1602);
nand U2449 (N_2449,N_1428,N_1669);
nand U2450 (N_2450,N_2271,N_1294);
and U2451 (N_2451,N_1788,N_2345);
and U2452 (N_2452,N_1068,N_1967);
nand U2453 (N_2453,N_2186,N_2353);
and U2454 (N_2454,In_477,N_2208);
or U2455 (N_2455,N_2393,N_2039);
nor U2456 (N_2456,N_2173,N_2291);
or U2457 (N_2457,N_2399,N_1508);
or U2458 (N_2458,N_1171,In_1349);
nand U2459 (N_2459,N_2368,N_2394);
nand U2460 (N_2460,N_2292,N_1826);
and U2461 (N_2461,N_2194,N_2389);
and U2462 (N_2462,N_2098,In_19);
or U2463 (N_2463,N_2094,N_1821);
nor U2464 (N_2464,N_2036,N_2195);
nor U2465 (N_2465,N_2323,In_2468);
nor U2466 (N_2466,N_2217,N_2025);
and U2467 (N_2467,In_2448,N_2298);
and U2468 (N_2468,N_261,N_1899);
nor U2469 (N_2469,N_2249,N_1847);
nand U2470 (N_2470,N_2267,N_2386);
and U2471 (N_2471,N_2062,In_2193);
xor U2472 (N_2472,N_1007,N_2328);
or U2473 (N_2473,N_1554,N_2366);
nand U2474 (N_2474,N_1817,N_696);
nand U2475 (N_2475,N_2288,N_942);
xor U2476 (N_2476,N_1951,N_1963);
xor U2477 (N_2477,N_1674,N_1423);
or U2478 (N_2478,N_2050,N_2344);
and U2479 (N_2479,N_809,N_1961);
or U2480 (N_2480,N_2207,N_490);
nor U2481 (N_2481,N_2257,N_2071);
nor U2482 (N_2482,N_2170,N_1965);
xnor U2483 (N_2483,N_1823,In_2198);
and U2484 (N_2484,N_2211,N_2214);
xnor U2485 (N_2485,N_319,N_2268);
and U2486 (N_2486,N_1320,In_1523);
nor U2487 (N_2487,In_2558,N_2280);
xor U2488 (N_2488,N_2276,N_2192);
nor U2489 (N_2489,N_2274,N_2290);
or U2490 (N_2490,N_1327,N_2219);
nand U2491 (N_2491,N_2263,N_1907);
and U2492 (N_2492,N_2283,In_1029);
xor U2493 (N_2493,In_1039,N_1306);
or U2494 (N_2494,In_1672,In_473);
nand U2495 (N_2495,N_2165,N_1209);
nand U2496 (N_2496,In_955,N_2277);
nor U2497 (N_2497,N_1872,N_310);
and U2498 (N_2498,N_2230,N_701);
xnor U2499 (N_2499,N_2202,N_1750);
nand U2500 (N_2500,N_2032,N_1727);
xor U2501 (N_2501,In_2639,N_1717);
or U2502 (N_2502,In_768,N_2201);
nor U2503 (N_2503,N_2300,N_234);
and U2504 (N_2504,N_2001,N_2332);
nand U2505 (N_2505,N_1580,N_2356);
or U2506 (N_2506,N_2279,N_1410);
nand U2507 (N_2507,N_2176,N_2239);
xnor U2508 (N_2508,N_2143,In_1836);
or U2509 (N_2509,N_42,N_2184);
and U2510 (N_2510,N_2273,N_1949);
nor U2511 (N_2511,N_179,N_2002);
or U2512 (N_2512,In_1645,N_2221);
or U2513 (N_2513,N_2253,N_1656);
and U2514 (N_2514,N_534,N_2130);
nand U2515 (N_2515,N_2043,N_2324);
xnor U2516 (N_2516,N_2387,N_1852);
nor U2517 (N_2517,N_1205,N_2397);
nor U2518 (N_2518,N_2065,N_1208);
nand U2519 (N_2519,N_1031,N_1625);
xor U2520 (N_2520,N_2085,N_2354);
or U2521 (N_2521,In_2858,N_1808);
nand U2522 (N_2522,N_2373,N_2382);
xor U2523 (N_2523,N_1814,In_1244);
or U2524 (N_2524,N_1059,In_2697);
or U2525 (N_2525,N_2045,N_1407);
and U2526 (N_2526,N_2361,N_2189);
xnor U2527 (N_2527,N_1780,N_2383);
xnor U2528 (N_2528,N_2337,N_1881);
and U2529 (N_2529,N_2379,N_1566);
or U2530 (N_2530,N_634,N_218);
and U2531 (N_2531,N_2321,In_912);
xnor U2532 (N_2532,N_120,In_212);
and U2533 (N_2533,N_2369,N_298);
nor U2534 (N_2534,In_2266,N_1470);
nand U2535 (N_2535,N_2364,N_2282);
or U2536 (N_2536,In_2890,N_2008);
and U2537 (N_2537,N_2302,N_2204);
nand U2538 (N_2538,N_2381,N_1863);
or U2539 (N_2539,N_2035,N_2151);
and U2540 (N_2540,N_2017,N_2331);
xnor U2541 (N_2541,In_2055,N_2081);
nor U2542 (N_2542,N_1954,N_2287);
nand U2543 (N_2543,N_2149,N_366);
or U2544 (N_2544,N_1911,N_1792);
and U2545 (N_2545,N_1372,N_661);
and U2546 (N_2546,N_2224,N_2363);
nand U2547 (N_2547,N_752,N_115);
nor U2548 (N_2548,N_2377,N_2022);
nand U2549 (N_2549,In_789,In_1180);
or U2550 (N_2550,N_1550,N_1526);
nand U2551 (N_2551,N_207,N_2258);
and U2552 (N_2552,N_747,N_2326);
xor U2553 (N_2553,N_2398,N_2297);
and U2554 (N_2554,N_2226,N_1783);
nor U2555 (N_2555,N_2048,N_2360);
nor U2556 (N_2556,N_1416,N_1897);
or U2557 (N_2557,N_2242,N_2203);
and U2558 (N_2558,N_1542,N_1981);
nor U2559 (N_2559,N_1975,In_1979);
xor U2560 (N_2560,N_2352,N_1464);
and U2561 (N_2561,In_1541,N_2030);
or U2562 (N_2562,N_2066,N_1822);
xnor U2563 (N_2563,N_2333,N_2104);
and U2564 (N_2564,N_2168,N_2355);
and U2565 (N_2565,N_2084,N_2052);
or U2566 (N_2566,N_1891,N_2295);
xnor U2567 (N_2567,N_2310,In_1530);
and U2568 (N_2568,N_1552,In_2827);
or U2569 (N_2569,In_2878,N_2251);
and U2570 (N_2570,N_1182,N_2340);
xnor U2571 (N_2571,N_2329,In_388);
nor U2572 (N_2572,N_852,N_2237);
xnor U2573 (N_2573,N_1997,In_926);
nand U2574 (N_2574,N_2193,N_1067);
xnor U2575 (N_2575,N_1853,N_1801);
or U2576 (N_2576,N_2132,N_1960);
and U2577 (N_2577,N_2375,N_2248);
nor U2578 (N_2578,N_2388,N_2245);
and U2579 (N_2579,N_2299,N_2307);
xnor U2580 (N_2580,N_351,N_2057);
nor U2581 (N_2581,N_1220,In_2964);
and U2582 (N_2582,N_1751,N_2392);
nor U2583 (N_2583,N_2265,N_2016);
nand U2584 (N_2584,N_2256,N_1465);
xor U2585 (N_2585,N_1694,N_1070);
and U2586 (N_2586,In_1267,N_2247);
and U2587 (N_2587,N_2308,In_2948);
nor U2588 (N_2588,In_469,N_1916);
nand U2589 (N_2589,N_2351,N_2152);
and U2590 (N_2590,N_2334,N_909);
nor U2591 (N_2591,N_2047,N_1962);
or U2592 (N_2592,N_1639,N_2395);
and U2593 (N_2593,N_2294,In_2051);
and U2594 (N_2594,N_2261,N_2114);
nor U2595 (N_2595,N_1771,N_1986);
nor U2596 (N_2596,N_2241,N_2238);
and U2597 (N_2597,In_1030,In_1438);
nand U2598 (N_2598,N_1992,N_993);
and U2599 (N_2599,N_1950,N_2157);
or U2600 (N_2600,N_2346,N_2512);
xnor U2601 (N_2601,N_2439,N_2412);
nor U2602 (N_2602,N_2421,N_2424);
or U2603 (N_2603,N_2566,N_706);
or U2604 (N_2604,N_2582,N_2550);
nor U2605 (N_2605,N_1876,N_2583);
xor U2606 (N_2606,N_2490,N_2322);
nand U2607 (N_2607,N_2416,N_1977);
nor U2608 (N_2608,N_1979,N_2486);
nand U2609 (N_2609,N_2589,N_2289);
or U2610 (N_2610,In_635,In_2417);
and U2611 (N_2611,N_2544,N_2469);
or U2612 (N_2612,In_2703,N_2485);
nand U2613 (N_2613,N_2461,N_2252);
nor U2614 (N_2614,N_2063,N_1100);
nand U2615 (N_2615,N_2451,N_1099);
nand U2616 (N_2616,N_2571,N_1058);
nand U2617 (N_2617,N_2404,N_2494);
nor U2618 (N_2618,N_2222,N_2452);
nand U2619 (N_2619,N_553,N_2575);
and U2620 (N_2620,In_1129,N_2538);
and U2621 (N_2621,N_2309,N_1930);
and U2622 (N_2622,N_2435,N_1737);
or U2623 (N_2623,N_2205,N_2489);
xor U2624 (N_2624,In_2,N_2422);
nand U2625 (N_2625,N_951,N_2338);
nand U2626 (N_2626,N_1993,N_2460);
nand U2627 (N_2627,N_2513,In_355);
nor U2628 (N_2628,N_2570,N_2519);
nand U2629 (N_2629,N_2445,N_2592);
xor U2630 (N_2630,N_1482,N_2335);
xor U2631 (N_2631,In_2879,N_2254);
nand U2632 (N_2632,In_266,N_2005);
nand U2633 (N_2633,N_2528,N_2095);
nor U2634 (N_2634,N_2407,N_2530);
or U2635 (N_2635,N_2484,N_1832);
xor U2636 (N_2636,In_186,N_1922);
nor U2637 (N_2637,N_2101,N_2285);
xor U2638 (N_2638,N_2171,N_844);
and U2639 (N_2639,N_2581,N_2413);
nor U2640 (N_2640,N_1532,N_2236);
nand U2641 (N_2641,N_2053,N_2505);
xnor U2642 (N_2642,N_2483,N_2558);
or U2643 (N_2643,N_2590,N_1637);
nor U2644 (N_2644,N_2464,N_2511);
nor U2645 (N_2645,N_2556,In_2007);
nand U2646 (N_2646,In_1598,N_2555);
xnor U2647 (N_2647,N_2467,N_2456);
and U2648 (N_2648,N_1601,N_2546);
or U2649 (N_2649,N_2465,N_2500);
and U2650 (N_2650,N_2330,N_2336);
and U2651 (N_2651,N_2508,N_2524);
nor U2652 (N_2652,In_2791,N_2430);
and U2653 (N_2653,N_2318,N_2499);
nor U2654 (N_2654,N_2419,N_2341);
or U2655 (N_2655,N_1501,N_524);
nand U2656 (N_2656,N_2437,N_2449);
nand U2657 (N_2657,N_1996,N_2438);
or U2658 (N_2658,N_2411,N_1940);
nand U2659 (N_2659,N_2199,N_2586);
or U2660 (N_2660,N_2121,In_1291);
nor U2661 (N_2661,N_2561,N_2301);
and U2662 (N_2662,N_2391,In_2453);
and U2663 (N_2663,In_569,N_2502);
nor U2664 (N_2664,N_2487,N_2434);
and U2665 (N_2665,N_2443,N_2547);
nor U2666 (N_2666,N_547,N_1474);
nand U2667 (N_2667,N_2343,N_2567);
xor U2668 (N_2668,N_1606,N_2218);
nor U2669 (N_2669,N_719,N_2028);
or U2670 (N_2670,N_2507,N_2266);
or U2671 (N_2671,In_2991,N_2410);
or U2672 (N_2672,N_2216,N_2573);
or U2673 (N_2673,N_2223,N_2501);
and U2674 (N_2674,N_2577,N_2594);
and U2675 (N_2675,N_2560,N_2517);
nand U2676 (N_2676,N_2540,N_2281);
and U2677 (N_2677,In_1061,N_903);
nand U2678 (N_2678,In_2945,N_2455);
or U2679 (N_2679,In_1642,N_2255);
xor U2680 (N_2680,N_2470,N_2339);
xnor U2681 (N_2681,N_920,N_2526);
and U2682 (N_2682,N_2212,N_795);
and U2683 (N_2683,N_2420,N_2415);
xor U2684 (N_2684,N_2140,N_2244);
nand U2685 (N_2685,N_2313,N_2529);
nand U2686 (N_2686,N_2262,N_2584);
xnor U2687 (N_2687,N_2559,N_1943);
or U2688 (N_2688,N_2006,N_2518);
or U2689 (N_2689,N_2429,N_2493);
nand U2690 (N_2690,N_1643,N_2385);
xor U2691 (N_2691,N_2478,N_2551);
nand U2692 (N_2692,N_2545,N_2510);
and U2693 (N_2693,N_2442,N_2003);
or U2694 (N_2694,N_2474,N_2491);
nor U2695 (N_2695,N_2246,N_2374);
and U2696 (N_2696,N_2396,N_2233);
and U2697 (N_2697,N_2093,N_1541);
nand U2698 (N_2698,N_2453,N_2319);
xor U2699 (N_2699,N_1573,In_726);
and U2700 (N_2700,N_1594,N_2516);
xnor U2701 (N_2701,N_2367,N_2563);
nand U2702 (N_2702,N_2286,N_2126);
nand U2703 (N_2703,N_2347,N_2553);
and U2704 (N_2704,N_1446,N_2549);
or U2705 (N_2705,N_2250,N_2471);
xor U2706 (N_2706,N_2096,N_2105);
or U2707 (N_2707,N_2174,N_2496);
and U2708 (N_2708,N_2523,N_1310);
xor U2709 (N_2709,N_2552,N_2428);
xnor U2710 (N_2710,N_2314,N_2440);
and U2711 (N_2711,N_2534,N_2542);
nand U2712 (N_2712,N_1415,N_749);
nor U2713 (N_2713,N_2405,N_2463);
nor U2714 (N_2714,N_2531,N_1206);
and U2715 (N_2715,N_2591,N_2515);
nand U2716 (N_2716,N_2520,N_2525);
nand U2717 (N_2717,N_1597,N_2488);
nand U2718 (N_2718,In_342,N_865);
nor U2719 (N_2719,N_2596,N_2535);
nor U2720 (N_2720,N_2564,N_2479);
nand U2721 (N_2721,N_1216,N_1679);
xor U2722 (N_2722,N_2587,In_526);
xor U2723 (N_2723,N_2444,N_2227);
xor U2724 (N_2724,N_2029,N_2433);
nand U2725 (N_2725,In_2612,In_2769);
xor U2726 (N_2726,N_2135,N_1280);
or U2727 (N_2727,N_2572,N_2588);
nand U2728 (N_2728,In_2363,N_2046);
or U2729 (N_2729,In_2529,N_2362);
nand U2730 (N_2730,N_2079,N_2495);
and U2731 (N_2731,N_2401,N_2459);
xor U2732 (N_2732,In_798,N_2070);
xnor U2733 (N_2733,N_2457,N_2597);
nor U2734 (N_2734,N_2432,N_2436);
or U2735 (N_2735,N_2585,N_2284);
and U2736 (N_2736,N_1918,N_2400);
nand U2737 (N_2737,N_2532,N_2358);
or U2738 (N_2738,N_2541,N_2303);
nand U2739 (N_2739,N_141,N_959);
and U2740 (N_2740,N_2475,N_2213);
nand U2741 (N_2741,N_2537,N_1270);
nor U2742 (N_2742,N_1763,N_2348);
nand U2743 (N_2743,N_2482,N_2580);
nor U2744 (N_2744,N_2305,In_2649);
nor U2745 (N_2745,N_2264,N_1757);
xnor U2746 (N_2746,N_2188,N_2568);
and U2747 (N_2747,N_2450,N_2315);
or U2748 (N_2748,N_1927,N_2514);
or U2749 (N_2749,N_2481,N_1328);
nor U2750 (N_2750,N_2492,N_2554);
and U2751 (N_2751,N_1330,In_2989);
xnor U2752 (N_2752,N_2406,N_2231);
or U2753 (N_2753,N_2409,N_2260);
xnor U2754 (N_2754,N_2064,N_2476);
nand U2755 (N_2755,N_2390,N_1842);
nand U2756 (N_2756,In_167,N_2593);
xnor U2757 (N_2757,N_2521,N_444);
nand U2758 (N_2758,N_1473,N_2498);
nor U2759 (N_2759,N_2349,N_2304);
or U2760 (N_2760,N_2503,N_2533);
nor U2761 (N_2761,N_2068,In_2195);
xnor U2762 (N_2762,N_2595,N_1631);
xnor U2763 (N_2763,N_2423,N_1735);
and U2764 (N_2764,N_2446,N_2473);
or U2765 (N_2765,N_2472,N_2598);
nand U2766 (N_2766,N_2466,N_2548);
nor U2767 (N_2767,In_626,N_2055);
xnor U2768 (N_2768,N_2058,N_2215);
and U2769 (N_2769,N_2038,N_2431);
xor U2770 (N_2770,N_2599,N_2408);
or U2771 (N_2771,N_2522,N_2209);
and U2772 (N_2772,N_2418,N_1985);
and U2773 (N_2773,In_1326,N_2370);
nand U2774 (N_2774,N_2506,N_2325);
nand U2775 (N_2775,N_2458,In_2493);
or U2776 (N_2776,N_2468,N_1755);
or U2777 (N_2777,N_2543,N_2569);
and U2778 (N_2778,N_2504,N_1509);
nand U2779 (N_2779,N_2579,N_2427);
or U2780 (N_2780,N_2477,N_1483);
nor U2781 (N_2781,N_2160,N_2536);
or U2782 (N_2782,N_1752,N_2425);
nor U2783 (N_2783,N_2565,N_2557);
and U2784 (N_2784,N_2539,N_2576);
xor U2785 (N_2785,N_2562,N_2447);
or U2786 (N_2786,N_2414,N_2206);
nor U2787 (N_2787,N_2480,N_2378);
or U2788 (N_2788,N_2225,N_2403);
or U2789 (N_2789,N_2229,N_2426);
or U2790 (N_2790,N_2574,N_2448);
nor U2791 (N_2791,N_2509,N_2497);
nor U2792 (N_2792,N_2270,N_2148);
nand U2793 (N_2793,N_2240,N_2232);
nand U2794 (N_2794,N_2527,N_2417);
xnor U2795 (N_2795,N_2372,N_1871);
and U2796 (N_2796,N_2162,N_2441);
nor U2797 (N_2797,N_2342,N_1363);
nor U2798 (N_2798,N_2578,N_2462);
nor U2799 (N_2799,N_2454,N_2402);
nand U2800 (N_2800,N_2709,N_2719);
and U2801 (N_2801,N_2684,N_2783);
or U2802 (N_2802,N_2677,N_2699);
and U2803 (N_2803,N_2713,N_2668);
or U2804 (N_2804,N_2718,N_2799);
or U2805 (N_2805,N_2639,N_2635);
or U2806 (N_2806,N_2728,N_2630);
or U2807 (N_2807,N_2647,N_2773);
nor U2808 (N_2808,N_2756,N_2735);
and U2809 (N_2809,N_2690,N_2696);
nand U2810 (N_2810,N_2765,N_2622);
nand U2811 (N_2811,N_2732,N_2664);
nor U2812 (N_2812,N_2620,N_2643);
or U2813 (N_2813,N_2753,N_2694);
nor U2814 (N_2814,N_2637,N_2663);
and U2815 (N_2815,N_2628,N_2623);
or U2816 (N_2816,N_2769,N_2665);
nor U2817 (N_2817,N_2605,N_2638);
nand U2818 (N_2818,N_2785,N_2767);
and U2819 (N_2819,N_2715,N_2727);
nand U2820 (N_2820,N_2680,N_2793);
and U2821 (N_2821,N_2698,N_2616);
nor U2822 (N_2822,N_2724,N_2776);
nand U2823 (N_2823,N_2688,N_2758);
nor U2824 (N_2824,N_2762,N_2611);
and U2825 (N_2825,N_2760,N_2786);
xor U2826 (N_2826,N_2681,N_2654);
or U2827 (N_2827,N_2743,N_2631);
xnor U2828 (N_2828,N_2657,N_2650);
and U2829 (N_2829,N_2703,N_2603);
and U2830 (N_2830,N_2777,N_2645);
nor U2831 (N_2831,N_2749,N_2775);
xnor U2832 (N_2832,N_2656,N_2619);
nor U2833 (N_2833,N_2658,N_2624);
nand U2834 (N_2834,N_2625,N_2636);
xnor U2835 (N_2835,N_2606,N_2738);
nor U2836 (N_2836,N_2771,N_2734);
nand U2837 (N_2837,N_2685,N_2669);
nor U2838 (N_2838,N_2692,N_2733);
nor U2839 (N_2839,N_2700,N_2644);
or U2840 (N_2840,N_2781,N_2655);
or U2841 (N_2841,N_2641,N_2748);
nor U2842 (N_2842,N_2780,N_2746);
nand U2843 (N_2843,N_2687,N_2774);
nor U2844 (N_2844,N_2798,N_2614);
and U2845 (N_2845,N_2676,N_2652);
xor U2846 (N_2846,N_2796,N_2744);
and U2847 (N_2847,N_2674,N_2768);
nand U2848 (N_2848,N_2626,N_2618);
nor U2849 (N_2849,N_2646,N_2686);
and U2850 (N_2850,N_2660,N_2717);
xor U2851 (N_2851,N_2742,N_2667);
nand U2852 (N_2852,N_2659,N_2731);
and U2853 (N_2853,N_2716,N_2615);
xor U2854 (N_2854,N_2633,N_2726);
xnor U2855 (N_2855,N_2705,N_2675);
and U2856 (N_2856,N_2601,N_2693);
nand U2857 (N_2857,N_2751,N_2683);
or U2858 (N_2858,N_2712,N_2662);
or U2859 (N_2859,N_2602,N_2792);
xnor U2860 (N_2860,N_2666,N_2609);
xor U2861 (N_2861,N_2782,N_2740);
nand U2862 (N_2862,N_2741,N_2607);
or U2863 (N_2863,N_2617,N_2629);
and U2864 (N_2864,N_2707,N_2691);
and U2865 (N_2865,N_2789,N_2621);
nand U2866 (N_2866,N_2640,N_2627);
nand U2867 (N_2867,N_2722,N_2737);
nor U2868 (N_2868,N_2610,N_2720);
xnor U2869 (N_2869,N_2600,N_2784);
xnor U2870 (N_2870,N_2711,N_2745);
and U2871 (N_2871,N_2770,N_2708);
nand U2872 (N_2872,N_2763,N_2797);
xnor U2873 (N_2873,N_2697,N_2642);
nand U2874 (N_2874,N_2604,N_2729);
xnor U2875 (N_2875,N_2747,N_2678);
and U2876 (N_2876,N_2723,N_2788);
nor U2877 (N_2877,N_2739,N_2766);
or U2878 (N_2878,N_2679,N_2701);
xnor U2879 (N_2879,N_2632,N_2649);
xor U2880 (N_2880,N_2653,N_2772);
and U2881 (N_2881,N_2759,N_2648);
or U2882 (N_2882,N_2671,N_2651);
and U2883 (N_2883,N_2778,N_2736);
nor U2884 (N_2884,N_2795,N_2682);
or U2885 (N_2885,N_2670,N_2752);
nor U2886 (N_2886,N_2672,N_2695);
and U2887 (N_2887,N_2613,N_2725);
nor U2888 (N_2888,N_2710,N_2714);
or U2889 (N_2889,N_2612,N_2794);
nand U2890 (N_2890,N_2761,N_2661);
nor U2891 (N_2891,N_2689,N_2721);
or U2892 (N_2892,N_2673,N_2791);
and U2893 (N_2893,N_2755,N_2702);
nand U2894 (N_2894,N_2787,N_2730);
nor U2895 (N_2895,N_2757,N_2704);
nand U2896 (N_2896,N_2764,N_2754);
xnor U2897 (N_2897,N_2750,N_2790);
or U2898 (N_2898,N_2608,N_2706);
or U2899 (N_2899,N_2634,N_2779);
nor U2900 (N_2900,N_2609,N_2630);
nand U2901 (N_2901,N_2682,N_2637);
nor U2902 (N_2902,N_2709,N_2624);
or U2903 (N_2903,N_2756,N_2614);
or U2904 (N_2904,N_2765,N_2796);
nand U2905 (N_2905,N_2671,N_2642);
nor U2906 (N_2906,N_2782,N_2757);
nand U2907 (N_2907,N_2796,N_2703);
nand U2908 (N_2908,N_2661,N_2694);
or U2909 (N_2909,N_2624,N_2682);
nor U2910 (N_2910,N_2643,N_2613);
nand U2911 (N_2911,N_2660,N_2637);
nor U2912 (N_2912,N_2787,N_2685);
or U2913 (N_2913,N_2702,N_2759);
nor U2914 (N_2914,N_2608,N_2746);
nand U2915 (N_2915,N_2771,N_2756);
nand U2916 (N_2916,N_2765,N_2682);
and U2917 (N_2917,N_2720,N_2601);
or U2918 (N_2918,N_2786,N_2622);
nand U2919 (N_2919,N_2765,N_2766);
and U2920 (N_2920,N_2704,N_2697);
nand U2921 (N_2921,N_2715,N_2734);
or U2922 (N_2922,N_2749,N_2788);
and U2923 (N_2923,N_2719,N_2740);
or U2924 (N_2924,N_2725,N_2779);
and U2925 (N_2925,N_2704,N_2637);
xnor U2926 (N_2926,N_2672,N_2776);
nor U2927 (N_2927,N_2604,N_2796);
xor U2928 (N_2928,N_2665,N_2733);
nor U2929 (N_2929,N_2667,N_2641);
nor U2930 (N_2930,N_2744,N_2606);
or U2931 (N_2931,N_2750,N_2644);
nand U2932 (N_2932,N_2737,N_2786);
xor U2933 (N_2933,N_2706,N_2723);
xnor U2934 (N_2934,N_2675,N_2763);
and U2935 (N_2935,N_2651,N_2678);
nor U2936 (N_2936,N_2686,N_2751);
nor U2937 (N_2937,N_2763,N_2667);
xor U2938 (N_2938,N_2784,N_2690);
or U2939 (N_2939,N_2648,N_2768);
or U2940 (N_2940,N_2792,N_2716);
or U2941 (N_2941,N_2722,N_2611);
or U2942 (N_2942,N_2763,N_2601);
nand U2943 (N_2943,N_2610,N_2736);
xnor U2944 (N_2944,N_2778,N_2641);
xnor U2945 (N_2945,N_2790,N_2740);
nand U2946 (N_2946,N_2723,N_2797);
or U2947 (N_2947,N_2687,N_2658);
and U2948 (N_2948,N_2789,N_2617);
nor U2949 (N_2949,N_2669,N_2624);
xor U2950 (N_2950,N_2670,N_2600);
or U2951 (N_2951,N_2781,N_2791);
nand U2952 (N_2952,N_2725,N_2734);
xnor U2953 (N_2953,N_2725,N_2681);
and U2954 (N_2954,N_2640,N_2723);
nand U2955 (N_2955,N_2746,N_2713);
or U2956 (N_2956,N_2757,N_2788);
or U2957 (N_2957,N_2637,N_2755);
xor U2958 (N_2958,N_2640,N_2762);
xnor U2959 (N_2959,N_2797,N_2639);
and U2960 (N_2960,N_2707,N_2775);
nor U2961 (N_2961,N_2796,N_2713);
nand U2962 (N_2962,N_2622,N_2728);
or U2963 (N_2963,N_2784,N_2789);
or U2964 (N_2964,N_2699,N_2619);
xnor U2965 (N_2965,N_2773,N_2680);
and U2966 (N_2966,N_2782,N_2734);
nand U2967 (N_2967,N_2750,N_2699);
nand U2968 (N_2968,N_2702,N_2677);
or U2969 (N_2969,N_2769,N_2742);
nor U2970 (N_2970,N_2615,N_2730);
nand U2971 (N_2971,N_2716,N_2703);
nor U2972 (N_2972,N_2604,N_2630);
nor U2973 (N_2973,N_2617,N_2725);
nand U2974 (N_2974,N_2611,N_2607);
or U2975 (N_2975,N_2664,N_2699);
nand U2976 (N_2976,N_2797,N_2726);
nand U2977 (N_2977,N_2608,N_2621);
or U2978 (N_2978,N_2726,N_2709);
nor U2979 (N_2979,N_2791,N_2676);
and U2980 (N_2980,N_2687,N_2739);
nor U2981 (N_2981,N_2790,N_2725);
or U2982 (N_2982,N_2655,N_2789);
or U2983 (N_2983,N_2632,N_2659);
nor U2984 (N_2984,N_2735,N_2796);
xnor U2985 (N_2985,N_2642,N_2767);
nor U2986 (N_2986,N_2704,N_2726);
xnor U2987 (N_2987,N_2619,N_2738);
nor U2988 (N_2988,N_2694,N_2645);
xnor U2989 (N_2989,N_2692,N_2735);
xor U2990 (N_2990,N_2663,N_2776);
nand U2991 (N_2991,N_2663,N_2750);
xor U2992 (N_2992,N_2663,N_2659);
nand U2993 (N_2993,N_2733,N_2734);
and U2994 (N_2994,N_2699,N_2679);
or U2995 (N_2995,N_2631,N_2600);
xor U2996 (N_2996,N_2605,N_2734);
nand U2997 (N_2997,N_2725,N_2787);
nand U2998 (N_2998,N_2658,N_2760);
or U2999 (N_2999,N_2606,N_2616);
nor U3000 (N_3000,N_2928,N_2825);
or U3001 (N_3001,N_2971,N_2830);
nor U3002 (N_3002,N_2887,N_2872);
nor U3003 (N_3003,N_2835,N_2803);
and U3004 (N_3004,N_2911,N_2921);
nand U3005 (N_3005,N_2805,N_2916);
and U3006 (N_3006,N_2960,N_2836);
xnor U3007 (N_3007,N_2972,N_2976);
nand U3008 (N_3008,N_2987,N_2854);
nand U3009 (N_3009,N_2858,N_2896);
nand U3010 (N_3010,N_2925,N_2938);
nor U3011 (N_3011,N_2945,N_2839);
or U3012 (N_3012,N_2885,N_2873);
and U3013 (N_3013,N_2826,N_2984);
and U3014 (N_3014,N_2841,N_2807);
nor U3015 (N_3015,N_2892,N_2943);
xor U3016 (N_3016,N_2821,N_2850);
and U3017 (N_3017,N_2931,N_2888);
and U3018 (N_3018,N_2894,N_2957);
or U3019 (N_3019,N_2920,N_2964);
or U3020 (N_3020,N_2950,N_2991);
and U3021 (N_3021,N_2905,N_2812);
or U3022 (N_3022,N_2901,N_2923);
nor U3023 (N_3023,N_2904,N_2862);
or U3024 (N_3024,N_2948,N_2910);
nor U3025 (N_3025,N_2927,N_2952);
nand U3026 (N_3026,N_2820,N_2906);
nand U3027 (N_3027,N_2809,N_2973);
or U3028 (N_3028,N_2818,N_2967);
and U3029 (N_3029,N_2875,N_2993);
and U3030 (N_3030,N_2840,N_2956);
or U3031 (N_3031,N_2986,N_2932);
nor U3032 (N_3032,N_2897,N_2893);
nor U3033 (N_3033,N_2823,N_2962);
nor U3034 (N_3034,N_2867,N_2937);
nand U3035 (N_3035,N_2969,N_2992);
or U3036 (N_3036,N_2856,N_2822);
nor U3037 (N_3037,N_2935,N_2814);
nand U3038 (N_3038,N_2806,N_2974);
or U3039 (N_3039,N_2870,N_2804);
and U3040 (N_3040,N_2908,N_2912);
nor U3041 (N_3041,N_2929,N_2918);
or U3042 (N_3042,N_2829,N_2847);
nor U3043 (N_3043,N_2878,N_2955);
nand U3044 (N_3044,N_2832,N_2917);
nand U3045 (N_3045,N_2919,N_2848);
nor U3046 (N_3046,N_2815,N_2977);
and U3047 (N_3047,N_2843,N_2801);
xnor U3048 (N_3048,N_2884,N_2936);
xor U3049 (N_3049,N_2869,N_2990);
nor U3050 (N_3050,N_2995,N_2914);
xor U3051 (N_3051,N_2933,N_2802);
nand U3052 (N_3052,N_2880,N_2819);
nand U3053 (N_3053,N_2842,N_2808);
and U3054 (N_3054,N_2865,N_2881);
xor U3055 (N_3055,N_2890,N_2999);
nor U3056 (N_3056,N_2926,N_2855);
or U3057 (N_3057,N_2951,N_2859);
and U3058 (N_3058,N_2970,N_2942);
nand U3059 (N_3059,N_2949,N_2982);
and U3060 (N_3060,N_2889,N_2898);
nand U3061 (N_3061,N_2810,N_2837);
nand U3062 (N_3062,N_2868,N_2980);
nor U3063 (N_3063,N_2874,N_2975);
nor U3064 (N_3064,N_2994,N_2909);
nand U3065 (N_3065,N_2891,N_2851);
nand U3066 (N_3066,N_2988,N_2834);
and U3067 (N_3067,N_2922,N_2954);
and U3068 (N_3068,N_2965,N_2939);
or U3069 (N_3069,N_2913,N_2981);
nand U3070 (N_3070,N_2966,N_2877);
xnor U3071 (N_3071,N_2940,N_2899);
and U3072 (N_3072,N_2866,N_2861);
nor U3073 (N_3073,N_2968,N_2852);
nand U3074 (N_3074,N_2998,N_2903);
and U3075 (N_3075,N_2816,N_2947);
and U3076 (N_3076,N_2963,N_2846);
or U3077 (N_3077,N_2882,N_2831);
and U3078 (N_3078,N_2857,N_2886);
and U3079 (N_3079,N_2863,N_2941);
and U3080 (N_3080,N_2883,N_2871);
xor U3081 (N_3081,N_2828,N_2983);
or U3082 (N_3082,N_2845,N_2979);
nor U3083 (N_3083,N_2985,N_2833);
nand U3084 (N_3084,N_2864,N_2879);
xnor U3085 (N_3085,N_2959,N_2876);
and U3086 (N_3086,N_2900,N_2849);
or U3087 (N_3087,N_2944,N_2930);
nor U3088 (N_3088,N_2958,N_2915);
nand U3089 (N_3089,N_2989,N_2895);
and U3090 (N_3090,N_2961,N_2907);
xor U3091 (N_3091,N_2817,N_2946);
nand U3092 (N_3092,N_2996,N_2953);
or U3093 (N_3093,N_2824,N_2838);
nand U3094 (N_3094,N_2813,N_2827);
nor U3095 (N_3095,N_2811,N_2844);
nand U3096 (N_3096,N_2902,N_2860);
or U3097 (N_3097,N_2800,N_2934);
and U3098 (N_3098,N_2997,N_2978);
xor U3099 (N_3099,N_2853,N_2924);
nor U3100 (N_3100,N_2980,N_2901);
xnor U3101 (N_3101,N_2919,N_2899);
and U3102 (N_3102,N_2917,N_2905);
nor U3103 (N_3103,N_2878,N_2880);
and U3104 (N_3104,N_2936,N_2964);
nor U3105 (N_3105,N_2909,N_2980);
xor U3106 (N_3106,N_2904,N_2822);
nor U3107 (N_3107,N_2886,N_2998);
and U3108 (N_3108,N_2901,N_2999);
nand U3109 (N_3109,N_2855,N_2882);
nor U3110 (N_3110,N_2828,N_2934);
nor U3111 (N_3111,N_2957,N_2945);
nand U3112 (N_3112,N_2833,N_2820);
nand U3113 (N_3113,N_2899,N_2903);
or U3114 (N_3114,N_2833,N_2897);
nand U3115 (N_3115,N_2914,N_2842);
and U3116 (N_3116,N_2962,N_2935);
nand U3117 (N_3117,N_2978,N_2923);
nand U3118 (N_3118,N_2802,N_2984);
nand U3119 (N_3119,N_2862,N_2893);
xor U3120 (N_3120,N_2840,N_2997);
nor U3121 (N_3121,N_2876,N_2828);
nor U3122 (N_3122,N_2992,N_2847);
nand U3123 (N_3123,N_2957,N_2885);
xnor U3124 (N_3124,N_2827,N_2853);
xor U3125 (N_3125,N_2888,N_2802);
nand U3126 (N_3126,N_2819,N_2876);
and U3127 (N_3127,N_2886,N_2928);
and U3128 (N_3128,N_2920,N_2817);
and U3129 (N_3129,N_2881,N_2927);
xor U3130 (N_3130,N_2934,N_2894);
and U3131 (N_3131,N_2918,N_2857);
nor U3132 (N_3132,N_2961,N_2918);
xnor U3133 (N_3133,N_2967,N_2903);
nand U3134 (N_3134,N_2830,N_2897);
nor U3135 (N_3135,N_2929,N_2994);
or U3136 (N_3136,N_2911,N_2940);
nor U3137 (N_3137,N_2979,N_2915);
or U3138 (N_3138,N_2870,N_2856);
nand U3139 (N_3139,N_2811,N_2987);
nand U3140 (N_3140,N_2900,N_2938);
and U3141 (N_3141,N_2825,N_2994);
and U3142 (N_3142,N_2911,N_2837);
nor U3143 (N_3143,N_2910,N_2946);
nand U3144 (N_3144,N_2923,N_2953);
or U3145 (N_3145,N_2865,N_2871);
xnor U3146 (N_3146,N_2878,N_2990);
or U3147 (N_3147,N_2927,N_2817);
xnor U3148 (N_3148,N_2957,N_2936);
nor U3149 (N_3149,N_2913,N_2955);
or U3150 (N_3150,N_2836,N_2864);
nand U3151 (N_3151,N_2924,N_2902);
and U3152 (N_3152,N_2918,N_2823);
or U3153 (N_3153,N_2826,N_2875);
or U3154 (N_3154,N_2951,N_2838);
or U3155 (N_3155,N_2940,N_2871);
xor U3156 (N_3156,N_2863,N_2957);
xnor U3157 (N_3157,N_2916,N_2966);
and U3158 (N_3158,N_2920,N_2992);
nor U3159 (N_3159,N_2907,N_2890);
and U3160 (N_3160,N_2935,N_2983);
nand U3161 (N_3161,N_2805,N_2949);
nand U3162 (N_3162,N_2950,N_2954);
nand U3163 (N_3163,N_2985,N_2848);
xor U3164 (N_3164,N_2820,N_2995);
or U3165 (N_3165,N_2837,N_2922);
nor U3166 (N_3166,N_2872,N_2971);
and U3167 (N_3167,N_2870,N_2886);
xnor U3168 (N_3168,N_2976,N_2845);
xor U3169 (N_3169,N_2869,N_2971);
nor U3170 (N_3170,N_2901,N_2825);
and U3171 (N_3171,N_2894,N_2886);
xnor U3172 (N_3172,N_2911,N_2998);
xnor U3173 (N_3173,N_2943,N_2824);
and U3174 (N_3174,N_2803,N_2878);
and U3175 (N_3175,N_2906,N_2989);
xnor U3176 (N_3176,N_2909,N_2974);
and U3177 (N_3177,N_2857,N_2882);
nor U3178 (N_3178,N_2939,N_2863);
or U3179 (N_3179,N_2896,N_2999);
or U3180 (N_3180,N_2927,N_2922);
xor U3181 (N_3181,N_2848,N_2872);
and U3182 (N_3182,N_2968,N_2974);
and U3183 (N_3183,N_2962,N_2910);
or U3184 (N_3184,N_2898,N_2920);
or U3185 (N_3185,N_2898,N_2934);
or U3186 (N_3186,N_2998,N_2910);
or U3187 (N_3187,N_2948,N_2958);
nand U3188 (N_3188,N_2824,N_2989);
nand U3189 (N_3189,N_2869,N_2812);
or U3190 (N_3190,N_2981,N_2848);
nand U3191 (N_3191,N_2926,N_2937);
nor U3192 (N_3192,N_2841,N_2933);
and U3193 (N_3193,N_2933,N_2986);
and U3194 (N_3194,N_2925,N_2869);
and U3195 (N_3195,N_2889,N_2984);
and U3196 (N_3196,N_2803,N_2998);
or U3197 (N_3197,N_2967,N_2969);
and U3198 (N_3198,N_2947,N_2884);
xor U3199 (N_3199,N_2882,N_2900);
nor U3200 (N_3200,N_3047,N_3133);
xor U3201 (N_3201,N_3007,N_3137);
or U3202 (N_3202,N_3129,N_3051);
or U3203 (N_3203,N_3166,N_3145);
xor U3204 (N_3204,N_3004,N_3013);
and U3205 (N_3205,N_3080,N_3075);
nand U3206 (N_3206,N_3082,N_3087);
and U3207 (N_3207,N_3054,N_3086);
nand U3208 (N_3208,N_3159,N_3117);
xor U3209 (N_3209,N_3027,N_3081);
xor U3210 (N_3210,N_3164,N_3084);
nand U3211 (N_3211,N_3008,N_3098);
and U3212 (N_3212,N_3128,N_3088);
nand U3213 (N_3213,N_3093,N_3114);
nor U3214 (N_3214,N_3123,N_3005);
nand U3215 (N_3215,N_3076,N_3132);
nand U3216 (N_3216,N_3192,N_3060);
xor U3217 (N_3217,N_3169,N_3174);
xnor U3218 (N_3218,N_3062,N_3110);
and U3219 (N_3219,N_3194,N_3101);
nor U3220 (N_3220,N_3085,N_3193);
xor U3221 (N_3221,N_3138,N_3154);
or U3222 (N_3222,N_3023,N_3028);
and U3223 (N_3223,N_3189,N_3002);
or U3224 (N_3224,N_3160,N_3172);
xnor U3225 (N_3225,N_3018,N_3183);
nor U3226 (N_3226,N_3000,N_3177);
and U3227 (N_3227,N_3178,N_3014);
nand U3228 (N_3228,N_3125,N_3141);
nand U3229 (N_3229,N_3115,N_3078);
or U3230 (N_3230,N_3040,N_3056);
and U3231 (N_3231,N_3171,N_3064);
nand U3232 (N_3232,N_3143,N_3030);
or U3233 (N_3233,N_3100,N_3197);
nand U3234 (N_3234,N_3144,N_3147);
xnor U3235 (N_3235,N_3130,N_3184);
xor U3236 (N_3236,N_3006,N_3071);
and U3237 (N_3237,N_3083,N_3079);
nor U3238 (N_3238,N_3161,N_3042);
or U3239 (N_3239,N_3155,N_3034);
or U3240 (N_3240,N_3150,N_3163);
xor U3241 (N_3241,N_3126,N_3070);
nor U3242 (N_3242,N_3066,N_3121);
or U3243 (N_3243,N_3022,N_3041);
nor U3244 (N_3244,N_3165,N_3103);
or U3245 (N_3245,N_3196,N_3118);
and U3246 (N_3246,N_3146,N_3190);
and U3247 (N_3247,N_3059,N_3127);
xnor U3248 (N_3248,N_3109,N_3020);
xnor U3249 (N_3249,N_3156,N_3122);
nor U3250 (N_3250,N_3046,N_3061);
and U3251 (N_3251,N_3116,N_3096);
nand U3252 (N_3252,N_3095,N_3058);
xor U3253 (N_3253,N_3072,N_3015);
nand U3254 (N_3254,N_3113,N_3199);
nand U3255 (N_3255,N_3037,N_3025);
nand U3256 (N_3256,N_3131,N_3175);
and U3257 (N_3257,N_3043,N_3050);
xor U3258 (N_3258,N_3182,N_3019);
and U3259 (N_3259,N_3011,N_3167);
or U3260 (N_3260,N_3111,N_3107);
and U3261 (N_3261,N_3057,N_3029);
and U3262 (N_3262,N_3135,N_3017);
nor U3263 (N_3263,N_3055,N_3038);
nand U3264 (N_3264,N_3136,N_3105);
nand U3265 (N_3265,N_3195,N_3024);
nand U3266 (N_3266,N_3089,N_3120);
xor U3267 (N_3267,N_3092,N_3010);
and U3268 (N_3268,N_3090,N_3067);
nor U3269 (N_3269,N_3104,N_3035);
or U3270 (N_3270,N_3162,N_3185);
or U3271 (N_3271,N_3012,N_3099);
nand U3272 (N_3272,N_3153,N_3097);
or U3273 (N_3273,N_3069,N_3026);
nor U3274 (N_3274,N_3049,N_3140);
xnor U3275 (N_3275,N_3108,N_3003);
xor U3276 (N_3276,N_3102,N_3170);
nor U3277 (N_3277,N_3045,N_3001);
nor U3278 (N_3278,N_3106,N_3091);
or U3279 (N_3279,N_3158,N_3181);
nand U3280 (N_3280,N_3074,N_3188);
nand U3281 (N_3281,N_3180,N_3009);
and U3282 (N_3282,N_3142,N_3063);
nor U3283 (N_3283,N_3053,N_3033);
xor U3284 (N_3284,N_3149,N_3186);
nor U3285 (N_3285,N_3191,N_3173);
xor U3286 (N_3286,N_3016,N_3065);
nor U3287 (N_3287,N_3148,N_3179);
or U3288 (N_3288,N_3139,N_3031);
xnor U3289 (N_3289,N_3073,N_3036);
and U3290 (N_3290,N_3198,N_3176);
and U3291 (N_3291,N_3021,N_3044);
or U3292 (N_3292,N_3039,N_3119);
nor U3293 (N_3293,N_3157,N_3094);
xor U3294 (N_3294,N_3134,N_3152);
nand U3295 (N_3295,N_3151,N_3048);
xor U3296 (N_3296,N_3187,N_3032);
nand U3297 (N_3297,N_3124,N_3168);
nor U3298 (N_3298,N_3068,N_3052);
nand U3299 (N_3299,N_3112,N_3077);
and U3300 (N_3300,N_3164,N_3135);
or U3301 (N_3301,N_3154,N_3028);
nand U3302 (N_3302,N_3166,N_3071);
or U3303 (N_3303,N_3134,N_3127);
or U3304 (N_3304,N_3067,N_3040);
and U3305 (N_3305,N_3002,N_3169);
xnor U3306 (N_3306,N_3016,N_3082);
and U3307 (N_3307,N_3036,N_3067);
nand U3308 (N_3308,N_3104,N_3126);
nand U3309 (N_3309,N_3169,N_3093);
nand U3310 (N_3310,N_3175,N_3156);
and U3311 (N_3311,N_3196,N_3150);
nand U3312 (N_3312,N_3098,N_3103);
nor U3313 (N_3313,N_3021,N_3050);
nor U3314 (N_3314,N_3030,N_3149);
and U3315 (N_3315,N_3073,N_3181);
and U3316 (N_3316,N_3008,N_3033);
nor U3317 (N_3317,N_3057,N_3091);
and U3318 (N_3318,N_3140,N_3098);
xor U3319 (N_3319,N_3190,N_3124);
nor U3320 (N_3320,N_3177,N_3065);
or U3321 (N_3321,N_3120,N_3180);
and U3322 (N_3322,N_3157,N_3051);
nor U3323 (N_3323,N_3184,N_3056);
xor U3324 (N_3324,N_3173,N_3107);
or U3325 (N_3325,N_3158,N_3198);
xor U3326 (N_3326,N_3122,N_3001);
nor U3327 (N_3327,N_3024,N_3101);
nand U3328 (N_3328,N_3108,N_3188);
nand U3329 (N_3329,N_3054,N_3049);
xnor U3330 (N_3330,N_3134,N_3089);
and U3331 (N_3331,N_3034,N_3028);
nor U3332 (N_3332,N_3169,N_3050);
or U3333 (N_3333,N_3044,N_3118);
and U3334 (N_3334,N_3059,N_3176);
and U3335 (N_3335,N_3024,N_3179);
and U3336 (N_3336,N_3059,N_3196);
xor U3337 (N_3337,N_3139,N_3142);
nand U3338 (N_3338,N_3157,N_3141);
xor U3339 (N_3339,N_3088,N_3042);
xor U3340 (N_3340,N_3147,N_3146);
xnor U3341 (N_3341,N_3008,N_3088);
nor U3342 (N_3342,N_3080,N_3131);
nand U3343 (N_3343,N_3032,N_3085);
and U3344 (N_3344,N_3143,N_3172);
or U3345 (N_3345,N_3183,N_3080);
nor U3346 (N_3346,N_3138,N_3195);
nor U3347 (N_3347,N_3033,N_3128);
xnor U3348 (N_3348,N_3045,N_3179);
xnor U3349 (N_3349,N_3158,N_3167);
and U3350 (N_3350,N_3035,N_3066);
nor U3351 (N_3351,N_3177,N_3109);
nor U3352 (N_3352,N_3194,N_3013);
xnor U3353 (N_3353,N_3186,N_3076);
nor U3354 (N_3354,N_3160,N_3175);
and U3355 (N_3355,N_3124,N_3021);
xnor U3356 (N_3356,N_3054,N_3148);
xnor U3357 (N_3357,N_3051,N_3087);
xor U3358 (N_3358,N_3102,N_3187);
or U3359 (N_3359,N_3067,N_3020);
and U3360 (N_3360,N_3046,N_3134);
nand U3361 (N_3361,N_3071,N_3050);
nand U3362 (N_3362,N_3181,N_3186);
xnor U3363 (N_3363,N_3113,N_3022);
xor U3364 (N_3364,N_3162,N_3078);
and U3365 (N_3365,N_3164,N_3001);
xor U3366 (N_3366,N_3178,N_3008);
nor U3367 (N_3367,N_3120,N_3175);
xor U3368 (N_3368,N_3103,N_3063);
xor U3369 (N_3369,N_3084,N_3016);
or U3370 (N_3370,N_3184,N_3010);
and U3371 (N_3371,N_3131,N_3181);
nor U3372 (N_3372,N_3108,N_3032);
xor U3373 (N_3373,N_3044,N_3183);
xor U3374 (N_3374,N_3120,N_3103);
nand U3375 (N_3375,N_3151,N_3001);
or U3376 (N_3376,N_3058,N_3129);
or U3377 (N_3377,N_3057,N_3030);
xnor U3378 (N_3378,N_3159,N_3039);
and U3379 (N_3379,N_3078,N_3158);
or U3380 (N_3380,N_3093,N_3132);
nand U3381 (N_3381,N_3164,N_3046);
or U3382 (N_3382,N_3025,N_3186);
xor U3383 (N_3383,N_3073,N_3100);
xnor U3384 (N_3384,N_3137,N_3027);
or U3385 (N_3385,N_3122,N_3137);
xor U3386 (N_3386,N_3042,N_3057);
nand U3387 (N_3387,N_3091,N_3135);
nand U3388 (N_3388,N_3139,N_3165);
nand U3389 (N_3389,N_3054,N_3152);
and U3390 (N_3390,N_3072,N_3064);
or U3391 (N_3391,N_3190,N_3182);
xor U3392 (N_3392,N_3097,N_3038);
and U3393 (N_3393,N_3197,N_3179);
nor U3394 (N_3394,N_3108,N_3157);
nor U3395 (N_3395,N_3046,N_3036);
and U3396 (N_3396,N_3176,N_3086);
or U3397 (N_3397,N_3001,N_3157);
and U3398 (N_3398,N_3168,N_3034);
xor U3399 (N_3399,N_3124,N_3071);
and U3400 (N_3400,N_3358,N_3209);
nand U3401 (N_3401,N_3266,N_3391);
nor U3402 (N_3402,N_3272,N_3331);
nor U3403 (N_3403,N_3367,N_3220);
or U3404 (N_3404,N_3216,N_3298);
xnor U3405 (N_3405,N_3218,N_3312);
nor U3406 (N_3406,N_3378,N_3265);
xnor U3407 (N_3407,N_3355,N_3339);
and U3408 (N_3408,N_3241,N_3305);
or U3409 (N_3409,N_3325,N_3307);
and U3410 (N_3410,N_3208,N_3222);
nor U3411 (N_3411,N_3205,N_3296);
nor U3412 (N_3412,N_3225,N_3233);
or U3413 (N_3413,N_3314,N_3224);
nand U3414 (N_3414,N_3267,N_3369);
nand U3415 (N_3415,N_3376,N_3246);
nor U3416 (N_3416,N_3277,N_3282);
and U3417 (N_3417,N_3235,N_3306);
xor U3418 (N_3418,N_3336,N_3219);
nor U3419 (N_3419,N_3395,N_3327);
xor U3420 (N_3420,N_3399,N_3291);
and U3421 (N_3421,N_3340,N_3288);
nand U3422 (N_3422,N_3384,N_3309);
nand U3423 (N_3423,N_3381,N_3351);
and U3424 (N_3424,N_3249,N_3210);
nor U3425 (N_3425,N_3337,N_3356);
xnor U3426 (N_3426,N_3290,N_3315);
and U3427 (N_3427,N_3281,N_3365);
xor U3428 (N_3428,N_3385,N_3343);
xor U3429 (N_3429,N_3338,N_3260);
or U3430 (N_3430,N_3389,N_3238);
nand U3431 (N_3431,N_3326,N_3375);
nand U3432 (N_3432,N_3251,N_3230);
nand U3433 (N_3433,N_3313,N_3371);
or U3434 (N_3434,N_3348,N_3239);
nor U3435 (N_3435,N_3259,N_3345);
nor U3436 (N_3436,N_3354,N_3333);
or U3437 (N_3437,N_3328,N_3254);
or U3438 (N_3438,N_3321,N_3357);
nand U3439 (N_3439,N_3329,N_3271);
and U3440 (N_3440,N_3317,N_3200);
or U3441 (N_3441,N_3289,N_3353);
nand U3442 (N_3442,N_3394,N_3300);
nand U3443 (N_3443,N_3203,N_3244);
and U3444 (N_3444,N_3373,N_3231);
and U3445 (N_3445,N_3202,N_3303);
or U3446 (N_3446,N_3372,N_3311);
and U3447 (N_3447,N_3279,N_3363);
or U3448 (N_3448,N_3269,N_3276);
nor U3449 (N_3449,N_3264,N_3212);
or U3450 (N_3450,N_3310,N_3280);
xnor U3451 (N_3451,N_3286,N_3390);
nor U3452 (N_3452,N_3293,N_3250);
nor U3453 (N_3453,N_3240,N_3302);
or U3454 (N_3454,N_3330,N_3334);
and U3455 (N_3455,N_3344,N_3262);
xnor U3456 (N_3456,N_3347,N_3253);
xnor U3457 (N_3457,N_3297,N_3226);
nor U3458 (N_3458,N_3304,N_3228);
and U3459 (N_3459,N_3227,N_3256);
nand U3460 (N_3460,N_3319,N_3287);
nor U3461 (N_3461,N_3215,N_3388);
or U3462 (N_3462,N_3229,N_3382);
nor U3463 (N_3463,N_3273,N_3285);
nor U3464 (N_3464,N_3350,N_3323);
nand U3465 (N_3465,N_3318,N_3361);
and U3466 (N_3466,N_3234,N_3379);
xor U3467 (N_3467,N_3362,N_3397);
or U3468 (N_3468,N_3346,N_3257);
or U3469 (N_3469,N_3268,N_3322);
nor U3470 (N_3470,N_3393,N_3324);
nor U3471 (N_3471,N_3217,N_3352);
and U3472 (N_3472,N_3242,N_3247);
nor U3473 (N_3473,N_3236,N_3275);
nor U3474 (N_3474,N_3335,N_3221);
nand U3475 (N_3475,N_3214,N_3243);
xor U3476 (N_3476,N_3255,N_3360);
xnor U3477 (N_3477,N_3301,N_3342);
xnor U3478 (N_3478,N_3223,N_3207);
xnor U3479 (N_3479,N_3349,N_3366);
or U3480 (N_3480,N_3232,N_3364);
and U3481 (N_3481,N_3341,N_3320);
nor U3482 (N_3482,N_3204,N_3211);
and U3483 (N_3483,N_3270,N_3374);
xor U3484 (N_3484,N_3308,N_3213);
or U3485 (N_3485,N_3377,N_3258);
xnor U3486 (N_3486,N_3294,N_3201);
nor U3487 (N_3487,N_3386,N_3206);
or U3488 (N_3488,N_3387,N_3396);
nor U3489 (N_3489,N_3359,N_3332);
nand U3490 (N_3490,N_3278,N_3283);
or U3491 (N_3491,N_3263,N_3248);
nor U3492 (N_3492,N_3261,N_3370);
xnor U3493 (N_3493,N_3368,N_3295);
or U3494 (N_3494,N_3398,N_3383);
nand U3495 (N_3495,N_3292,N_3299);
nand U3496 (N_3496,N_3274,N_3237);
nor U3497 (N_3497,N_3392,N_3245);
nand U3498 (N_3498,N_3380,N_3316);
or U3499 (N_3499,N_3252,N_3284);
or U3500 (N_3500,N_3232,N_3213);
and U3501 (N_3501,N_3393,N_3314);
and U3502 (N_3502,N_3366,N_3398);
xor U3503 (N_3503,N_3282,N_3241);
nand U3504 (N_3504,N_3207,N_3290);
or U3505 (N_3505,N_3387,N_3331);
or U3506 (N_3506,N_3205,N_3209);
or U3507 (N_3507,N_3385,N_3244);
and U3508 (N_3508,N_3235,N_3381);
nor U3509 (N_3509,N_3310,N_3266);
nor U3510 (N_3510,N_3232,N_3224);
xor U3511 (N_3511,N_3281,N_3321);
nand U3512 (N_3512,N_3362,N_3357);
nor U3513 (N_3513,N_3398,N_3265);
and U3514 (N_3514,N_3302,N_3281);
nor U3515 (N_3515,N_3310,N_3311);
nor U3516 (N_3516,N_3254,N_3318);
and U3517 (N_3517,N_3236,N_3387);
and U3518 (N_3518,N_3338,N_3311);
or U3519 (N_3519,N_3216,N_3338);
nor U3520 (N_3520,N_3338,N_3278);
nor U3521 (N_3521,N_3281,N_3398);
xnor U3522 (N_3522,N_3287,N_3326);
nand U3523 (N_3523,N_3217,N_3364);
nor U3524 (N_3524,N_3257,N_3254);
nor U3525 (N_3525,N_3258,N_3227);
nand U3526 (N_3526,N_3382,N_3364);
nor U3527 (N_3527,N_3231,N_3337);
nand U3528 (N_3528,N_3302,N_3381);
xnor U3529 (N_3529,N_3207,N_3200);
xor U3530 (N_3530,N_3335,N_3204);
and U3531 (N_3531,N_3359,N_3341);
or U3532 (N_3532,N_3276,N_3277);
or U3533 (N_3533,N_3238,N_3321);
and U3534 (N_3534,N_3377,N_3331);
xor U3535 (N_3535,N_3256,N_3365);
nand U3536 (N_3536,N_3226,N_3247);
nand U3537 (N_3537,N_3267,N_3213);
nand U3538 (N_3538,N_3361,N_3227);
nor U3539 (N_3539,N_3318,N_3267);
or U3540 (N_3540,N_3341,N_3228);
and U3541 (N_3541,N_3244,N_3283);
xnor U3542 (N_3542,N_3317,N_3260);
or U3543 (N_3543,N_3364,N_3271);
and U3544 (N_3544,N_3390,N_3361);
xnor U3545 (N_3545,N_3265,N_3260);
nand U3546 (N_3546,N_3353,N_3317);
and U3547 (N_3547,N_3323,N_3228);
or U3548 (N_3548,N_3234,N_3347);
or U3549 (N_3549,N_3212,N_3331);
or U3550 (N_3550,N_3221,N_3289);
xnor U3551 (N_3551,N_3391,N_3339);
nand U3552 (N_3552,N_3225,N_3300);
and U3553 (N_3553,N_3276,N_3319);
xnor U3554 (N_3554,N_3230,N_3359);
nand U3555 (N_3555,N_3225,N_3264);
and U3556 (N_3556,N_3275,N_3306);
and U3557 (N_3557,N_3294,N_3245);
or U3558 (N_3558,N_3381,N_3236);
and U3559 (N_3559,N_3305,N_3301);
xnor U3560 (N_3560,N_3265,N_3376);
xor U3561 (N_3561,N_3223,N_3397);
xor U3562 (N_3562,N_3300,N_3377);
xor U3563 (N_3563,N_3394,N_3329);
or U3564 (N_3564,N_3244,N_3358);
nand U3565 (N_3565,N_3312,N_3327);
nand U3566 (N_3566,N_3346,N_3246);
nand U3567 (N_3567,N_3328,N_3349);
nand U3568 (N_3568,N_3275,N_3276);
or U3569 (N_3569,N_3225,N_3396);
or U3570 (N_3570,N_3385,N_3381);
nand U3571 (N_3571,N_3345,N_3265);
or U3572 (N_3572,N_3244,N_3351);
nand U3573 (N_3573,N_3213,N_3275);
or U3574 (N_3574,N_3390,N_3395);
or U3575 (N_3575,N_3223,N_3283);
or U3576 (N_3576,N_3252,N_3215);
or U3577 (N_3577,N_3200,N_3361);
nor U3578 (N_3578,N_3291,N_3323);
nor U3579 (N_3579,N_3392,N_3223);
nor U3580 (N_3580,N_3316,N_3347);
nor U3581 (N_3581,N_3206,N_3362);
xor U3582 (N_3582,N_3329,N_3380);
or U3583 (N_3583,N_3262,N_3391);
and U3584 (N_3584,N_3329,N_3213);
nor U3585 (N_3585,N_3393,N_3209);
nand U3586 (N_3586,N_3382,N_3390);
or U3587 (N_3587,N_3314,N_3310);
or U3588 (N_3588,N_3360,N_3264);
or U3589 (N_3589,N_3364,N_3365);
xor U3590 (N_3590,N_3350,N_3249);
or U3591 (N_3591,N_3361,N_3248);
nand U3592 (N_3592,N_3285,N_3395);
nand U3593 (N_3593,N_3334,N_3393);
xnor U3594 (N_3594,N_3219,N_3397);
or U3595 (N_3595,N_3331,N_3333);
and U3596 (N_3596,N_3316,N_3202);
and U3597 (N_3597,N_3324,N_3360);
nor U3598 (N_3598,N_3331,N_3203);
nor U3599 (N_3599,N_3228,N_3289);
nor U3600 (N_3600,N_3577,N_3460);
nand U3601 (N_3601,N_3424,N_3403);
nand U3602 (N_3602,N_3492,N_3401);
xnor U3603 (N_3603,N_3407,N_3428);
nor U3604 (N_3604,N_3525,N_3469);
nand U3605 (N_3605,N_3514,N_3489);
nand U3606 (N_3606,N_3464,N_3593);
or U3607 (N_3607,N_3473,N_3420);
or U3608 (N_3608,N_3459,N_3440);
nor U3609 (N_3609,N_3470,N_3505);
nand U3610 (N_3610,N_3538,N_3481);
xnor U3611 (N_3611,N_3565,N_3432);
or U3612 (N_3612,N_3485,N_3591);
nor U3613 (N_3613,N_3445,N_3595);
and U3614 (N_3614,N_3461,N_3465);
xor U3615 (N_3615,N_3524,N_3587);
and U3616 (N_3616,N_3497,N_3520);
xnor U3617 (N_3617,N_3521,N_3433);
xor U3618 (N_3618,N_3430,N_3502);
nor U3619 (N_3619,N_3567,N_3418);
xnor U3620 (N_3620,N_3496,N_3490);
and U3621 (N_3621,N_3527,N_3478);
or U3622 (N_3622,N_3541,N_3531);
nor U3623 (N_3623,N_3457,N_3536);
nor U3624 (N_3624,N_3439,N_3406);
and U3625 (N_3625,N_3471,N_3443);
nand U3626 (N_3626,N_3426,N_3556);
and U3627 (N_3627,N_3557,N_3472);
nor U3628 (N_3628,N_3411,N_3421);
nor U3629 (N_3629,N_3571,N_3451);
or U3630 (N_3630,N_3408,N_3437);
nand U3631 (N_3631,N_3599,N_3419);
nor U3632 (N_3632,N_3572,N_3503);
xor U3633 (N_3633,N_3512,N_3410);
xnor U3634 (N_3634,N_3530,N_3491);
nand U3635 (N_3635,N_3546,N_3553);
and U3636 (N_3636,N_3441,N_3523);
or U3637 (N_3637,N_3494,N_3518);
nor U3638 (N_3638,N_3549,N_3559);
xor U3639 (N_3639,N_3533,N_3542);
and U3640 (N_3640,N_3581,N_3598);
nor U3641 (N_3641,N_3551,N_3462);
nand U3642 (N_3642,N_3509,N_3574);
or U3643 (N_3643,N_3501,N_3522);
xor U3644 (N_3644,N_3402,N_3414);
and U3645 (N_3645,N_3575,N_3488);
xor U3646 (N_3646,N_3422,N_3544);
nand U3647 (N_3647,N_3539,N_3586);
and U3648 (N_3648,N_3526,N_3555);
and U3649 (N_3649,N_3409,N_3429);
nand U3650 (N_3650,N_3467,N_3552);
xor U3651 (N_3651,N_3561,N_3540);
or U3652 (N_3652,N_3436,N_3550);
xor U3653 (N_3653,N_3589,N_3417);
xnor U3654 (N_3654,N_3579,N_3435);
and U3655 (N_3655,N_3506,N_3534);
and U3656 (N_3656,N_3442,N_3529);
nor U3657 (N_3657,N_3583,N_3573);
or U3658 (N_3658,N_3519,N_3570);
and U3659 (N_3659,N_3596,N_3486);
nor U3660 (N_3660,N_3484,N_3427);
xor U3661 (N_3661,N_3498,N_3569);
xnor U3662 (N_3662,N_3483,N_3588);
nand U3663 (N_3663,N_3590,N_3558);
nand U3664 (N_3664,N_3476,N_3532);
and U3665 (N_3665,N_3480,N_3515);
nor U3666 (N_3666,N_3463,N_3444);
and U3667 (N_3667,N_3563,N_3450);
or U3668 (N_3668,N_3511,N_3487);
xor U3669 (N_3669,N_3431,N_3425);
nor U3670 (N_3670,N_3517,N_3400);
nand U3671 (N_3671,N_3415,N_3477);
nand U3672 (N_3672,N_3499,N_3447);
nor U3673 (N_3673,N_3543,N_3438);
nor U3674 (N_3674,N_3547,N_3566);
and U3675 (N_3675,N_3548,N_3453);
nand U3676 (N_3676,N_3452,N_3592);
and U3677 (N_3677,N_3597,N_3448);
nor U3678 (N_3678,N_3585,N_3560);
xor U3679 (N_3679,N_3510,N_3413);
and U3680 (N_3680,N_3562,N_3564);
and U3681 (N_3681,N_3423,N_3456);
nor U3682 (N_3682,N_3535,N_3454);
xor U3683 (N_3683,N_3449,N_3537);
or U3684 (N_3684,N_3495,N_3493);
nor U3685 (N_3685,N_3458,N_3578);
xnor U3686 (N_3686,N_3504,N_3568);
nand U3687 (N_3687,N_3479,N_3584);
nand U3688 (N_3688,N_3405,N_3446);
xor U3689 (N_3689,N_3404,N_3455);
nor U3690 (N_3690,N_3528,N_3412);
xnor U3691 (N_3691,N_3554,N_3468);
xor U3692 (N_3692,N_3466,N_3516);
nor U3693 (N_3693,N_3434,N_3594);
or U3694 (N_3694,N_3507,N_3416);
and U3695 (N_3695,N_3580,N_3582);
or U3696 (N_3696,N_3513,N_3475);
nand U3697 (N_3697,N_3576,N_3545);
or U3698 (N_3698,N_3474,N_3500);
nor U3699 (N_3699,N_3508,N_3482);
and U3700 (N_3700,N_3577,N_3403);
nor U3701 (N_3701,N_3531,N_3459);
or U3702 (N_3702,N_3445,N_3404);
or U3703 (N_3703,N_3597,N_3574);
xor U3704 (N_3704,N_3430,N_3401);
nand U3705 (N_3705,N_3422,N_3452);
nor U3706 (N_3706,N_3494,N_3504);
nor U3707 (N_3707,N_3426,N_3598);
and U3708 (N_3708,N_3584,N_3564);
or U3709 (N_3709,N_3551,N_3578);
or U3710 (N_3710,N_3582,N_3405);
nor U3711 (N_3711,N_3415,N_3502);
xnor U3712 (N_3712,N_3553,N_3427);
nand U3713 (N_3713,N_3576,N_3500);
and U3714 (N_3714,N_3407,N_3435);
nand U3715 (N_3715,N_3584,N_3556);
xor U3716 (N_3716,N_3419,N_3441);
nand U3717 (N_3717,N_3429,N_3572);
nand U3718 (N_3718,N_3593,N_3566);
and U3719 (N_3719,N_3406,N_3515);
and U3720 (N_3720,N_3463,N_3483);
xnor U3721 (N_3721,N_3549,N_3447);
xnor U3722 (N_3722,N_3530,N_3582);
xor U3723 (N_3723,N_3517,N_3557);
and U3724 (N_3724,N_3568,N_3597);
and U3725 (N_3725,N_3509,N_3402);
nand U3726 (N_3726,N_3587,N_3412);
xor U3727 (N_3727,N_3545,N_3458);
xor U3728 (N_3728,N_3565,N_3474);
and U3729 (N_3729,N_3569,N_3422);
nand U3730 (N_3730,N_3413,N_3564);
and U3731 (N_3731,N_3485,N_3548);
and U3732 (N_3732,N_3453,N_3470);
or U3733 (N_3733,N_3506,N_3465);
and U3734 (N_3734,N_3511,N_3593);
nand U3735 (N_3735,N_3588,N_3469);
nand U3736 (N_3736,N_3575,N_3518);
and U3737 (N_3737,N_3564,N_3426);
nand U3738 (N_3738,N_3564,N_3585);
and U3739 (N_3739,N_3560,N_3579);
nand U3740 (N_3740,N_3471,N_3557);
or U3741 (N_3741,N_3480,N_3421);
xor U3742 (N_3742,N_3574,N_3515);
xnor U3743 (N_3743,N_3545,N_3592);
nand U3744 (N_3744,N_3591,N_3447);
nor U3745 (N_3745,N_3501,N_3499);
and U3746 (N_3746,N_3468,N_3455);
nor U3747 (N_3747,N_3558,N_3553);
nor U3748 (N_3748,N_3408,N_3529);
or U3749 (N_3749,N_3452,N_3457);
and U3750 (N_3750,N_3456,N_3584);
nor U3751 (N_3751,N_3473,N_3556);
nor U3752 (N_3752,N_3520,N_3493);
or U3753 (N_3753,N_3537,N_3487);
and U3754 (N_3754,N_3539,N_3546);
or U3755 (N_3755,N_3448,N_3440);
and U3756 (N_3756,N_3470,N_3401);
and U3757 (N_3757,N_3470,N_3528);
nand U3758 (N_3758,N_3574,N_3583);
nor U3759 (N_3759,N_3512,N_3579);
nand U3760 (N_3760,N_3451,N_3523);
or U3761 (N_3761,N_3480,N_3511);
nor U3762 (N_3762,N_3514,N_3471);
and U3763 (N_3763,N_3496,N_3578);
nand U3764 (N_3764,N_3454,N_3475);
nand U3765 (N_3765,N_3508,N_3406);
nor U3766 (N_3766,N_3592,N_3402);
nand U3767 (N_3767,N_3557,N_3503);
nor U3768 (N_3768,N_3577,N_3525);
nand U3769 (N_3769,N_3458,N_3481);
xnor U3770 (N_3770,N_3525,N_3430);
nand U3771 (N_3771,N_3435,N_3452);
and U3772 (N_3772,N_3479,N_3483);
and U3773 (N_3773,N_3427,N_3527);
and U3774 (N_3774,N_3468,N_3551);
xor U3775 (N_3775,N_3461,N_3594);
or U3776 (N_3776,N_3549,N_3581);
or U3777 (N_3777,N_3534,N_3591);
or U3778 (N_3778,N_3411,N_3552);
xnor U3779 (N_3779,N_3599,N_3511);
nor U3780 (N_3780,N_3456,N_3480);
nand U3781 (N_3781,N_3547,N_3440);
or U3782 (N_3782,N_3486,N_3512);
and U3783 (N_3783,N_3551,N_3491);
and U3784 (N_3784,N_3444,N_3573);
and U3785 (N_3785,N_3545,N_3507);
nor U3786 (N_3786,N_3569,N_3597);
or U3787 (N_3787,N_3474,N_3564);
or U3788 (N_3788,N_3490,N_3582);
nor U3789 (N_3789,N_3459,N_3434);
xnor U3790 (N_3790,N_3535,N_3478);
and U3791 (N_3791,N_3570,N_3558);
and U3792 (N_3792,N_3550,N_3592);
nor U3793 (N_3793,N_3503,N_3402);
xor U3794 (N_3794,N_3576,N_3429);
nor U3795 (N_3795,N_3498,N_3445);
or U3796 (N_3796,N_3551,N_3466);
nor U3797 (N_3797,N_3584,N_3587);
or U3798 (N_3798,N_3416,N_3527);
xor U3799 (N_3799,N_3526,N_3569);
nand U3800 (N_3800,N_3712,N_3635);
and U3801 (N_3801,N_3778,N_3759);
nor U3802 (N_3802,N_3659,N_3715);
or U3803 (N_3803,N_3647,N_3682);
and U3804 (N_3804,N_3783,N_3733);
xor U3805 (N_3805,N_3771,N_3741);
or U3806 (N_3806,N_3615,N_3745);
or U3807 (N_3807,N_3793,N_3725);
nand U3808 (N_3808,N_3625,N_3760);
nand U3809 (N_3809,N_3763,N_3652);
nor U3810 (N_3810,N_3604,N_3797);
nor U3811 (N_3811,N_3665,N_3617);
xnor U3812 (N_3812,N_3714,N_3799);
or U3813 (N_3813,N_3656,N_3641);
xor U3814 (N_3814,N_3710,N_3628);
xor U3815 (N_3815,N_3614,N_3609);
nand U3816 (N_3816,N_3700,N_3648);
nand U3817 (N_3817,N_3692,N_3705);
and U3818 (N_3818,N_3776,N_3798);
or U3819 (N_3819,N_3777,N_3764);
nor U3820 (N_3820,N_3790,N_3761);
and U3821 (N_3821,N_3717,N_3616);
nor U3822 (N_3822,N_3681,N_3750);
or U3823 (N_3823,N_3689,N_3608);
or U3824 (N_3824,N_3758,N_3662);
or U3825 (N_3825,N_3651,N_3735);
nor U3826 (N_3826,N_3774,N_3637);
nor U3827 (N_3827,N_3630,N_3664);
xor U3828 (N_3828,N_3737,N_3785);
nand U3829 (N_3829,N_3698,N_3743);
xnor U3830 (N_3830,N_3666,N_3711);
nand U3831 (N_3831,N_3718,N_3685);
and U3832 (N_3832,N_3674,N_3749);
or U3833 (N_3833,N_3618,N_3694);
and U3834 (N_3834,N_3719,N_3629);
xor U3835 (N_3835,N_3697,N_3627);
or U3836 (N_3836,N_3748,N_3723);
nand U3837 (N_3837,N_3600,N_3732);
or U3838 (N_3838,N_3684,N_3702);
or U3839 (N_3839,N_3691,N_3730);
and U3840 (N_3840,N_3686,N_3706);
nor U3841 (N_3841,N_3756,N_3736);
and U3842 (N_3842,N_3680,N_3739);
or U3843 (N_3843,N_3645,N_3786);
nor U3844 (N_3844,N_3653,N_3727);
and U3845 (N_3845,N_3713,N_3738);
and U3846 (N_3846,N_3796,N_3678);
xor U3847 (N_3847,N_3658,N_3670);
nor U3848 (N_3848,N_3746,N_3729);
xnor U3849 (N_3849,N_3787,N_3757);
nor U3850 (N_3850,N_3636,N_3644);
xnor U3851 (N_3851,N_3650,N_3709);
or U3852 (N_3852,N_3769,N_3782);
and U3853 (N_3853,N_3649,N_3696);
nor U3854 (N_3854,N_3780,N_3695);
or U3855 (N_3855,N_3669,N_3707);
nand U3856 (N_3856,N_3671,N_3688);
and U3857 (N_3857,N_3704,N_3703);
nand U3858 (N_3858,N_3767,N_3667);
and U3859 (N_3859,N_3623,N_3701);
nand U3860 (N_3860,N_3765,N_3742);
nor U3861 (N_3861,N_3643,N_3744);
and U3862 (N_3862,N_3642,N_3753);
or U3863 (N_3863,N_3734,N_3654);
and U3864 (N_3864,N_3632,N_3721);
nor U3865 (N_3865,N_3646,N_3661);
or U3866 (N_3866,N_3601,N_3708);
nor U3867 (N_3867,N_3754,N_3775);
nor U3868 (N_3868,N_3794,N_3676);
nand U3869 (N_3869,N_3690,N_3619);
and U3870 (N_3870,N_3747,N_3766);
nand U3871 (N_3871,N_3795,N_3607);
nand U3872 (N_3872,N_3675,N_3687);
and U3873 (N_3873,N_3655,N_3621);
nand U3874 (N_3874,N_3626,N_3657);
xor U3875 (N_3875,N_3631,N_3699);
xor U3876 (N_3876,N_3693,N_3788);
and U3877 (N_3877,N_3603,N_3779);
and U3878 (N_3878,N_3639,N_3728);
and U3879 (N_3879,N_3622,N_3663);
and U3880 (N_3880,N_3740,N_3605);
and U3881 (N_3881,N_3731,N_3762);
or U3882 (N_3882,N_3724,N_3668);
nand U3883 (N_3883,N_3768,N_3640);
and U3884 (N_3884,N_3792,N_3716);
xnor U3885 (N_3885,N_3784,N_3770);
nand U3886 (N_3886,N_3755,N_3679);
and U3887 (N_3887,N_3751,N_3722);
xor U3888 (N_3888,N_3660,N_3606);
and U3889 (N_3889,N_3752,N_3683);
nand U3890 (N_3890,N_3613,N_3610);
nand U3891 (N_3891,N_3726,N_3624);
nand U3892 (N_3892,N_3677,N_3720);
or U3893 (N_3893,N_3772,N_3611);
or U3894 (N_3894,N_3620,N_3638);
nor U3895 (N_3895,N_3773,N_3673);
nor U3896 (N_3896,N_3633,N_3789);
nor U3897 (N_3897,N_3634,N_3781);
xnor U3898 (N_3898,N_3612,N_3672);
xnor U3899 (N_3899,N_3791,N_3602);
or U3900 (N_3900,N_3605,N_3627);
nor U3901 (N_3901,N_3690,N_3634);
nand U3902 (N_3902,N_3651,N_3682);
or U3903 (N_3903,N_3645,N_3725);
and U3904 (N_3904,N_3672,N_3794);
nand U3905 (N_3905,N_3623,N_3762);
xnor U3906 (N_3906,N_3770,N_3760);
nor U3907 (N_3907,N_3799,N_3726);
and U3908 (N_3908,N_3686,N_3637);
nor U3909 (N_3909,N_3656,N_3671);
or U3910 (N_3910,N_3648,N_3738);
xor U3911 (N_3911,N_3708,N_3685);
or U3912 (N_3912,N_3652,N_3630);
nand U3913 (N_3913,N_3634,N_3662);
and U3914 (N_3914,N_3693,N_3620);
and U3915 (N_3915,N_3652,N_3657);
xnor U3916 (N_3916,N_3645,N_3721);
or U3917 (N_3917,N_3714,N_3602);
nor U3918 (N_3918,N_3659,N_3649);
nand U3919 (N_3919,N_3733,N_3781);
nor U3920 (N_3920,N_3722,N_3784);
or U3921 (N_3921,N_3696,N_3746);
nand U3922 (N_3922,N_3795,N_3793);
or U3923 (N_3923,N_3797,N_3728);
and U3924 (N_3924,N_3677,N_3746);
nor U3925 (N_3925,N_3638,N_3696);
nand U3926 (N_3926,N_3695,N_3674);
nor U3927 (N_3927,N_3758,N_3608);
and U3928 (N_3928,N_3619,N_3665);
nand U3929 (N_3929,N_3606,N_3772);
nor U3930 (N_3930,N_3697,N_3720);
xnor U3931 (N_3931,N_3729,N_3624);
or U3932 (N_3932,N_3740,N_3766);
nand U3933 (N_3933,N_3683,N_3623);
nand U3934 (N_3934,N_3787,N_3797);
nor U3935 (N_3935,N_3672,N_3644);
or U3936 (N_3936,N_3627,N_3696);
or U3937 (N_3937,N_3693,N_3678);
and U3938 (N_3938,N_3762,N_3670);
or U3939 (N_3939,N_3665,N_3644);
and U3940 (N_3940,N_3638,N_3799);
nand U3941 (N_3941,N_3725,N_3651);
xor U3942 (N_3942,N_3795,N_3608);
and U3943 (N_3943,N_3763,N_3676);
nand U3944 (N_3944,N_3633,N_3765);
nand U3945 (N_3945,N_3726,N_3741);
or U3946 (N_3946,N_3651,N_3653);
nor U3947 (N_3947,N_3688,N_3669);
and U3948 (N_3948,N_3717,N_3649);
nand U3949 (N_3949,N_3632,N_3733);
nor U3950 (N_3950,N_3638,N_3628);
nand U3951 (N_3951,N_3619,N_3739);
nand U3952 (N_3952,N_3692,N_3778);
nand U3953 (N_3953,N_3799,N_3793);
nor U3954 (N_3954,N_3716,N_3715);
xnor U3955 (N_3955,N_3715,N_3790);
and U3956 (N_3956,N_3620,N_3661);
nand U3957 (N_3957,N_3702,N_3778);
nor U3958 (N_3958,N_3758,N_3711);
or U3959 (N_3959,N_3717,N_3709);
or U3960 (N_3960,N_3672,N_3662);
nor U3961 (N_3961,N_3631,N_3798);
xor U3962 (N_3962,N_3792,N_3656);
nand U3963 (N_3963,N_3746,N_3763);
xnor U3964 (N_3964,N_3797,N_3660);
nand U3965 (N_3965,N_3603,N_3772);
and U3966 (N_3966,N_3601,N_3765);
nor U3967 (N_3967,N_3670,N_3797);
nor U3968 (N_3968,N_3684,N_3676);
nand U3969 (N_3969,N_3609,N_3661);
or U3970 (N_3970,N_3775,N_3773);
or U3971 (N_3971,N_3649,N_3738);
and U3972 (N_3972,N_3702,N_3784);
nor U3973 (N_3973,N_3657,N_3628);
xnor U3974 (N_3974,N_3602,N_3752);
or U3975 (N_3975,N_3632,N_3628);
and U3976 (N_3976,N_3781,N_3629);
or U3977 (N_3977,N_3684,N_3628);
nor U3978 (N_3978,N_3683,N_3780);
xor U3979 (N_3979,N_3649,N_3628);
nand U3980 (N_3980,N_3731,N_3795);
and U3981 (N_3981,N_3683,N_3791);
xnor U3982 (N_3982,N_3774,N_3674);
or U3983 (N_3983,N_3610,N_3791);
nand U3984 (N_3984,N_3608,N_3708);
nor U3985 (N_3985,N_3700,N_3798);
and U3986 (N_3986,N_3636,N_3761);
nor U3987 (N_3987,N_3771,N_3680);
or U3988 (N_3988,N_3652,N_3626);
nor U3989 (N_3989,N_3726,N_3703);
or U3990 (N_3990,N_3734,N_3681);
xor U3991 (N_3991,N_3629,N_3732);
and U3992 (N_3992,N_3791,N_3666);
nor U3993 (N_3993,N_3765,N_3764);
xor U3994 (N_3994,N_3637,N_3723);
or U3995 (N_3995,N_3609,N_3788);
nand U3996 (N_3996,N_3645,N_3638);
nand U3997 (N_3997,N_3743,N_3711);
xnor U3998 (N_3998,N_3747,N_3635);
and U3999 (N_3999,N_3775,N_3684);
xor U4000 (N_4000,N_3834,N_3924);
nor U4001 (N_4001,N_3951,N_3848);
nor U4002 (N_4002,N_3965,N_3850);
and U4003 (N_4003,N_3856,N_3824);
and U4004 (N_4004,N_3933,N_3847);
nor U4005 (N_4005,N_3873,N_3859);
xnor U4006 (N_4006,N_3949,N_3872);
or U4007 (N_4007,N_3958,N_3808);
xor U4008 (N_4008,N_3820,N_3925);
or U4009 (N_4009,N_3912,N_3876);
nand U4010 (N_4010,N_3800,N_3815);
or U4011 (N_4011,N_3950,N_3962);
or U4012 (N_4012,N_3904,N_3978);
or U4013 (N_4013,N_3863,N_3897);
nor U4014 (N_4014,N_3898,N_3982);
nor U4015 (N_4015,N_3845,N_3999);
nor U4016 (N_4016,N_3987,N_3967);
nand U4017 (N_4017,N_3854,N_3988);
or U4018 (N_4018,N_3869,N_3959);
nor U4019 (N_4019,N_3915,N_3833);
xnor U4020 (N_4020,N_3812,N_3909);
nor U4021 (N_4021,N_3805,N_3953);
and U4022 (N_4022,N_3851,N_3963);
xor U4023 (N_4023,N_3899,N_3816);
xor U4024 (N_4024,N_3857,N_3846);
xor U4025 (N_4025,N_3998,N_3841);
or U4026 (N_4026,N_3893,N_3921);
xor U4027 (N_4027,N_3908,N_3989);
nor U4028 (N_4028,N_3985,N_3969);
xnor U4029 (N_4029,N_3906,N_3984);
xor U4030 (N_4030,N_3922,N_3870);
nand U4031 (N_4031,N_3896,N_3954);
nor U4032 (N_4032,N_3914,N_3943);
or U4033 (N_4033,N_3977,N_3844);
xnor U4034 (N_4034,N_3817,N_3952);
xnor U4035 (N_4035,N_3852,N_3849);
nor U4036 (N_4036,N_3973,N_3941);
or U4037 (N_4037,N_3936,N_3993);
nor U4038 (N_4038,N_3971,N_3990);
nor U4039 (N_4039,N_3911,N_3866);
nor U4040 (N_4040,N_3860,N_3884);
and U4041 (N_4041,N_3831,N_3992);
or U4042 (N_4042,N_3940,N_3858);
or U4043 (N_4043,N_3837,N_3995);
xor U4044 (N_4044,N_3881,N_3862);
xnor U4045 (N_4045,N_3901,N_3807);
xnor U4046 (N_4046,N_3835,N_3806);
nand U4047 (N_4047,N_3894,N_3905);
nor U4048 (N_4048,N_3916,N_3891);
nand U4049 (N_4049,N_3970,N_3811);
xor U4050 (N_4050,N_3827,N_3928);
nand U4051 (N_4051,N_3853,N_3926);
nand U4052 (N_4052,N_3983,N_3929);
nor U4053 (N_4053,N_3829,N_3980);
and U4054 (N_4054,N_3956,N_3828);
or U4055 (N_4055,N_3919,N_3935);
or U4056 (N_4056,N_3974,N_3875);
nand U4057 (N_4057,N_3832,N_3960);
xor U4058 (N_4058,N_3947,N_3887);
nor U4059 (N_4059,N_3937,N_3930);
or U4060 (N_4060,N_3920,N_3944);
xnor U4061 (N_4061,N_3902,N_3968);
nand U4062 (N_4062,N_3945,N_3927);
and U4063 (N_4063,N_3913,N_3810);
xor U4064 (N_4064,N_3839,N_3889);
nor U4065 (N_4065,N_3801,N_3964);
and U4066 (N_4066,N_3955,N_3886);
or U4067 (N_4067,N_3838,N_3809);
nand U4068 (N_4068,N_3802,N_3986);
nor U4069 (N_4069,N_3961,N_3907);
xor U4070 (N_4070,N_3991,N_3892);
and U4071 (N_4071,N_3934,N_3900);
xor U4072 (N_4072,N_3910,N_3877);
or U4073 (N_4073,N_3883,N_3903);
or U4074 (N_4074,N_3836,N_3996);
nor U4075 (N_4075,N_3868,N_3918);
nor U4076 (N_4076,N_3931,N_3994);
and U4077 (N_4077,N_3840,N_3979);
nor U4078 (N_4078,N_3946,N_3821);
or U4079 (N_4079,N_3923,N_3864);
and U4080 (N_4080,N_3972,N_3830);
or U4081 (N_4081,N_3938,N_3880);
nor U4082 (N_4082,N_3975,N_3890);
xnor U4083 (N_4083,N_3885,N_3976);
and U4084 (N_4084,N_3861,N_3855);
or U4085 (N_4085,N_3842,N_3867);
and U4086 (N_4086,N_3822,N_3843);
or U4087 (N_4087,N_3948,N_3957);
xor U4088 (N_4088,N_3814,N_3818);
nand U4089 (N_4089,N_3871,N_3997);
xnor U4090 (N_4090,N_3895,N_3826);
xor U4091 (N_4091,N_3888,N_3813);
and U4092 (N_4092,N_3804,N_3865);
nand U4093 (N_4093,N_3825,N_3981);
xor U4094 (N_4094,N_3878,N_3882);
or U4095 (N_4095,N_3966,N_3874);
xor U4096 (N_4096,N_3879,N_3917);
nor U4097 (N_4097,N_3823,N_3942);
xor U4098 (N_4098,N_3803,N_3819);
and U4099 (N_4099,N_3939,N_3932);
and U4100 (N_4100,N_3860,N_3875);
or U4101 (N_4101,N_3828,N_3973);
nor U4102 (N_4102,N_3910,N_3920);
xnor U4103 (N_4103,N_3984,N_3853);
or U4104 (N_4104,N_3833,N_3853);
nor U4105 (N_4105,N_3894,N_3878);
and U4106 (N_4106,N_3946,N_3847);
nand U4107 (N_4107,N_3880,N_3990);
and U4108 (N_4108,N_3960,N_3927);
nor U4109 (N_4109,N_3876,N_3832);
or U4110 (N_4110,N_3918,N_3858);
nand U4111 (N_4111,N_3858,N_3990);
nor U4112 (N_4112,N_3858,N_3959);
or U4113 (N_4113,N_3915,N_3800);
nand U4114 (N_4114,N_3971,N_3912);
nand U4115 (N_4115,N_3934,N_3992);
xor U4116 (N_4116,N_3959,N_3829);
nand U4117 (N_4117,N_3870,N_3843);
nor U4118 (N_4118,N_3833,N_3992);
nand U4119 (N_4119,N_3967,N_3860);
or U4120 (N_4120,N_3827,N_3854);
xor U4121 (N_4121,N_3935,N_3924);
xnor U4122 (N_4122,N_3921,N_3945);
and U4123 (N_4123,N_3836,N_3869);
or U4124 (N_4124,N_3900,N_3983);
and U4125 (N_4125,N_3816,N_3916);
nor U4126 (N_4126,N_3920,N_3876);
or U4127 (N_4127,N_3983,N_3906);
nor U4128 (N_4128,N_3836,N_3811);
nor U4129 (N_4129,N_3861,N_3825);
nor U4130 (N_4130,N_3875,N_3924);
or U4131 (N_4131,N_3839,N_3946);
or U4132 (N_4132,N_3896,N_3871);
and U4133 (N_4133,N_3924,N_3891);
or U4134 (N_4134,N_3969,N_3875);
or U4135 (N_4135,N_3867,N_3955);
nand U4136 (N_4136,N_3827,N_3817);
nor U4137 (N_4137,N_3876,N_3805);
and U4138 (N_4138,N_3880,N_3848);
nor U4139 (N_4139,N_3839,N_3903);
nand U4140 (N_4140,N_3842,N_3837);
or U4141 (N_4141,N_3909,N_3963);
xnor U4142 (N_4142,N_3876,N_3906);
nand U4143 (N_4143,N_3920,N_3837);
nand U4144 (N_4144,N_3865,N_3908);
nor U4145 (N_4145,N_3876,N_3999);
nor U4146 (N_4146,N_3839,N_3842);
nor U4147 (N_4147,N_3802,N_3999);
or U4148 (N_4148,N_3829,N_3988);
and U4149 (N_4149,N_3949,N_3839);
nor U4150 (N_4150,N_3896,N_3876);
nand U4151 (N_4151,N_3970,N_3827);
nor U4152 (N_4152,N_3883,N_3860);
nor U4153 (N_4153,N_3881,N_3816);
xnor U4154 (N_4154,N_3975,N_3982);
and U4155 (N_4155,N_3841,N_3840);
xor U4156 (N_4156,N_3966,N_3979);
xor U4157 (N_4157,N_3988,N_3825);
nor U4158 (N_4158,N_3905,N_3832);
or U4159 (N_4159,N_3919,N_3869);
nor U4160 (N_4160,N_3835,N_3983);
or U4161 (N_4161,N_3938,N_3851);
xor U4162 (N_4162,N_3847,N_3835);
or U4163 (N_4163,N_3800,N_3943);
xnor U4164 (N_4164,N_3888,N_3934);
or U4165 (N_4165,N_3891,N_3935);
xor U4166 (N_4166,N_3817,N_3847);
and U4167 (N_4167,N_3835,N_3845);
and U4168 (N_4168,N_3976,N_3982);
nand U4169 (N_4169,N_3960,N_3995);
or U4170 (N_4170,N_3923,N_3993);
nand U4171 (N_4171,N_3896,N_3826);
and U4172 (N_4172,N_3858,N_3873);
or U4173 (N_4173,N_3893,N_3915);
or U4174 (N_4174,N_3997,N_3848);
xor U4175 (N_4175,N_3941,N_3923);
and U4176 (N_4176,N_3878,N_3935);
nand U4177 (N_4177,N_3881,N_3833);
nand U4178 (N_4178,N_3907,N_3900);
nor U4179 (N_4179,N_3858,N_3899);
nand U4180 (N_4180,N_3886,N_3823);
or U4181 (N_4181,N_3830,N_3968);
or U4182 (N_4182,N_3828,N_3949);
nand U4183 (N_4183,N_3846,N_3900);
or U4184 (N_4184,N_3803,N_3844);
nor U4185 (N_4185,N_3950,N_3805);
and U4186 (N_4186,N_3850,N_3984);
nor U4187 (N_4187,N_3896,N_3811);
xor U4188 (N_4188,N_3874,N_3945);
or U4189 (N_4189,N_3929,N_3938);
nand U4190 (N_4190,N_3967,N_3946);
nand U4191 (N_4191,N_3830,N_3977);
or U4192 (N_4192,N_3949,N_3986);
or U4193 (N_4193,N_3996,N_3986);
nor U4194 (N_4194,N_3901,N_3903);
nor U4195 (N_4195,N_3987,N_3990);
or U4196 (N_4196,N_3893,N_3931);
and U4197 (N_4197,N_3970,N_3847);
nor U4198 (N_4198,N_3862,N_3934);
xor U4199 (N_4199,N_3993,N_3880);
xnor U4200 (N_4200,N_4124,N_4188);
nand U4201 (N_4201,N_4134,N_4015);
nor U4202 (N_4202,N_4114,N_4049);
and U4203 (N_4203,N_4141,N_4166);
or U4204 (N_4204,N_4099,N_4098);
nand U4205 (N_4205,N_4061,N_4018);
nor U4206 (N_4206,N_4131,N_4145);
or U4207 (N_4207,N_4170,N_4169);
nand U4208 (N_4208,N_4168,N_4122);
nand U4209 (N_4209,N_4123,N_4075);
or U4210 (N_4210,N_4133,N_4156);
nor U4211 (N_4211,N_4062,N_4160);
xor U4212 (N_4212,N_4086,N_4077);
xnor U4213 (N_4213,N_4095,N_4130);
nand U4214 (N_4214,N_4029,N_4017);
or U4215 (N_4215,N_4147,N_4157);
or U4216 (N_4216,N_4172,N_4076);
nand U4217 (N_4217,N_4078,N_4022);
and U4218 (N_4218,N_4135,N_4041);
nor U4219 (N_4219,N_4126,N_4071);
nand U4220 (N_4220,N_4033,N_4034);
nor U4221 (N_4221,N_4199,N_4132);
and U4222 (N_4222,N_4107,N_4092);
nand U4223 (N_4223,N_4119,N_4009);
and U4224 (N_4224,N_4084,N_4103);
and U4225 (N_4225,N_4091,N_4138);
and U4226 (N_4226,N_4043,N_4198);
or U4227 (N_4227,N_4026,N_4180);
or U4228 (N_4228,N_4111,N_4035);
xor U4229 (N_4229,N_4096,N_4072);
or U4230 (N_4230,N_4105,N_4008);
nand U4231 (N_4231,N_4151,N_4193);
xor U4232 (N_4232,N_4142,N_4044);
or U4233 (N_4233,N_4149,N_4000);
xnor U4234 (N_4234,N_4176,N_4191);
xnor U4235 (N_4235,N_4177,N_4150);
nand U4236 (N_4236,N_4113,N_4056);
or U4237 (N_4237,N_4154,N_4004);
or U4238 (N_4238,N_4137,N_4182);
xnor U4239 (N_4239,N_4139,N_4031);
xor U4240 (N_4240,N_4070,N_4187);
nand U4241 (N_4241,N_4185,N_4047);
or U4242 (N_4242,N_4059,N_4081);
nand U4243 (N_4243,N_4128,N_4069);
xnor U4244 (N_4244,N_4010,N_4073);
xor U4245 (N_4245,N_4067,N_4194);
and U4246 (N_4246,N_4163,N_4184);
nor U4247 (N_4247,N_4014,N_4110);
xnor U4248 (N_4248,N_4055,N_4115);
nand U4249 (N_4249,N_4129,N_4020);
and U4250 (N_4250,N_4016,N_4087);
or U4251 (N_4251,N_4167,N_4097);
nor U4252 (N_4252,N_4025,N_4165);
or U4253 (N_4253,N_4024,N_4012);
xor U4254 (N_4254,N_4053,N_4011);
nand U4255 (N_4255,N_4036,N_4100);
nor U4256 (N_4256,N_4155,N_4195);
nand U4257 (N_4257,N_4040,N_4117);
xnor U4258 (N_4258,N_4052,N_4063);
or U4259 (N_4259,N_4136,N_4179);
and U4260 (N_4260,N_4183,N_4125);
nand U4261 (N_4261,N_4046,N_4102);
or U4262 (N_4262,N_4007,N_4057);
and U4263 (N_4263,N_4197,N_4003);
nor U4264 (N_4264,N_4094,N_4083);
or U4265 (N_4265,N_4032,N_4152);
and U4266 (N_4266,N_4173,N_4048);
or U4267 (N_4267,N_4108,N_4112);
nor U4268 (N_4268,N_4101,N_4079);
xnor U4269 (N_4269,N_4190,N_4181);
xor U4270 (N_4270,N_4002,N_4064);
xnor U4271 (N_4271,N_4192,N_4085);
or U4272 (N_4272,N_4065,N_4058);
and U4273 (N_4273,N_4127,N_4178);
nand U4274 (N_4274,N_4045,N_4189);
or U4275 (N_4275,N_4120,N_4104);
or U4276 (N_4276,N_4143,N_4001);
xor U4277 (N_4277,N_4066,N_4196);
or U4278 (N_4278,N_4121,N_4038);
xnor U4279 (N_4279,N_4023,N_4148);
nor U4280 (N_4280,N_4116,N_4164);
nor U4281 (N_4281,N_4118,N_4042);
or U4282 (N_4282,N_4060,N_4021);
xnor U4283 (N_4283,N_4090,N_4186);
nor U4284 (N_4284,N_4089,N_4039);
xor U4285 (N_4285,N_4037,N_4005);
nor U4286 (N_4286,N_4082,N_4074);
nand U4287 (N_4287,N_4159,N_4068);
or U4288 (N_4288,N_4028,N_4175);
or U4289 (N_4289,N_4027,N_4106);
nand U4290 (N_4290,N_4019,N_4161);
nor U4291 (N_4291,N_4171,N_4013);
or U4292 (N_4292,N_4174,N_4054);
and U4293 (N_4293,N_4109,N_4162);
xor U4294 (N_4294,N_4030,N_4088);
and U4295 (N_4295,N_4158,N_4051);
xor U4296 (N_4296,N_4050,N_4140);
or U4297 (N_4297,N_4080,N_4153);
nand U4298 (N_4298,N_4006,N_4144);
nor U4299 (N_4299,N_4093,N_4146);
xor U4300 (N_4300,N_4065,N_4106);
or U4301 (N_4301,N_4027,N_4192);
or U4302 (N_4302,N_4010,N_4128);
and U4303 (N_4303,N_4013,N_4022);
or U4304 (N_4304,N_4048,N_4077);
and U4305 (N_4305,N_4188,N_4076);
xor U4306 (N_4306,N_4045,N_4095);
xnor U4307 (N_4307,N_4080,N_4012);
nor U4308 (N_4308,N_4070,N_4167);
and U4309 (N_4309,N_4195,N_4145);
nand U4310 (N_4310,N_4171,N_4184);
nand U4311 (N_4311,N_4145,N_4130);
nor U4312 (N_4312,N_4013,N_4001);
xnor U4313 (N_4313,N_4178,N_4126);
and U4314 (N_4314,N_4092,N_4088);
and U4315 (N_4315,N_4041,N_4195);
nor U4316 (N_4316,N_4038,N_4189);
and U4317 (N_4317,N_4125,N_4190);
and U4318 (N_4318,N_4189,N_4057);
or U4319 (N_4319,N_4055,N_4060);
xnor U4320 (N_4320,N_4093,N_4074);
nand U4321 (N_4321,N_4166,N_4061);
or U4322 (N_4322,N_4009,N_4162);
or U4323 (N_4323,N_4192,N_4196);
and U4324 (N_4324,N_4120,N_4168);
nand U4325 (N_4325,N_4163,N_4054);
xor U4326 (N_4326,N_4165,N_4008);
xor U4327 (N_4327,N_4191,N_4097);
xnor U4328 (N_4328,N_4080,N_4077);
nand U4329 (N_4329,N_4018,N_4121);
or U4330 (N_4330,N_4082,N_4142);
nand U4331 (N_4331,N_4116,N_4100);
nor U4332 (N_4332,N_4174,N_4104);
and U4333 (N_4333,N_4145,N_4108);
and U4334 (N_4334,N_4081,N_4020);
nor U4335 (N_4335,N_4122,N_4162);
nor U4336 (N_4336,N_4167,N_4058);
nand U4337 (N_4337,N_4095,N_4149);
and U4338 (N_4338,N_4113,N_4061);
xor U4339 (N_4339,N_4181,N_4031);
or U4340 (N_4340,N_4002,N_4074);
nor U4341 (N_4341,N_4083,N_4072);
xnor U4342 (N_4342,N_4068,N_4081);
nand U4343 (N_4343,N_4084,N_4066);
or U4344 (N_4344,N_4066,N_4187);
xor U4345 (N_4345,N_4163,N_4090);
xor U4346 (N_4346,N_4171,N_4172);
xnor U4347 (N_4347,N_4113,N_4006);
and U4348 (N_4348,N_4169,N_4047);
xor U4349 (N_4349,N_4021,N_4124);
nor U4350 (N_4350,N_4182,N_4092);
and U4351 (N_4351,N_4019,N_4040);
xor U4352 (N_4352,N_4183,N_4059);
nor U4353 (N_4353,N_4014,N_4048);
or U4354 (N_4354,N_4044,N_4138);
xor U4355 (N_4355,N_4040,N_4070);
nor U4356 (N_4356,N_4048,N_4178);
and U4357 (N_4357,N_4019,N_4192);
and U4358 (N_4358,N_4196,N_4005);
xor U4359 (N_4359,N_4109,N_4065);
nand U4360 (N_4360,N_4048,N_4065);
nand U4361 (N_4361,N_4120,N_4190);
or U4362 (N_4362,N_4148,N_4099);
nand U4363 (N_4363,N_4094,N_4086);
nand U4364 (N_4364,N_4024,N_4090);
nor U4365 (N_4365,N_4006,N_4022);
and U4366 (N_4366,N_4197,N_4014);
and U4367 (N_4367,N_4171,N_4127);
and U4368 (N_4368,N_4079,N_4075);
xor U4369 (N_4369,N_4120,N_4024);
xnor U4370 (N_4370,N_4024,N_4151);
and U4371 (N_4371,N_4024,N_4133);
xnor U4372 (N_4372,N_4077,N_4144);
or U4373 (N_4373,N_4027,N_4061);
nand U4374 (N_4374,N_4141,N_4129);
and U4375 (N_4375,N_4174,N_4180);
nand U4376 (N_4376,N_4178,N_4009);
xnor U4377 (N_4377,N_4102,N_4180);
or U4378 (N_4378,N_4115,N_4117);
nand U4379 (N_4379,N_4122,N_4115);
and U4380 (N_4380,N_4096,N_4111);
nand U4381 (N_4381,N_4130,N_4115);
nand U4382 (N_4382,N_4137,N_4156);
nand U4383 (N_4383,N_4088,N_4135);
nand U4384 (N_4384,N_4007,N_4109);
or U4385 (N_4385,N_4185,N_4118);
nor U4386 (N_4386,N_4114,N_4014);
and U4387 (N_4387,N_4117,N_4041);
nor U4388 (N_4388,N_4061,N_4194);
xnor U4389 (N_4389,N_4144,N_4053);
xor U4390 (N_4390,N_4191,N_4196);
and U4391 (N_4391,N_4165,N_4075);
nand U4392 (N_4392,N_4121,N_4167);
nand U4393 (N_4393,N_4162,N_4176);
nand U4394 (N_4394,N_4132,N_4120);
or U4395 (N_4395,N_4139,N_4083);
nor U4396 (N_4396,N_4142,N_4181);
xnor U4397 (N_4397,N_4049,N_4019);
or U4398 (N_4398,N_4054,N_4001);
nand U4399 (N_4399,N_4082,N_4009);
xnor U4400 (N_4400,N_4327,N_4323);
and U4401 (N_4401,N_4289,N_4380);
or U4402 (N_4402,N_4347,N_4311);
nand U4403 (N_4403,N_4325,N_4271);
xor U4404 (N_4404,N_4256,N_4317);
and U4405 (N_4405,N_4268,N_4227);
nor U4406 (N_4406,N_4370,N_4288);
or U4407 (N_4407,N_4331,N_4388);
and U4408 (N_4408,N_4368,N_4326);
nand U4409 (N_4409,N_4304,N_4374);
nand U4410 (N_4410,N_4309,N_4366);
nand U4411 (N_4411,N_4228,N_4232);
nand U4412 (N_4412,N_4329,N_4299);
or U4413 (N_4413,N_4298,N_4343);
xnor U4414 (N_4414,N_4348,N_4360);
and U4415 (N_4415,N_4395,N_4376);
or U4416 (N_4416,N_4259,N_4276);
and U4417 (N_4417,N_4332,N_4242);
nor U4418 (N_4418,N_4231,N_4245);
xnor U4419 (N_4419,N_4350,N_4312);
nand U4420 (N_4420,N_4291,N_4226);
or U4421 (N_4421,N_4212,N_4274);
xnor U4422 (N_4422,N_4210,N_4377);
nand U4423 (N_4423,N_4363,N_4253);
and U4424 (N_4424,N_4303,N_4292);
and U4425 (N_4425,N_4225,N_4319);
nor U4426 (N_4426,N_4270,N_4398);
nor U4427 (N_4427,N_4254,N_4399);
xor U4428 (N_4428,N_4364,N_4346);
nor U4429 (N_4429,N_4279,N_4387);
and U4430 (N_4430,N_4344,N_4273);
and U4431 (N_4431,N_4248,N_4308);
nor U4432 (N_4432,N_4310,N_4294);
or U4433 (N_4433,N_4251,N_4320);
xnor U4434 (N_4434,N_4287,N_4204);
or U4435 (N_4435,N_4339,N_4391);
or U4436 (N_4436,N_4240,N_4397);
nor U4437 (N_4437,N_4338,N_4223);
or U4438 (N_4438,N_4229,N_4283);
nor U4439 (N_4439,N_4324,N_4306);
and U4440 (N_4440,N_4355,N_4341);
xnor U4441 (N_4441,N_4238,N_4255);
nor U4442 (N_4442,N_4384,N_4373);
nor U4443 (N_4443,N_4237,N_4233);
or U4444 (N_4444,N_4284,N_4278);
nand U4445 (N_4445,N_4342,N_4390);
or U4446 (N_4446,N_4275,N_4205);
and U4447 (N_4447,N_4266,N_4315);
nand U4448 (N_4448,N_4379,N_4285);
nor U4449 (N_4449,N_4215,N_4230);
or U4450 (N_4450,N_4345,N_4280);
nand U4451 (N_4451,N_4220,N_4356);
or U4452 (N_4452,N_4260,N_4200);
or U4453 (N_4453,N_4206,N_4293);
nor U4454 (N_4454,N_4297,N_4241);
and U4455 (N_4455,N_4396,N_4265);
nand U4456 (N_4456,N_4340,N_4333);
nand U4457 (N_4457,N_4336,N_4239);
or U4458 (N_4458,N_4357,N_4316);
xnor U4459 (N_4459,N_4282,N_4286);
xor U4460 (N_4460,N_4349,N_4330);
nor U4461 (N_4461,N_4321,N_4246);
xor U4462 (N_4462,N_4257,N_4381);
or U4463 (N_4463,N_4378,N_4362);
xnor U4464 (N_4464,N_4337,N_4249);
and U4465 (N_4465,N_4277,N_4263);
or U4466 (N_4466,N_4328,N_4236);
or U4467 (N_4467,N_4361,N_4234);
xor U4468 (N_4468,N_4371,N_4353);
nand U4469 (N_4469,N_4258,N_4267);
or U4470 (N_4470,N_4208,N_4252);
and U4471 (N_4471,N_4217,N_4243);
nand U4472 (N_4472,N_4375,N_4365);
xor U4473 (N_4473,N_4367,N_4358);
and U4474 (N_4474,N_4269,N_4209);
and U4475 (N_4475,N_4392,N_4305);
xnor U4476 (N_4476,N_4302,N_4313);
or U4477 (N_4477,N_4222,N_4221);
and U4478 (N_4478,N_4322,N_4264);
and U4479 (N_4479,N_4383,N_4207);
nor U4480 (N_4480,N_4295,N_4261);
nand U4481 (N_4481,N_4213,N_4250);
or U4482 (N_4482,N_4334,N_4262);
xor U4483 (N_4483,N_4218,N_4352);
and U4484 (N_4484,N_4394,N_4318);
nor U4485 (N_4485,N_4385,N_4281);
xor U4486 (N_4486,N_4211,N_4389);
and U4487 (N_4487,N_4301,N_4372);
nand U4488 (N_4488,N_4202,N_4386);
nor U4489 (N_4489,N_4235,N_4351);
or U4490 (N_4490,N_4314,N_4247);
xnor U4491 (N_4491,N_4201,N_4354);
nand U4492 (N_4492,N_4300,N_4296);
nor U4493 (N_4493,N_4369,N_4290);
or U4494 (N_4494,N_4244,N_4393);
and U4495 (N_4495,N_4307,N_4203);
xor U4496 (N_4496,N_4214,N_4219);
nor U4497 (N_4497,N_4359,N_4224);
xor U4498 (N_4498,N_4216,N_4382);
and U4499 (N_4499,N_4335,N_4272);
xnor U4500 (N_4500,N_4377,N_4248);
nand U4501 (N_4501,N_4227,N_4250);
nor U4502 (N_4502,N_4309,N_4350);
xor U4503 (N_4503,N_4248,N_4224);
and U4504 (N_4504,N_4356,N_4286);
and U4505 (N_4505,N_4311,N_4255);
nand U4506 (N_4506,N_4249,N_4242);
xor U4507 (N_4507,N_4363,N_4316);
or U4508 (N_4508,N_4383,N_4235);
and U4509 (N_4509,N_4241,N_4201);
and U4510 (N_4510,N_4250,N_4284);
nand U4511 (N_4511,N_4331,N_4307);
nor U4512 (N_4512,N_4207,N_4386);
nor U4513 (N_4513,N_4339,N_4241);
and U4514 (N_4514,N_4371,N_4332);
or U4515 (N_4515,N_4383,N_4294);
and U4516 (N_4516,N_4236,N_4362);
nor U4517 (N_4517,N_4225,N_4310);
or U4518 (N_4518,N_4220,N_4202);
and U4519 (N_4519,N_4224,N_4382);
or U4520 (N_4520,N_4225,N_4328);
or U4521 (N_4521,N_4386,N_4281);
nor U4522 (N_4522,N_4369,N_4391);
or U4523 (N_4523,N_4299,N_4390);
or U4524 (N_4524,N_4350,N_4261);
nand U4525 (N_4525,N_4208,N_4329);
or U4526 (N_4526,N_4204,N_4264);
xor U4527 (N_4527,N_4231,N_4267);
xor U4528 (N_4528,N_4264,N_4368);
and U4529 (N_4529,N_4393,N_4346);
nand U4530 (N_4530,N_4214,N_4244);
nor U4531 (N_4531,N_4320,N_4344);
xor U4532 (N_4532,N_4309,N_4267);
and U4533 (N_4533,N_4399,N_4369);
and U4534 (N_4534,N_4234,N_4388);
nor U4535 (N_4535,N_4277,N_4369);
nand U4536 (N_4536,N_4236,N_4293);
and U4537 (N_4537,N_4272,N_4249);
nand U4538 (N_4538,N_4332,N_4359);
or U4539 (N_4539,N_4237,N_4219);
nand U4540 (N_4540,N_4370,N_4248);
nand U4541 (N_4541,N_4341,N_4390);
xor U4542 (N_4542,N_4374,N_4256);
nor U4543 (N_4543,N_4305,N_4317);
xnor U4544 (N_4544,N_4397,N_4224);
xnor U4545 (N_4545,N_4248,N_4331);
nand U4546 (N_4546,N_4335,N_4396);
and U4547 (N_4547,N_4219,N_4343);
xor U4548 (N_4548,N_4233,N_4375);
or U4549 (N_4549,N_4272,N_4228);
xor U4550 (N_4550,N_4314,N_4387);
nand U4551 (N_4551,N_4398,N_4314);
and U4552 (N_4552,N_4301,N_4365);
nand U4553 (N_4553,N_4342,N_4297);
xor U4554 (N_4554,N_4302,N_4299);
nor U4555 (N_4555,N_4223,N_4323);
xnor U4556 (N_4556,N_4265,N_4373);
or U4557 (N_4557,N_4338,N_4302);
and U4558 (N_4558,N_4292,N_4250);
xnor U4559 (N_4559,N_4229,N_4375);
or U4560 (N_4560,N_4282,N_4258);
nor U4561 (N_4561,N_4225,N_4366);
xnor U4562 (N_4562,N_4344,N_4294);
nand U4563 (N_4563,N_4277,N_4345);
xnor U4564 (N_4564,N_4310,N_4296);
nand U4565 (N_4565,N_4320,N_4306);
xnor U4566 (N_4566,N_4240,N_4390);
nor U4567 (N_4567,N_4225,N_4270);
or U4568 (N_4568,N_4372,N_4398);
or U4569 (N_4569,N_4204,N_4340);
nor U4570 (N_4570,N_4319,N_4257);
nor U4571 (N_4571,N_4265,N_4366);
or U4572 (N_4572,N_4270,N_4396);
xnor U4573 (N_4573,N_4297,N_4380);
xor U4574 (N_4574,N_4270,N_4325);
xor U4575 (N_4575,N_4397,N_4266);
nand U4576 (N_4576,N_4285,N_4385);
nor U4577 (N_4577,N_4373,N_4335);
or U4578 (N_4578,N_4225,N_4239);
or U4579 (N_4579,N_4382,N_4325);
nor U4580 (N_4580,N_4314,N_4351);
or U4581 (N_4581,N_4228,N_4282);
and U4582 (N_4582,N_4364,N_4347);
and U4583 (N_4583,N_4349,N_4245);
nand U4584 (N_4584,N_4253,N_4202);
or U4585 (N_4585,N_4275,N_4294);
xor U4586 (N_4586,N_4247,N_4347);
nand U4587 (N_4587,N_4242,N_4213);
xnor U4588 (N_4588,N_4329,N_4281);
or U4589 (N_4589,N_4207,N_4232);
nand U4590 (N_4590,N_4380,N_4326);
nor U4591 (N_4591,N_4354,N_4267);
xor U4592 (N_4592,N_4335,N_4345);
and U4593 (N_4593,N_4226,N_4300);
and U4594 (N_4594,N_4237,N_4298);
nor U4595 (N_4595,N_4303,N_4250);
nand U4596 (N_4596,N_4371,N_4220);
and U4597 (N_4597,N_4359,N_4312);
xor U4598 (N_4598,N_4287,N_4357);
and U4599 (N_4599,N_4320,N_4378);
or U4600 (N_4600,N_4442,N_4445);
and U4601 (N_4601,N_4583,N_4546);
nand U4602 (N_4602,N_4475,N_4540);
xor U4603 (N_4603,N_4531,N_4432);
nor U4604 (N_4604,N_4434,N_4514);
and U4605 (N_4605,N_4482,N_4408);
or U4606 (N_4606,N_4576,N_4456);
xnor U4607 (N_4607,N_4595,N_4566);
and U4608 (N_4608,N_4509,N_4458);
or U4609 (N_4609,N_4452,N_4515);
nand U4610 (N_4610,N_4589,N_4469);
and U4611 (N_4611,N_4429,N_4501);
nor U4612 (N_4612,N_4507,N_4426);
and U4613 (N_4613,N_4460,N_4544);
or U4614 (N_4614,N_4403,N_4559);
and U4615 (N_4615,N_4440,N_4573);
or U4616 (N_4616,N_4499,N_4543);
xor U4617 (N_4617,N_4541,N_4539);
nor U4618 (N_4618,N_4565,N_4579);
nor U4619 (N_4619,N_4532,N_4560);
and U4620 (N_4620,N_4570,N_4446);
nand U4621 (N_4621,N_4506,N_4520);
nand U4622 (N_4622,N_4451,N_4468);
and U4623 (N_4623,N_4585,N_4465);
or U4624 (N_4624,N_4530,N_4455);
nor U4625 (N_4625,N_4572,N_4502);
and U4626 (N_4626,N_4419,N_4400);
xor U4627 (N_4627,N_4487,N_4443);
xnor U4628 (N_4628,N_4441,N_4587);
nor U4629 (N_4629,N_4497,N_4527);
nand U4630 (N_4630,N_4417,N_4411);
or U4631 (N_4631,N_4597,N_4479);
and U4632 (N_4632,N_4554,N_4457);
nand U4633 (N_4633,N_4553,N_4427);
xnor U4634 (N_4634,N_4536,N_4568);
xnor U4635 (N_4635,N_4563,N_4519);
xor U4636 (N_4636,N_4537,N_4581);
or U4637 (N_4637,N_4569,N_4490);
xor U4638 (N_4638,N_4409,N_4438);
nor U4639 (N_4639,N_4462,N_4582);
or U4640 (N_4640,N_4418,N_4511);
and U4641 (N_4641,N_4454,N_4574);
nand U4642 (N_4642,N_4447,N_4557);
nor U4643 (N_4643,N_4421,N_4464);
nand U4644 (N_4644,N_4472,N_4406);
and U4645 (N_4645,N_4513,N_4430);
nor U4646 (N_4646,N_4594,N_4584);
or U4647 (N_4647,N_4538,N_4503);
nand U4648 (N_4648,N_4521,N_4550);
nand U4649 (N_4649,N_4575,N_4510);
or U4650 (N_4650,N_4470,N_4598);
nor U4651 (N_4651,N_4486,N_4410);
xnor U4652 (N_4652,N_4593,N_4422);
and U4653 (N_4653,N_4552,N_4525);
nand U4654 (N_4654,N_4562,N_4523);
and U4655 (N_4655,N_4590,N_4596);
nor U4656 (N_4656,N_4444,N_4526);
nand U4657 (N_4657,N_4558,N_4498);
or U4658 (N_4658,N_4548,N_4413);
and U4659 (N_4659,N_4533,N_4555);
and U4660 (N_4660,N_4453,N_4588);
and U4661 (N_4661,N_4571,N_4524);
nand U4662 (N_4662,N_4450,N_4578);
nand U4663 (N_4663,N_4528,N_4437);
xor U4664 (N_4664,N_4476,N_4481);
xor U4665 (N_4665,N_4489,N_4529);
nor U4666 (N_4666,N_4478,N_4549);
nor U4667 (N_4667,N_4488,N_4477);
xnor U4668 (N_4668,N_4586,N_4404);
and U4669 (N_4669,N_4547,N_4480);
xnor U4670 (N_4670,N_4551,N_4577);
and U4671 (N_4671,N_4580,N_4518);
nor U4672 (N_4672,N_4431,N_4407);
and U4673 (N_4673,N_4491,N_4415);
nor U4674 (N_4674,N_4504,N_4401);
nor U4675 (N_4675,N_4516,N_4599);
or U4676 (N_4676,N_4428,N_4500);
nand U4677 (N_4677,N_4436,N_4591);
or U4678 (N_4678,N_4423,N_4414);
xnor U4679 (N_4679,N_4485,N_4412);
or U4680 (N_4680,N_4534,N_4435);
nor U4681 (N_4681,N_4512,N_4439);
and U4682 (N_4682,N_4561,N_4466);
or U4683 (N_4683,N_4433,N_4473);
nor U4684 (N_4684,N_4492,N_4420);
or U4685 (N_4685,N_4493,N_4424);
and U4686 (N_4686,N_4517,N_4564);
xnor U4687 (N_4687,N_4495,N_4449);
or U4688 (N_4688,N_4467,N_4545);
xnor U4689 (N_4689,N_4463,N_4484);
or U4690 (N_4690,N_4461,N_4416);
nand U4691 (N_4691,N_4505,N_4448);
nor U4692 (N_4692,N_4459,N_4483);
or U4693 (N_4693,N_4508,N_4556);
or U4694 (N_4694,N_4535,N_4471);
and U4695 (N_4695,N_4425,N_4542);
nor U4696 (N_4696,N_4522,N_4405);
or U4697 (N_4697,N_4474,N_4494);
or U4698 (N_4698,N_4592,N_4496);
nor U4699 (N_4699,N_4567,N_4402);
nor U4700 (N_4700,N_4450,N_4423);
nor U4701 (N_4701,N_4565,N_4513);
and U4702 (N_4702,N_4522,N_4447);
xor U4703 (N_4703,N_4461,N_4578);
or U4704 (N_4704,N_4477,N_4588);
or U4705 (N_4705,N_4522,N_4472);
nor U4706 (N_4706,N_4527,N_4496);
nand U4707 (N_4707,N_4490,N_4548);
nor U4708 (N_4708,N_4599,N_4532);
nand U4709 (N_4709,N_4544,N_4487);
nand U4710 (N_4710,N_4510,N_4451);
or U4711 (N_4711,N_4579,N_4401);
and U4712 (N_4712,N_4520,N_4507);
nor U4713 (N_4713,N_4457,N_4517);
nor U4714 (N_4714,N_4439,N_4567);
and U4715 (N_4715,N_4570,N_4502);
nand U4716 (N_4716,N_4425,N_4448);
nor U4717 (N_4717,N_4426,N_4577);
nand U4718 (N_4718,N_4582,N_4551);
or U4719 (N_4719,N_4515,N_4527);
xor U4720 (N_4720,N_4584,N_4492);
xor U4721 (N_4721,N_4457,N_4598);
xor U4722 (N_4722,N_4426,N_4405);
and U4723 (N_4723,N_4547,N_4453);
nand U4724 (N_4724,N_4464,N_4572);
nand U4725 (N_4725,N_4486,N_4415);
xor U4726 (N_4726,N_4442,N_4561);
xnor U4727 (N_4727,N_4463,N_4578);
nor U4728 (N_4728,N_4494,N_4408);
or U4729 (N_4729,N_4527,N_4548);
nor U4730 (N_4730,N_4402,N_4563);
or U4731 (N_4731,N_4517,N_4430);
or U4732 (N_4732,N_4483,N_4570);
or U4733 (N_4733,N_4447,N_4520);
and U4734 (N_4734,N_4559,N_4591);
nand U4735 (N_4735,N_4416,N_4470);
nand U4736 (N_4736,N_4571,N_4554);
or U4737 (N_4737,N_4424,N_4454);
nand U4738 (N_4738,N_4589,N_4596);
xnor U4739 (N_4739,N_4561,N_4488);
nand U4740 (N_4740,N_4414,N_4528);
and U4741 (N_4741,N_4449,N_4417);
or U4742 (N_4742,N_4501,N_4404);
or U4743 (N_4743,N_4571,N_4429);
or U4744 (N_4744,N_4547,N_4437);
nand U4745 (N_4745,N_4505,N_4581);
xnor U4746 (N_4746,N_4401,N_4428);
nand U4747 (N_4747,N_4462,N_4481);
or U4748 (N_4748,N_4540,N_4570);
xor U4749 (N_4749,N_4404,N_4419);
nand U4750 (N_4750,N_4540,N_4585);
and U4751 (N_4751,N_4517,N_4516);
and U4752 (N_4752,N_4502,N_4552);
nand U4753 (N_4753,N_4480,N_4430);
xor U4754 (N_4754,N_4545,N_4490);
nand U4755 (N_4755,N_4543,N_4557);
or U4756 (N_4756,N_4496,N_4462);
nand U4757 (N_4757,N_4487,N_4457);
nor U4758 (N_4758,N_4518,N_4543);
and U4759 (N_4759,N_4434,N_4453);
and U4760 (N_4760,N_4529,N_4493);
and U4761 (N_4761,N_4472,N_4518);
or U4762 (N_4762,N_4561,N_4492);
and U4763 (N_4763,N_4443,N_4545);
xnor U4764 (N_4764,N_4572,N_4562);
nand U4765 (N_4765,N_4411,N_4439);
nand U4766 (N_4766,N_4447,N_4598);
nor U4767 (N_4767,N_4436,N_4485);
nand U4768 (N_4768,N_4568,N_4479);
nor U4769 (N_4769,N_4451,N_4431);
nor U4770 (N_4770,N_4599,N_4556);
and U4771 (N_4771,N_4446,N_4528);
nand U4772 (N_4772,N_4483,N_4405);
nand U4773 (N_4773,N_4581,N_4466);
nor U4774 (N_4774,N_4409,N_4467);
nand U4775 (N_4775,N_4586,N_4412);
and U4776 (N_4776,N_4415,N_4420);
or U4777 (N_4777,N_4552,N_4444);
nor U4778 (N_4778,N_4470,N_4551);
nor U4779 (N_4779,N_4591,N_4427);
nor U4780 (N_4780,N_4435,N_4583);
nand U4781 (N_4781,N_4489,N_4443);
and U4782 (N_4782,N_4546,N_4433);
nand U4783 (N_4783,N_4529,N_4597);
and U4784 (N_4784,N_4439,N_4417);
and U4785 (N_4785,N_4564,N_4440);
nand U4786 (N_4786,N_4445,N_4500);
or U4787 (N_4787,N_4526,N_4579);
or U4788 (N_4788,N_4520,N_4564);
nor U4789 (N_4789,N_4488,N_4530);
and U4790 (N_4790,N_4490,N_4599);
nor U4791 (N_4791,N_4434,N_4592);
and U4792 (N_4792,N_4529,N_4592);
xnor U4793 (N_4793,N_4442,N_4492);
xor U4794 (N_4794,N_4448,N_4591);
nor U4795 (N_4795,N_4511,N_4599);
nor U4796 (N_4796,N_4574,N_4516);
or U4797 (N_4797,N_4477,N_4505);
and U4798 (N_4798,N_4409,N_4578);
nor U4799 (N_4799,N_4473,N_4588);
nor U4800 (N_4800,N_4686,N_4652);
and U4801 (N_4801,N_4656,N_4753);
nand U4802 (N_4802,N_4712,N_4761);
or U4803 (N_4803,N_4737,N_4710);
xnor U4804 (N_4804,N_4650,N_4731);
nand U4805 (N_4805,N_4697,N_4741);
nor U4806 (N_4806,N_4759,N_4640);
and U4807 (N_4807,N_4718,N_4784);
or U4808 (N_4808,N_4627,N_4701);
xor U4809 (N_4809,N_4680,N_4653);
xor U4810 (N_4810,N_4657,N_4654);
or U4811 (N_4811,N_4704,N_4622);
nor U4812 (N_4812,N_4764,N_4698);
nor U4813 (N_4813,N_4715,N_4744);
xor U4814 (N_4814,N_4736,N_4687);
xor U4815 (N_4815,N_4688,N_4706);
xor U4816 (N_4816,N_4695,N_4658);
nand U4817 (N_4817,N_4766,N_4732);
nor U4818 (N_4818,N_4790,N_4614);
and U4819 (N_4819,N_4748,N_4689);
and U4820 (N_4820,N_4740,N_4711);
xor U4821 (N_4821,N_4683,N_4625);
and U4822 (N_4822,N_4705,N_4608);
xor U4823 (N_4823,N_4708,N_4660);
or U4824 (N_4824,N_4783,N_4756);
xor U4825 (N_4825,N_4716,N_4649);
xnor U4826 (N_4826,N_4621,N_4671);
xor U4827 (N_4827,N_4779,N_4643);
or U4828 (N_4828,N_4601,N_4796);
or U4829 (N_4829,N_4624,N_4677);
xnor U4830 (N_4830,N_4612,N_4738);
and U4831 (N_4831,N_4763,N_4728);
or U4832 (N_4832,N_4709,N_4691);
xnor U4833 (N_4833,N_4629,N_4786);
and U4834 (N_4834,N_4757,N_4678);
nand U4835 (N_4835,N_4610,N_4762);
nand U4836 (N_4836,N_4722,N_4604);
or U4837 (N_4837,N_4747,N_4672);
or U4838 (N_4838,N_4735,N_4615);
or U4839 (N_4839,N_4659,N_4631);
xnor U4840 (N_4840,N_4662,N_4664);
nand U4841 (N_4841,N_4618,N_4647);
nand U4842 (N_4842,N_4645,N_4690);
or U4843 (N_4843,N_4787,N_4776);
and U4844 (N_4844,N_4758,N_4720);
nor U4845 (N_4845,N_4768,N_4693);
nor U4846 (N_4846,N_4794,N_4770);
nor U4847 (N_4847,N_4743,N_4772);
nor U4848 (N_4848,N_4623,N_4775);
nor U4849 (N_4849,N_4639,N_4634);
nor U4850 (N_4850,N_4773,N_4745);
or U4851 (N_4851,N_4651,N_4670);
xnor U4852 (N_4852,N_4724,N_4609);
nor U4853 (N_4853,N_4788,N_4754);
and U4854 (N_4854,N_4752,N_4730);
nand U4855 (N_4855,N_4798,N_4714);
nor U4856 (N_4856,N_4605,N_4694);
and U4857 (N_4857,N_4792,N_4637);
nand U4858 (N_4858,N_4638,N_4603);
and U4859 (N_4859,N_4644,N_4727);
or U4860 (N_4860,N_4789,N_4646);
nand U4861 (N_4861,N_4751,N_4696);
xnor U4862 (N_4862,N_4655,N_4674);
nand U4863 (N_4863,N_4725,N_4717);
and U4864 (N_4864,N_4666,N_4667);
nand U4865 (N_4865,N_4785,N_4739);
nand U4866 (N_4866,N_4765,N_4777);
and U4867 (N_4867,N_4681,N_4606);
nand U4868 (N_4868,N_4733,N_4682);
nor U4869 (N_4869,N_4749,N_4692);
and U4870 (N_4870,N_4702,N_4742);
or U4871 (N_4871,N_4755,N_4746);
or U4872 (N_4872,N_4633,N_4676);
and U4873 (N_4873,N_4721,N_4632);
xnor U4874 (N_4874,N_4648,N_4760);
nor U4875 (N_4875,N_4750,N_4617);
or U4876 (N_4876,N_4707,N_4607);
or U4877 (N_4877,N_4791,N_4641);
nand U4878 (N_4878,N_4600,N_4769);
xnor U4879 (N_4879,N_4726,N_4616);
xor U4880 (N_4880,N_4635,N_4781);
xnor U4881 (N_4881,N_4793,N_4602);
nor U4882 (N_4882,N_4665,N_4780);
nand U4883 (N_4883,N_4729,N_4626);
xor U4884 (N_4884,N_4668,N_4673);
nor U4885 (N_4885,N_4669,N_4767);
nand U4886 (N_4886,N_4703,N_4630);
xor U4887 (N_4887,N_4799,N_4700);
nand U4888 (N_4888,N_4719,N_4663);
nand U4889 (N_4889,N_4774,N_4619);
nand U4890 (N_4890,N_4679,N_4613);
xor U4891 (N_4891,N_4661,N_4795);
xnor U4892 (N_4892,N_4684,N_4797);
nor U4893 (N_4893,N_4734,N_4620);
nor U4894 (N_4894,N_4642,N_4628);
or U4895 (N_4895,N_4723,N_4778);
and U4896 (N_4896,N_4771,N_4699);
or U4897 (N_4897,N_4685,N_4636);
and U4898 (N_4898,N_4782,N_4675);
or U4899 (N_4899,N_4611,N_4713);
or U4900 (N_4900,N_4604,N_4744);
nand U4901 (N_4901,N_4631,N_4744);
or U4902 (N_4902,N_4673,N_4651);
nand U4903 (N_4903,N_4684,N_4680);
and U4904 (N_4904,N_4623,N_4750);
nor U4905 (N_4905,N_4742,N_4604);
and U4906 (N_4906,N_4626,N_4605);
or U4907 (N_4907,N_4742,N_4606);
nor U4908 (N_4908,N_4721,N_4627);
xor U4909 (N_4909,N_4779,N_4793);
nand U4910 (N_4910,N_4640,N_4726);
xor U4911 (N_4911,N_4782,N_4718);
or U4912 (N_4912,N_4738,N_4604);
xor U4913 (N_4913,N_4774,N_4712);
or U4914 (N_4914,N_4791,N_4690);
nor U4915 (N_4915,N_4624,N_4790);
or U4916 (N_4916,N_4695,N_4719);
and U4917 (N_4917,N_4791,N_4737);
and U4918 (N_4918,N_4753,N_4644);
nor U4919 (N_4919,N_4654,N_4737);
nand U4920 (N_4920,N_4611,N_4783);
and U4921 (N_4921,N_4751,N_4669);
nand U4922 (N_4922,N_4655,N_4742);
or U4923 (N_4923,N_4777,N_4652);
or U4924 (N_4924,N_4646,N_4714);
nor U4925 (N_4925,N_4610,N_4644);
and U4926 (N_4926,N_4673,N_4727);
or U4927 (N_4927,N_4709,N_4642);
or U4928 (N_4928,N_4798,N_4686);
or U4929 (N_4929,N_4733,N_4627);
xnor U4930 (N_4930,N_4788,N_4766);
nand U4931 (N_4931,N_4629,N_4794);
nand U4932 (N_4932,N_4757,N_4755);
nand U4933 (N_4933,N_4670,N_4672);
nand U4934 (N_4934,N_4779,N_4636);
xnor U4935 (N_4935,N_4648,N_4716);
nor U4936 (N_4936,N_4763,N_4695);
nor U4937 (N_4937,N_4683,N_4749);
or U4938 (N_4938,N_4798,N_4666);
and U4939 (N_4939,N_4728,N_4796);
and U4940 (N_4940,N_4747,N_4709);
nand U4941 (N_4941,N_4630,N_4614);
and U4942 (N_4942,N_4712,N_4623);
xnor U4943 (N_4943,N_4662,N_4607);
nand U4944 (N_4944,N_4720,N_4791);
or U4945 (N_4945,N_4652,N_4647);
nand U4946 (N_4946,N_4726,N_4777);
xor U4947 (N_4947,N_4635,N_4737);
or U4948 (N_4948,N_4674,N_4691);
xnor U4949 (N_4949,N_4649,N_4710);
and U4950 (N_4950,N_4616,N_4719);
or U4951 (N_4951,N_4664,N_4772);
or U4952 (N_4952,N_4668,N_4615);
and U4953 (N_4953,N_4620,N_4778);
nor U4954 (N_4954,N_4782,N_4707);
and U4955 (N_4955,N_4741,N_4771);
nand U4956 (N_4956,N_4648,N_4659);
nor U4957 (N_4957,N_4625,N_4788);
nor U4958 (N_4958,N_4667,N_4702);
nor U4959 (N_4959,N_4632,N_4735);
or U4960 (N_4960,N_4655,N_4625);
and U4961 (N_4961,N_4616,N_4607);
and U4962 (N_4962,N_4743,N_4693);
or U4963 (N_4963,N_4660,N_4790);
or U4964 (N_4964,N_4730,N_4672);
nand U4965 (N_4965,N_4729,N_4650);
and U4966 (N_4966,N_4622,N_4628);
xor U4967 (N_4967,N_4656,N_4659);
nor U4968 (N_4968,N_4787,N_4671);
or U4969 (N_4969,N_4761,N_4654);
or U4970 (N_4970,N_4670,N_4780);
nand U4971 (N_4971,N_4755,N_4732);
nand U4972 (N_4972,N_4787,N_4683);
xnor U4973 (N_4973,N_4757,N_4638);
nand U4974 (N_4974,N_4718,N_4687);
xnor U4975 (N_4975,N_4635,N_4700);
or U4976 (N_4976,N_4742,N_4638);
and U4977 (N_4977,N_4786,N_4760);
and U4978 (N_4978,N_4615,N_4774);
nand U4979 (N_4979,N_4600,N_4639);
nand U4980 (N_4980,N_4671,N_4777);
nor U4981 (N_4981,N_4628,N_4681);
nand U4982 (N_4982,N_4737,N_4691);
and U4983 (N_4983,N_4638,N_4615);
and U4984 (N_4984,N_4698,N_4669);
xnor U4985 (N_4985,N_4684,N_4729);
xnor U4986 (N_4986,N_4715,N_4608);
or U4987 (N_4987,N_4696,N_4666);
and U4988 (N_4988,N_4644,N_4704);
nand U4989 (N_4989,N_4740,N_4724);
xnor U4990 (N_4990,N_4727,N_4692);
and U4991 (N_4991,N_4629,N_4654);
nand U4992 (N_4992,N_4785,N_4771);
and U4993 (N_4993,N_4620,N_4664);
xor U4994 (N_4994,N_4735,N_4612);
and U4995 (N_4995,N_4655,N_4762);
nor U4996 (N_4996,N_4658,N_4783);
nand U4997 (N_4997,N_4619,N_4699);
and U4998 (N_4998,N_4605,N_4723);
nor U4999 (N_4999,N_4742,N_4668);
xor U5000 (N_5000,N_4873,N_4858);
xor U5001 (N_5001,N_4864,N_4924);
nor U5002 (N_5002,N_4981,N_4991);
or U5003 (N_5003,N_4952,N_4819);
and U5004 (N_5004,N_4853,N_4972);
or U5005 (N_5005,N_4856,N_4802);
nor U5006 (N_5006,N_4838,N_4938);
nand U5007 (N_5007,N_4886,N_4898);
nor U5008 (N_5008,N_4909,N_4840);
and U5009 (N_5009,N_4891,N_4863);
xor U5010 (N_5010,N_4892,N_4903);
nor U5011 (N_5011,N_4806,N_4948);
nor U5012 (N_5012,N_4859,N_4975);
xnor U5013 (N_5013,N_4967,N_4922);
xnor U5014 (N_5014,N_4917,N_4932);
xnor U5015 (N_5015,N_4887,N_4827);
nand U5016 (N_5016,N_4990,N_4977);
and U5017 (N_5017,N_4823,N_4973);
nand U5018 (N_5018,N_4843,N_4996);
or U5019 (N_5019,N_4835,N_4986);
and U5020 (N_5020,N_4916,N_4867);
nand U5021 (N_5021,N_4900,N_4880);
nor U5022 (N_5022,N_4934,N_4974);
nand U5023 (N_5023,N_4800,N_4937);
or U5024 (N_5024,N_4866,N_4978);
and U5025 (N_5025,N_4889,N_4885);
nand U5026 (N_5026,N_4923,N_4879);
nor U5027 (N_5027,N_4931,N_4965);
and U5028 (N_5028,N_4933,N_4921);
and U5029 (N_5029,N_4822,N_4824);
xor U5030 (N_5030,N_4888,N_4820);
nand U5031 (N_5031,N_4808,N_4812);
xnor U5032 (N_5032,N_4979,N_4998);
xor U5033 (N_5033,N_4901,N_4964);
or U5034 (N_5034,N_4970,N_4956);
nand U5035 (N_5035,N_4907,N_4814);
or U5036 (N_5036,N_4944,N_4946);
or U5037 (N_5037,N_4955,N_4941);
xnor U5038 (N_5038,N_4983,N_4926);
and U5039 (N_5039,N_4953,N_4947);
nand U5040 (N_5040,N_4945,N_4828);
and U5041 (N_5041,N_4989,N_4831);
and U5042 (N_5042,N_4833,N_4813);
xor U5043 (N_5043,N_4861,N_4875);
xnor U5044 (N_5044,N_4988,N_4980);
or U5045 (N_5045,N_4837,N_4925);
xnor U5046 (N_5046,N_4915,N_4817);
nand U5047 (N_5047,N_4816,N_4855);
xnor U5048 (N_5048,N_4811,N_4845);
or U5049 (N_5049,N_4834,N_4874);
and U5050 (N_5050,N_4890,N_4999);
nor U5051 (N_5051,N_4920,N_4857);
xnor U5052 (N_5052,N_4954,N_4995);
and U5053 (N_5053,N_4930,N_4818);
or U5054 (N_5054,N_4897,N_4804);
xnor U5055 (N_5055,N_4911,N_4905);
nand U5056 (N_5056,N_4884,N_4868);
nor U5057 (N_5057,N_4936,N_4877);
nand U5058 (N_5058,N_4997,N_4842);
nand U5059 (N_5059,N_4846,N_4850);
or U5060 (N_5060,N_4848,N_4896);
and U5061 (N_5061,N_4919,N_4815);
and U5062 (N_5062,N_4987,N_4935);
and U5063 (N_5063,N_4865,N_4962);
and U5064 (N_5064,N_4810,N_4825);
and U5065 (N_5065,N_4910,N_4906);
nor U5066 (N_5066,N_4801,N_4870);
nor U5067 (N_5067,N_4963,N_4958);
or U5068 (N_5068,N_4904,N_4872);
nor U5069 (N_5069,N_4830,N_4992);
and U5070 (N_5070,N_4982,N_4908);
nor U5071 (N_5071,N_4957,N_4847);
xor U5072 (N_5072,N_4829,N_4940);
or U5073 (N_5073,N_4807,N_4968);
nor U5074 (N_5074,N_4994,N_4826);
nand U5075 (N_5075,N_4993,N_4913);
nand U5076 (N_5076,N_4985,N_4893);
nor U5077 (N_5077,N_4882,N_4899);
and U5078 (N_5078,N_4950,N_4852);
nor U5079 (N_5079,N_4951,N_4894);
xor U5080 (N_5080,N_4851,N_4961);
nand U5081 (N_5081,N_4878,N_4927);
or U5082 (N_5082,N_4862,N_4809);
nor U5083 (N_5083,N_4883,N_4849);
xnor U5084 (N_5084,N_4969,N_4839);
xor U5085 (N_5085,N_4895,N_4881);
and U5086 (N_5086,N_4902,N_4871);
xnor U5087 (N_5087,N_4942,N_4971);
xnor U5088 (N_5088,N_4984,N_4844);
xnor U5089 (N_5089,N_4841,N_4949);
nand U5090 (N_5090,N_4860,N_4939);
nor U5091 (N_5091,N_4943,N_4959);
xnor U5092 (N_5092,N_4912,N_4966);
nand U5093 (N_5093,N_4914,N_4918);
nor U5094 (N_5094,N_4928,N_4869);
nor U5095 (N_5095,N_4960,N_4803);
nand U5096 (N_5096,N_4836,N_4929);
and U5097 (N_5097,N_4821,N_4854);
nor U5098 (N_5098,N_4832,N_4876);
nand U5099 (N_5099,N_4805,N_4976);
and U5100 (N_5100,N_4930,N_4862);
nor U5101 (N_5101,N_4851,N_4902);
nor U5102 (N_5102,N_4807,N_4999);
nand U5103 (N_5103,N_4873,N_4933);
or U5104 (N_5104,N_4840,N_4940);
nor U5105 (N_5105,N_4913,N_4996);
nor U5106 (N_5106,N_4922,N_4839);
or U5107 (N_5107,N_4814,N_4878);
and U5108 (N_5108,N_4936,N_4869);
nand U5109 (N_5109,N_4918,N_4844);
nor U5110 (N_5110,N_4919,N_4861);
xor U5111 (N_5111,N_4900,N_4840);
or U5112 (N_5112,N_4807,N_4993);
and U5113 (N_5113,N_4823,N_4835);
nand U5114 (N_5114,N_4908,N_4856);
or U5115 (N_5115,N_4933,N_4876);
nor U5116 (N_5116,N_4910,N_4897);
and U5117 (N_5117,N_4853,N_4910);
nand U5118 (N_5118,N_4912,N_4928);
xnor U5119 (N_5119,N_4803,N_4850);
or U5120 (N_5120,N_4935,N_4998);
or U5121 (N_5121,N_4982,N_4839);
or U5122 (N_5122,N_4810,N_4926);
nand U5123 (N_5123,N_4860,N_4854);
nand U5124 (N_5124,N_4934,N_4937);
and U5125 (N_5125,N_4993,N_4931);
xnor U5126 (N_5126,N_4891,N_4956);
nand U5127 (N_5127,N_4915,N_4921);
nor U5128 (N_5128,N_4850,N_4953);
or U5129 (N_5129,N_4816,N_4880);
nor U5130 (N_5130,N_4824,N_4974);
and U5131 (N_5131,N_4833,N_4899);
xnor U5132 (N_5132,N_4839,N_4829);
or U5133 (N_5133,N_4865,N_4845);
nor U5134 (N_5134,N_4814,N_4901);
nand U5135 (N_5135,N_4855,N_4957);
nand U5136 (N_5136,N_4951,N_4882);
and U5137 (N_5137,N_4924,N_4979);
nor U5138 (N_5138,N_4994,N_4975);
and U5139 (N_5139,N_4890,N_4979);
and U5140 (N_5140,N_4973,N_4871);
nand U5141 (N_5141,N_4993,N_4914);
xnor U5142 (N_5142,N_4941,N_4827);
nand U5143 (N_5143,N_4970,N_4983);
nor U5144 (N_5144,N_4812,N_4983);
xor U5145 (N_5145,N_4847,N_4989);
and U5146 (N_5146,N_4987,N_4992);
xor U5147 (N_5147,N_4925,N_4852);
xnor U5148 (N_5148,N_4931,N_4887);
and U5149 (N_5149,N_4910,N_4997);
and U5150 (N_5150,N_4904,N_4917);
and U5151 (N_5151,N_4876,N_4918);
or U5152 (N_5152,N_4818,N_4879);
nand U5153 (N_5153,N_4908,N_4983);
xor U5154 (N_5154,N_4984,N_4806);
or U5155 (N_5155,N_4950,N_4934);
and U5156 (N_5156,N_4862,N_4878);
nand U5157 (N_5157,N_4807,N_4845);
nand U5158 (N_5158,N_4813,N_4847);
nor U5159 (N_5159,N_4816,N_4918);
and U5160 (N_5160,N_4882,N_4959);
or U5161 (N_5161,N_4985,N_4945);
nor U5162 (N_5162,N_4980,N_4870);
or U5163 (N_5163,N_4917,N_4947);
or U5164 (N_5164,N_4960,N_4856);
or U5165 (N_5165,N_4959,N_4949);
nor U5166 (N_5166,N_4847,N_4829);
nand U5167 (N_5167,N_4916,N_4811);
and U5168 (N_5168,N_4816,N_4883);
xor U5169 (N_5169,N_4871,N_4899);
or U5170 (N_5170,N_4944,N_4985);
and U5171 (N_5171,N_4883,N_4937);
and U5172 (N_5172,N_4805,N_4871);
and U5173 (N_5173,N_4970,N_4842);
nand U5174 (N_5174,N_4975,N_4965);
nand U5175 (N_5175,N_4815,N_4852);
nor U5176 (N_5176,N_4947,N_4929);
xor U5177 (N_5177,N_4898,N_4847);
xnor U5178 (N_5178,N_4815,N_4839);
or U5179 (N_5179,N_4938,N_4960);
and U5180 (N_5180,N_4949,N_4850);
or U5181 (N_5181,N_4949,N_4873);
nand U5182 (N_5182,N_4853,N_4887);
and U5183 (N_5183,N_4903,N_4915);
or U5184 (N_5184,N_4982,N_4940);
nor U5185 (N_5185,N_4850,N_4899);
xnor U5186 (N_5186,N_4867,N_4907);
nand U5187 (N_5187,N_4914,N_4851);
nand U5188 (N_5188,N_4817,N_4852);
xnor U5189 (N_5189,N_4906,N_4822);
nor U5190 (N_5190,N_4835,N_4809);
nand U5191 (N_5191,N_4943,N_4956);
or U5192 (N_5192,N_4935,N_4938);
nand U5193 (N_5193,N_4893,N_4864);
nand U5194 (N_5194,N_4836,N_4943);
and U5195 (N_5195,N_4942,N_4862);
and U5196 (N_5196,N_4812,N_4998);
or U5197 (N_5197,N_4936,N_4824);
xnor U5198 (N_5198,N_4972,N_4942);
or U5199 (N_5199,N_4904,N_4956);
or U5200 (N_5200,N_5059,N_5094);
xnor U5201 (N_5201,N_5198,N_5154);
and U5202 (N_5202,N_5184,N_5179);
xnor U5203 (N_5203,N_5122,N_5159);
nor U5204 (N_5204,N_5197,N_5067);
and U5205 (N_5205,N_5049,N_5167);
nor U5206 (N_5206,N_5110,N_5089);
and U5207 (N_5207,N_5011,N_5058);
and U5208 (N_5208,N_5187,N_5051);
nor U5209 (N_5209,N_5071,N_5101);
xor U5210 (N_5210,N_5139,N_5075);
and U5211 (N_5211,N_5090,N_5019);
nor U5212 (N_5212,N_5032,N_5123);
and U5213 (N_5213,N_5102,N_5006);
nor U5214 (N_5214,N_5168,N_5120);
and U5215 (N_5215,N_5104,N_5156);
xnor U5216 (N_5216,N_5063,N_5162);
nor U5217 (N_5217,N_5065,N_5017);
and U5218 (N_5218,N_5093,N_5060);
or U5219 (N_5219,N_5066,N_5112);
and U5220 (N_5220,N_5082,N_5143);
xnor U5221 (N_5221,N_5009,N_5074);
nand U5222 (N_5222,N_5044,N_5107);
nand U5223 (N_5223,N_5170,N_5158);
nand U5224 (N_5224,N_5163,N_5057);
nor U5225 (N_5225,N_5173,N_5152);
and U5226 (N_5226,N_5099,N_5190);
nand U5227 (N_5227,N_5177,N_5108);
or U5228 (N_5228,N_5157,N_5174);
nor U5229 (N_5229,N_5026,N_5161);
xnor U5230 (N_5230,N_5015,N_5048);
xor U5231 (N_5231,N_5041,N_5151);
nand U5232 (N_5232,N_5091,N_5037);
xor U5233 (N_5233,N_5047,N_5046);
xor U5234 (N_5234,N_5155,N_5118);
nand U5235 (N_5235,N_5133,N_5181);
and U5236 (N_5236,N_5195,N_5175);
and U5237 (N_5237,N_5146,N_5130);
or U5238 (N_5238,N_5160,N_5196);
or U5239 (N_5239,N_5052,N_5115);
nor U5240 (N_5240,N_5081,N_5192);
or U5241 (N_5241,N_5088,N_5148);
xnor U5242 (N_5242,N_5153,N_5126);
and U5243 (N_5243,N_5042,N_5125);
or U5244 (N_5244,N_5064,N_5189);
nand U5245 (N_5245,N_5020,N_5188);
or U5246 (N_5246,N_5109,N_5165);
or U5247 (N_5247,N_5003,N_5073);
nor U5248 (N_5248,N_5069,N_5194);
xor U5249 (N_5249,N_5116,N_5014);
and U5250 (N_5250,N_5117,N_5033);
and U5251 (N_5251,N_5013,N_5055);
nor U5252 (N_5252,N_5022,N_5135);
or U5253 (N_5253,N_5035,N_5053);
and U5254 (N_5254,N_5005,N_5199);
and U5255 (N_5255,N_5147,N_5136);
nor U5256 (N_5256,N_5039,N_5085);
and U5257 (N_5257,N_5128,N_5018);
xnor U5258 (N_5258,N_5138,N_5176);
xor U5259 (N_5259,N_5103,N_5098);
nor U5260 (N_5260,N_5043,N_5097);
xnor U5261 (N_5261,N_5183,N_5023);
or U5262 (N_5262,N_5087,N_5024);
and U5263 (N_5263,N_5054,N_5129);
nor U5264 (N_5264,N_5132,N_5106);
and U5265 (N_5265,N_5027,N_5114);
nor U5266 (N_5266,N_5172,N_5149);
xor U5267 (N_5267,N_5025,N_5164);
xnor U5268 (N_5268,N_5186,N_5077);
nand U5269 (N_5269,N_5016,N_5137);
and U5270 (N_5270,N_5080,N_5002);
and U5271 (N_5271,N_5036,N_5096);
nor U5272 (N_5272,N_5100,N_5072);
nand U5273 (N_5273,N_5070,N_5119);
or U5274 (N_5274,N_5105,N_5021);
nor U5275 (N_5275,N_5144,N_5062);
nor U5276 (N_5276,N_5121,N_5145);
or U5277 (N_5277,N_5095,N_5185);
nor U5278 (N_5278,N_5141,N_5079);
or U5279 (N_5279,N_5084,N_5191);
or U5280 (N_5280,N_5169,N_5004);
nor U5281 (N_5281,N_5028,N_5142);
or U5282 (N_5282,N_5076,N_5178);
nor U5283 (N_5283,N_5061,N_5031);
xor U5284 (N_5284,N_5040,N_5166);
and U5285 (N_5285,N_5029,N_5127);
nor U5286 (N_5286,N_5134,N_5193);
or U5287 (N_5287,N_5038,N_5092);
nor U5288 (N_5288,N_5068,N_5045);
or U5289 (N_5289,N_5078,N_5007);
xnor U5290 (N_5290,N_5034,N_5050);
or U5291 (N_5291,N_5171,N_5086);
and U5292 (N_5292,N_5000,N_5140);
nor U5293 (N_5293,N_5001,N_5111);
xor U5294 (N_5294,N_5030,N_5056);
nand U5295 (N_5295,N_5124,N_5113);
or U5296 (N_5296,N_5008,N_5182);
nor U5297 (N_5297,N_5131,N_5012);
and U5298 (N_5298,N_5180,N_5010);
or U5299 (N_5299,N_5083,N_5150);
nor U5300 (N_5300,N_5021,N_5118);
and U5301 (N_5301,N_5044,N_5192);
xor U5302 (N_5302,N_5071,N_5136);
nand U5303 (N_5303,N_5101,N_5050);
xnor U5304 (N_5304,N_5086,N_5081);
nor U5305 (N_5305,N_5051,N_5174);
or U5306 (N_5306,N_5039,N_5188);
and U5307 (N_5307,N_5185,N_5193);
or U5308 (N_5308,N_5091,N_5065);
xor U5309 (N_5309,N_5085,N_5169);
xnor U5310 (N_5310,N_5011,N_5145);
nand U5311 (N_5311,N_5191,N_5117);
nand U5312 (N_5312,N_5110,N_5127);
xor U5313 (N_5313,N_5067,N_5094);
or U5314 (N_5314,N_5053,N_5062);
and U5315 (N_5315,N_5011,N_5178);
nand U5316 (N_5316,N_5195,N_5185);
and U5317 (N_5317,N_5114,N_5092);
nand U5318 (N_5318,N_5038,N_5199);
or U5319 (N_5319,N_5120,N_5011);
and U5320 (N_5320,N_5088,N_5139);
or U5321 (N_5321,N_5068,N_5055);
nor U5322 (N_5322,N_5067,N_5049);
and U5323 (N_5323,N_5137,N_5059);
nor U5324 (N_5324,N_5041,N_5040);
nor U5325 (N_5325,N_5191,N_5170);
nand U5326 (N_5326,N_5123,N_5164);
or U5327 (N_5327,N_5036,N_5133);
or U5328 (N_5328,N_5007,N_5024);
xnor U5329 (N_5329,N_5033,N_5052);
and U5330 (N_5330,N_5105,N_5073);
nor U5331 (N_5331,N_5168,N_5092);
or U5332 (N_5332,N_5093,N_5065);
xor U5333 (N_5333,N_5026,N_5012);
nor U5334 (N_5334,N_5137,N_5063);
or U5335 (N_5335,N_5085,N_5145);
and U5336 (N_5336,N_5196,N_5095);
nand U5337 (N_5337,N_5017,N_5143);
nand U5338 (N_5338,N_5143,N_5094);
nand U5339 (N_5339,N_5046,N_5061);
xnor U5340 (N_5340,N_5111,N_5148);
or U5341 (N_5341,N_5097,N_5155);
nand U5342 (N_5342,N_5067,N_5119);
nand U5343 (N_5343,N_5183,N_5176);
and U5344 (N_5344,N_5110,N_5054);
nand U5345 (N_5345,N_5179,N_5108);
nand U5346 (N_5346,N_5068,N_5145);
nor U5347 (N_5347,N_5188,N_5010);
nor U5348 (N_5348,N_5059,N_5005);
xnor U5349 (N_5349,N_5129,N_5071);
nor U5350 (N_5350,N_5167,N_5196);
or U5351 (N_5351,N_5097,N_5166);
nor U5352 (N_5352,N_5177,N_5056);
nand U5353 (N_5353,N_5142,N_5185);
xnor U5354 (N_5354,N_5027,N_5028);
xor U5355 (N_5355,N_5121,N_5088);
xor U5356 (N_5356,N_5148,N_5132);
xor U5357 (N_5357,N_5109,N_5103);
nor U5358 (N_5358,N_5186,N_5035);
nand U5359 (N_5359,N_5023,N_5184);
and U5360 (N_5360,N_5144,N_5126);
or U5361 (N_5361,N_5103,N_5066);
nor U5362 (N_5362,N_5044,N_5110);
xnor U5363 (N_5363,N_5036,N_5183);
nand U5364 (N_5364,N_5126,N_5111);
and U5365 (N_5365,N_5062,N_5066);
nor U5366 (N_5366,N_5185,N_5033);
xnor U5367 (N_5367,N_5063,N_5066);
xor U5368 (N_5368,N_5102,N_5169);
or U5369 (N_5369,N_5038,N_5141);
nand U5370 (N_5370,N_5010,N_5019);
or U5371 (N_5371,N_5166,N_5106);
or U5372 (N_5372,N_5046,N_5178);
or U5373 (N_5373,N_5127,N_5005);
xor U5374 (N_5374,N_5063,N_5183);
and U5375 (N_5375,N_5176,N_5035);
nor U5376 (N_5376,N_5070,N_5004);
nor U5377 (N_5377,N_5148,N_5032);
xnor U5378 (N_5378,N_5156,N_5169);
nand U5379 (N_5379,N_5107,N_5097);
nand U5380 (N_5380,N_5093,N_5103);
and U5381 (N_5381,N_5046,N_5037);
or U5382 (N_5382,N_5046,N_5192);
nor U5383 (N_5383,N_5028,N_5152);
nand U5384 (N_5384,N_5013,N_5100);
nor U5385 (N_5385,N_5059,N_5120);
nand U5386 (N_5386,N_5156,N_5035);
xnor U5387 (N_5387,N_5117,N_5111);
and U5388 (N_5388,N_5113,N_5183);
or U5389 (N_5389,N_5136,N_5016);
or U5390 (N_5390,N_5113,N_5060);
nor U5391 (N_5391,N_5168,N_5040);
nand U5392 (N_5392,N_5127,N_5060);
nor U5393 (N_5393,N_5029,N_5120);
xor U5394 (N_5394,N_5036,N_5171);
xnor U5395 (N_5395,N_5159,N_5044);
and U5396 (N_5396,N_5033,N_5118);
or U5397 (N_5397,N_5194,N_5198);
or U5398 (N_5398,N_5098,N_5193);
xor U5399 (N_5399,N_5015,N_5068);
or U5400 (N_5400,N_5336,N_5353);
nor U5401 (N_5401,N_5320,N_5226);
and U5402 (N_5402,N_5237,N_5339);
nand U5403 (N_5403,N_5321,N_5366);
nand U5404 (N_5404,N_5221,N_5322);
nand U5405 (N_5405,N_5241,N_5248);
or U5406 (N_5406,N_5211,N_5252);
nor U5407 (N_5407,N_5259,N_5265);
and U5408 (N_5408,N_5388,N_5206);
xnor U5409 (N_5409,N_5247,N_5251);
nand U5410 (N_5410,N_5332,N_5340);
and U5411 (N_5411,N_5234,N_5217);
and U5412 (N_5412,N_5271,N_5278);
nor U5413 (N_5413,N_5394,N_5311);
or U5414 (N_5414,N_5242,N_5210);
nand U5415 (N_5415,N_5325,N_5371);
or U5416 (N_5416,N_5239,N_5273);
xor U5417 (N_5417,N_5395,N_5246);
and U5418 (N_5418,N_5370,N_5244);
nor U5419 (N_5419,N_5346,N_5367);
nand U5420 (N_5420,N_5208,N_5203);
and U5421 (N_5421,N_5345,N_5357);
nand U5422 (N_5422,N_5213,N_5362);
nand U5423 (N_5423,N_5232,N_5308);
or U5424 (N_5424,N_5304,N_5397);
xor U5425 (N_5425,N_5352,N_5282);
nor U5426 (N_5426,N_5379,N_5399);
or U5427 (N_5427,N_5205,N_5287);
and U5428 (N_5428,N_5391,N_5316);
nand U5429 (N_5429,N_5269,N_5218);
or U5430 (N_5430,N_5348,N_5342);
nand U5431 (N_5431,N_5364,N_5295);
xor U5432 (N_5432,N_5262,N_5343);
or U5433 (N_5433,N_5292,N_5272);
or U5434 (N_5434,N_5297,N_5337);
and U5435 (N_5435,N_5341,N_5326);
xor U5436 (N_5436,N_5245,N_5298);
and U5437 (N_5437,N_5233,N_5214);
nor U5438 (N_5438,N_5314,N_5305);
and U5439 (N_5439,N_5301,N_5277);
or U5440 (N_5440,N_5331,N_5312);
xnor U5441 (N_5441,N_5286,N_5275);
or U5442 (N_5442,N_5220,N_5238);
and U5443 (N_5443,N_5288,N_5378);
and U5444 (N_5444,N_5284,N_5329);
xor U5445 (N_5445,N_5293,N_5257);
nand U5446 (N_5446,N_5317,N_5363);
or U5447 (N_5447,N_5310,N_5347);
xor U5448 (N_5448,N_5385,N_5349);
nand U5449 (N_5449,N_5254,N_5338);
nor U5450 (N_5450,N_5324,N_5276);
or U5451 (N_5451,N_5300,N_5250);
and U5452 (N_5452,N_5376,N_5204);
or U5453 (N_5453,N_5260,N_5296);
xnor U5454 (N_5454,N_5381,N_5303);
xor U5455 (N_5455,N_5313,N_5207);
xor U5456 (N_5456,N_5231,N_5258);
nor U5457 (N_5457,N_5228,N_5219);
nor U5458 (N_5458,N_5383,N_5369);
and U5459 (N_5459,N_5264,N_5229);
nor U5460 (N_5460,N_5253,N_5267);
nor U5461 (N_5461,N_5255,N_5372);
and U5462 (N_5462,N_5209,N_5279);
nand U5463 (N_5463,N_5382,N_5212);
or U5464 (N_5464,N_5291,N_5330);
nor U5465 (N_5465,N_5307,N_5361);
or U5466 (N_5466,N_5222,N_5333);
nor U5467 (N_5467,N_5274,N_5299);
xnor U5468 (N_5468,N_5356,N_5266);
nor U5469 (N_5469,N_5223,N_5359);
nand U5470 (N_5470,N_5354,N_5365);
or U5471 (N_5471,N_5368,N_5386);
and U5472 (N_5472,N_5350,N_5235);
or U5473 (N_5473,N_5315,N_5268);
nand U5474 (N_5474,N_5373,N_5306);
xor U5475 (N_5475,N_5289,N_5309);
and U5476 (N_5476,N_5225,N_5355);
nor U5477 (N_5477,N_5387,N_5256);
xor U5478 (N_5478,N_5200,N_5396);
or U5479 (N_5479,N_5327,N_5224);
and U5480 (N_5480,N_5302,N_5249);
and U5481 (N_5481,N_5351,N_5390);
nor U5482 (N_5482,N_5202,N_5360);
or U5483 (N_5483,N_5398,N_5374);
and U5484 (N_5484,N_5230,N_5294);
and U5485 (N_5485,N_5270,N_5201);
and U5486 (N_5486,N_5243,N_5328);
and U5487 (N_5487,N_5215,N_5335);
xnor U5488 (N_5488,N_5227,N_5280);
and U5489 (N_5489,N_5323,N_5290);
nand U5490 (N_5490,N_5380,N_5375);
and U5491 (N_5491,N_5281,N_5344);
nor U5492 (N_5492,N_5240,N_5283);
xor U5493 (N_5493,N_5334,N_5285);
or U5494 (N_5494,N_5263,N_5236);
or U5495 (N_5495,N_5384,N_5358);
nand U5496 (N_5496,N_5319,N_5377);
nor U5497 (N_5497,N_5393,N_5389);
nor U5498 (N_5498,N_5261,N_5216);
and U5499 (N_5499,N_5392,N_5318);
nand U5500 (N_5500,N_5303,N_5312);
and U5501 (N_5501,N_5253,N_5260);
nand U5502 (N_5502,N_5250,N_5227);
xor U5503 (N_5503,N_5352,N_5254);
xnor U5504 (N_5504,N_5352,N_5215);
nand U5505 (N_5505,N_5241,N_5201);
or U5506 (N_5506,N_5285,N_5315);
and U5507 (N_5507,N_5214,N_5322);
xnor U5508 (N_5508,N_5273,N_5207);
and U5509 (N_5509,N_5200,N_5337);
and U5510 (N_5510,N_5354,N_5214);
nor U5511 (N_5511,N_5315,N_5255);
nand U5512 (N_5512,N_5240,N_5344);
xnor U5513 (N_5513,N_5339,N_5369);
nor U5514 (N_5514,N_5208,N_5302);
and U5515 (N_5515,N_5398,N_5392);
nor U5516 (N_5516,N_5215,N_5210);
and U5517 (N_5517,N_5324,N_5381);
xnor U5518 (N_5518,N_5374,N_5336);
and U5519 (N_5519,N_5263,N_5224);
nand U5520 (N_5520,N_5367,N_5224);
and U5521 (N_5521,N_5255,N_5228);
xnor U5522 (N_5522,N_5350,N_5210);
nor U5523 (N_5523,N_5256,N_5206);
and U5524 (N_5524,N_5267,N_5338);
or U5525 (N_5525,N_5226,N_5230);
and U5526 (N_5526,N_5251,N_5375);
nand U5527 (N_5527,N_5360,N_5348);
xnor U5528 (N_5528,N_5373,N_5331);
xor U5529 (N_5529,N_5288,N_5244);
nor U5530 (N_5530,N_5256,N_5254);
nand U5531 (N_5531,N_5332,N_5382);
xor U5532 (N_5532,N_5377,N_5217);
xnor U5533 (N_5533,N_5273,N_5360);
or U5534 (N_5534,N_5312,N_5330);
xor U5535 (N_5535,N_5355,N_5257);
nor U5536 (N_5536,N_5304,N_5288);
or U5537 (N_5537,N_5284,N_5292);
nor U5538 (N_5538,N_5378,N_5205);
nand U5539 (N_5539,N_5209,N_5356);
nand U5540 (N_5540,N_5321,N_5326);
nand U5541 (N_5541,N_5372,N_5212);
xnor U5542 (N_5542,N_5273,N_5284);
and U5543 (N_5543,N_5223,N_5394);
nand U5544 (N_5544,N_5294,N_5384);
nor U5545 (N_5545,N_5208,N_5361);
xnor U5546 (N_5546,N_5321,N_5369);
or U5547 (N_5547,N_5212,N_5357);
nor U5548 (N_5548,N_5326,N_5345);
nor U5549 (N_5549,N_5333,N_5332);
nand U5550 (N_5550,N_5231,N_5357);
nor U5551 (N_5551,N_5397,N_5285);
or U5552 (N_5552,N_5251,N_5349);
and U5553 (N_5553,N_5295,N_5370);
and U5554 (N_5554,N_5386,N_5224);
and U5555 (N_5555,N_5382,N_5229);
nand U5556 (N_5556,N_5375,N_5214);
xor U5557 (N_5557,N_5397,N_5260);
nand U5558 (N_5558,N_5271,N_5203);
and U5559 (N_5559,N_5212,N_5312);
and U5560 (N_5560,N_5378,N_5327);
or U5561 (N_5561,N_5309,N_5216);
xnor U5562 (N_5562,N_5211,N_5345);
or U5563 (N_5563,N_5392,N_5369);
nor U5564 (N_5564,N_5380,N_5223);
xnor U5565 (N_5565,N_5306,N_5280);
and U5566 (N_5566,N_5308,N_5260);
nand U5567 (N_5567,N_5303,N_5338);
xor U5568 (N_5568,N_5342,N_5242);
and U5569 (N_5569,N_5333,N_5322);
and U5570 (N_5570,N_5350,N_5353);
nand U5571 (N_5571,N_5207,N_5333);
nand U5572 (N_5572,N_5267,N_5344);
or U5573 (N_5573,N_5334,N_5287);
or U5574 (N_5574,N_5206,N_5277);
xnor U5575 (N_5575,N_5386,N_5263);
and U5576 (N_5576,N_5324,N_5292);
and U5577 (N_5577,N_5285,N_5201);
and U5578 (N_5578,N_5275,N_5274);
or U5579 (N_5579,N_5383,N_5285);
nand U5580 (N_5580,N_5248,N_5318);
xnor U5581 (N_5581,N_5388,N_5319);
nor U5582 (N_5582,N_5244,N_5290);
or U5583 (N_5583,N_5358,N_5340);
and U5584 (N_5584,N_5317,N_5265);
and U5585 (N_5585,N_5386,N_5219);
xor U5586 (N_5586,N_5212,N_5348);
nor U5587 (N_5587,N_5235,N_5243);
nor U5588 (N_5588,N_5316,N_5266);
xnor U5589 (N_5589,N_5361,N_5278);
and U5590 (N_5590,N_5291,N_5221);
nor U5591 (N_5591,N_5323,N_5214);
nor U5592 (N_5592,N_5238,N_5211);
xor U5593 (N_5593,N_5242,N_5224);
xor U5594 (N_5594,N_5258,N_5391);
and U5595 (N_5595,N_5272,N_5238);
or U5596 (N_5596,N_5393,N_5269);
nand U5597 (N_5597,N_5241,N_5208);
xor U5598 (N_5598,N_5294,N_5397);
nor U5599 (N_5599,N_5283,N_5263);
nor U5600 (N_5600,N_5561,N_5442);
nand U5601 (N_5601,N_5554,N_5589);
xor U5602 (N_5602,N_5533,N_5429);
and U5603 (N_5603,N_5492,N_5490);
xnor U5604 (N_5604,N_5423,N_5560);
nand U5605 (N_5605,N_5476,N_5588);
nor U5606 (N_5606,N_5566,N_5449);
xor U5607 (N_5607,N_5537,N_5438);
or U5608 (N_5608,N_5412,N_5462);
nand U5609 (N_5609,N_5559,N_5427);
and U5610 (N_5610,N_5435,N_5482);
xnor U5611 (N_5611,N_5568,N_5456);
or U5612 (N_5612,N_5461,N_5453);
nor U5613 (N_5613,N_5584,N_5549);
and U5614 (N_5614,N_5421,N_5466);
xor U5615 (N_5615,N_5485,N_5570);
and U5616 (N_5616,N_5530,N_5504);
nor U5617 (N_5617,N_5477,N_5571);
xnor U5618 (N_5618,N_5437,N_5593);
nand U5619 (N_5619,N_5599,N_5590);
and U5620 (N_5620,N_5440,N_5410);
nand U5621 (N_5621,N_5544,N_5527);
or U5622 (N_5622,N_5404,N_5407);
or U5623 (N_5623,N_5509,N_5596);
nor U5624 (N_5624,N_5460,N_5553);
or U5625 (N_5625,N_5434,N_5441);
xnor U5626 (N_5626,N_5415,N_5489);
nand U5627 (N_5627,N_5558,N_5542);
xnor U5628 (N_5628,N_5524,N_5487);
xor U5629 (N_5629,N_5400,N_5592);
or U5630 (N_5630,N_5432,N_5416);
nor U5631 (N_5631,N_5496,N_5480);
nor U5632 (N_5632,N_5468,N_5595);
xor U5633 (N_5633,N_5497,N_5548);
and U5634 (N_5634,N_5479,N_5591);
or U5635 (N_5635,N_5406,N_5522);
or U5636 (N_5636,N_5557,N_5563);
or U5637 (N_5637,N_5538,N_5578);
xor U5638 (N_5638,N_5414,N_5539);
nor U5639 (N_5639,N_5488,N_5574);
nor U5640 (N_5640,N_5505,N_5495);
and U5641 (N_5641,N_5580,N_5587);
xnor U5642 (N_5642,N_5511,N_5597);
nor U5643 (N_5643,N_5551,N_5469);
nand U5644 (N_5644,N_5535,N_5443);
xnor U5645 (N_5645,N_5426,N_5439);
and U5646 (N_5646,N_5541,N_5543);
xnor U5647 (N_5647,N_5491,N_5425);
nor U5648 (N_5648,N_5446,N_5576);
or U5649 (N_5649,N_5467,N_5512);
nor U5650 (N_5650,N_5545,N_5401);
nor U5651 (N_5651,N_5517,N_5454);
or U5652 (N_5652,N_5455,N_5452);
or U5653 (N_5653,N_5471,N_5420);
xor U5654 (N_5654,N_5499,N_5408);
nor U5655 (N_5655,N_5478,N_5564);
xor U5656 (N_5656,N_5457,N_5556);
nand U5657 (N_5657,N_5519,N_5508);
and U5658 (N_5658,N_5546,N_5507);
and U5659 (N_5659,N_5532,N_5575);
nor U5660 (N_5660,N_5459,N_5419);
or U5661 (N_5661,N_5534,N_5422);
nor U5662 (N_5662,N_5565,N_5433);
and U5663 (N_5663,N_5418,N_5585);
xnor U5664 (N_5664,N_5510,N_5498);
xor U5665 (N_5665,N_5555,N_5424);
nand U5666 (N_5666,N_5493,N_5486);
or U5667 (N_5667,N_5463,N_5562);
and U5668 (N_5668,N_5430,N_5451);
nand U5669 (N_5669,N_5583,N_5514);
nand U5670 (N_5670,N_5531,N_5515);
nand U5671 (N_5671,N_5448,N_5402);
nor U5672 (N_5672,N_5413,N_5465);
and U5673 (N_5673,N_5523,N_5444);
or U5674 (N_5674,N_5431,N_5502);
or U5675 (N_5675,N_5550,N_5581);
xor U5676 (N_5676,N_5582,N_5569);
nor U5677 (N_5677,N_5572,N_5526);
and U5678 (N_5678,N_5501,N_5494);
xor U5679 (N_5679,N_5436,N_5540);
and U5680 (N_5680,N_5529,N_5567);
or U5681 (N_5681,N_5458,N_5577);
or U5682 (N_5682,N_5573,N_5520);
and U5683 (N_5683,N_5500,N_5447);
and U5684 (N_5684,N_5450,N_5579);
nor U5685 (N_5685,N_5536,N_5598);
nor U5686 (N_5686,N_5528,N_5411);
and U5687 (N_5687,N_5473,N_5472);
or U5688 (N_5688,N_5470,N_5445);
or U5689 (N_5689,N_5586,N_5594);
nor U5690 (N_5690,N_5518,N_5484);
or U5691 (N_5691,N_5403,N_5503);
nand U5692 (N_5692,N_5428,N_5475);
or U5693 (N_5693,N_5516,N_5474);
nand U5694 (N_5694,N_5483,N_5525);
xnor U5695 (N_5695,N_5552,N_5409);
nand U5696 (N_5696,N_5417,N_5513);
and U5697 (N_5697,N_5521,N_5547);
nand U5698 (N_5698,N_5481,N_5405);
xor U5699 (N_5699,N_5464,N_5506);
nor U5700 (N_5700,N_5440,N_5502);
xnor U5701 (N_5701,N_5451,N_5557);
or U5702 (N_5702,N_5531,N_5591);
nor U5703 (N_5703,N_5409,N_5446);
nand U5704 (N_5704,N_5521,N_5561);
and U5705 (N_5705,N_5561,N_5513);
xnor U5706 (N_5706,N_5486,N_5597);
and U5707 (N_5707,N_5560,N_5545);
or U5708 (N_5708,N_5444,N_5404);
nor U5709 (N_5709,N_5484,N_5550);
or U5710 (N_5710,N_5409,N_5474);
or U5711 (N_5711,N_5598,N_5511);
and U5712 (N_5712,N_5426,N_5555);
nand U5713 (N_5713,N_5498,N_5565);
nor U5714 (N_5714,N_5413,N_5506);
or U5715 (N_5715,N_5574,N_5455);
nand U5716 (N_5716,N_5466,N_5489);
nand U5717 (N_5717,N_5423,N_5553);
nor U5718 (N_5718,N_5582,N_5449);
or U5719 (N_5719,N_5530,N_5547);
and U5720 (N_5720,N_5563,N_5490);
and U5721 (N_5721,N_5531,N_5511);
xnor U5722 (N_5722,N_5431,N_5527);
nand U5723 (N_5723,N_5440,N_5402);
xor U5724 (N_5724,N_5499,N_5430);
nand U5725 (N_5725,N_5483,N_5585);
xnor U5726 (N_5726,N_5409,N_5458);
xor U5727 (N_5727,N_5595,N_5593);
or U5728 (N_5728,N_5468,N_5441);
nand U5729 (N_5729,N_5580,N_5497);
nor U5730 (N_5730,N_5521,N_5579);
xor U5731 (N_5731,N_5456,N_5563);
nand U5732 (N_5732,N_5441,N_5485);
and U5733 (N_5733,N_5456,N_5509);
xor U5734 (N_5734,N_5453,N_5523);
and U5735 (N_5735,N_5552,N_5514);
xnor U5736 (N_5736,N_5429,N_5511);
or U5737 (N_5737,N_5531,N_5583);
or U5738 (N_5738,N_5575,N_5459);
and U5739 (N_5739,N_5441,N_5464);
nand U5740 (N_5740,N_5591,N_5521);
xor U5741 (N_5741,N_5460,N_5515);
nor U5742 (N_5742,N_5591,N_5518);
and U5743 (N_5743,N_5491,N_5565);
xor U5744 (N_5744,N_5424,N_5473);
and U5745 (N_5745,N_5463,N_5470);
or U5746 (N_5746,N_5480,N_5498);
xor U5747 (N_5747,N_5465,N_5442);
xor U5748 (N_5748,N_5523,N_5483);
nor U5749 (N_5749,N_5567,N_5512);
xor U5750 (N_5750,N_5511,N_5596);
and U5751 (N_5751,N_5557,N_5580);
or U5752 (N_5752,N_5457,N_5507);
or U5753 (N_5753,N_5588,N_5440);
nand U5754 (N_5754,N_5536,N_5478);
xor U5755 (N_5755,N_5401,N_5550);
and U5756 (N_5756,N_5460,N_5431);
xor U5757 (N_5757,N_5478,N_5435);
nor U5758 (N_5758,N_5404,N_5437);
or U5759 (N_5759,N_5494,N_5423);
nand U5760 (N_5760,N_5502,N_5462);
xnor U5761 (N_5761,N_5502,N_5595);
and U5762 (N_5762,N_5508,N_5549);
or U5763 (N_5763,N_5594,N_5535);
or U5764 (N_5764,N_5549,N_5510);
or U5765 (N_5765,N_5499,N_5434);
nor U5766 (N_5766,N_5512,N_5574);
xnor U5767 (N_5767,N_5472,N_5495);
or U5768 (N_5768,N_5524,N_5543);
and U5769 (N_5769,N_5418,N_5581);
nor U5770 (N_5770,N_5572,N_5417);
nor U5771 (N_5771,N_5526,N_5569);
and U5772 (N_5772,N_5444,N_5576);
nand U5773 (N_5773,N_5570,N_5471);
nand U5774 (N_5774,N_5463,N_5573);
xor U5775 (N_5775,N_5573,N_5431);
or U5776 (N_5776,N_5598,N_5541);
nand U5777 (N_5777,N_5583,N_5472);
nor U5778 (N_5778,N_5428,N_5555);
nor U5779 (N_5779,N_5572,N_5564);
nand U5780 (N_5780,N_5579,N_5411);
or U5781 (N_5781,N_5428,N_5565);
xnor U5782 (N_5782,N_5503,N_5480);
xor U5783 (N_5783,N_5477,N_5462);
nand U5784 (N_5784,N_5488,N_5463);
nand U5785 (N_5785,N_5437,N_5424);
and U5786 (N_5786,N_5495,N_5477);
or U5787 (N_5787,N_5528,N_5594);
xor U5788 (N_5788,N_5430,N_5454);
nand U5789 (N_5789,N_5551,N_5453);
nand U5790 (N_5790,N_5421,N_5567);
nand U5791 (N_5791,N_5561,N_5409);
nor U5792 (N_5792,N_5556,N_5414);
nand U5793 (N_5793,N_5455,N_5448);
or U5794 (N_5794,N_5523,N_5446);
or U5795 (N_5795,N_5438,N_5486);
nand U5796 (N_5796,N_5489,N_5539);
and U5797 (N_5797,N_5586,N_5555);
xor U5798 (N_5798,N_5548,N_5494);
and U5799 (N_5799,N_5512,N_5416);
nand U5800 (N_5800,N_5788,N_5697);
xnor U5801 (N_5801,N_5762,N_5755);
nand U5802 (N_5802,N_5688,N_5651);
nor U5803 (N_5803,N_5620,N_5747);
nor U5804 (N_5804,N_5708,N_5639);
nor U5805 (N_5805,N_5763,N_5775);
or U5806 (N_5806,N_5710,N_5640);
xor U5807 (N_5807,N_5777,N_5718);
or U5808 (N_5808,N_5634,N_5655);
xor U5809 (N_5809,N_5605,N_5624);
nand U5810 (N_5810,N_5692,N_5613);
or U5811 (N_5811,N_5623,N_5673);
or U5812 (N_5812,N_5733,N_5695);
or U5813 (N_5813,N_5721,N_5606);
or U5814 (N_5814,N_5676,N_5659);
nor U5815 (N_5815,N_5772,N_5770);
nand U5816 (N_5816,N_5736,N_5783);
nand U5817 (N_5817,N_5722,N_5671);
or U5818 (N_5818,N_5678,N_5675);
or U5819 (N_5819,N_5654,N_5715);
nor U5820 (N_5820,N_5608,N_5734);
or U5821 (N_5821,N_5668,N_5699);
and U5822 (N_5822,N_5682,N_5744);
nor U5823 (N_5823,N_5662,N_5751);
or U5824 (N_5824,N_5709,N_5694);
and U5825 (N_5825,N_5773,N_5680);
nand U5826 (N_5826,N_5661,N_5667);
and U5827 (N_5827,N_5626,N_5740);
xnor U5828 (N_5828,N_5732,N_5792);
nor U5829 (N_5829,N_5707,N_5630);
xor U5830 (N_5830,N_5713,N_5700);
or U5831 (N_5831,N_5689,N_5614);
or U5832 (N_5832,N_5632,N_5723);
and U5833 (N_5833,N_5728,N_5696);
nor U5834 (N_5834,N_5690,N_5650);
or U5835 (N_5835,N_5769,N_5797);
and U5836 (N_5836,N_5617,N_5693);
nor U5837 (N_5837,N_5658,N_5759);
and U5838 (N_5838,N_5714,N_5616);
or U5839 (N_5839,N_5635,N_5717);
xor U5840 (N_5840,N_5766,N_5648);
xor U5841 (N_5841,N_5646,N_5704);
and U5842 (N_5842,N_5745,N_5603);
or U5843 (N_5843,N_5643,N_5701);
or U5844 (N_5844,N_5794,N_5679);
or U5845 (N_5845,N_5685,N_5637);
and U5846 (N_5846,N_5622,N_5621);
nand U5847 (N_5847,N_5666,N_5750);
nor U5848 (N_5848,N_5672,N_5785);
nor U5849 (N_5849,N_5735,N_5647);
and U5850 (N_5850,N_5765,N_5706);
xnor U5851 (N_5851,N_5610,N_5698);
nand U5852 (N_5852,N_5600,N_5776);
xor U5853 (N_5853,N_5645,N_5757);
xnor U5854 (N_5854,N_5771,N_5741);
nand U5855 (N_5855,N_5758,N_5674);
xor U5856 (N_5856,N_5656,N_5636);
or U5857 (N_5857,N_5793,N_5652);
nor U5858 (N_5858,N_5738,N_5782);
and U5859 (N_5859,N_5615,N_5711);
or U5860 (N_5860,N_5649,N_5754);
or U5861 (N_5861,N_5739,N_5726);
nand U5862 (N_5862,N_5719,N_5787);
and U5863 (N_5863,N_5798,N_5602);
xor U5864 (N_5864,N_5653,N_5609);
and U5865 (N_5865,N_5607,N_5691);
nor U5866 (N_5866,N_5768,N_5778);
and U5867 (N_5867,N_5629,N_5752);
nand U5868 (N_5868,N_5799,N_5641);
and U5869 (N_5869,N_5724,N_5731);
nand U5870 (N_5870,N_5795,N_5705);
xnor U5871 (N_5871,N_5774,N_5791);
xnor U5872 (N_5872,N_5725,N_5677);
and U5873 (N_5873,N_5749,N_5611);
or U5874 (N_5874,N_5657,N_5670);
xnor U5875 (N_5875,N_5702,N_5664);
xor U5876 (N_5876,N_5742,N_5746);
nor U5877 (N_5877,N_5786,N_5796);
xnor U5878 (N_5878,N_5730,N_5761);
xor U5879 (N_5879,N_5716,N_5665);
xor U5880 (N_5880,N_5644,N_5625);
nor U5881 (N_5881,N_5764,N_5627);
nand U5882 (N_5882,N_5604,N_5743);
xnor U5883 (N_5883,N_5642,N_5631);
and U5884 (N_5884,N_5638,N_5703);
xor U5885 (N_5885,N_5720,N_5618);
and U5886 (N_5886,N_5712,N_5686);
and U5887 (N_5887,N_5619,N_5789);
and U5888 (N_5888,N_5684,N_5681);
nor U5889 (N_5889,N_5683,N_5737);
and U5890 (N_5890,N_5660,N_5729);
nor U5891 (N_5891,N_5687,N_5727);
xnor U5892 (N_5892,N_5784,N_5767);
and U5893 (N_5893,N_5628,N_5780);
nand U5894 (N_5894,N_5601,N_5633);
or U5895 (N_5895,N_5779,N_5748);
or U5896 (N_5896,N_5612,N_5669);
nor U5897 (N_5897,N_5753,N_5663);
nor U5898 (N_5898,N_5756,N_5760);
nand U5899 (N_5899,N_5790,N_5781);
nor U5900 (N_5900,N_5791,N_5700);
nor U5901 (N_5901,N_5615,N_5743);
nor U5902 (N_5902,N_5674,N_5608);
and U5903 (N_5903,N_5639,N_5797);
xnor U5904 (N_5904,N_5797,N_5667);
or U5905 (N_5905,N_5637,N_5795);
or U5906 (N_5906,N_5747,N_5603);
xor U5907 (N_5907,N_5785,N_5790);
and U5908 (N_5908,N_5628,N_5799);
nor U5909 (N_5909,N_5713,N_5662);
and U5910 (N_5910,N_5630,N_5662);
xnor U5911 (N_5911,N_5791,N_5635);
nor U5912 (N_5912,N_5710,N_5788);
xnor U5913 (N_5913,N_5762,N_5731);
xor U5914 (N_5914,N_5780,N_5614);
nand U5915 (N_5915,N_5746,N_5687);
nor U5916 (N_5916,N_5748,N_5657);
and U5917 (N_5917,N_5625,N_5749);
or U5918 (N_5918,N_5794,N_5695);
nor U5919 (N_5919,N_5761,N_5615);
or U5920 (N_5920,N_5653,N_5600);
nand U5921 (N_5921,N_5629,N_5775);
xnor U5922 (N_5922,N_5789,N_5621);
xnor U5923 (N_5923,N_5754,N_5759);
or U5924 (N_5924,N_5704,N_5765);
nor U5925 (N_5925,N_5741,N_5663);
or U5926 (N_5926,N_5739,N_5755);
nand U5927 (N_5927,N_5759,N_5771);
and U5928 (N_5928,N_5746,N_5704);
nand U5929 (N_5929,N_5678,N_5762);
nand U5930 (N_5930,N_5636,N_5777);
and U5931 (N_5931,N_5737,N_5754);
and U5932 (N_5932,N_5615,N_5782);
nor U5933 (N_5933,N_5761,N_5704);
xnor U5934 (N_5934,N_5650,N_5691);
or U5935 (N_5935,N_5665,N_5756);
nand U5936 (N_5936,N_5711,N_5716);
xnor U5937 (N_5937,N_5742,N_5644);
nor U5938 (N_5938,N_5628,N_5665);
nor U5939 (N_5939,N_5746,N_5664);
and U5940 (N_5940,N_5740,N_5710);
or U5941 (N_5941,N_5633,N_5773);
or U5942 (N_5942,N_5666,N_5691);
xor U5943 (N_5943,N_5783,N_5790);
nand U5944 (N_5944,N_5611,N_5680);
xor U5945 (N_5945,N_5618,N_5712);
nor U5946 (N_5946,N_5778,N_5766);
or U5947 (N_5947,N_5718,N_5781);
and U5948 (N_5948,N_5725,N_5628);
nand U5949 (N_5949,N_5653,N_5606);
and U5950 (N_5950,N_5667,N_5673);
nand U5951 (N_5951,N_5754,N_5752);
nor U5952 (N_5952,N_5652,N_5607);
nand U5953 (N_5953,N_5781,N_5752);
xnor U5954 (N_5954,N_5634,N_5601);
xor U5955 (N_5955,N_5632,N_5750);
or U5956 (N_5956,N_5676,N_5713);
nand U5957 (N_5957,N_5632,N_5793);
nand U5958 (N_5958,N_5626,N_5785);
or U5959 (N_5959,N_5712,N_5611);
and U5960 (N_5960,N_5650,N_5607);
nand U5961 (N_5961,N_5656,N_5642);
nor U5962 (N_5962,N_5761,N_5795);
nand U5963 (N_5963,N_5718,N_5746);
and U5964 (N_5964,N_5600,N_5618);
xor U5965 (N_5965,N_5701,N_5671);
and U5966 (N_5966,N_5632,N_5790);
nand U5967 (N_5967,N_5744,N_5740);
and U5968 (N_5968,N_5624,N_5633);
or U5969 (N_5969,N_5728,N_5638);
nand U5970 (N_5970,N_5633,N_5740);
xor U5971 (N_5971,N_5661,N_5708);
xor U5972 (N_5972,N_5689,N_5671);
nor U5973 (N_5973,N_5605,N_5638);
nor U5974 (N_5974,N_5767,N_5659);
and U5975 (N_5975,N_5683,N_5625);
nand U5976 (N_5976,N_5609,N_5691);
nor U5977 (N_5977,N_5770,N_5629);
and U5978 (N_5978,N_5795,N_5718);
nor U5979 (N_5979,N_5781,N_5697);
and U5980 (N_5980,N_5619,N_5730);
xor U5981 (N_5981,N_5644,N_5684);
or U5982 (N_5982,N_5606,N_5712);
nor U5983 (N_5983,N_5601,N_5738);
xor U5984 (N_5984,N_5736,N_5798);
nand U5985 (N_5985,N_5656,N_5671);
xnor U5986 (N_5986,N_5634,N_5680);
xnor U5987 (N_5987,N_5692,N_5604);
or U5988 (N_5988,N_5742,N_5652);
nor U5989 (N_5989,N_5751,N_5690);
or U5990 (N_5990,N_5762,N_5727);
nand U5991 (N_5991,N_5732,N_5735);
and U5992 (N_5992,N_5748,N_5745);
nand U5993 (N_5993,N_5632,N_5718);
nor U5994 (N_5994,N_5619,N_5701);
or U5995 (N_5995,N_5771,N_5691);
nor U5996 (N_5996,N_5629,N_5626);
and U5997 (N_5997,N_5748,N_5755);
nand U5998 (N_5998,N_5637,N_5666);
nor U5999 (N_5999,N_5794,N_5624);
nor U6000 (N_6000,N_5994,N_5952);
and U6001 (N_6001,N_5831,N_5967);
and U6002 (N_6002,N_5872,N_5867);
nand U6003 (N_6003,N_5855,N_5822);
nand U6004 (N_6004,N_5826,N_5815);
nor U6005 (N_6005,N_5887,N_5974);
nor U6006 (N_6006,N_5889,N_5847);
xnor U6007 (N_6007,N_5892,N_5875);
nand U6008 (N_6008,N_5921,N_5869);
xnor U6009 (N_6009,N_5836,N_5806);
and U6010 (N_6010,N_5947,N_5945);
nand U6011 (N_6011,N_5807,N_5919);
or U6012 (N_6012,N_5981,N_5810);
nor U6013 (N_6013,N_5963,N_5949);
or U6014 (N_6014,N_5844,N_5969);
and U6015 (N_6015,N_5894,N_5876);
nand U6016 (N_6016,N_5843,N_5902);
and U6017 (N_6017,N_5958,N_5828);
nor U6018 (N_6018,N_5837,N_5939);
nor U6019 (N_6019,N_5948,N_5870);
or U6020 (N_6020,N_5864,N_5917);
xor U6021 (N_6021,N_5951,N_5895);
or U6022 (N_6022,N_5931,N_5805);
or U6023 (N_6023,N_5907,N_5854);
nor U6024 (N_6024,N_5941,N_5922);
nor U6025 (N_6025,N_5834,N_5988);
nand U6026 (N_6026,N_5935,N_5818);
nor U6027 (N_6027,N_5842,N_5937);
nand U6028 (N_6028,N_5996,N_5986);
xor U6029 (N_6029,N_5962,N_5801);
and U6030 (N_6030,N_5804,N_5976);
nor U6031 (N_6031,N_5802,N_5888);
and U6032 (N_6032,N_5903,N_5874);
xor U6033 (N_6033,N_5978,N_5882);
xnor U6034 (N_6034,N_5929,N_5835);
nor U6035 (N_6035,N_5816,N_5954);
nand U6036 (N_6036,N_5838,N_5808);
nand U6037 (N_6037,N_5979,N_5860);
or U6038 (N_6038,N_5964,N_5823);
or U6039 (N_6039,N_5830,N_5977);
nand U6040 (N_6040,N_5857,N_5879);
or U6041 (N_6041,N_5925,N_5862);
and U6042 (N_6042,N_5944,N_5960);
xor U6043 (N_6043,N_5966,N_5881);
nor U6044 (N_6044,N_5914,N_5961);
xor U6045 (N_6045,N_5858,N_5953);
nand U6046 (N_6046,N_5871,N_5968);
xor U6047 (N_6047,N_5936,N_5861);
nor U6048 (N_6048,N_5908,N_5841);
nand U6049 (N_6049,N_5846,N_5965);
nor U6050 (N_6050,N_5800,N_5928);
or U6051 (N_6051,N_5901,N_5878);
xnor U6052 (N_6052,N_5814,N_5820);
or U6053 (N_6053,N_5900,N_5910);
or U6054 (N_6054,N_5918,N_5911);
or U6055 (N_6055,N_5856,N_5848);
or U6056 (N_6056,N_5817,N_5923);
xor U6057 (N_6057,N_5885,N_5975);
nor U6058 (N_6058,N_5859,N_5821);
or U6059 (N_6059,N_5991,N_5950);
or U6060 (N_6060,N_5896,N_5829);
xor U6061 (N_6061,N_5877,N_5956);
and U6062 (N_6062,N_5880,N_5839);
or U6063 (N_6063,N_5833,N_5970);
nand U6064 (N_6064,N_5819,N_5943);
nor U6065 (N_6065,N_5890,N_5825);
nand U6066 (N_6066,N_5811,N_5926);
or U6067 (N_6067,N_5930,N_5989);
xor U6068 (N_6068,N_5973,N_5924);
or U6069 (N_6069,N_5868,N_5985);
and U6070 (N_6070,N_5851,N_5997);
xnor U6071 (N_6071,N_5992,N_5852);
xor U6072 (N_6072,N_5809,N_5995);
nand U6073 (N_6073,N_5972,N_5840);
and U6074 (N_6074,N_5946,N_5942);
and U6075 (N_6075,N_5803,N_5933);
nor U6076 (N_6076,N_5827,N_5915);
or U6077 (N_6077,N_5980,N_5932);
nand U6078 (N_6078,N_5812,N_5916);
and U6079 (N_6079,N_5909,N_5883);
or U6080 (N_6080,N_5897,N_5959);
xor U6081 (N_6081,N_5866,N_5999);
xnor U6082 (N_6082,N_5853,N_5849);
and U6083 (N_6083,N_5993,N_5990);
and U6084 (N_6084,N_5845,N_5984);
or U6085 (N_6085,N_5955,N_5873);
or U6086 (N_6086,N_5983,N_5904);
xnor U6087 (N_6087,N_5927,N_5886);
xnor U6088 (N_6088,N_5905,N_5832);
and U6089 (N_6089,N_5899,N_5884);
xor U6090 (N_6090,N_5893,N_5934);
nor U6091 (N_6091,N_5998,N_5912);
or U6092 (N_6092,N_5824,N_5971);
nor U6093 (N_6093,N_5850,N_5987);
nor U6094 (N_6094,N_5913,N_5891);
xor U6095 (N_6095,N_5906,N_5865);
nand U6096 (N_6096,N_5813,N_5938);
and U6097 (N_6097,N_5863,N_5940);
and U6098 (N_6098,N_5957,N_5920);
or U6099 (N_6099,N_5982,N_5898);
nand U6100 (N_6100,N_5878,N_5945);
xnor U6101 (N_6101,N_5980,N_5960);
or U6102 (N_6102,N_5832,N_5840);
and U6103 (N_6103,N_5959,N_5961);
xnor U6104 (N_6104,N_5942,N_5906);
or U6105 (N_6105,N_5895,N_5875);
and U6106 (N_6106,N_5916,N_5962);
nand U6107 (N_6107,N_5861,N_5949);
or U6108 (N_6108,N_5801,N_5840);
or U6109 (N_6109,N_5982,N_5850);
nor U6110 (N_6110,N_5805,N_5824);
or U6111 (N_6111,N_5874,N_5996);
xor U6112 (N_6112,N_5960,N_5924);
and U6113 (N_6113,N_5938,N_5831);
nand U6114 (N_6114,N_5883,N_5856);
or U6115 (N_6115,N_5885,N_5812);
nor U6116 (N_6116,N_5951,N_5937);
nor U6117 (N_6117,N_5959,N_5819);
nand U6118 (N_6118,N_5878,N_5835);
or U6119 (N_6119,N_5826,N_5996);
or U6120 (N_6120,N_5870,N_5961);
and U6121 (N_6121,N_5924,N_5832);
nand U6122 (N_6122,N_5925,N_5921);
xnor U6123 (N_6123,N_5869,N_5955);
nand U6124 (N_6124,N_5899,N_5997);
nand U6125 (N_6125,N_5836,N_5809);
xnor U6126 (N_6126,N_5847,N_5863);
and U6127 (N_6127,N_5807,N_5834);
xnor U6128 (N_6128,N_5877,N_5998);
xor U6129 (N_6129,N_5924,N_5911);
xnor U6130 (N_6130,N_5942,N_5974);
and U6131 (N_6131,N_5958,N_5995);
xor U6132 (N_6132,N_5899,N_5875);
nand U6133 (N_6133,N_5869,N_5884);
or U6134 (N_6134,N_5878,N_5883);
nor U6135 (N_6135,N_5914,N_5990);
nand U6136 (N_6136,N_5930,N_5941);
and U6137 (N_6137,N_5925,N_5970);
nor U6138 (N_6138,N_5948,N_5802);
nor U6139 (N_6139,N_5884,N_5883);
and U6140 (N_6140,N_5978,N_5819);
and U6141 (N_6141,N_5849,N_5866);
nor U6142 (N_6142,N_5969,N_5965);
nand U6143 (N_6143,N_5906,N_5883);
or U6144 (N_6144,N_5966,N_5814);
xor U6145 (N_6145,N_5906,N_5987);
and U6146 (N_6146,N_5871,N_5903);
xor U6147 (N_6147,N_5867,N_5964);
or U6148 (N_6148,N_5980,N_5985);
xnor U6149 (N_6149,N_5951,N_5938);
and U6150 (N_6150,N_5952,N_5829);
and U6151 (N_6151,N_5931,N_5851);
xnor U6152 (N_6152,N_5845,N_5915);
and U6153 (N_6153,N_5950,N_5965);
nor U6154 (N_6154,N_5924,N_5895);
or U6155 (N_6155,N_5868,N_5973);
nor U6156 (N_6156,N_5961,N_5905);
and U6157 (N_6157,N_5944,N_5979);
and U6158 (N_6158,N_5878,N_5895);
or U6159 (N_6159,N_5988,N_5887);
and U6160 (N_6160,N_5946,N_5912);
nor U6161 (N_6161,N_5920,N_5871);
xnor U6162 (N_6162,N_5842,N_5800);
nor U6163 (N_6163,N_5894,N_5854);
nand U6164 (N_6164,N_5818,N_5937);
xnor U6165 (N_6165,N_5872,N_5974);
or U6166 (N_6166,N_5999,N_5921);
xnor U6167 (N_6167,N_5957,N_5922);
xnor U6168 (N_6168,N_5854,N_5944);
xor U6169 (N_6169,N_5838,N_5802);
nand U6170 (N_6170,N_5815,N_5821);
and U6171 (N_6171,N_5964,N_5955);
and U6172 (N_6172,N_5942,N_5858);
xnor U6173 (N_6173,N_5824,N_5801);
or U6174 (N_6174,N_5906,N_5837);
nor U6175 (N_6175,N_5952,N_5979);
xor U6176 (N_6176,N_5923,N_5879);
xor U6177 (N_6177,N_5981,N_5905);
nand U6178 (N_6178,N_5950,N_5879);
nor U6179 (N_6179,N_5802,N_5839);
or U6180 (N_6180,N_5932,N_5921);
or U6181 (N_6181,N_5835,N_5887);
nor U6182 (N_6182,N_5815,N_5832);
and U6183 (N_6183,N_5936,N_5871);
and U6184 (N_6184,N_5874,N_5843);
and U6185 (N_6185,N_5895,N_5954);
nand U6186 (N_6186,N_5876,N_5962);
xor U6187 (N_6187,N_5937,N_5919);
xnor U6188 (N_6188,N_5873,N_5989);
nor U6189 (N_6189,N_5942,N_5903);
xor U6190 (N_6190,N_5880,N_5844);
and U6191 (N_6191,N_5842,N_5910);
xnor U6192 (N_6192,N_5933,N_5970);
nand U6193 (N_6193,N_5808,N_5839);
xnor U6194 (N_6194,N_5905,N_5997);
nand U6195 (N_6195,N_5996,N_5959);
or U6196 (N_6196,N_5976,N_5863);
and U6197 (N_6197,N_5954,N_5958);
xnor U6198 (N_6198,N_5817,N_5965);
xnor U6199 (N_6199,N_5958,N_5939);
nand U6200 (N_6200,N_6113,N_6151);
xnor U6201 (N_6201,N_6178,N_6131);
nand U6202 (N_6202,N_6017,N_6195);
nor U6203 (N_6203,N_6123,N_6008);
nor U6204 (N_6204,N_6175,N_6191);
and U6205 (N_6205,N_6058,N_6062);
nor U6206 (N_6206,N_6009,N_6045);
or U6207 (N_6207,N_6019,N_6124);
nor U6208 (N_6208,N_6037,N_6091);
and U6209 (N_6209,N_6070,N_6032);
nor U6210 (N_6210,N_6159,N_6156);
and U6211 (N_6211,N_6161,N_6100);
nor U6212 (N_6212,N_6135,N_6134);
and U6213 (N_6213,N_6196,N_6075);
or U6214 (N_6214,N_6077,N_6160);
nand U6215 (N_6215,N_6104,N_6105);
nor U6216 (N_6216,N_6099,N_6038);
and U6217 (N_6217,N_6090,N_6164);
or U6218 (N_6218,N_6093,N_6048);
nand U6219 (N_6219,N_6116,N_6073);
nor U6220 (N_6220,N_6112,N_6013);
and U6221 (N_6221,N_6181,N_6106);
and U6222 (N_6222,N_6060,N_6173);
nand U6223 (N_6223,N_6168,N_6194);
xnor U6224 (N_6224,N_6051,N_6003);
or U6225 (N_6225,N_6197,N_6133);
nor U6226 (N_6226,N_6056,N_6170);
and U6227 (N_6227,N_6021,N_6001);
nand U6228 (N_6228,N_6066,N_6154);
xor U6229 (N_6229,N_6166,N_6057);
or U6230 (N_6230,N_6082,N_6031);
nor U6231 (N_6231,N_6087,N_6147);
or U6232 (N_6232,N_6030,N_6040);
nand U6233 (N_6233,N_6130,N_6086);
nor U6234 (N_6234,N_6169,N_6094);
nor U6235 (N_6235,N_6153,N_6046);
and U6236 (N_6236,N_6138,N_6177);
or U6237 (N_6237,N_6150,N_6121);
nand U6238 (N_6238,N_6149,N_6018);
and U6239 (N_6239,N_6050,N_6067);
or U6240 (N_6240,N_6182,N_6061);
nand U6241 (N_6241,N_6085,N_6127);
nand U6242 (N_6242,N_6010,N_6089);
or U6243 (N_6243,N_6141,N_6155);
nand U6244 (N_6244,N_6024,N_6176);
nand U6245 (N_6245,N_6078,N_6080);
xor U6246 (N_6246,N_6041,N_6006);
or U6247 (N_6247,N_6096,N_6126);
or U6248 (N_6248,N_6137,N_6110);
or U6249 (N_6249,N_6072,N_6083);
and U6250 (N_6250,N_6023,N_6095);
nor U6251 (N_6251,N_6068,N_6071);
nand U6252 (N_6252,N_6047,N_6189);
xnor U6253 (N_6253,N_6052,N_6199);
and U6254 (N_6254,N_6179,N_6055);
and U6255 (N_6255,N_6049,N_6117);
nor U6256 (N_6256,N_6042,N_6165);
nand U6257 (N_6257,N_6039,N_6102);
nand U6258 (N_6258,N_6184,N_6098);
and U6259 (N_6259,N_6188,N_6136);
nor U6260 (N_6260,N_6107,N_6081);
nand U6261 (N_6261,N_6064,N_6044);
and U6262 (N_6262,N_6174,N_6059);
or U6263 (N_6263,N_6092,N_6043);
and U6264 (N_6264,N_6016,N_6183);
xor U6265 (N_6265,N_6119,N_6022);
and U6266 (N_6266,N_6180,N_6146);
xor U6267 (N_6267,N_6012,N_6004);
xnor U6268 (N_6268,N_6167,N_6084);
nor U6269 (N_6269,N_6005,N_6109);
xnor U6270 (N_6270,N_6097,N_6139);
nand U6271 (N_6271,N_6114,N_6033);
and U6272 (N_6272,N_6198,N_6036);
nand U6273 (N_6273,N_6140,N_6088);
and U6274 (N_6274,N_6069,N_6035);
xnor U6275 (N_6275,N_6079,N_6186);
nand U6276 (N_6276,N_6108,N_6027);
or U6277 (N_6277,N_6193,N_6162);
and U6278 (N_6278,N_6128,N_6101);
and U6279 (N_6279,N_6007,N_6002);
nand U6280 (N_6280,N_6000,N_6025);
xor U6281 (N_6281,N_6163,N_6029);
nor U6282 (N_6282,N_6028,N_6158);
nand U6283 (N_6283,N_6063,N_6015);
nand U6284 (N_6284,N_6145,N_6011);
nor U6285 (N_6285,N_6122,N_6120);
and U6286 (N_6286,N_6103,N_6142);
xnor U6287 (N_6287,N_6115,N_6026);
xnor U6288 (N_6288,N_6034,N_6111);
nand U6289 (N_6289,N_6132,N_6125);
nor U6290 (N_6290,N_6190,N_6187);
xor U6291 (N_6291,N_6144,N_6171);
nor U6292 (N_6292,N_6192,N_6065);
xor U6293 (N_6293,N_6152,N_6054);
and U6294 (N_6294,N_6129,N_6014);
xnor U6295 (N_6295,N_6074,N_6076);
nor U6296 (N_6296,N_6185,N_6020);
and U6297 (N_6297,N_6143,N_6172);
nor U6298 (N_6298,N_6157,N_6053);
nand U6299 (N_6299,N_6148,N_6118);
and U6300 (N_6300,N_6071,N_6070);
or U6301 (N_6301,N_6046,N_6126);
xor U6302 (N_6302,N_6091,N_6056);
or U6303 (N_6303,N_6147,N_6054);
and U6304 (N_6304,N_6026,N_6053);
nor U6305 (N_6305,N_6074,N_6103);
and U6306 (N_6306,N_6073,N_6095);
xor U6307 (N_6307,N_6082,N_6129);
and U6308 (N_6308,N_6025,N_6122);
nand U6309 (N_6309,N_6183,N_6163);
nor U6310 (N_6310,N_6117,N_6064);
xor U6311 (N_6311,N_6177,N_6096);
and U6312 (N_6312,N_6083,N_6165);
xor U6313 (N_6313,N_6136,N_6012);
nor U6314 (N_6314,N_6184,N_6196);
nor U6315 (N_6315,N_6144,N_6083);
or U6316 (N_6316,N_6160,N_6125);
nand U6317 (N_6317,N_6017,N_6100);
nor U6318 (N_6318,N_6166,N_6086);
nor U6319 (N_6319,N_6032,N_6046);
or U6320 (N_6320,N_6049,N_6177);
nor U6321 (N_6321,N_6053,N_6149);
and U6322 (N_6322,N_6058,N_6102);
nand U6323 (N_6323,N_6123,N_6178);
nor U6324 (N_6324,N_6152,N_6032);
nand U6325 (N_6325,N_6012,N_6165);
nor U6326 (N_6326,N_6042,N_6144);
nor U6327 (N_6327,N_6013,N_6031);
and U6328 (N_6328,N_6190,N_6051);
nor U6329 (N_6329,N_6089,N_6189);
and U6330 (N_6330,N_6199,N_6097);
nand U6331 (N_6331,N_6000,N_6086);
or U6332 (N_6332,N_6110,N_6177);
or U6333 (N_6333,N_6070,N_6069);
or U6334 (N_6334,N_6016,N_6145);
or U6335 (N_6335,N_6191,N_6187);
nor U6336 (N_6336,N_6149,N_6190);
xor U6337 (N_6337,N_6188,N_6036);
nand U6338 (N_6338,N_6135,N_6138);
nand U6339 (N_6339,N_6182,N_6183);
and U6340 (N_6340,N_6038,N_6001);
nor U6341 (N_6341,N_6040,N_6025);
or U6342 (N_6342,N_6190,N_6113);
and U6343 (N_6343,N_6019,N_6132);
or U6344 (N_6344,N_6054,N_6174);
nand U6345 (N_6345,N_6019,N_6174);
or U6346 (N_6346,N_6175,N_6092);
nor U6347 (N_6347,N_6068,N_6014);
xor U6348 (N_6348,N_6197,N_6056);
nor U6349 (N_6349,N_6143,N_6128);
nand U6350 (N_6350,N_6143,N_6119);
or U6351 (N_6351,N_6159,N_6058);
nand U6352 (N_6352,N_6080,N_6164);
xor U6353 (N_6353,N_6022,N_6061);
nor U6354 (N_6354,N_6035,N_6002);
nand U6355 (N_6355,N_6000,N_6103);
nand U6356 (N_6356,N_6062,N_6037);
xor U6357 (N_6357,N_6047,N_6155);
nor U6358 (N_6358,N_6069,N_6118);
or U6359 (N_6359,N_6042,N_6189);
or U6360 (N_6360,N_6102,N_6135);
xnor U6361 (N_6361,N_6094,N_6119);
nor U6362 (N_6362,N_6038,N_6170);
xnor U6363 (N_6363,N_6133,N_6189);
or U6364 (N_6364,N_6090,N_6163);
nor U6365 (N_6365,N_6047,N_6091);
nor U6366 (N_6366,N_6084,N_6061);
xnor U6367 (N_6367,N_6065,N_6144);
nor U6368 (N_6368,N_6129,N_6093);
xor U6369 (N_6369,N_6144,N_6020);
xor U6370 (N_6370,N_6063,N_6199);
nand U6371 (N_6371,N_6144,N_6103);
and U6372 (N_6372,N_6059,N_6019);
and U6373 (N_6373,N_6060,N_6050);
and U6374 (N_6374,N_6150,N_6088);
or U6375 (N_6375,N_6104,N_6078);
nor U6376 (N_6376,N_6193,N_6025);
nor U6377 (N_6377,N_6179,N_6029);
or U6378 (N_6378,N_6196,N_6174);
xnor U6379 (N_6379,N_6136,N_6016);
or U6380 (N_6380,N_6155,N_6006);
or U6381 (N_6381,N_6036,N_6006);
or U6382 (N_6382,N_6049,N_6005);
nor U6383 (N_6383,N_6116,N_6049);
or U6384 (N_6384,N_6196,N_6050);
or U6385 (N_6385,N_6155,N_6044);
or U6386 (N_6386,N_6005,N_6146);
nand U6387 (N_6387,N_6041,N_6102);
nor U6388 (N_6388,N_6021,N_6003);
nor U6389 (N_6389,N_6141,N_6072);
and U6390 (N_6390,N_6127,N_6011);
and U6391 (N_6391,N_6169,N_6051);
and U6392 (N_6392,N_6145,N_6074);
or U6393 (N_6393,N_6058,N_6017);
xor U6394 (N_6394,N_6178,N_6124);
and U6395 (N_6395,N_6084,N_6023);
and U6396 (N_6396,N_6164,N_6177);
xor U6397 (N_6397,N_6029,N_6189);
and U6398 (N_6398,N_6112,N_6000);
and U6399 (N_6399,N_6071,N_6089);
xnor U6400 (N_6400,N_6280,N_6319);
nand U6401 (N_6401,N_6251,N_6262);
nor U6402 (N_6402,N_6352,N_6382);
and U6403 (N_6403,N_6227,N_6293);
nor U6404 (N_6404,N_6397,N_6351);
and U6405 (N_6405,N_6266,N_6278);
or U6406 (N_6406,N_6252,N_6288);
and U6407 (N_6407,N_6313,N_6222);
nand U6408 (N_6408,N_6249,N_6343);
nand U6409 (N_6409,N_6215,N_6205);
xor U6410 (N_6410,N_6396,N_6250);
and U6411 (N_6411,N_6289,N_6349);
or U6412 (N_6412,N_6243,N_6208);
xor U6413 (N_6413,N_6388,N_6223);
nand U6414 (N_6414,N_6314,N_6360);
nand U6415 (N_6415,N_6300,N_6338);
nand U6416 (N_6416,N_6342,N_6204);
and U6417 (N_6417,N_6332,N_6391);
nand U6418 (N_6418,N_6380,N_6206);
nor U6419 (N_6419,N_6221,N_6274);
xnor U6420 (N_6420,N_6202,N_6261);
and U6421 (N_6421,N_6348,N_6375);
nand U6422 (N_6422,N_6372,N_6231);
nor U6423 (N_6423,N_6290,N_6269);
and U6424 (N_6424,N_6233,N_6350);
or U6425 (N_6425,N_6385,N_6246);
or U6426 (N_6426,N_6329,N_6253);
nand U6427 (N_6427,N_6307,N_6347);
nand U6428 (N_6428,N_6317,N_6230);
nor U6429 (N_6429,N_6209,N_6239);
or U6430 (N_6430,N_6341,N_6268);
xor U6431 (N_6431,N_6257,N_6229);
xnor U6432 (N_6432,N_6273,N_6379);
xor U6433 (N_6433,N_6287,N_6285);
or U6434 (N_6434,N_6294,N_6308);
and U6435 (N_6435,N_6245,N_6299);
or U6436 (N_6436,N_6399,N_6366);
or U6437 (N_6437,N_6258,N_6217);
and U6438 (N_6438,N_6296,N_6345);
nand U6439 (N_6439,N_6241,N_6256);
xor U6440 (N_6440,N_6331,N_6359);
nor U6441 (N_6441,N_6254,N_6364);
xor U6442 (N_6442,N_6376,N_6298);
nor U6443 (N_6443,N_6395,N_6270);
or U6444 (N_6444,N_6235,N_6312);
nand U6445 (N_6445,N_6301,N_6377);
and U6446 (N_6446,N_6276,N_6327);
xor U6447 (N_6447,N_6247,N_6295);
and U6448 (N_6448,N_6219,N_6302);
and U6449 (N_6449,N_6369,N_6212);
and U6450 (N_6450,N_6333,N_6381);
nand U6451 (N_6451,N_6207,N_6303);
xor U6452 (N_6452,N_6218,N_6267);
nor U6453 (N_6453,N_6226,N_6330);
xnor U6454 (N_6454,N_6390,N_6370);
or U6455 (N_6455,N_6322,N_6200);
xnor U6456 (N_6456,N_6255,N_6335);
nor U6457 (N_6457,N_6384,N_6292);
xor U6458 (N_6458,N_6281,N_6387);
nand U6459 (N_6459,N_6318,N_6225);
and U6460 (N_6460,N_6279,N_6311);
nand U6461 (N_6461,N_6236,N_6220);
nor U6462 (N_6462,N_6373,N_6260);
or U6463 (N_6463,N_6357,N_6284);
xnor U6464 (N_6464,N_6326,N_6334);
or U6465 (N_6465,N_6328,N_6392);
nor U6466 (N_6466,N_6201,N_6323);
and U6467 (N_6467,N_6356,N_6378);
and U6468 (N_6468,N_6363,N_6367);
nand U6469 (N_6469,N_6259,N_6358);
nand U6470 (N_6470,N_6232,N_6337);
and U6471 (N_6471,N_6310,N_6271);
nand U6472 (N_6472,N_6210,N_6216);
or U6473 (N_6473,N_6316,N_6354);
xor U6474 (N_6474,N_6211,N_6365);
nor U6475 (N_6475,N_6355,N_6304);
nor U6476 (N_6476,N_6265,N_6306);
nand U6477 (N_6477,N_6240,N_6393);
or U6478 (N_6478,N_6234,N_6321);
nand U6479 (N_6479,N_6368,N_6346);
nand U6480 (N_6480,N_6325,N_6336);
and U6481 (N_6481,N_6353,N_6248);
nor U6482 (N_6482,N_6228,N_6242);
xnor U6483 (N_6483,N_6320,N_6339);
and U6484 (N_6484,N_6275,N_6291);
nand U6485 (N_6485,N_6224,N_6383);
xnor U6486 (N_6486,N_6386,N_6374);
and U6487 (N_6487,N_6237,N_6315);
xnor U6488 (N_6488,N_6309,N_6244);
and U6489 (N_6489,N_6297,N_6340);
xor U6490 (N_6490,N_6282,N_6394);
xor U6491 (N_6491,N_6203,N_6214);
nor U6492 (N_6492,N_6263,N_6389);
nand U6493 (N_6493,N_6213,N_6305);
nand U6494 (N_6494,N_6362,N_6361);
nand U6495 (N_6495,N_6272,N_6324);
nand U6496 (N_6496,N_6238,N_6371);
or U6497 (N_6497,N_6398,N_6283);
or U6498 (N_6498,N_6344,N_6277);
and U6499 (N_6499,N_6264,N_6286);
and U6500 (N_6500,N_6383,N_6262);
nor U6501 (N_6501,N_6258,N_6389);
and U6502 (N_6502,N_6377,N_6388);
xor U6503 (N_6503,N_6266,N_6296);
nand U6504 (N_6504,N_6234,N_6242);
xnor U6505 (N_6505,N_6282,N_6379);
xor U6506 (N_6506,N_6305,N_6389);
nand U6507 (N_6507,N_6356,N_6264);
or U6508 (N_6508,N_6224,N_6359);
or U6509 (N_6509,N_6367,N_6249);
xor U6510 (N_6510,N_6252,N_6345);
and U6511 (N_6511,N_6293,N_6325);
xor U6512 (N_6512,N_6220,N_6267);
and U6513 (N_6513,N_6204,N_6218);
or U6514 (N_6514,N_6305,N_6216);
nand U6515 (N_6515,N_6329,N_6394);
nor U6516 (N_6516,N_6308,N_6255);
nand U6517 (N_6517,N_6202,N_6391);
nor U6518 (N_6518,N_6273,N_6251);
nand U6519 (N_6519,N_6332,N_6288);
or U6520 (N_6520,N_6269,N_6340);
nand U6521 (N_6521,N_6377,N_6290);
nor U6522 (N_6522,N_6287,N_6335);
xor U6523 (N_6523,N_6238,N_6237);
and U6524 (N_6524,N_6203,N_6385);
nor U6525 (N_6525,N_6258,N_6247);
nor U6526 (N_6526,N_6299,N_6395);
nor U6527 (N_6527,N_6357,N_6216);
nor U6528 (N_6528,N_6304,N_6311);
nor U6529 (N_6529,N_6241,N_6324);
xnor U6530 (N_6530,N_6373,N_6355);
nand U6531 (N_6531,N_6226,N_6249);
nand U6532 (N_6532,N_6281,N_6299);
and U6533 (N_6533,N_6370,N_6330);
or U6534 (N_6534,N_6314,N_6384);
nand U6535 (N_6535,N_6397,N_6264);
xnor U6536 (N_6536,N_6280,N_6203);
nor U6537 (N_6537,N_6263,N_6313);
xnor U6538 (N_6538,N_6299,N_6340);
nand U6539 (N_6539,N_6237,N_6301);
xnor U6540 (N_6540,N_6244,N_6242);
nand U6541 (N_6541,N_6298,N_6310);
nor U6542 (N_6542,N_6353,N_6355);
or U6543 (N_6543,N_6364,N_6325);
nor U6544 (N_6544,N_6315,N_6338);
or U6545 (N_6545,N_6308,N_6324);
or U6546 (N_6546,N_6222,N_6203);
nor U6547 (N_6547,N_6251,N_6310);
nand U6548 (N_6548,N_6280,N_6317);
and U6549 (N_6549,N_6319,N_6323);
or U6550 (N_6550,N_6292,N_6210);
and U6551 (N_6551,N_6246,N_6337);
or U6552 (N_6552,N_6351,N_6337);
nor U6553 (N_6553,N_6220,N_6264);
nor U6554 (N_6554,N_6352,N_6240);
nor U6555 (N_6555,N_6380,N_6347);
and U6556 (N_6556,N_6289,N_6219);
nor U6557 (N_6557,N_6313,N_6334);
and U6558 (N_6558,N_6361,N_6374);
nand U6559 (N_6559,N_6233,N_6223);
nand U6560 (N_6560,N_6325,N_6275);
or U6561 (N_6561,N_6282,N_6375);
xor U6562 (N_6562,N_6350,N_6322);
nand U6563 (N_6563,N_6208,N_6235);
and U6564 (N_6564,N_6223,N_6358);
nand U6565 (N_6565,N_6251,N_6386);
and U6566 (N_6566,N_6228,N_6371);
xor U6567 (N_6567,N_6223,N_6361);
nand U6568 (N_6568,N_6207,N_6298);
and U6569 (N_6569,N_6243,N_6382);
xor U6570 (N_6570,N_6229,N_6296);
or U6571 (N_6571,N_6272,N_6363);
or U6572 (N_6572,N_6219,N_6331);
xor U6573 (N_6573,N_6325,N_6366);
nor U6574 (N_6574,N_6205,N_6397);
xor U6575 (N_6575,N_6251,N_6256);
xnor U6576 (N_6576,N_6327,N_6207);
nor U6577 (N_6577,N_6292,N_6345);
xnor U6578 (N_6578,N_6270,N_6358);
or U6579 (N_6579,N_6350,N_6263);
or U6580 (N_6580,N_6236,N_6345);
or U6581 (N_6581,N_6335,N_6390);
nor U6582 (N_6582,N_6265,N_6336);
nand U6583 (N_6583,N_6358,N_6249);
or U6584 (N_6584,N_6262,N_6212);
nand U6585 (N_6585,N_6297,N_6319);
and U6586 (N_6586,N_6303,N_6240);
or U6587 (N_6587,N_6276,N_6347);
nand U6588 (N_6588,N_6347,N_6363);
or U6589 (N_6589,N_6344,N_6332);
xor U6590 (N_6590,N_6354,N_6372);
xnor U6591 (N_6591,N_6284,N_6347);
or U6592 (N_6592,N_6231,N_6281);
or U6593 (N_6593,N_6352,N_6262);
xnor U6594 (N_6594,N_6204,N_6341);
nand U6595 (N_6595,N_6396,N_6293);
nand U6596 (N_6596,N_6368,N_6264);
and U6597 (N_6597,N_6211,N_6389);
xor U6598 (N_6598,N_6373,N_6364);
and U6599 (N_6599,N_6260,N_6366);
or U6600 (N_6600,N_6416,N_6559);
nand U6601 (N_6601,N_6440,N_6545);
xor U6602 (N_6602,N_6422,N_6549);
nand U6603 (N_6603,N_6448,N_6496);
xor U6604 (N_6604,N_6513,N_6443);
nand U6605 (N_6605,N_6522,N_6525);
xnor U6606 (N_6606,N_6578,N_6592);
nand U6607 (N_6607,N_6480,N_6433);
xor U6608 (N_6608,N_6573,N_6519);
xor U6609 (N_6609,N_6420,N_6451);
nand U6610 (N_6610,N_6555,N_6491);
nor U6611 (N_6611,N_6537,N_6521);
nor U6612 (N_6612,N_6450,N_6484);
nor U6613 (N_6613,N_6591,N_6483);
xor U6614 (N_6614,N_6517,N_6575);
xnor U6615 (N_6615,N_6438,N_6577);
nand U6616 (N_6616,N_6539,N_6447);
nor U6617 (N_6617,N_6427,N_6572);
nand U6618 (N_6618,N_6586,N_6479);
xnor U6619 (N_6619,N_6478,N_6583);
or U6620 (N_6620,N_6538,N_6401);
or U6621 (N_6621,N_6454,N_6404);
and U6622 (N_6622,N_6441,N_6528);
and U6623 (N_6623,N_6520,N_6518);
nand U6624 (N_6624,N_6400,N_6485);
or U6625 (N_6625,N_6547,N_6426);
nand U6626 (N_6626,N_6506,N_6557);
nor U6627 (N_6627,N_6511,N_6567);
nor U6628 (N_6628,N_6501,N_6482);
xor U6629 (N_6629,N_6546,N_6424);
and U6630 (N_6630,N_6411,N_6526);
nor U6631 (N_6631,N_6588,N_6507);
nor U6632 (N_6632,N_6468,N_6428);
nand U6633 (N_6633,N_6530,N_6524);
and U6634 (N_6634,N_6434,N_6498);
nor U6635 (N_6635,N_6556,N_6599);
nand U6636 (N_6636,N_6534,N_6477);
nand U6637 (N_6637,N_6446,N_6500);
and U6638 (N_6638,N_6488,N_6475);
nand U6639 (N_6639,N_6492,N_6445);
or U6640 (N_6640,N_6570,N_6565);
or U6641 (N_6641,N_6571,N_6579);
or U6642 (N_6642,N_6505,N_6429);
xnor U6643 (N_6643,N_6412,N_6514);
or U6644 (N_6644,N_6452,N_6512);
xnor U6645 (N_6645,N_6435,N_6541);
or U6646 (N_6646,N_6405,N_6561);
and U6647 (N_6647,N_6402,N_6408);
nor U6648 (N_6648,N_6563,N_6516);
nand U6649 (N_6649,N_6499,N_6403);
nor U6650 (N_6650,N_6457,N_6407);
nor U6651 (N_6651,N_6535,N_6533);
or U6652 (N_6652,N_6560,N_6470);
or U6653 (N_6653,N_6585,N_6410);
nor U6654 (N_6654,N_6504,N_6460);
or U6655 (N_6655,N_6596,N_6423);
xor U6656 (N_6656,N_6473,N_6487);
or U6657 (N_6657,N_6515,N_6406);
nor U6658 (N_6658,N_6439,N_6471);
nor U6659 (N_6659,N_6493,N_6510);
or U6660 (N_6660,N_6432,N_6568);
xor U6661 (N_6661,N_6464,N_6414);
xor U6662 (N_6662,N_6574,N_6540);
nand U6663 (N_6663,N_6474,N_6497);
and U6664 (N_6664,N_6461,N_6564);
nand U6665 (N_6665,N_6542,N_6436);
xor U6666 (N_6666,N_6589,N_6430);
xnor U6667 (N_6667,N_6467,N_6503);
xor U6668 (N_6668,N_6544,N_6466);
xor U6669 (N_6669,N_6486,N_6459);
xor U6670 (N_6670,N_6529,N_6469);
nor U6671 (N_6671,N_6417,N_6431);
xnor U6672 (N_6672,N_6550,N_6508);
nor U6673 (N_6673,N_6581,N_6598);
nor U6674 (N_6674,N_6543,N_6553);
nand U6675 (N_6675,N_6409,N_6595);
and U6676 (N_6676,N_6523,N_6593);
nor U6677 (N_6677,N_6548,N_6421);
and U6678 (N_6678,N_6554,N_6536);
nand U6679 (N_6679,N_6456,N_6444);
nand U6680 (N_6680,N_6552,N_6415);
nor U6681 (N_6681,N_6476,N_6495);
nor U6682 (N_6682,N_6437,N_6442);
nor U6683 (N_6683,N_6413,N_6558);
or U6684 (N_6684,N_6590,N_6582);
nor U6685 (N_6685,N_6472,N_6566);
nand U6686 (N_6686,N_6453,N_6458);
nor U6687 (N_6687,N_6465,N_6481);
xnor U6688 (N_6688,N_6449,N_6419);
nor U6689 (N_6689,N_6594,N_6597);
and U6690 (N_6690,N_6490,N_6455);
nand U6691 (N_6691,N_6562,N_6502);
nor U6692 (N_6692,N_6532,N_6551);
and U6693 (N_6693,N_6584,N_6494);
xor U6694 (N_6694,N_6509,N_6418);
or U6695 (N_6695,N_6462,N_6576);
xnor U6696 (N_6696,N_6527,N_6489);
and U6697 (N_6697,N_6587,N_6463);
nor U6698 (N_6698,N_6425,N_6569);
nor U6699 (N_6699,N_6580,N_6531);
nor U6700 (N_6700,N_6544,N_6478);
nor U6701 (N_6701,N_6442,N_6592);
xor U6702 (N_6702,N_6463,N_6593);
xnor U6703 (N_6703,N_6577,N_6495);
or U6704 (N_6704,N_6419,N_6414);
nor U6705 (N_6705,N_6456,N_6539);
and U6706 (N_6706,N_6465,N_6417);
or U6707 (N_6707,N_6539,N_6469);
nor U6708 (N_6708,N_6405,N_6594);
nand U6709 (N_6709,N_6571,N_6432);
and U6710 (N_6710,N_6491,N_6424);
xnor U6711 (N_6711,N_6490,N_6405);
nor U6712 (N_6712,N_6430,N_6572);
or U6713 (N_6713,N_6538,N_6593);
and U6714 (N_6714,N_6573,N_6452);
and U6715 (N_6715,N_6449,N_6590);
and U6716 (N_6716,N_6513,N_6570);
nor U6717 (N_6717,N_6403,N_6468);
or U6718 (N_6718,N_6437,N_6405);
nor U6719 (N_6719,N_6525,N_6419);
or U6720 (N_6720,N_6559,N_6583);
and U6721 (N_6721,N_6427,N_6458);
xor U6722 (N_6722,N_6535,N_6434);
and U6723 (N_6723,N_6426,N_6574);
nor U6724 (N_6724,N_6515,N_6577);
nor U6725 (N_6725,N_6496,N_6454);
or U6726 (N_6726,N_6447,N_6513);
and U6727 (N_6727,N_6545,N_6429);
or U6728 (N_6728,N_6483,N_6508);
or U6729 (N_6729,N_6451,N_6433);
or U6730 (N_6730,N_6516,N_6583);
nand U6731 (N_6731,N_6423,N_6537);
nor U6732 (N_6732,N_6427,N_6448);
and U6733 (N_6733,N_6524,N_6401);
nand U6734 (N_6734,N_6573,N_6492);
nor U6735 (N_6735,N_6565,N_6422);
or U6736 (N_6736,N_6573,N_6461);
xnor U6737 (N_6737,N_6440,N_6573);
nand U6738 (N_6738,N_6426,N_6464);
nand U6739 (N_6739,N_6586,N_6492);
or U6740 (N_6740,N_6474,N_6565);
nor U6741 (N_6741,N_6425,N_6528);
nor U6742 (N_6742,N_6509,N_6535);
nand U6743 (N_6743,N_6516,N_6512);
xnor U6744 (N_6744,N_6466,N_6546);
nand U6745 (N_6745,N_6573,N_6403);
nor U6746 (N_6746,N_6458,N_6404);
and U6747 (N_6747,N_6447,N_6419);
nand U6748 (N_6748,N_6553,N_6540);
nand U6749 (N_6749,N_6450,N_6589);
nand U6750 (N_6750,N_6440,N_6492);
xor U6751 (N_6751,N_6410,N_6589);
and U6752 (N_6752,N_6492,N_6469);
nor U6753 (N_6753,N_6566,N_6401);
nor U6754 (N_6754,N_6541,N_6544);
or U6755 (N_6755,N_6461,N_6551);
or U6756 (N_6756,N_6471,N_6487);
nor U6757 (N_6757,N_6532,N_6412);
or U6758 (N_6758,N_6488,N_6410);
xnor U6759 (N_6759,N_6541,N_6566);
nand U6760 (N_6760,N_6463,N_6415);
nand U6761 (N_6761,N_6568,N_6464);
or U6762 (N_6762,N_6435,N_6462);
or U6763 (N_6763,N_6432,N_6539);
xnor U6764 (N_6764,N_6426,N_6541);
nand U6765 (N_6765,N_6581,N_6521);
xnor U6766 (N_6766,N_6469,N_6561);
nand U6767 (N_6767,N_6597,N_6482);
nand U6768 (N_6768,N_6483,N_6422);
xor U6769 (N_6769,N_6564,N_6574);
nor U6770 (N_6770,N_6555,N_6559);
xnor U6771 (N_6771,N_6493,N_6492);
nor U6772 (N_6772,N_6508,N_6461);
or U6773 (N_6773,N_6453,N_6466);
xnor U6774 (N_6774,N_6466,N_6419);
or U6775 (N_6775,N_6595,N_6530);
nand U6776 (N_6776,N_6465,N_6489);
xnor U6777 (N_6777,N_6546,N_6501);
or U6778 (N_6778,N_6502,N_6465);
and U6779 (N_6779,N_6555,N_6472);
or U6780 (N_6780,N_6520,N_6410);
nor U6781 (N_6781,N_6586,N_6429);
xor U6782 (N_6782,N_6547,N_6596);
nor U6783 (N_6783,N_6440,N_6455);
and U6784 (N_6784,N_6408,N_6559);
nor U6785 (N_6785,N_6527,N_6417);
or U6786 (N_6786,N_6490,N_6565);
xor U6787 (N_6787,N_6414,N_6448);
and U6788 (N_6788,N_6410,N_6534);
or U6789 (N_6789,N_6579,N_6500);
xnor U6790 (N_6790,N_6500,N_6582);
nor U6791 (N_6791,N_6584,N_6462);
nor U6792 (N_6792,N_6510,N_6547);
xnor U6793 (N_6793,N_6445,N_6433);
and U6794 (N_6794,N_6412,N_6513);
nor U6795 (N_6795,N_6425,N_6538);
or U6796 (N_6796,N_6546,N_6547);
and U6797 (N_6797,N_6492,N_6520);
nand U6798 (N_6798,N_6481,N_6539);
and U6799 (N_6799,N_6527,N_6524);
xnor U6800 (N_6800,N_6682,N_6768);
nand U6801 (N_6801,N_6631,N_6688);
and U6802 (N_6802,N_6755,N_6794);
and U6803 (N_6803,N_6616,N_6767);
and U6804 (N_6804,N_6704,N_6729);
nand U6805 (N_6805,N_6748,N_6732);
and U6806 (N_6806,N_6776,N_6617);
nand U6807 (N_6807,N_6698,N_6774);
nor U6808 (N_6808,N_6654,N_6670);
nor U6809 (N_6809,N_6763,N_6797);
xor U6810 (N_6810,N_6653,N_6675);
and U6811 (N_6811,N_6745,N_6714);
nor U6812 (N_6812,N_6666,N_6657);
xnor U6813 (N_6813,N_6671,N_6697);
nand U6814 (N_6814,N_6636,N_6790);
xnor U6815 (N_6815,N_6798,N_6614);
nor U6816 (N_6816,N_6681,N_6601);
or U6817 (N_6817,N_6751,N_6730);
xor U6818 (N_6818,N_6652,N_6679);
xnor U6819 (N_6819,N_6620,N_6693);
xor U6820 (N_6820,N_6765,N_6735);
and U6821 (N_6821,N_6695,N_6685);
xnor U6822 (N_6822,N_6626,N_6749);
and U6823 (N_6823,N_6739,N_6660);
and U6824 (N_6824,N_6773,N_6750);
xor U6825 (N_6825,N_6686,N_6766);
or U6826 (N_6826,N_6761,N_6771);
and U6827 (N_6827,N_6702,N_6658);
and U6828 (N_6828,N_6721,N_6689);
xnor U6829 (N_6829,N_6613,N_6777);
xnor U6830 (N_6830,N_6646,N_6612);
nand U6831 (N_6831,N_6703,N_6677);
nand U6832 (N_6832,N_6605,N_6788);
nor U6833 (N_6833,N_6778,N_6651);
or U6834 (N_6834,N_6673,N_6785);
or U6835 (N_6835,N_6710,N_6661);
nor U6836 (N_6836,N_6608,N_6764);
and U6837 (N_6837,N_6705,N_6731);
or U6838 (N_6838,N_6604,N_6784);
xor U6839 (N_6839,N_6602,N_6726);
or U6840 (N_6840,N_6725,N_6779);
and U6841 (N_6841,N_6753,N_6734);
nand U6842 (N_6842,N_6722,N_6648);
xor U6843 (N_6843,N_6706,N_6647);
xor U6844 (N_6844,N_6700,N_6793);
or U6845 (N_6845,N_6720,N_6772);
and U6846 (N_6846,N_6629,N_6709);
nor U6847 (N_6847,N_6684,N_6775);
xor U6848 (N_6848,N_6638,N_6787);
and U6849 (N_6849,N_6611,N_6633);
xor U6850 (N_6850,N_6667,N_6759);
or U6851 (N_6851,N_6719,N_6795);
or U6852 (N_6852,N_6770,N_6786);
and U6853 (N_6853,N_6740,N_6606);
xnor U6854 (N_6854,N_6643,N_6712);
nor U6855 (N_6855,N_6783,N_6746);
nor U6856 (N_6856,N_6644,N_6780);
and U6857 (N_6857,N_6758,N_6760);
nor U6858 (N_6858,N_6727,N_6649);
xnor U6859 (N_6859,N_6799,N_6756);
or U6860 (N_6860,N_6610,N_6639);
xnor U6861 (N_6861,N_6607,N_6630);
xor U6862 (N_6862,N_6669,N_6680);
nand U6863 (N_6863,N_6792,N_6628);
xor U6864 (N_6864,N_6664,N_6694);
or U6865 (N_6865,N_6713,N_6736);
or U6866 (N_6866,N_6641,N_6665);
and U6867 (N_6867,N_6747,N_6627);
nor U6868 (N_6868,N_6662,N_6623);
nand U6869 (N_6869,N_6655,N_6621);
nor U6870 (N_6870,N_6796,N_6656);
or U6871 (N_6871,N_6782,N_6738);
nand U6872 (N_6872,N_6741,N_6687);
nand U6873 (N_6873,N_6659,N_6691);
xnor U6874 (N_6874,N_6615,N_6622);
nand U6875 (N_6875,N_6692,N_6690);
or U6876 (N_6876,N_6625,N_6603);
and U6877 (N_6877,N_6737,N_6733);
or U6878 (N_6878,N_6619,N_6663);
or U6879 (N_6879,N_6683,N_6716);
nand U6880 (N_6880,N_6743,N_6781);
nand U6881 (N_6881,N_6637,N_6600);
nand U6882 (N_6882,N_6618,N_6717);
xnor U6883 (N_6883,N_6645,N_6676);
nor U6884 (N_6884,N_6752,N_6744);
or U6885 (N_6885,N_6668,N_6715);
nor U6886 (N_6886,N_6707,N_6757);
or U6887 (N_6887,N_6789,N_6699);
and U6888 (N_6888,N_6672,N_6708);
and U6889 (N_6889,N_6724,N_6718);
xnor U6890 (N_6890,N_6650,N_6728);
nor U6891 (N_6891,N_6635,N_6609);
xor U6892 (N_6892,N_6754,N_6632);
nand U6893 (N_6893,N_6696,N_6640);
xor U6894 (N_6894,N_6624,N_6791);
nor U6895 (N_6895,N_6701,N_6742);
xnor U6896 (N_6896,N_6678,N_6723);
or U6897 (N_6897,N_6762,N_6642);
xor U6898 (N_6898,N_6769,N_6634);
nor U6899 (N_6899,N_6711,N_6674);
nand U6900 (N_6900,N_6734,N_6789);
and U6901 (N_6901,N_6605,N_6765);
and U6902 (N_6902,N_6762,N_6739);
nor U6903 (N_6903,N_6731,N_6631);
nor U6904 (N_6904,N_6746,N_6734);
nand U6905 (N_6905,N_6623,N_6729);
and U6906 (N_6906,N_6632,N_6782);
xor U6907 (N_6907,N_6717,N_6749);
or U6908 (N_6908,N_6759,N_6668);
xor U6909 (N_6909,N_6690,N_6714);
or U6910 (N_6910,N_6703,N_6788);
nand U6911 (N_6911,N_6675,N_6710);
or U6912 (N_6912,N_6654,N_6774);
nand U6913 (N_6913,N_6784,N_6699);
xnor U6914 (N_6914,N_6627,N_6601);
and U6915 (N_6915,N_6798,N_6700);
and U6916 (N_6916,N_6738,N_6713);
nor U6917 (N_6917,N_6700,N_6671);
nor U6918 (N_6918,N_6686,N_6779);
nand U6919 (N_6919,N_6738,N_6652);
or U6920 (N_6920,N_6614,N_6725);
or U6921 (N_6921,N_6635,N_6641);
xnor U6922 (N_6922,N_6651,N_6694);
or U6923 (N_6923,N_6757,N_6621);
and U6924 (N_6924,N_6720,N_6736);
nand U6925 (N_6925,N_6672,N_6610);
and U6926 (N_6926,N_6757,N_6620);
nor U6927 (N_6927,N_6659,N_6776);
xor U6928 (N_6928,N_6685,N_6772);
xor U6929 (N_6929,N_6731,N_6748);
nand U6930 (N_6930,N_6690,N_6740);
and U6931 (N_6931,N_6782,N_6787);
nand U6932 (N_6932,N_6728,N_6780);
xnor U6933 (N_6933,N_6646,N_6651);
or U6934 (N_6934,N_6681,N_6690);
nand U6935 (N_6935,N_6638,N_6620);
nand U6936 (N_6936,N_6644,N_6683);
nand U6937 (N_6937,N_6643,N_6753);
and U6938 (N_6938,N_6720,N_6604);
xnor U6939 (N_6939,N_6713,N_6711);
nand U6940 (N_6940,N_6762,N_6682);
and U6941 (N_6941,N_6655,N_6657);
nor U6942 (N_6942,N_6651,N_6747);
nor U6943 (N_6943,N_6635,N_6704);
nand U6944 (N_6944,N_6687,N_6615);
nor U6945 (N_6945,N_6646,N_6680);
nand U6946 (N_6946,N_6740,N_6628);
nor U6947 (N_6947,N_6646,N_6762);
or U6948 (N_6948,N_6717,N_6728);
nand U6949 (N_6949,N_6772,N_6631);
nand U6950 (N_6950,N_6714,N_6782);
xor U6951 (N_6951,N_6747,N_6742);
nand U6952 (N_6952,N_6648,N_6667);
nor U6953 (N_6953,N_6624,N_6710);
nor U6954 (N_6954,N_6689,N_6736);
nor U6955 (N_6955,N_6617,N_6736);
xnor U6956 (N_6956,N_6710,N_6789);
or U6957 (N_6957,N_6654,N_6792);
and U6958 (N_6958,N_6734,N_6682);
xor U6959 (N_6959,N_6751,N_6676);
xnor U6960 (N_6960,N_6744,N_6689);
xor U6961 (N_6961,N_6676,N_6607);
and U6962 (N_6962,N_6618,N_6767);
and U6963 (N_6963,N_6723,N_6674);
or U6964 (N_6964,N_6676,N_6620);
nor U6965 (N_6965,N_6623,N_6695);
and U6966 (N_6966,N_6701,N_6625);
nand U6967 (N_6967,N_6778,N_6683);
xnor U6968 (N_6968,N_6740,N_6764);
nand U6969 (N_6969,N_6733,N_6694);
or U6970 (N_6970,N_6700,N_6763);
xnor U6971 (N_6971,N_6626,N_6691);
nor U6972 (N_6972,N_6742,N_6620);
xnor U6973 (N_6973,N_6616,N_6681);
and U6974 (N_6974,N_6621,N_6669);
or U6975 (N_6975,N_6623,N_6639);
nor U6976 (N_6976,N_6677,N_6790);
xor U6977 (N_6977,N_6686,N_6673);
or U6978 (N_6978,N_6682,N_6796);
xnor U6979 (N_6979,N_6722,N_6692);
nor U6980 (N_6980,N_6795,N_6703);
nor U6981 (N_6981,N_6719,N_6683);
nor U6982 (N_6982,N_6797,N_6764);
or U6983 (N_6983,N_6704,N_6642);
xnor U6984 (N_6984,N_6640,N_6738);
nor U6985 (N_6985,N_6680,N_6769);
or U6986 (N_6986,N_6696,N_6631);
and U6987 (N_6987,N_6761,N_6719);
nand U6988 (N_6988,N_6611,N_6678);
nor U6989 (N_6989,N_6726,N_6770);
and U6990 (N_6990,N_6642,N_6744);
nand U6991 (N_6991,N_6640,N_6695);
and U6992 (N_6992,N_6654,N_6649);
and U6993 (N_6993,N_6735,N_6621);
nand U6994 (N_6994,N_6686,N_6791);
or U6995 (N_6995,N_6621,N_6642);
xor U6996 (N_6996,N_6738,N_6726);
or U6997 (N_6997,N_6768,N_6750);
nor U6998 (N_6998,N_6618,N_6620);
and U6999 (N_6999,N_6706,N_6702);
nand U7000 (N_7000,N_6938,N_6926);
xor U7001 (N_7001,N_6937,N_6941);
nand U7002 (N_7002,N_6971,N_6898);
xnor U7003 (N_7003,N_6914,N_6963);
xor U7004 (N_7004,N_6882,N_6862);
nand U7005 (N_7005,N_6990,N_6968);
nor U7006 (N_7006,N_6906,N_6839);
xnor U7007 (N_7007,N_6805,N_6864);
nor U7008 (N_7008,N_6959,N_6944);
nor U7009 (N_7009,N_6913,N_6917);
nor U7010 (N_7010,N_6854,N_6909);
and U7011 (N_7011,N_6949,N_6988);
nor U7012 (N_7012,N_6936,N_6922);
xnor U7013 (N_7013,N_6973,N_6800);
xor U7014 (N_7014,N_6933,N_6902);
xor U7015 (N_7015,N_6974,N_6833);
nor U7016 (N_7016,N_6908,N_6916);
xor U7017 (N_7017,N_6993,N_6896);
xor U7018 (N_7018,N_6829,N_6994);
xor U7019 (N_7019,N_6984,N_6983);
and U7020 (N_7020,N_6856,N_6817);
nand U7021 (N_7021,N_6901,N_6960);
or U7022 (N_7022,N_6934,N_6905);
or U7023 (N_7023,N_6848,N_6821);
xor U7024 (N_7024,N_6883,N_6953);
nor U7025 (N_7025,N_6932,N_6807);
nor U7026 (N_7026,N_6834,N_6801);
or U7027 (N_7027,N_6989,N_6921);
and U7028 (N_7028,N_6952,N_6928);
or U7029 (N_7029,N_6894,N_6970);
nand U7030 (N_7030,N_6955,N_6965);
nor U7031 (N_7031,N_6840,N_6868);
and U7032 (N_7032,N_6930,N_6806);
nand U7033 (N_7033,N_6886,N_6890);
or U7034 (N_7034,N_6962,N_6948);
xor U7035 (N_7035,N_6857,N_6977);
xor U7036 (N_7036,N_6838,N_6925);
nor U7037 (N_7037,N_6855,N_6811);
or U7038 (N_7038,N_6810,N_6849);
nor U7039 (N_7039,N_6809,N_6825);
nand U7040 (N_7040,N_6995,N_6981);
nor U7041 (N_7041,N_6877,N_6845);
or U7042 (N_7042,N_6853,N_6912);
nand U7043 (N_7043,N_6987,N_6876);
nor U7044 (N_7044,N_6957,N_6803);
or U7045 (N_7045,N_6820,N_6920);
xor U7046 (N_7046,N_6844,N_6818);
and U7047 (N_7047,N_6978,N_6832);
nand U7048 (N_7048,N_6982,N_6824);
xnor U7049 (N_7049,N_6954,N_6900);
xor U7050 (N_7050,N_6804,N_6802);
xor U7051 (N_7051,N_6998,N_6992);
and U7052 (N_7052,N_6942,N_6892);
xor U7053 (N_7053,N_6836,N_6851);
xnor U7054 (N_7054,N_6852,N_6870);
xnor U7055 (N_7055,N_6843,N_6879);
nand U7056 (N_7056,N_6958,N_6891);
or U7057 (N_7057,N_6945,N_6915);
xor U7058 (N_7058,N_6888,N_6808);
nand U7059 (N_7059,N_6815,N_6923);
nor U7060 (N_7060,N_6904,N_6979);
nand U7061 (N_7061,N_6865,N_6860);
xnor U7062 (N_7062,N_6911,N_6859);
xor U7063 (N_7063,N_6903,N_6985);
nor U7064 (N_7064,N_6967,N_6918);
and U7065 (N_7065,N_6895,N_6881);
and U7066 (N_7066,N_6826,N_6880);
and U7067 (N_7067,N_6837,N_6822);
nor U7068 (N_7068,N_6927,N_6842);
and U7069 (N_7069,N_6885,N_6867);
nand U7070 (N_7070,N_6871,N_6893);
or U7071 (N_7071,N_6875,N_6878);
xor U7072 (N_7072,N_6969,N_6863);
or U7073 (N_7073,N_6999,N_6889);
or U7074 (N_7074,N_6869,N_6850);
or U7075 (N_7075,N_6835,N_6961);
or U7076 (N_7076,N_6940,N_6910);
nor U7077 (N_7077,N_6873,N_6846);
xnor U7078 (N_7078,N_6874,N_6939);
xnor U7079 (N_7079,N_6966,N_6847);
or U7080 (N_7080,N_6943,N_6964);
or U7081 (N_7081,N_6950,N_6972);
xnor U7082 (N_7082,N_6899,N_6997);
or U7083 (N_7083,N_6897,N_6980);
or U7084 (N_7084,N_6991,N_6887);
xor U7085 (N_7085,N_6812,N_6935);
xor U7086 (N_7086,N_6931,N_6884);
nor U7087 (N_7087,N_6976,N_6924);
nor U7088 (N_7088,N_6946,N_6816);
nand U7089 (N_7089,N_6841,N_6956);
nand U7090 (N_7090,N_6866,N_6919);
xnor U7091 (N_7091,N_6951,N_6947);
nand U7092 (N_7092,N_6872,N_6929);
xor U7093 (N_7093,N_6907,N_6830);
nor U7094 (N_7094,N_6831,N_6986);
xnor U7095 (N_7095,N_6813,N_6823);
or U7096 (N_7096,N_6827,N_6975);
xor U7097 (N_7097,N_6814,N_6828);
and U7098 (N_7098,N_6996,N_6858);
or U7099 (N_7099,N_6819,N_6861);
or U7100 (N_7100,N_6900,N_6816);
or U7101 (N_7101,N_6854,N_6996);
nand U7102 (N_7102,N_6935,N_6972);
nor U7103 (N_7103,N_6903,N_6942);
nor U7104 (N_7104,N_6968,N_6900);
xor U7105 (N_7105,N_6931,N_6912);
nand U7106 (N_7106,N_6848,N_6893);
xnor U7107 (N_7107,N_6972,N_6944);
and U7108 (N_7108,N_6919,N_6907);
nand U7109 (N_7109,N_6903,N_6807);
nand U7110 (N_7110,N_6960,N_6995);
xnor U7111 (N_7111,N_6997,N_6866);
nand U7112 (N_7112,N_6931,N_6824);
or U7113 (N_7113,N_6817,N_6819);
xor U7114 (N_7114,N_6957,N_6833);
and U7115 (N_7115,N_6844,N_6983);
nor U7116 (N_7116,N_6895,N_6835);
xnor U7117 (N_7117,N_6860,N_6884);
xor U7118 (N_7118,N_6931,N_6953);
nor U7119 (N_7119,N_6983,N_6817);
nor U7120 (N_7120,N_6971,N_6991);
nand U7121 (N_7121,N_6919,N_6878);
xor U7122 (N_7122,N_6909,N_6862);
nand U7123 (N_7123,N_6839,N_6805);
nand U7124 (N_7124,N_6933,N_6831);
xnor U7125 (N_7125,N_6869,N_6988);
xnor U7126 (N_7126,N_6930,N_6804);
or U7127 (N_7127,N_6831,N_6999);
nor U7128 (N_7128,N_6813,N_6837);
xor U7129 (N_7129,N_6842,N_6950);
nor U7130 (N_7130,N_6846,N_6951);
xnor U7131 (N_7131,N_6975,N_6986);
xor U7132 (N_7132,N_6852,N_6810);
nand U7133 (N_7133,N_6928,N_6919);
and U7134 (N_7134,N_6861,N_6977);
or U7135 (N_7135,N_6947,N_6965);
xor U7136 (N_7136,N_6864,N_6853);
nor U7137 (N_7137,N_6924,N_6816);
or U7138 (N_7138,N_6873,N_6910);
xnor U7139 (N_7139,N_6962,N_6896);
and U7140 (N_7140,N_6804,N_6928);
nand U7141 (N_7141,N_6951,N_6957);
or U7142 (N_7142,N_6913,N_6957);
nor U7143 (N_7143,N_6897,N_6893);
or U7144 (N_7144,N_6966,N_6824);
nand U7145 (N_7145,N_6853,N_6987);
nor U7146 (N_7146,N_6900,N_6959);
nor U7147 (N_7147,N_6817,N_6827);
xor U7148 (N_7148,N_6968,N_6885);
and U7149 (N_7149,N_6918,N_6990);
nor U7150 (N_7150,N_6904,N_6839);
and U7151 (N_7151,N_6811,N_6850);
or U7152 (N_7152,N_6877,N_6871);
and U7153 (N_7153,N_6847,N_6830);
nor U7154 (N_7154,N_6865,N_6914);
and U7155 (N_7155,N_6872,N_6921);
nor U7156 (N_7156,N_6996,N_6963);
and U7157 (N_7157,N_6870,N_6954);
and U7158 (N_7158,N_6898,N_6800);
xor U7159 (N_7159,N_6814,N_6857);
nand U7160 (N_7160,N_6989,N_6828);
xnor U7161 (N_7161,N_6953,N_6830);
nand U7162 (N_7162,N_6937,N_6853);
or U7163 (N_7163,N_6824,N_6943);
or U7164 (N_7164,N_6854,N_6859);
nand U7165 (N_7165,N_6895,N_6991);
nand U7166 (N_7166,N_6858,N_6874);
and U7167 (N_7167,N_6886,N_6880);
nor U7168 (N_7168,N_6863,N_6880);
nand U7169 (N_7169,N_6977,N_6870);
and U7170 (N_7170,N_6992,N_6906);
nor U7171 (N_7171,N_6878,N_6883);
nor U7172 (N_7172,N_6816,N_6860);
or U7173 (N_7173,N_6980,N_6916);
nand U7174 (N_7174,N_6809,N_6855);
or U7175 (N_7175,N_6972,N_6833);
or U7176 (N_7176,N_6927,N_6917);
nor U7177 (N_7177,N_6996,N_6948);
nand U7178 (N_7178,N_6866,N_6942);
or U7179 (N_7179,N_6838,N_6865);
xor U7180 (N_7180,N_6876,N_6992);
nand U7181 (N_7181,N_6806,N_6859);
or U7182 (N_7182,N_6980,N_6842);
and U7183 (N_7183,N_6841,N_6801);
nor U7184 (N_7184,N_6902,N_6960);
xnor U7185 (N_7185,N_6900,N_6912);
xor U7186 (N_7186,N_6810,N_6953);
nand U7187 (N_7187,N_6809,N_6911);
nand U7188 (N_7188,N_6896,N_6936);
and U7189 (N_7189,N_6947,N_6922);
and U7190 (N_7190,N_6910,N_6892);
nor U7191 (N_7191,N_6872,N_6814);
or U7192 (N_7192,N_6857,N_6926);
nand U7193 (N_7193,N_6905,N_6854);
nor U7194 (N_7194,N_6985,N_6916);
nor U7195 (N_7195,N_6885,N_6805);
nor U7196 (N_7196,N_6973,N_6986);
nor U7197 (N_7197,N_6836,N_6912);
and U7198 (N_7198,N_6849,N_6876);
xnor U7199 (N_7199,N_6825,N_6995);
or U7200 (N_7200,N_7144,N_7159);
nor U7201 (N_7201,N_7105,N_7068);
or U7202 (N_7202,N_7194,N_7002);
nor U7203 (N_7203,N_7182,N_7087);
xnor U7204 (N_7204,N_7037,N_7130);
nand U7205 (N_7205,N_7098,N_7143);
and U7206 (N_7206,N_7027,N_7170);
and U7207 (N_7207,N_7111,N_7031);
nand U7208 (N_7208,N_7119,N_7042);
and U7209 (N_7209,N_7125,N_7133);
nor U7210 (N_7210,N_7184,N_7021);
nand U7211 (N_7211,N_7050,N_7011);
xor U7212 (N_7212,N_7040,N_7036);
or U7213 (N_7213,N_7085,N_7145);
and U7214 (N_7214,N_7053,N_7058);
nand U7215 (N_7215,N_7175,N_7044);
and U7216 (N_7216,N_7008,N_7101);
and U7217 (N_7217,N_7001,N_7134);
and U7218 (N_7218,N_7158,N_7157);
xor U7219 (N_7219,N_7007,N_7173);
or U7220 (N_7220,N_7060,N_7198);
nor U7221 (N_7221,N_7128,N_7110);
xor U7222 (N_7222,N_7057,N_7108);
nor U7223 (N_7223,N_7035,N_7014);
nand U7224 (N_7224,N_7112,N_7181);
and U7225 (N_7225,N_7041,N_7048);
xor U7226 (N_7226,N_7043,N_7077);
xnor U7227 (N_7227,N_7047,N_7154);
xnor U7228 (N_7228,N_7074,N_7121);
or U7229 (N_7229,N_7033,N_7148);
nand U7230 (N_7230,N_7038,N_7034);
or U7231 (N_7231,N_7005,N_7045);
and U7232 (N_7232,N_7080,N_7131);
nor U7233 (N_7233,N_7165,N_7106);
nand U7234 (N_7234,N_7150,N_7089);
nor U7235 (N_7235,N_7117,N_7003);
xnor U7236 (N_7236,N_7188,N_7046);
nor U7237 (N_7237,N_7174,N_7123);
or U7238 (N_7238,N_7083,N_7063);
nor U7239 (N_7239,N_7103,N_7016);
and U7240 (N_7240,N_7006,N_7025);
or U7241 (N_7241,N_7090,N_7061);
or U7242 (N_7242,N_7114,N_7091);
or U7243 (N_7243,N_7024,N_7104);
nand U7244 (N_7244,N_7151,N_7116);
and U7245 (N_7245,N_7136,N_7012);
or U7246 (N_7246,N_7096,N_7192);
or U7247 (N_7247,N_7164,N_7095);
nand U7248 (N_7248,N_7019,N_7013);
or U7249 (N_7249,N_7177,N_7132);
nor U7250 (N_7250,N_7097,N_7029);
nand U7251 (N_7251,N_7113,N_7179);
xnor U7252 (N_7252,N_7139,N_7078);
and U7253 (N_7253,N_7082,N_7169);
and U7254 (N_7254,N_7018,N_7064);
xor U7255 (N_7255,N_7055,N_7065);
and U7256 (N_7256,N_7183,N_7191);
nor U7257 (N_7257,N_7156,N_7100);
nor U7258 (N_7258,N_7004,N_7168);
or U7259 (N_7259,N_7124,N_7028);
xnor U7260 (N_7260,N_7086,N_7023);
and U7261 (N_7261,N_7070,N_7010);
nand U7262 (N_7262,N_7196,N_7084);
nor U7263 (N_7263,N_7071,N_7138);
nor U7264 (N_7264,N_7185,N_7020);
nor U7265 (N_7265,N_7067,N_7122);
or U7266 (N_7266,N_7163,N_7000);
or U7267 (N_7267,N_7017,N_7102);
nand U7268 (N_7268,N_7039,N_7066);
nand U7269 (N_7269,N_7197,N_7146);
nand U7270 (N_7270,N_7187,N_7137);
and U7271 (N_7271,N_7180,N_7126);
xnor U7272 (N_7272,N_7081,N_7030);
nand U7273 (N_7273,N_7099,N_7147);
nor U7274 (N_7274,N_7161,N_7075);
and U7275 (N_7275,N_7141,N_7079);
or U7276 (N_7276,N_7051,N_7142);
and U7277 (N_7277,N_7120,N_7052);
xor U7278 (N_7278,N_7009,N_7199);
xnor U7279 (N_7279,N_7088,N_7073);
xnor U7280 (N_7280,N_7094,N_7186);
and U7281 (N_7281,N_7049,N_7172);
or U7282 (N_7282,N_7195,N_7176);
nor U7283 (N_7283,N_7189,N_7056);
or U7284 (N_7284,N_7171,N_7093);
or U7285 (N_7285,N_7140,N_7072);
and U7286 (N_7286,N_7076,N_7190);
and U7287 (N_7287,N_7022,N_7115);
xor U7288 (N_7288,N_7160,N_7092);
or U7289 (N_7289,N_7135,N_7153);
and U7290 (N_7290,N_7166,N_7107);
nand U7291 (N_7291,N_7109,N_7062);
or U7292 (N_7292,N_7193,N_7178);
xor U7293 (N_7293,N_7155,N_7054);
and U7294 (N_7294,N_7162,N_7152);
or U7295 (N_7295,N_7015,N_7149);
nor U7296 (N_7296,N_7127,N_7167);
nor U7297 (N_7297,N_7129,N_7118);
and U7298 (N_7298,N_7059,N_7026);
nor U7299 (N_7299,N_7069,N_7032);
and U7300 (N_7300,N_7147,N_7113);
nor U7301 (N_7301,N_7155,N_7016);
and U7302 (N_7302,N_7177,N_7157);
nor U7303 (N_7303,N_7044,N_7124);
xor U7304 (N_7304,N_7097,N_7082);
xor U7305 (N_7305,N_7148,N_7061);
nand U7306 (N_7306,N_7152,N_7168);
or U7307 (N_7307,N_7146,N_7040);
or U7308 (N_7308,N_7142,N_7138);
and U7309 (N_7309,N_7112,N_7160);
nor U7310 (N_7310,N_7155,N_7024);
nor U7311 (N_7311,N_7046,N_7170);
nand U7312 (N_7312,N_7174,N_7109);
nand U7313 (N_7313,N_7087,N_7017);
or U7314 (N_7314,N_7149,N_7007);
or U7315 (N_7315,N_7189,N_7116);
nor U7316 (N_7316,N_7054,N_7070);
xor U7317 (N_7317,N_7078,N_7140);
xnor U7318 (N_7318,N_7181,N_7070);
nand U7319 (N_7319,N_7113,N_7114);
nor U7320 (N_7320,N_7091,N_7093);
and U7321 (N_7321,N_7028,N_7062);
nand U7322 (N_7322,N_7119,N_7110);
nor U7323 (N_7323,N_7021,N_7196);
or U7324 (N_7324,N_7094,N_7072);
nand U7325 (N_7325,N_7156,N_7098);
nor U7326 (N_7326,N_7034,N_7195);
nor U7327 (N_7327,N_7031,N_7129);
and U7328 (N_7328,N_7043,N_7131);
xor U7329 (N_7329,N_7018,N_7129);
and U7330 (N_7330,N_7098,N_7199);
xnor U7331 (N_7331,N_7030,N_7071);
nor U7332 (N_7332,N_7131,N_7056);
or U7333 (N_7333,N_7182,N_7177);
nor U7334 (N_7334,N_7101,N_7139);
nor U7335 (N_7335,N_7150,N_7010);
nor U7336 (N_7336,N_7095,N_7022);
or U7337 (N_7337,N_7134,N_7193);
xor U7338 (N_7338,N_7198,N_7030);
nand U7339 (N_7339,N_7162,N_7128);
nor U7340 (N_7340,N_7173,N_7145);
and U7341 (N_7341,N_7002,N_7100);
nand U7342 (N_7342,N_7131,N_7053);
nand U7343 (N_7343,N_7142,N_7180);
or U7344 (N_7344,N_7155,N_7012);
nand U7345 (N_7345,N_7079,N_7097);
or U7346 (N_7346,N_7072,N_7118);
or U7347 (N_7347,N_7085,N_7173);
nand U7348 (N_7348,N_7182,N_7076);
and U7349 (N_7349,N_7003,N_7010);
xor U7350 (N_7350,N_7112,N_7043);
or U7351 (N_7351,N_7093,N_7042);
nor U7352 (N_7352,N_7122,N_7039);
or U7353 (N_7353,N_7179,N_7166);
and U7354 (N_7354,N_7181,N_7131);
or U7355 (N_7355,N_7095,N_7053);
or U7356 (N_7356,N_7178,N_7084);
nand U7357 (N_7357,N_7040,N_7126);
or U7358 (N_7358,N_7089,N_7154);
nor U7359 (N_7359,N_7143,N_7136);
xnor U7360 (N_7360,N_7045,N_7026);
xnor U7361 (N_7361,N_7154,N_7157);
nor U7362 (N_7362,N_7060,N_7004);
xor U7363 (N_7363,N_7150,N_7196);
nand U7364 (N_7364,N_7111,N_7159);
xnor U7365 (N_7365,N_7041,N_7051);
and U7366 (N_7366,N_7057,N_7153);
nor U7367 (N_7367,N_7121,N_7017);
or U7368 (N_7368,N_7168,N_7199);
and U7369 (N_7369,N_7100,N_7133);
and U7370 (N_7370,N_7141,N_7174);
or U7371 (N_7371,N_7162,N_7070);
or U7372 (N_7372,N_7110,N_7066);
xor U7373 (N_7373,N_7098,N_7018);
xnor U7374 (N_7374,N_7196,N_7168);
xor U7375 (N_7375,N_7149,N_7193);
or U7376 (N_7376,N_7028,N_7088);
nor U7377 (N_7377,N_7157,N_7190);
nor U7378 (N_7378,N_7008,N_7135);
xnor U7379 (N_7379,N_7032,N_7050);
xnor U7380 (N_7380,N_7136,N_7002);
nor U7381 (N_7381,N_7110,N_7135);
nor U7382 (N_7382,N_7019,N_7002);
nor U7383 (N_7383,N_7003,N_7131);
nor U7384 (N_7384,N_7007,N_7056);
nor U7385 (N_7385,N_7047,N_7095);
nor U7386 (N_7386,N_7192,N_7082);
xnor U7387 (N_7387,N_7165,N_7085);
nand U7388 (N_7388,N_7127,N_7002);
and U7389 (N_7389,N_7068,N_7174);
xor U7390 (N_7390,N_7053,N_7182);
nor U7391 (N_7391,N_7130,N_7099);
or U7392 (N_7392,N_7180,N_7149);
xor U7393 (N_7393,N_7124,N_7122);
or U7394 (N_7394,N_7151,N_7067);
nor U7395 (N_7395,N_7035,N_7012);
nand U7396 (N_7396,N_7135,N_7168);
nor U7397 (N_7397,N_7063,N_7111);
and U7398 (N_7398,N_7157,N_7025);
nand U7399 (N_7399,N_7162,N_7167);
xnor U7400 (N_7400,N_7227,N_7332);
nand U7401 (N_7401,N_7201,N_7316);
xnor U7402 (N_7402,N_7210,N_7240);
xnor U7403 (N_7403,N_7248,N_7285);
xnor U7404 (N_7404,N_7250,N_7360);
or U7405 (N_7405,N_7321,N_7219);
xnor U7406 (N_7406,N_7306,N_7302);
xnor U7407 (N_7407,N_7315,N_7322);
xor U7408 (N_7408,N_7331,N_7323);
or U7409 (N_7409,N_7356,N_7258);
and U7410 (N_7410,N_7252,N_7267);
nor U7411 (N_7411,N_7355,N_7231);
and U7412 (N_7412,N_7290,N_7212);
xor U7413 (N_7413,N_7353,N_7372);
nand U7414 (N_7414,N_7394,N_7270);
nor U7415 (N_7415,N_7349,N_7271);
and U7416 (N_7416,N_7329,N_7273);
nand U7417 (N_7417,N_7225,N_7217);
and U7418 (N_7418,N_7251,N_7284);
xor U7419 (N_7419,N_7341,N_7357);
or U7420 (N_7420,N_7289,N_7202);
xor U7421 (N_7421,N_7208,N_7260);
and U7422 (N_7422,N_7390,N_7314);
or U7423 (N_7423,N_7264,N_7375);
nor U7424 (N_7424,N_7268,N_7253);
xnor U7425 (N_7425,N_7343,N_7377);
and U7426 (N_7426,N_7230,N_7373);
nand U7427 (N_7427,N_7358,N_7241);
nor U7428 (N_7428,N_7278,N_7311);
nand U7429 (N_7429,N_7348,N_7393);
nor U7430 (N_7430,N_7342,N_7336);
nand U7431 (N_7431,N_7370,N_7203);
nand U7432 (N_7432,N_7381,N_7216);
or U7433 (N_7433,N_7274,N_7294);
and U7434 (N_7434,N_7256,N_7337);
or U7435 (N_7435,N_7281,N_7269);
or U7436 (N_7436,N_7395,N_7277);
and U7437 (N_7437,N_7378,N_7214);
nor U7438 (N_7438,N_7213,N_7310);
nor U7439 (N_7439,N_7220,N_7215);
and U7440 (N_7440,N_7364,N_7325);
or U7441 (N_7441,N_7317,N_7304);
xnor U7442 (N_7442,N_7369,N_7338);
and U7443 (N_7443,N_7303,N_7229);
nand U7444 (N_7444,N_7300,N_7243);
xor U7445 (N_7445,N_7218,N_7297);
or U7446 (N_7446,N_7295,N_7235);
nor U7447 (N_7447,N_7396,N_7261);
or U7448 (N_7448,N_7205,N_7388);
nor U7449 (N_7449,N_7262,N_7339);
or U7450 (N_7450,N_7263,N_7293);
xnor U7451 (N_7451,N_7224,N_7391);
or U7452 (N_7452,N_7376,N_7366);
nand U7453 (N_7453,N_7379,N_7207);
nor U7454 (N_7454,N_7362,N_7318);
and U7455 (N_7455,N_7398,N_7313);
nor U7456 (N_7456,N_7382,N_7222);
nand U7457 (N_7457,N_7280,N_7299);
nand U7458 (N_7458,N_7334,N_7383);
nor U7459 (N_7459,N_7239,N_7272);
and U7460 (N_7460,N_7328,N_7347);
nand U7461 (N_7461,N_7234,N_7352);
and U7462 (N_7462,N_7363,N_7221);
xnor U7463 (N_7463,N_7320,N_7324);
and U7464 (N_7464,N_7249,N_7232);
nand U7465 (N_7465,N_7333,N_7309);
nand U7466 (N_7466,N_7345,N_7308);
or U7467 (N_7467,N_7340,N_7226);
and U7468 (N_7468,N_7327,N_7228);
nand U7469 (N_7469,N_7296,N_7330);
and U7470 (N_7470,N_7371,N_7266);
nand U7471 (N_7471,N_7384,N_7206);
nor U7472 (N_7472,N_7292,N_7319);
and U7473 (N_7473,N_7211,N_7283);
nand U7474 (N_7474,N_7335,N_7244);
nor U7475 (N_7475,N_7259,N_7385);
and U7476 (N_7476,N_7374,N_7276);
nor U7477 (N_7477,N_7380,N_7397);
nor U7478 (N_7478,N_7344,N_7350);
and U7479 (N_7479,N_7399,N_7298);
nand U7480 (N_7480,N_7351,N_7254);
nor U7481 (N_7481,N_7291,N_7286);
nand U7482 (N_7482,N_7392,N_7368);
xnor U7483 (N_7483,N_7386,N_7238);
xor U7484 (N_7484,N_7301,N_7237);
and U7485 (N_7485,N_7242,N_7257);
nor U7486 (N_7486,N_7204,N_7305);
nor U7487 (N_7487,N_7275,N_7255);
xnor U7488 (N_7488,N_7223,N_7245);
nand U7489 (N_7489,N_7247,N_7282);
xor U7490 (N_7490,N_7279,N_7365);
nand U7491 (N_7491,N_7307,N_7389);
xnor U7492 (N_7492,N_7287,N_7359);
and U7493 (N_7493,N_7200,N_7209);
nor U7494 (N_7494,N_7387,N_7312);
xnor U7495 (N_7495,N_7367,N_7354);
nand U7496 (N_7496,N_7233,N_7236);
xnor U7497 (N_7497,N_7326,N_7288);
nand U7498 (N_7498,N_7361,N_7246);
nand U7499 (N_7499,N_7346,N_7265);
or U7500 (N_7500,N_7314,N_7232);
nand U7501 (N_7501,N_7275,N_7371);
or U7502 (N_7502,N_7277,N_7380);
nor U7503 (N_7503,N_7385,N_7348);
or U7504 (N_7504,N_7296,N_7338);
xnor U7505 (N_7505,N_7212,N_7224);
or U7506 (N_7506,N_7298,N_7355);
and U7507 (N_7507,N_7346,N_7219);
and U7508 (N_7508,N_7396,N_7224);
xnor U7509 (N_7509,N_7332,N_7308);
nand U7510 (N_7510,N_7369,N_7249);
nand U7511 (N_7511,N_7202,N_7270);
and U7512 (N_7512,N_7335,N_7365);
nand U7513 (N_7513,N_7326,N_7295);
xnor U7514 (N_7514,N_7366,N_7266);
xnor U7515 (N_7515,N_7253,N_7352);
and U7516 (N_7516,N_7274,N_7397);
nor U7517 (N_7517,N_7395,N_7339);
nor U7518 (N_7518,N_7241,N_7311);
nor U7519 (N_7519,N_7305,N_7369);
and U7520 (N_7520,N_7205,N_7294);
nor U7521 (N_7521,N_7304,N_7288);
or U7522 (N_7522,N_7353,N_7317);
and U7523 (N_7523,N_7319,N_7360);
nand U7524 (N_7524,N_7293,N_7239);
nor U7525 (N_7525,N_7209,N_7232);
xnor U7526 (N_7526,N_7382,N_7214);
xor U7527 (N_7527,N_7331,N_7317);
and U7528 (N_7528,N_7237,N_7328);
nor U7529 (N_7529,N_7382,N_7373);
or U7530 (N_7530,N_7213,N_7380);
or U7531 (N_7531,N_7272,N_7234);
nor U7532 (N_7532,N_7252,N_7341);
nand U7533 (N_7533,N_7239,N_7228);
and U7534 (N_7534,N_7369,N_7200);
or U7535 (N_7535,N_7251,N_7304);
nor U7536 (N_7536,N_7259,N_7372);
nor U7537 (N_7537,N_7397,N_7375);
xnor U7538 (N_7538,N_7260,N_7341);
xnor U7539 (N_7539,N_7243,N_7270);
xor U7540 (N_7540,N_7282,N_7366);
nand U7541 (N_7541,N_7229,N_7256);
and U7542 (N_7542,N_7398,N_7324);
and U7543 (N_7543,N_7209,N_7247);
or U7544 (N_7544,N_7341,N_7304);
nor U7545 (N_7545,N_7393,N_7337);
nand U7546 (N_7546,N_7283,N_7338);
or U7547 (N_7547,N_7227,N_7223);
or U7548 (N_7548,N_7229,N_7375);
xor U7549 (N_7549,N_7214,N_7305);
nor U7550 (N_7550,N_7330,N_7323);
nand U7551 (N_7551,N_7315,N_7222);
and U7552 (N_7552,N_7399,N_7356);
xnor U7553 (N_7553,N_7274,N_7379);
and U7554 (N_7554,N_7303,N_7318);
and U7555 (N_7555,N_7295,N_7234);
nor U7556 (N_7556,N_7235,N_7259);
or U7557 (N_7557,N_7343,N_7245);
and U7558 (N_7558,N_7344,N_7288);
nor U7559 (N_7559,N_7364,N_7340);
nor U7560 (N_7560,N_7310,N_7335);
and U7561 (N_7561,N_7205,N_7281);
xnor U7562 (N_7562,N_7223,N_7363);
xor U7563 (N_7563,N_7211,N_7320);
nand U7564 (N_7564,N_7324,N_7272);
and U7565 (N_7565,N_7385,N_7349);
and U7566 (N_7566,N_7299,N_7216);
xnor U7567 (N_7567,N_7261,N_7332);
or U7568 (N_7568,N_7328,N_7350);
nor U7569 (N_7569,N_7369,N_7283);
nor U7570 (N_7570,N_7340,N_7363);
nor U7571 (N_7571,N_7363,N_7359);
nor U7572 (N_7572,N_7242,N_7336);
xor U7573 (N_7573,N_7365,N_7205);
nand U7574 (N_7574,N_7217,N_7310);
or U7575 (N_7575,N_7358,N_7239);
nand U7576 (N_7576,N_7232,N_7238);
nand U7577 (N_7577,N_7233,N_7384);
nand U7578 (N_7578,N_7233,N_7377);
or U7579 (N_7579,N_7259,N_7251);
nor U7580 (N_7580,N_7370,N_7226);
and U7581 (N_7581,N_7322,N_7314);
or U7582 (N_7582,N_7382,N_7350);
xnor U7583 (N_7583,N_7220,N_7348);
nand U7584 (N_7584,N_7337,N_7249);
nor U7585 (N_7585,N_7244,N_7270);
and U7586 (N_7586,N_7216,N_7298);
xnor U7587 (N_7587,N_7341,N_7335);
or U7588 (N_7588,N_7276,N_7293);
nor U7589 (N_7589,N_7279,N_7341);
and U7590 (N_7590,N_7310,N_7248);
and U7591 (N_7591,N_7321,N_7290);
xnor U7592 (N_7592,N_7206,N_7382);
xnor U7593 (N_7593,N_7391,N_7240);
xnor U7594 (N_7594,N_7263,N_7388);
nand U7595 (N_7595,N_7336,N_7299);
or U7596 (N_7596,N_7353,N_7233);
and U7597 (N_7597,N_7216,N_7245);
nor U7598 (N_7598,N_7373,N_7258);
xor U7599 (N_7599,N_7219,N_7240);
or U7600 (N_7600,N_7408,N_7501);
or U7601 (N_7601,N_7490,N_7578);
nand U7602 (N_7602,N_7448,N_7436);
xor U7603 (N_7603,N_7491,N_7405);
or U7604 (N_7604,N_7461,N_7510);
and U7605 (N_7605,N_7532,N_7512);
or U7606 (N_7606,N_7494,N_7585);
and U7607 (N_7607,N_7425,N_7438);
and U7608 (N_7608,N_7479,N_7483);
xor U7609 (N_7609,N_7450,N_7435);
and U7610 (N_7610,N_7567,N_7487);
xor U7611 (N_7611,N_7553,N_7582);
nand U7612 (N_7612,N_7498,N_7440);
or U7613 (N_7613,N_7492,N_7449);
and U7614 (N_7614,N_7441,N_7592);
nand U7615 (N_7615,N_7576,N_7533);
nand U7616 (N_7616,N_7515,N_7456);
nand U7617 (N_7617,N_7555,N_7443);
xor U7618 (N_7618,N_7542,N_7548);
nand U7619 (N_7619,N_7423,N_7442);
or U7620 (N_7620,N_7412,N_7526);
xnor U7621 (N_7621,N_7588,N_7473);
xnor U7622 (N_7622,N_7429,N_7531);
nand U7623 (N_7623,N_7453,N_7572);
xnor U7624 (N_7624,N_7559,N_7458);
or U7625 (N_7625,N_7554,N_7562);
xor U7626 (N_7626,N_7566,N_7444);
nand U7627 (N_7627,N_7577,N_7482);
nand U7628 (N_7628,N_7421,N_7537);
nor U7629 (N_7629,N_7424,N_7426);
xor U7630 (N_7630,N_7541,N_7475);
or U7631 (N_7631,N_7573,N_7500);
and U7632 (N_7632,N_7481,N_7570);
xnor U7633 (N_7633,N_7459,N_7469);
and U7634 (N_7634,N_7506,N_7489);
xnor U7635 (N_7635,N_7595,N_7536);
nor U7636 (N_7636,N_7556,N_7579);
nor U7637 (N_7637,N_7552,N_7594);
xnor U7638 (N_7638,N_7513,N_7511);
or U7639 (N_7639,N_7466,N_7560);
nor U7640 (N_7640,N_7587,N_7563);
xnor U7641 (N_7641,N_7472,N_7464);
nand U7642 (N_7642,N_7583,N_7514);
nor U7643 (N_7643,N_7462,N_7455);
xor U7644 (N_7644,N_7452,N_7460);
xnor U7645 (N_7645,N_7519,N_7516);
and U7646 (N_7646,N_7427,N_7530);
and U7647 (N_7647,N_7546,N_7529);
nor U7648 (N_7648,N_7584,N_7463);
and U7649 (N_7649,N_7589,N_7538);
xnor U7650 (N_7650,N_7540,N_7418);
nand U7651 (N_7651,N_7598,N_7571);
xor U7652 (N_7652,N_7565,N_7525);
and U7653 (N_7653,N_7596,N_7557);
nor U7654 (N_7654,N_7432,N_7439);
nor U7655 (N_7655,N_7454,N_7451);
and U7656 (N_7656,N_7591,N_7569);
or U7657 (N_7657,N_7597,N_7545);
nor U7658 (N_7658,N_7496,N_7476);
and U7659 (N_7659,N_7404,N_7465);
nor U7660 (N_7660,N_7504,N_7543);
and U7661 (N_7661,N_7457,N_7401);
xor U7662 (N_7662,N_7586,N_7550);
xnor U7663 (N_7663,N_7508,N_7470);
nand U7664 (N_7664,N_7402,N_7580);
or U7665 (N_7665,N_7437,N_7518);
nand U7666 (N_7666,N_7517,N_7485);
nand U7667 (N_7667,N_7406,N_7446);
and U7668 (N_7668,N_7522,N_7484);
and U7669 (N_7669,N_7551,N_7599);
xor U7670 (N_7670,N_7564,N_7549);
nor U7671 (N_7671,N_7474,N_7471);
and U7672 (N_7672,N_7509,N_7581);
nand U7673 (N_7673,N_7575,N_7413);
and U7674 (N_7674,N_7414,N_7422);
and U7675 (N_7675,N_7416,N_7574);
and U7676 (N_7676,N_7410,N_7568);
and U7677 (N_7677,N_7497,N_7527);
or U7678 (N_7678,N_7415,N_7411);
nand U7679 (N_7679,N_7558,N_7520);
xor U7680 (N_7680,N_7499,N_7488);
xor U7681 (N_7681,N_7502,N_7445);
nand U7682 (N_7682,N_7428,N_7503);
nor U7683 (N_7683,N_7486,N_7478);
xor U7684 (N_7684,N_7521,N_7407);
and U7685 (N_7685,N_7409,N_7480);
and U7686 (N_7686,N_7420,N_7468);
or U7687 (N_7687,N_7539,N_7534);
and U7688 (N_7688,N_7434,N_7535);
nor U7689 (N_7689,N_7544,N_7547);
xor U7690 (N_7690,N_7528,N_7523);
and U7691 (N_7691,N_7495,N_7431);
nor U7692 (N_7692,N_7505,N_7467);
and U7693 (N_7693,N_7593,N_7477);
nand U7694 (N_7694,N_7493,N_7433);
nor U7695 (N_7695,N_7403,N_7417);
xnor U7696 (N_7696,N_7507,N_7524);
or U7697 (N_7697,N_7561,N_7430);
or U7698 (N_7698,N_7590,N_7400);
xor U7699 (N_7699,N_7419,N_7447);
xnor U7700 (N_7700,N_7425,N_7593);
nor U7701 (N_7701,N_7572,N_7461);
xnor U7702 (N_7702,N_7590,N_7527);
and U7703 (N_7703,N_7506,N_7528);
xor U7704 (N_7704,N_7423,N_7469);
nand U7705 (N_7705,N_7493,N_7418);
and U7706 (N_7706,N_7566,N_7501);
nand U7707 (N_7707,N_7489,N_7522);
and U7708 (N_7708,N_7494,N_7477);
xnor U7709 (N_7709,N_7469,N_7453);
nor U7710 (N_7710,N_7559,N_7422);
xnor U7711 (N_7711,N_7424,N_7418);
and U7712 (N_7712,N_7578,N_7513);
or U7713 (N_7713,N_7521,N_7420);
nor U7714 (N_7714,N_7483,N_7505);
and U7715 (N_7715,N_7504,N_7551);
or U7716 (N_7716,N_7424,N_7577);
or U7717 (N_7717,N_7494,N_7496);
xnor U7718 (N_7718,N_7466,N_7501);
nor U7719 (N_7719,N_7506,N_7484);
xnor U7720 (N_7720,N_7472,N_7582);
and U7721 (N_7721,N_7409,N_7483);
xnor U7722 (N_7722,N_7534,N_7537);
xnor U7723 (N_7723,N_7586,N_7543);
nor U7724 (N_7724,N_7410,N_7457);
nand U7725 (N_7725,N_7455,N_7582);
xor U7726 (N_7726,N_7557,N_7511);
xnor U7727 (N_7727,N_7553,N_7475);
nor U7728 (N_7728,N_7513,N_7478);
xor U7729 (N_7729,N_7417,N_7495);
and U7730 (N_7730,N_7442,N_7580);
and U7731 (N_7731,N_7580,N_7587);
or U7732 (N_7732,N_7408,N_7530);
xnor U7733 (N_7733,N_7497,N_7541);
nor U7734 (N_7734,N_7406,N_7589);
and U7735 (N_7735,N_7473,N_7587);
and U7736 (N_7736,N_7513,N_7518);
or U7737 (N_7737,N_7425,N_7495);
xor U7738 (N_7738,N_7470,N_7466);
xnor U7739 (N_7739,N_7579,N_7408);
nand U7740 (N_7740,N_7413,N_7492);
nor U7741 (N_7741,N_7533,N_7553);
or U7742 (N_7742,N_7457,N_7585);
or U7743 (N_7743,N_7549,N_7504);
nor U7744 (N_7744,N_7474,N_7590);
nor U7745 (N_7745,N_7569,N_7447);
nor U7746 (N_7746,N_7539,N_7491);
or U7747 (N_7747,N_7549,N_7456);
and U7748 (N_7748,N_7495,N_7460);
and U7749 (N_7749,N_7591,N_7451);
or U7750 (N_7750,N_7482,N_7420);
nand U7751 (N_7751,N_7497,N_7414);
or U7752 (N_7752,N_7512,N_7506);
or U7753 (N_7753,N_7410,N_7474);
or U7754 (N_7754,N_7564,N_7456);
xor U7755 (N_7755,N_7411,N_7447);
xnor U7756 (N_7756,N_7527,N_7563);
nor U7757 (N_7757,N_7540,N_7588);
nor U7758 (N_7758,N_7478,N_7533);
xor U7759 (N_7759,N_7492,N_7419);
and U7760 (N_7760,N_7425,N_7446);
nand U7761 (N_7761,N_7452,N_7408);
and U7762 (N_7762,N_7484,N_7558);
xnor U7763 (N_7763,N_7574,N_7560);
xor U7764 (N_7764,N_7565,N_7527);
nand U7765 (N_7765,N_7470,N_7431);
nand U7766 (N_7766,N_7474,N_7426);
nand U7767 (N_7767,N_7466,N_7554);
nand U7768 (N_7768,N_7585,N_7507);
nand U7769 (N_7769,N_7583,N_7554);
nor U7770 (N_7770,N_7404,N_7493);
nor U7771 (N_7771,N_7599,N_7500);
xor U7772 (N_7772,N_7433,N_7555);
nand U7773 (N_7773,N_7580,N_7447);
or U7774 (N_7774,N_7433,N_7488);
xor U7775 (N_7775,N_7469,N_7506);
nand U7776 (N_7776,N_7529,N_7465);
nor U7777 (N_7777,N_7440,N_7447);
or U7778 (N_7778,N_7577,N_7495);
nand U7779 (N_7779,N_7551,N_7420);
nor U7780 (N_7780,N_7556,N_7401);
and U7781 (N_7781,N_7517,N_7542);
nor U7782 (N_7782,N_7408,N_7455);
or U7783 (N_7783,N_7459,N_7541);
xnor U7784 (N_7784,N_7465,N_7478);
or U7785 (N_7785,N_7506,N_7476);
and U7786 (N_7786,N_7473,N_7517);
nand U7787 (N_7787,N_7408,N_7598);
and U7788 (N_7788,N_7433,N_7566);
or U7789 (N_7789,N_7450,N_7469);
nor U7790 (N_7790,N_7488,N_7468);
or U7791 (N_7791,N_7549,N_7423);
nand U7792 (N_7792,N_7406,N_7485);
nand U7793 (N_7793,N_7564,N_7508);
nor U7794 (N_7794,N_7445,N_7562);
or U7795 (N_7795,N_7512,N_7535);
xnor U7796 (N_7796,N_7530,N_7486);
or U7797 (N_7797,N_7580,N_7401);
and U7798 (N_7798,N_7447,N_7409);
xnor U7799 (N_7799,N_7457,N_7535);
or U7800 (N_7800,N_7760,N_7629);
nand U7801 (N_7801,N_7638,N_7612);
and U7802 (N_7802,N_7646,N_7793);
nor U7803 (N_7803,N_7672,N_7726);
xnor U7804 (N_7804,N_7603,N_7781);
nor U7805 (N_7805,N_7727,N_7758);
and U7806 (N_7806,N_7604,N_7644);
nand U7807 (N_7807,N_7670,N_7645);
xor U7808 (N_7808,N_7729,N_7624);
or U7809 (N_7809,N_7634,N_7734);
nand U7810 (N_7810,N_7723,N_7632);
nor U7811 (N_7811,N_7621,N_7707);
or U7812 (N_7812,N_7657,N_7768);
and U7813 (N_7813,N_7666,N_7724);
or U7814 (N_7814,N_7628,N_7671);
xnor U7815 (N_7815,N_7709,N_7610);
nand U7816 (N_7816,N_7688,N_7679);
xnor U7817 (N_7817,N_7792,N_7627);
nand U7818 (N_7818,N_7761,N_7746);
or U7819 (N_7819,N_7751,N_7696);
xor U7820 (N_7820,N_7722,N_7630);
nand U7821 (N_7821,N_7772,N_7795);
xnor U7822 (N_7822,N_7663,N_7625);
nand U7823 (N_7823,N_7736,N_7704);
nand U7824 (N_7824,N_7797,N_7782);
and U7825 (N_7825,N_7665,N_7698);
nand U7826 (N_7826,N_7659,N_7749);
xnor U7827 (N_7827,N_7778,N_7770);
nor U7828 (N_7828,N_7676,N_7668);
and U7829 (N_7829,N_7690,N_7733);
and U7830 (N_7830,N_7790,N_7623);
or U7831 (N_7831,N_7613,N_7667);
or U7832 (N_7832,N_7701,N_7615);
and U7833 (N_7833,N_7673,N_7675);
nand U7834 (N_7834,N_7677,N_7681);
nor U7835 (N_7835,N_7753,N_7757);
nor U7836 (N_7836,N_7641,N_7687);
and U7837 (N_7837,N_7614,N_7682);
or U7838 (N_7838,N_7739,N_7703);
xnor U7839 (N_7839,N_7654,N_7784);
nand U7840 (N_7840,N_7622,N_7741);
or U7841 (N_7841,N_7611,N_7650);
nor U7842 (N_7842,N_7637,N_7743);
nor U7843 (N_7843,N_7785,N_7652);
and U7844 (N_7844,N_7780,N_7602);
nor U7845 (N_7845,N_7725,N_7694);
xnor U7846 (N_7846,N_7789,N_7752);
nor U7847 (N_7847,N_7636,N_7740);
nand U7848 (N_7848,N_7619,N_7783);
nand U7849 (N_7849,N_7647,N_7773);
and U7850 (N_7850,N_7718,N_7769);
xor U7851 (N_7851,N_7745,N_7748);
nor U7852 (N_7852,N_7779,N_7765);
and U7853 (N_7853,N_7787,N_7691);
and U7854 (N_7854,N_7786,N_7617);
nor U7855 (N_7855,N_7762,N_7633);
or U7856 (N_7856,N_7699,N_7750);
or U7857 (N_7857,N_7656,N_7719);
or U7858 (N_7858,N_7683,N_7730);
nor U7859 (N_7859,N_7735,N_7643);
and U7860 (N_7860,N_7642,N_7754);
and U7861 (N_7861,N_7664,N_7744);
xnor U7862 (N_7862,N_7732,N_7686);
or U7863 (N_7863,N_7708,N_7639);
nand U7864 (N_7864,N_7640,N_7731);
or U7865 (N_7865,N_7607,N_7618);
or U7866 (N_7866,N_7712,N_7794);
nand U7867 (N_7867,N_7692,N_7777);
or U7868 (N_7868,N_7674,N_7775);
nand U7869 (N_7869,N_7774,N_7626);
nor U7870 (N_7870,N_7742,N_7756);
nor U7871 (N_7871,N_7705,N_7685);
xnor U7872 (N_7872,N_7713,N_7721);
or U7873 (N_7873,N_7678,N_7714);
nor U7874 (N_7874,N_7648,N_7716);
xor U7875 (N_7875,N_7695,N_7717);
or U7876 (N_7876,N_7655,N_7711);
nand U7877 (N_7877,N_7609,N_7771);
xnor U7878 (N_7878,N_7684,N_7669);
nor U7879 (N_7879,N_7737,N_7680);
nand U7880 (N_7880,N_7689,N_7616);
or U7881 (N_7881,N_7766,N_7631);
or U7882 (N_7882,N_7661,N_7658);
nand U7883 (N_7883,N_7798,N_7660);
nand U7884 (N_7884,N_7693,N_7653);
nor U7885 (N_7885,N_7662,N_7764);
xnor U7886 (N_7886,N_7796,N_7715);
xnor U7887 (N_7887,N_7767,N_7606);
nand U7888 (N_7888,N_7700,N_7697);
nand U7889 (N_7889,N_7738,N_7710);
nor U7890 (N_7890,N_7620,N_7601);
nand U7891 (N_7891,N_7799,N_7728);
xor U7892 (N_7892,N_7791,N_7605);
nor U7893 (N_7893,N_7759,N_7747);
xnor U7894 (N_7894,N_7788,N_7600);
xor U7895 (N_7895,N_7649,N_7702);
xnor U7896 (N_7896,N_7651,N_7763);
and U7897 (N_7897,N_7720,N_7755);
nand U7898 (N_7898,N_7608,N_7776);
nand U7899 (N_7899,N_7635,N_7706);
nor U7900 (N_7900,N_7633,N_7790);
and U7901 (N_7901,N_7795,N_7603);
and U7902 (N_7902,N_7733,N_7762);
nor U7903 (N_7903,N_7643,N_7743);
nand U7904 (N_7904,N_7663,N_7737);
nand U7905 (N_7905,N_7733,N_7667);
nand U7906 (N_7906,N_7759,N_7709);
xor U7907 (N_7907,N_7760,N_7706);
nor U7908 (N_7908,N_7623,N_7693);
xnor U7909 (N_7909,N_7639,N_7750);
xor U7910 (N_7910,N_7760,N_7654);
and U7911 (N_7911,N_7642,N_7778);
nand U7912 (N_7912,N_7759,N_7666);
xnor U7913 (N_7913,N_7758,N_7639);
nor U7914 (N_7914,N_7726,N_7627);
and U7915 (N_7915,N_7734,N_7667);
xnor U7916 (N_7916,N_7699,N_7714);
nor U7917 (N_7917,N_7735,N_7604);
nor U7918 (N_7918,N_7711,N_7682);
or U7919 (N_7919,N_7763,N_7712);
xor U7920 (N_7920,N_7768,N_7789);
xnor U7921 (N_7921,N_7622,N_7725);
xor U7922 (N_7922,N_7605,N_7668);
nand U7923 (N_7923,N_7768,N_7680);
nor U7924 (N_7924,N_7607,N_7790);
and U7925 (N_7925,N_7768,N_7622);
nand U7926 (N_7926,N_7656,N_7770);
and U7927 (N_7927,N_7667,N_7721);
and U7928 (N_7928,N_7682,N_7683);
nand U7929 (N_7929,N_7799,N_7775);
and U7930 (N_7930,N_7775,N_7761);
and U7931 (N_7931,N_7768,N_7733);
nand U7932 (N_7932,N_7763,N_7724);
nor U7933 (N_7933,N_7678,N_7783);
or U7934 (N_7934,N_7697,N_7600);
nor U7935 (N_7935,N_7715,N_7792);
nand U7936 (N_7936,N_7688,N_7700);
nor U7937 (N_7937,N_7692,N_7784);
or U7938 (N_7938,N_7794,N_7719);
xnor U7939 (N_7939,N_7679,N_7658);
and U7940 (N_7940,N_7751,N_7722);
and U7941 (N_7941,N_7727,N_7628);
xor U7942 (N_7942,N_7784,N_7691);
nand U7943 (N_7943,N_7727,N_7621);
nand U7944 (N_7944,N_7636,N_7668);
and U7945 (N_7945,N_7625,N_7601);
xor U7946 (N_7946,N_7715,N_7770);
xor U7947 (N_7947,N_7721,N_7626);
nand U7948 (N_7948,N_7686,N_7634);
or U7949 (N_7949,N_7607,N_7793);
and U7950 (N_7950,N_7772,N_7720);
or U7951 (N_7951,N_7652,N_7665);
xnor U7952 (N_7952,N_7774,N_7797);
or U7953 (N_7953,N_7728,N_7619);
and U7954 (N_7954,N_7667,N_7778);
or U7955 (N_7955,N_7649,N_7739);
xnor U7956 (N_7956,N_7670,N_7678);
or U7957 (N_7957,N_7618,N_7726);
and U7958 (N_7958,N_7608,N_7791);
and U7959 (N_7959,N_7717,N_7679);
nor U7960 (N_7960,N_7783,N_7750);
nand U7961 (N_7961,N_7617,N_7650);
nor U7962 (N_7962,N_7794,N_7758);
xnor U7963 (N_7963,N_7674,N_7692);
nor U7964 (N_7964,N_7731,N_7617);
nand U7965 (N_7965,N_7729,N_7703);
and U7966 (N_7966,N_7649,N_7656);
xnor U7967 (N_7967,N_7692,N_7650);
and U7968 (N_7968,N_7707,N_7695);
xnor U7969 (N_7969,N_7796,N_7665);
nor U7970 (N_7970,N_7673,N_7604);
or U7971 (N_7971,N_7727,N_7792);
or U7972 (N_7972,N_7680,N_7678);
and U7973 (N_7973,N_7624,N_7704);
nor U7974 (N_7974,N_7602,N_7746);
nand U7975 (N_7975,N_7776,N_7688);
and U7976 (N_7976,N_7622,N_7696);
or U7977 (N_7977,N_7739,N_7779);
nand U7978 (N_7978,N_7621,N_7659);
and U7979 (N_7979,N_7697,N_7663);
nor U7980 (N_7980,N_7629,N_7722);
nor U7981 (N_7981,N_7736,N_7780);
nor U7982 (N_7982,N_7788,N_7677);
and U7983 (N_7983,N_7666,N_7779);
and U7984 (N_7984,N_7692,N_7734);
xnor U7985 (N_7985,N_7652,N_7791);
or U7986 (N_7986,N_7671,N_7623);
xnor U7987 (N_7987,N_7660,N_7751);
or U7988 (N_7988,N_7677,N_7686);
nor U7989 (N_7989,N_7614,N_7727);
nor U7990 (N_7990,N_7789,N_7702);
nand U7991 (N_7991,N_7695,N_7708);
nor U7992 (N_7992,N_7641,N_7740);
nand U7993 (N_7993,N_7726,N_7772);
xor U7994 (N_7994,N_7620,N_7710);
nand U7995 (N_7995,N_7756,N_7667);
nand U7996 (N_7996,N_7702,N_7782);
or U7997 (N_7997,N_7740,N_7644);
nand U7998 (N_7998,N_7648,N_7640);
and U7999 (N_7999,N_7671,N_7780);
xor U8000 (N_8000,N_7822,N_7954);
nand U8001 (N_8001,N_7872,N_7987);
or U8002 (N_8002,N_7900,N_7887);
and U8003 (N_8003,N_7895,N_7858);
and U8004 (N_8004,N_7964,N_7871);
or U8005 (N_8005,N_7912,N_7849);
nor U8006 (N_8006,N_7970,N_7991);
and U8007 (N_8007,N_7807,N_7921);
or U8008 (N_8008,N_7853,N_7962);
nor U8009 (N_8009,N_7841,N_7878);
xnor U8010 (N_8010,N_7833,N_7832);
or U8011 (N_8011,N_7974,N_7862);
and U8012 (N_8012,N_7901,N_7930);
or U8013 (N_8013,N_7910,N_7886);
nand U8014 (N_8014,N_7811,N_7857);
or U8015 (N_8015,N_7920,N_7993);
or U8016 (N_8016,N_7927,N_7821);
xnor U8017 (N_8017,N_7983,N_7814);
nor U8018 (N_8018,N_7928,N_7976);
and U8019 (N_8019,N_7942,N_7864);
and U8020 (N_8020,N_7972,N_7997);
xnor U8021 (N_8021,N_7875,N_7968);
xor U8022 (N_8022,N_7955,N_7836);
and U8023 (N_8023,N_7916,N_7838);
xor U8024 (N_8024,N_7820,N_7933);
xor U8025 (N_8025,N_7937,N_7852);
and U8026 (N_8026,N_7996,N_7800);
nor U8027 (N_8027,N_7902,N_7881);
xnor U8028 (N_8028,N_7860,N_7845);
nor U8029 (N_8029,N_7948,N_7870);
and U8030 (N_8030,N_7950,N_7869);
and U8031 (N_8031,N_7868,N_7919);
or U8032 (N_8032,N_7911,N_7810);
xnor U8033 (N_8033,N_7913,N_7896);
xnor U8034 (N_8034,N_7889,N_7859);
and U8035 (N_8035,N_7877,N_7943);
and U8036 (N_8036,N_7961,N_7829);
nand U8037 (N_8037,N_7865,N_7866);
xor U8038 (N_8038,N_7893,N_7917);
or U8039 (N_8039,N_7844,N_7957);
nor U8040 (N_8040,N_7940,N_7932);
or U8041 (N_8041,N_7969,N_7978);
xor U8042 (N_8042,N_7922,N_7894);
nand U8043 (N_8043,N_7803,N_7817);
nor U8044 (N_8044,N_7826,N_7924);
and U8045 (N_8045,N_7890,N_7973);
nor U8046 (N_8046,N_7825,N_7882);
and U8047 (N_8047,N_7994,N_7958);
nor U8048 (N_8048,N_7952,N_7989);
nor U8049 (N_8049,N_7819,N_7876);
nand U8050 (N_8050,N_7884,N_7938);
nor U8051 (N_8051,N_7808,N_7984);
xnor U8052 (N_8052,N_7805,N_7986);
nand U8053 (N_8053,N_7963,N_7947);
and U8054 (N_8054,N_7892,N_7979);
or U8055 (N_8055,N_7944,N_7975);
nor U8056 (N_8056,N_7843,N_7899);
or U8057 (N_8057,N_7823,N_7966);
and U8058 (N_8058,N_7802,N_7846);
xor U8059 (N_8059,N_7842,N_7945);
nand U8060 (N_8060,N_7946,N_7809);
nor U8061 (N_8061,N_7813,N_7971);
nand U8062 (N_8062,N_7988,N_7831);
and U8063 (N_8063,N_7908,N_7873);
nor U8064 (N_8064,N_7982,N_7999);
xor U8065 (N_8065,N_7960,N_7804);
nor U8066 (N_8066,N_7941,N_7935);
and U8067 (N_8067,N_7897,N_7816);
and U8068 (N_8068,N_7830,N_7827);
and U8069 (N_8069,N_7981,N_7879);
nand U8070 (N_8070,N_7909,N_7874);
xnor U8071 (N_8071,N_7906,N_7848);
and U8072 (N_8072,N_7907,N_7939);
xor U8073 (N_8073,N_7936,N_7925);
nor U8074 (N_8074,N_7965,N_7905);
and U8075 (N_8075,N_7861,N_7835);
nor U8076 (N_8076,N_7904,N_7898);
nand U8077 (N_8077,N_7926,N_7918);
nor U8078 (N_8078,N_7923,N_7992);
xor U8079 (N_8079,N_7856,N_7998);
nor U8080 (N_8080,N_7914,N_7990);
and U8081 (N_8081,N_7847,N_7915);
nor U8082 (N_8082,N_7929,N_7959);
and U8083 (N_8083,N_7967,N_7812);
or U8084 (N_8084,N_7828,N_7806);
nand U8085 (N_8085,N_7888,N_7837);
nand U8086 (N_8086,N_7980,N_7977);
nand U8087 (N_8087,N_7891,N_7855);
nor U8088 (N_8088,N_7801,N_7839);
or U8089 (N_8089,N_7995,N_7818);
nor U8090 (N_8090,N_7931,N_7834);
nor U8091 (N_8091,N_7956,N_7854);
and U8092 (N_8092,N_7903,N_7985);
xor U8093 (N_8093,N_7953,N_7883);
nand U8094 (N_8094,N_7863,N_7880);
nor U8095 (N_8095,N_7951,N_7851);
nor U8096 (N_8096,N_7885,N_7824);
nand U8097 (N_8097,N_7949,N_7867);
xor U8098 (N_8098,N_7850,N_7815);
and U8099 (N_8099,N_7840,N_7934);
or U8100 (N_8100,N_7812,N_7996);
xor U8101 (N_8101,N_7906,N_7810);
and U8102 (N_8102,N_7971,N_7860);
nor U8103 (N_8103,N_7928,N_7875);
nor U8104 (N_8104,N_7937,N_7985);
xor U8105 (N_8105,N_7867,N_7807);
or U8106 (N_8106,N_7949,N_7857);
nor U8107 (N_8107,N_7863,N_7984);
nor U8108 (N_8108,N_7800,N_7859);
and U8109 (N_8109,N_7931,N_7952);
or U8110 (N_8110,N_7920,N_7888);
or U8111 (N_8111,N_7996,N_7910);
nor U8112 (N_8112,N_7880,N_7903);
and U8113 (N_8113,N_7958,N_7917);
and U8114 (N_8114,N_7840,N_7952);
nand U8115 (N_8115,N_7949,N_7879);
nor U8116 (N_8116,N_7891,N_7939);
nor U8117 (N_8117,N_7850,N_7946);
and U8118 (N_8118,N_7959,N_7992);
nand U8119 (N_8119,N_7862,N_7942);
nand U8120 (N_8120,N_7948,N_7982);
or U8121 (N_8121,N_7837,N_7868);
and U8122 (N_8122,N_7894,N_7815);
or U8123 (N_8123,N_7812,N_7893);
nand U8124 (N_8124,N_7961,N_7908);
xnor U8125 (N_8125,N_7963,N_7859);
xor U8126 (N_8126,N_7895,N_7876);
and U8127 (N_8127,N_7883,N_7875);
and U8128 (N_8128,N_7982,N_7847);
nor U8129 (N_8129,N_7931,N_7833);
and U8130 (N_8130,N_7980,N_7829);
or U8131 (N_8131,N_7966,N_7933);
xor U8132 (N_8132,N_7906,N_7815);
nand U8133 (N_8133,N_7901,N_7813);
nand U8134 (N_8134,N_7898,N_7916);
xor U8135 (N_8135,N_7815,N_7801);
nor U8136 (N_8136,N_7904,N_7837);
xor U8137 (N_8137,N_7818,N_7896);
or U8138 (N_8138,N_7872,N_7808);
nand U8139 (N_8139,N_7815,N_7948);
and U8140 (N_8140,N_7994,N_7944);
xnor U8141 (N_8141,N_7991,N_7897);
xnor U8142 (N_8142,N_7963,N_7804);
xnor U8143 (N_8143,N_7838,N_7851);
or U8144 (N_8144,N_7933,N_7821);
nand U8145 (N_8145,N_7820,N_7909);
xor U8146 (N_8146,N_7882,N_7953);
or U8147 (N_8147,N_7885,N_7997);
or U8148 (N_8148,N_7919,N_7952);
nand U8149 (N_8149,N_7967,N_7859);
or U8150 (N_8150,N_7845,N_7962);
xor U8151 (N_8151,N_7994,N_7826);
or U8152 (N_8152,N_7992,N_7859);
and U8153 (N_8153,N_7875,N_7817);
or U8154 (N_8154,N_7836,N_7933);
nor U8155 (N_8155,N_7805,N_7965);
nand U8156 (N_8156,N_7860,N_7949);
or U8157 (N_8157,N_7865,N_7848);
nand U8158 (N_8158,N_7991,N_7837);
xnor U8159 (N_8159,N_7865,N_7993);
nor U8160 (N_8160,N_7952,N_7903);
and U8161 (N_8161,N_7897,N_7804);
xor U8162 (N_8162,N_7804,N_7947);
and U8163 (N_8163,N_7815,N_7858);
nand U8164 (N_8164,N_7955,N_7871);
xor U8165 (N_8165,N_7855,N_7933);
or U8166 (N_8166,N_7977,N_7918);
and U8167 (N_8167,N_7857,N_7819);
nand U8168 (N_8168,N_7970,N_7886);
xor U8169 (N_8169,N_7842,N_7874);
nor U8170 (N_8170,N_7912,N_7802);
nand U8171 (N_8171,N_7978,N_7873);
nor U8172 (N_8172,N_7841,N_7965);
nand U8173 (N_8173,N_7859,N_7916);
and U8174 (N_8174,N_7960,N_7911);
nand U8175 (N_8175,N_7831,N_7973);
and U8176 (N_8176,N_7976,N_7990);
xnor U8177 (N_8177,N_7985,N_7954);
nor U8178 (N_8178,N_7980,N_7964);
xor U8179 (N_8179,N_7863,N_7928);
or U8180 (N_8180,N_7849,N_7929);
nor U8181 (N_8181,N_7986,N_7866);
or U8182 (N_8182,N_7881,N_7958);
xor U8183 (N_8183,N_7994,N_7910);
xor U8184 (N_8184,N_7833,N_7944);
nand U8185 (N_8185,N_7913,N_7902);
xor U8186 (N_8186,N_7841,N_7806);
or U8187 (N_8187,N_7959,N_7961);
and U8188 (N_8188,N_7860,N_7863);
nor U8189 (N_8189,N_7888,N_7891);
and U8190 (N_8190,N_7839,N_7867);
nor U8191 (N_8191,N_7842,N_7917);
and U8192 (N_8192,N_7950,N_7976);
xnor U8193 (N_8193,N_7894,N_7999);
nand U8194 (N_8194,N_7897,N_7859);
or U8195 (N_8195,N_7800,N_7821);
nand U8196 (N_8196,N_7893,N_7933);
and U8197 (N_8197,N_7832,N_7869);
nand U8198 (N_8198,N_7844,N_7984);
and U8199 (N_8199,N_7824,N_7844);
and U8200 (N_8200,N_8165,N_8031);
nor U8201 (N_8201,N_8037,N_8026);
nand U8202 (N_8202,N_8027,N_8196);
and U8203 (N_8203,N_8181,N_8113);
nand U8204 (N_8204,N_8016,N_8099);
and U8205 (N_8205,N_8182,N_8096);
xnor U8206 (N_8206,N_8043,N_8151);
or U8207 (N_8207,N_8140,N_8020);
xnor U8208 (N_8208,N_8157,N_8064);
xor U8209 (N_8209,N_8084,N_8105);
or U8210 (N_8210,N_8118,N_8090);
nand U8211 (N_8211,N_8056,N_8126);
or U8212 (N_8212,N_8022,N_8061);
nand U8213 (N_8213,N_8047,N_8005);
nor U8214 (N_8214,N_8039,N_8139);
and U8215 (N_8215,N_8094,N_8191);
and U8216 (N_8216,N_8193,N_8083);
and U8217 (N_8217,N_8173,N_8128);
or U8218 (N_8218,N_8018,N_8065);
or U8219 (N_8219,N_8098,N_8102);
and U8220 (N_8220,N_8198,N_8123);
or U8221 (N_8221,N_8058,N_8127);
or U8222 (N_8222,N_8046,N_8070);
nor U8223 (N_8223,N_8017,N_8186);
nand U8224 (N_8224,N_8121,N_8171);
nand U8225 (N_8225,N_8156,N_8132);
xor U8226 (N_8226,N_8095,N_8003);
and U8227 (N_8227,N_8066,N_8042);
nand U8228 (N_8228,N_8009,N_8142);
nand U8229 (N_8229,N_8041,N_8000);
nand U8230 (N_8230,N_8068,N_8082);
nand U8231 (N_8231,N_8073,N_8057);
and U8232 (N_8232,N_8115,N_8035);
and U8233 (N_8233,N_8010,N_8032);
or U8234 (N_8234,N_8087,N_8021);
xnor U8235 (N_8235,N_8122,N_8185);
xnor U8236 (N_8236,N_8166,N_8133);
and U8237 (N_8237,N_8164,N_8050);
nor U8238 (N_8238,N_8184,N_8081);
or U8239 (N_8239,N_8177,N_8153);
and U8240 (N_8240,N_8143,N_8135);
xor U8241 (N_8241,N_8008,N_8145);
and U8242 (N_8242,N_8012,N_8174);
nor U8243 (N_8243,N_8125,N_8036);
nor U8244 (N_8244,N_8108,N_8045);
nor U8245 (N_8245,N_8011,N_8162);
and U8246 (N_8246,N_8052,N_8188);
nor U8247 (N_8247,N_8054,N_8148);
or U8248 (N_8248,N_8024,N_8152);
and U8249 (N_8249,N_8110,N_8167);
and U8250 (N_8250,N_8030,N_8169);
xnor U8251 (N_8251,N_8100,N_8172);
nand U8252 (N_8252,N_8044,N_8154);
nor U8253 (N_8253,N_8025,N_8134);
xnor U8254 (N_8254,N_8116,N_8002);
or U8255 (N_8255,N_8195,N_8144);
nor U8256 (N_8256,N_8136,N_8161);
xor U8257 (N_8257,N_8120,N_8137);
and U8258 (N_8258,N_8138,N_8155);
nand U8259 (N_8259,N_8101,N_8053);
xnor U8260 (N_8260,N_8117,N_8033);
xnor U8261 (N_8261,N_8189,N_8063);
and U8262 (N_8262,N_8014,N_8075);
xnor U8263 (N_8263,N_8129,N_8176);
nand U8264 (N_8264,N_8006,N_8124);
nor U8265 (N_8265,N_8091,N_8158);
nor U8266 (N_8266,N_8079,N_8168);
xnor U8267 (N_8267,N_8106,N_8060);
or U8268 (N_8268,N_8114,N_8059);
or U8269 (N_8269,N_8112,N_8072);
nand U8270 (N_8270,N_8175,N_8170);
or U8271 (N_8271,N_8131,N_8055);
nand U8272 (N_8272,N_8004,N_8192);
or U8273 (N_8273,N_8062,N_8150);
xor U8274 (N_8274,N_8190,N_8104);
nand U8275 (N_8275,N_8147,N_8103);
nand U8276 (N_8276,N_8038,N_8141);
nand U8277 (N_8277,N_8092,N_8074);
and U8278 (N_8278,N_8160,N_8178);
and U8279 (N_8279,N_8159,N_8130);
or U8280 (N_8280,N_8048,N_8163);
nor U8281 (N_8281,N_8049,N_8076);
nand U8282 (N_8282,N_8109,N_8040);
or U8283 (N_8283,N_8107,N_8183);
nor U8284 (N_8284,N_8088,N_8051);
nor U8285 (N_8285,N_8199,N_8029);
and U8286 (N_8286,N_8019,N_8111);
and U8287 (N_8287,N_8007,N_8028);
nand U8288 (N_8288,N_8194,N_8078);
nor U8289 (N_8289,N_8093,N_8069);
xnor U8290 (N_8290,N_8197,N_8001);
nand U8291 (N_8291,N_8085,N_8089);
nor U8292 (N_8292,N_8013,N_8146);
or U8293 (N_8293,N_8097,N_8015);
and U8294 (N_8294,N_8119,N_8067);
xnor U8295 (N_8295,N_8034,N_8149);
nand U8296 (N_8296,N_8180,N_8071);
or U8297 (N_8297,N_8086,N_8023);
and U8298 (N_8298,N_8077,N_8179);
nand U8299 (N_8299,N_8187,N_8080);
and U8300 (N_8300,N_8034,N_8117);
nor U8301 (N_8301,N_8098,N_8125);
or U8302 (N_8302,N_8174,N_8002);
xor U8303 (N_8303,N_8084,N_8051);
nand U8304 (N_8304,N_8122,N_8190);
and U8305 (N_8305,N_8056,N_8157);
nor U8306 (N_8306,N_8106,N_8000);
or U8307 (N_8307,N_8115,N_8143);
nor U8308 (N_8308,N_8108,N_8093);
xor U8309 (N_8309,N_8115,N_8104);
nor U8310 (N_8310,N_8054,N_8034);
and U8311 (N_8311,N_8079,N_8148);
nand U8312 (N_8312,N_8156,N_8196);
and U8313 (N_8313,N_8142,N_8044);
xor U8314 (N_8314,N_8184,N_8015);
or U8315 (N_8315,N_8083,N_8136);
and U8316 (N_8316,N_8004,N_8105);
xnor U8317 (N_8317,N_8143,N_8136);
nor U8318 (N_8318,N_8169,N_8124);
and U8319 (N_8319,N_8082,N_8190);
nand U8320 (N_8320,N_8171,N_8070);
nor U8321 (N_8321,N_8141,N_8000);
nor U8322 (N_8322,N_8146,N_8047);
or U8323 (N_8323,N_8197,N_8158);
nand U8324 (N_8324,N_8180,N_8150);
or U8325 (N_8325,N_8052,N_8056);
xnor U8326 (N_8326,N_8150,N_8133);
and U8327 (N_8327,N_8179,N_8116);
nor U8328 (N_8328,N_8081,N_8098);
xor U8329 (N_8329,N_8023,N_8166);
or U8330 (N_8330,N_8022,N_8070);
nand U8331 (N_8331,N_8136,N_8016);
xor U8332 (N_8332,N_8197,N_8190);
nor U8333 (N_8333,N_8156,N_8138);
and U8334 (N_8334,N_8044,N_8144);
nor U8335 (N_8335,N_8036,N_8017);
or U8336 (N_8336,N_8027,N_8180);
nand U8337 (N_8337,N_8173,N_8123);
nand U8338 (N_8338,N_8085,N_8071);
nor U8339 (N_8339,N_8135,N_8149);
nand U8340 (N_8340,N_8113,N_8175);
or U8341 (N_8341,N_8110,N_8008);
nand U8342 (N_8342,N_8024,N_8193);
or U8343 (N_8343,N_8121,N_8001);
nor U8344 (N_8344,N_8106,N_8027);
or U8345 (N_8345,N_8096,N_8125);
xnor U8346 (N_8346,N_8048,N_8164);
nand U8347 (N_8347,N_8189,N_8131);
nand U8348 (N_8348,N_8101,N_8120);
nand U8349 (N_8349,N_8155,N_8157);
nand U8350 (N_8350,N_8053,N_8001);
or U8351 (N_8351,N_8009,N_8096);
nor U8352 (N_8352,N_8039,N_8010);
nand U8353 (N_8353,N_8162,N_8145);
nor U8354 (N_8354,N_8101,N_8158);
xor U8355 (N_8355,N_8177,N_8023);
xnor U8356 (N_8356,N_8196,N_8070);
and U8357 (N_8357,N_8070,N_8167);
nand U8358 (N_8358,N_8063,N_8030);
and U8359 (N_8359,N_8033,N_8069);
and U8360 (N_8360,N_8008,N_8100);
nor U8361 (N_8361,N_8053,N_8116);
nor U8362 (N_8362,N_8189,N_8029);
xor U8363 (N_8363,N_8068,N_8072);
xnor U8364 (N_8364,N_8167,N_8108);
xor U8365 (N_8365,N_8010,N_8158);
or U8366 (N_8366,N_8180,N_8123);
nor U8367 (N_8367,N_8098,N_8042);
nand U8368 (N_8368,N_8028,N_8117);
nand U8369 (N_8369,N_8153,N_8070);
or U8370 (N_8370,N_8061,N_8109);
xnor U8371 (N_8371,N_8147,N_8119);
and U8372 (N_8372,N_8115,N_8141);
xnor U8373 (N_8373,N_8046,N_8022);
xor U8374 (N_8374,N_8177,N_8192);
or U8375 (N_8375,N_8047,N_8089);
nand U8376 (N_8376,N_8152,N_8194);
xor U8377 (N_8377,N_8019,N_8131);
or U8378 (N_8378,N_8089,N_8155);
and U8379 (N_8379,N_8168,N_8123);
nand U8380 (N_8380,N_8045,N_8113);
or U8381 (N_8381,N_8007,N_8153);
and U8382 (N_8382,N_8182,N_8192);
or U8383 (N_8383,N_8090,N_8107);
and U8384 (N_8384,N_8105,N_8139);
nor U8385 (N_8385,N_8034,N_8051);
nand U8386 (N_8386,N_8113,N_8023);
and U8387 (N_8387,N_8085,N_8126);
xnor U8388 (N_8388,N_8183,N_8169);
nor U8389 (N_8389,N_8101,N_8079);
nand U8390 (N_8390,N_8055,N_8108);
nand U8391 (N_8391,N_8071,N_8069);
xor U8392 (N_8392,N_8137,N_8141);
xnor U8393 (N_8393,N_8079,N_8080);
xor U8394 (N_8394,N_8078,N_8108);
xnor U8395 (N_8395,N_8154,N_8199);
nor U8396 (N_8396,N_8070,N_8198);
and U8397 (N_8397,N_8107,N_8197);
or U8398 (N_8398,N_8049,N_8005);
nor U8399 (N_8399,N_8132,N_8166);
nand U8400 (N_8400,N_8308,N_8220);
or U8401 (N_8401,N_8242,N_8365);
xnor U8402 (N_8402,N_8265,N_8328);
nand U8403 (N_8403,N_8344,N_8299);
xor U8404 (N_8404,N_8288,N_8310);
and U8405 (N_8405,N_8259,N_8213);
nor U8406 (N_8406,N_8315,N_8227);
or U8407 (N_8407,N_8396,N_8290);
xor U8408 (N_8408,N_8364,N_8331);
nand U8409 (N_8409,N_8380,N_8292);
nor U8410 (N_8410,N_8234,N_8203);
and U8411 (N_8411,N_8267,N_8313);
nor U8412 (N_8412,N_8384,N_8352);
and U8413 (N_8413,N_8363,N_8230);
nor U8414 (N_8414,N_8258,N_8362);
or U8415 (N_8415,N_8266,N_8335);
and U8416 (N_8416,N_8272,N_8371);
nand U8417 (N_8417,N_8249,N_8302);
or U8418 (N_8418,N_8238,N_8314);
xnor U8419 (N_8419,N_8337,N_8354);
xor U8420 (N_8420,N_8255,N_8205);
xnor U8421 (N_8421,N_8274,N_8260);
xor U8422 (N_8422,N_8296,N_8221);
or U8423 (N_8423,N_8253,N_8254);
xor U8424 (N_8424,N_8357,N_8273);
nor U8425 (N_8425,N_8211,N_8316);
xnor U8426 (N_8426,N_8360,N_8386);
xnor U8427 (N_8427,N_8324,N_8368);
xor U8428 (N_8428,N_8398,N_8372);
or U8429 (N_8429,N_8370,N_8291);
or U8430 (N_8430,N_8226,N_8341);
nor U8431 (N_8431,N_8275,N_8224);
or U8432 (N_8432,N_8228,N_8252);
or U8433 (N_8433,N_8369,N_8319);
nand U8434 (N_8434,N_8340,N_8367);
xor U8435 (N_8435,N_8209,N_8350);
nand U8436 (N_8436,N_8235,N_8218);
xor U8437 (N_8437,N_8347,N_8378);
and U8438 (N_8438,N_8321,N_8358);
xnor U8439 (N_8439,N_8286,N_8373);
xor U8440 (N_8440,N_8217,N_8387);
xor U8441 (N_8441,N_8293,N_8216);
and U8442 (N_8442,N_8261,N_8222);
and U8443 (N_8443,N_8244,N_8332);
or U8444 (N_8444,N_8317,N_8379);
and U8445 (N_8445,N_8377,N_8200);
nor U8446 (N_8446,N_8338,N_8279);
xnor U8447 (N_8447,N_8329,N_8283);
and U8448 (N_8448,N_8382,N_8393);
and U8449 (N_8449,N_8256,N_8241);
nand U8450 (N_8450,N_8269,N_8355);
and U8451 (N_8451,N_8215,N_8278);
nand U8452 (N_8452,N_8246,N_8305);
nor U8453 (N_8453,N_8229,N_8351);
nand U8454 (N_8454,N_8298,N_8207);
nand U8455 (N_8455,N_8346,N_8281);
and U8456 (N_8456,N_8276,N_8223);
xor U8457 (N_8457,N_8326,N_8202);
nor U8458 (N_8458,N_8348,N_8243);
and U8459 (N_8459,N_8270,N_8320);
or U8460 (N_8460,N_8214,N_8312);
xnor U8461 (N_8461,N_8233,N_8376);
or U8462 (N_8462,N_8389,N_8264);
or U8463 (N_8463,N_8394,N_8277);
nor U8464 (N_8464,N_8391,N_8271);
or U8465 (N_8465,N_8322,N_8353);
nor U8466 (N_8466,N_8388,N_8250);
nor U8467 (N_8467,N_8232,N_8361);
xnor U8468 (N_8468,N_8301,N_8300);
xor U8469 (N_8469,N_8306,N_8383);
or U8470 (N_8470,N_8311,N_8297);
xnor U8471 (N_8471,N_8206,N_8374);
xor U8472 (N_8472,N_8231,N_8289);
nand U8473 (N_8473,N_8294,N_8240);
nor U8474 (N_8474,N_8304,N_8247);
and U8475 (N_8475,N_8345,N_8257);
xnor U8476 (N_8476,N_8236,N_8263);
or U8477 (N_8477,N_8339,N_8295);
nand U8478 (N_8478,N_8284,N_8208);
nor U8479 (N_8479,N_8325,N_8285);
xnor U8480 (N_8480,N_8323,N_8334);
nand U8481 (N_8481,N_8333,N_8280);
nand U8482 (N_8482,N_8366,N_8330);
xor U8483 (N_8483,N_8239,N_8307);
nand U8484 (N_8484,N_8210,N_8262);
nor U8485 (N_8485,N_8342,N_8381);
or U8486 (N_8486,N_8309,N_8399);
or U8487 (N_8487,N_8219,N_8356);
xnor U8488 (N_8488,N_8375,N_8251);
and U8489 (N_8489,N_8397,N_8359);
and U8490 (N_8490,N_8390,N_8343);
xnor U8491 (N_8491,N_8204,N_8201);
nor U8492 (N_8492,N_8282,N_8385);
xor U8493 (N_8493,N_8248,N_8268);
nor U8494 (N_8494,N_8392,N_8237);
nand U8495 (N_8495,N_8349,N_8395);
or U8496 (N_8496,N_8303,N_8318);
or U8497 (N_8497,N_8336,N_8287);
or U8498 (N_8498,N_8225,N_8327);
xor U8499 (N_8499,N_8212,N_8245);
nor U8500 (N_8500,N_8281,N_8227);
nor U8501 (N_8501,N_8253,N_8350);
nand U8502 (N_8502,N_8291,N_8334);
or U8503 (N_8503,N_8356,N_8245);
or U8504 (N_8504,N_8382,N_8352);
nand U8505 (N_8505,N_8349,N_8302);
nand U8506 (N_8506,N_8266,N_8374);
or U8507 (N_8507,N_8316,N_8376);
xnor U8508 (N_8508,N_8371,N_8257);
and U8509 (N_8509,N_8227,N_8286);
nand U8510 (N_8510,N_8282,N_8291);
nand U8511 (N_8511,N_8214,N_8389);
or U8512 (N_8512,N_8322,N_8220);
nand U8513 (N_8513,N_8358,N_8285);
or U8514 (N_8514,N_8308,N_8321);
nand U8515 (N_8515,N_8239,N_8295);
xor U8516 (N_8516,N_8355,N_8322);
nor U8517 (N_8517,N_8360,N_8272);
xor U8518 (N_8518,N_8238,N_8274);
xnor U8519 (N_8519,N_8271,N_8277);
xnor U8520 (N_8520,N_8340,N_8225);
and U8521 (N_8521,N_8380,N_8225);
and U8522 (N_8522,N_8266,N_8249);
nor U8523 (N_8523,N_8380,N_8228);
or U8524 (N_8524,N_8237,N_8243);
and U8525 (N_8525,N_8210,N_8213);
and U8526 (N_8526,N_8345,N_8367);
nand U8527 (N_8527,N_8292,N_8382);
or U8528 (N_8528,N_8314,N_8269);
xnor U8529 (N_8529,N_8254,N_8290);
nor U8530 (N_8530,N_8390,N_8268);
xnor U8531 (N_8531,N_8253,N_8219);
and U8532 (N_8532,N_8318,N_8291);
nor U8533 (N_8533,N_8202,N_8205);
nor U8534 (N_8534,N_8289,N_8277);
and U8535 (N_8535,N_8353,N_8385);
and U8536 (N_8536,N_8201,N_8271);
nor U8537 (N_8537,N_8262,N_8269);
nor U8538 (N_8538,N_8252,N_8283);
nand U8539 (N_8539,N_8270,N_8272);
nor U8540 (N_8540,N_8325,N_8383);
xnor U8541 (N_8541,N_8230,N_8239);
xor U8542 (N_8542,N_8207,N_8299);
xnor U8543 (N_8543,N_8350,N_8240);
and U8544 (N_8544,N_8346,N_8378);
or U8545 (N_8545,N_8377,N_8395);
and U8546 (N_8546,N_8371,N_8275);
nand U8547 (N_8547,N_8368,N_8358);
or U8548 (N_8548,N_8342,N_8254);
or U8549 (N_8549,N_8211,N_8268);
nand U8550 (N_8550,N_8388,N_8277);
or U8551 (N_8551,N_8223,N_8362);
nor U8552 (N_8552,N_8229,N_8336);
xor U8553 (N_8553,N_8362,N_8284);
or U8554 (N_8554,N_8212,N_8333);
and U8555 (N_8555,N_8306,N_8295);
and U8556 (N_8556,N_8288,N_8359);
nand U8557 (N_8557,N_8359,N_8341);
nand U8558 (N_8558,N_8286,N_8355);
nand U8559 (N_8559,N_8263,N_8299);
and U8560 (N_8560,N_8379,N_8304);
nand U8561 (N_8561,N_8289,N_8389);
xor U8562 (N_8562,N_8282,N_8328);
xnor U8563 (N_8563,N_8357,N_8291);
nor U8564 (N_8564,N_8271,N_8317);
nand U8565 (N_8565,N_8221,N_8397);
nor U8566 (N_8566,N_8319,N_8314);
and U8567 (N_8567,N_8200,N_8239);
xnor U8568 (N_8568,N_8220,N_8329);
xnor U8569 (N_8569,N_8242,N_8318);
nand U8570 (N_8570,N_8328,N_8235);
nor U8571 (N_8571,N_8358,N_8355);
and U8572 (N_8572,N_8222,N_8308);
or U8573 (N_8573,N_8263,N_8261);
xnor U8574 (N_8574,N_8322,N_8258);
nand U8575 (N_8575,N_8386,N_8374);
nand U8576 (N_8576,N_8221,N_8279);
nand U8577 (N_8577,N_8359,N_8223);
xnor U8578 (N_8578,N_8310,N_8238);
xnor U8579 (N_8579,N_8258,N_8265);
or U8580 (N_8580,N_8379,N_8345);
and U8581 (N_8581,N_8307,N_8387);
and U8582 (N_8582,N_8231,N_8273);
nor U8583 (N_8583,N_8270,N_8221);
and U8584 (N_8584,N_8333,N_8343);
nor U8585 (N_8585,N_8395,N_8266);
or U8586 (N_8586,N_8365,N_8360);
nand U8587 (N_8587,N_8309,N_8249);
nand U8588 (N_8588,N_8300,N_8252);
xnor U8589 (N_8589,N_8208,N_8211);
nor U8590 (N_8590,N_8338,N_8395);
or U8591 (N_8591,N_8394,N_8249);
or U8592 (N_8592,N_8204,N_8288);
or U8593 (N_8593,N_8303,N_8397);
or U8594 (N_8594,N_8381,N_8324);
or U8595 (N_8595,N_8297,N_8326);
xnor U8596 (N_8596,N_8380,N_8224);
nor U8597 (N_8597,N_8214,N_8358);
xor U8598 (N_8598,N_8226,N_8274);
and U8599 (N_8599,N_8363,N_8350);
nand U8600 (N_8600,N_8591,N_8429);
or U8601 (N_8601,N_8515,N_8478);
xnor U8602 (N_8602,N_8483,N_8406);
or U8603 (N_8603,N_8400,N_8412);
nand U8604 (N_8604,N_8596,N_8566);
nand U8605 (N_8605,N_8492,N_8595);
xor U8606 (N_8606,N_8403,N_8507);
nand U8607 (N_8607,N_8580,N_8466);
xnor U8608 (N_8608,N_8567,N_8484);
xnor U8609 (N_8609,N_8474,N_8442);
nor U8610 (N_8610,N_8405,N_8565);
nand U8611 (N_8611,N_8419,N_8527);
nand U8612 (N_8612,N_8417,N_8531);
xor U8613 (N_8613,N_8587,N_8488);
nor U8614 (N_8614,N_8582,N_8509);
and U8615 (N_8615,N_8516,N_8409);
xnor U8616 (N_8616,N_8577,N_8413);
nand U8617 (N_8617,N_8575,N_8514);
nand U8618 (N_8618,N_8557,N_8414);
or U8619 (N_8619,N_8511,N_8501);
nand U8620 (N_8620,N_8598,N_8599);
nor U8621 (N_8621,N_8467,N_8505);
and U8622 (N_8622,N_8427,N_8537);
xnor U8623 (N_8623,N_8446,N_8506);
or U8624 (N_8624,N_8482,N_8435);
nand U8625 (N_8625,N_8408,N_8451);
or U8626 (N_8626,N_8593,N_8562);
and U8627 (N_8627,N_8493,N_8533);
nor U8628 (N_8628,N_8545,N_8581);
and U8629 (N_8629,N_8401,N_8423);
nor U8630 (N_8630,N_8463,N_8495);
nand U8631 (N_8631,N_8473,N_8535);
nand U8632 (N_8632,N_8512,N_8592);
nor U8633 (N_8633,N_8547,N_8583);
nand U8634 (N_8634,N_8458,N_8444);
nor U8635 (N_8635,N_8540,N_8447);
nor U8636 (N_8636,N_8574,N_8499);
nand U8637 (N_8637,N_8550,N_8510);
nor U8638 (N_8638,N_8569,N_8472);
nor U8639 (N_8639,N_8420,N_8462);
nor U8640 (N_8640,N_8411,N_8520);
and U8641 (N_8641,N_8441,N_8498);
nor U8642 (N_8642,N_8572,N_8448);
or U8643 (N_8643,N_8502,N_8486);
and U8644 (N_8644,N_8496,N_8563);
or U8645 (N_8645,N_8439,N_8558);
nor U8646 (N_8646,N_8404,N_8469);
and U8647 (N_8647,N_8489,N_8526);
xnor U8648 (N_8648,N_8454,N_8544);
nand U8649 (N_8649,N_8437,N_8538);
and U8650 (N_8650,N_8559,N_8443);
xnor U8651 (N_8651,N_8532,N_8530);
and U8652 (N_8652,N_8428,N_8543);
xnor U8653 (N_8653,N_8534,N_8546);
or U8654 (N_8654,N_8578,N_8571);
xor U8655 (N_8655,N_8433,N_8576);
nand U8656 (N_8656,N_8480,N_8518);
and U8657 (N_8657,N_8457,N_8584);
and U8658 (N_8658,N_8568,N_8471);
and U8659 (N_8659,N_8553,N_8468);
nand U8660 (N_8660,N_8524,N_8453);
nand U8661 (N_8661,N_8438,N_8497);
nor U8662 (N_8662,N_8551,N_8464);
xnor U8663 (N_8663,N_8589,N_8561);
xor U8664 (N_8664,N_8449,N_8426);
nor U8665 (N_8665,N_8432,N_8421);
nor U8666 (N_8666,N_8564,N_8586);
or U8667 (N_8667,N_8536,N_8475);
nand U8668 (N_8668,N_8477,N_8523);
nor U8669 (N_8669,N_8422,N_8425);
and U8670 (N_8670,N_8415,N_8542);
nor U8671 (N_8671,N_8500,N_8430);
and U8672 (N_8672,N_8487,N_8424);
nand U8673 (N_8673,N_8445,N_8560);
and U8674 (N_8674,N_8456,N_8416);
nor U8675 (N_8675,N_8418,N_8555);
or U8676 (N_8676,N_8490,N_8573);
or U8677 (N_8677,N_8450,N_8597);
nand U8678 (N_8678,N_8552,N_8556);
nor U8679 (N_8679,N_8594,N_8579);
and U8680 (N_8680,N_8407,N_8479);
nand U8681 (N_8681,N_8476,N_8402);
and U8682 (N_8682,N_8548,N_8460);
xor U8683 (N_8683,N_8541,N_8461);
nor U8684 (N_8684,N_8522,N_8491);
or U8685 (N_8685,N_8434,N_8554);
and U8686 (N_8686,N_8539,N_8590);
and U8687 (N_8687,N_8517,N_8481);
nor U8688 (N_8688,N_8494,N_8508);
or U8689 (N_8689,N_8519,N_8513);
xor U8690 (N_8690,N_8585,N_8504);
and U8691 (N_8691,N_8410,N_8570);
xnor U8692 (N_8692,N_8588,N_8440);
nand U8693 (N_8693,N_8529,N_8549);
or U8694 (N_8694,N_8525,N_8465);
xnor U8695 (N_8695,N_8521,N_8470);
xor U8696 (N_8696,N_8485,N_8503);
or U8697 (N_8697,N_8431,N_8436);
nand U8698 (N_8698,N_8528,N_8455);
nand U8699 (N_8699,N_8452,N_8459);
nand U8700 (N_8700,N_8522,N_8599);
xor U8701 (N_8701,N_8599,N_8442);
nand U8702 (N_8702,N_8472,N_8511);
nor U8703 (N_8703,N_8472,N_8471);
and U8704 (N_8704,N_8414,N_8507);
nor U8705 (N_8705,N_8579,N_8592);
and U8706 (N_8706,N_8572,N_8436);
or U8707 (N_8707,N_8540,N_8549);
or U8708 (N_8708,N_8578,N_8594);
nand U8709 (N_8709,N_8462,N_8537);
xor U8710 (N_8710,N_8523,N_8414);
or U8711 (N_8711,N_8454,N_8596);
xnor U8712 (N_8712,N_8533,N_8582);
nand U8713 (N_8713,N_8570,N_8492);
nand U8714 (N_8714,N_8439,N_8433);
xor U8715 (N_8715,N_8422,N_8488);
nor U8716 (N_8716,N_8591,N_8454);
and U8717 (N_8717,N_8534,N_8472);
nor U8718 (N_8718,N_8437,N_8400);
and U8719 (N_8719,N_8405,N_8587);
nand U8720 (N_8720,N_8542,N_8432);
nor U8721 (N_8721,N_8461,N_8531);
and U8722 (N_8722,N_8560,N_8490);
xnor U8723 (N_8723,N_8435,N_8501);
and U8724 (N_8724,N_8417,N_8480);
nor U8725 (N_8725,N_8501,N_8554);
or U8726 (N_8726,N_8495,N_8571);
and U8727 (N_8727,N_8596,N_8589);
nor U8728 (N_8728,N_8441,N_8474);
xor U8729 (N_8729,N_8500,N_8453);
or U8730 (N_8730,N_8519,N_8457);
xnor U8731 (N_8731,N_8570,N_8416);
nor U8732 (N_8732,N_8404,N_8491);
nor U8733 (N_8733,N_8486,N_8568);
or U8734 (N_8734,N_8557,N_8408);
or U8735 (N_8735,N_8458,N_8566);
and U8736 (N_8736,N_8471,N_8597);
xor U8737 (N_8737,N_8452,N_8479);
and U8738 (N_8738,N_8460,N_8520);
xor U8739 (N_8739,N_8560,N_8419);
nor U8740 (N_8740,N_8445,N_8589);
and U8741 (N_8741,N_8515,N_8503);
nand U8742 (N_8742,N_8564,N_8528);
xnor U8743 (N_8743,N_8403,N_8485);
or U8744 (N_8744,N_8569,N_8578);
xor U8745 (N_8745,N_8538,N_8431);
nand U8746 (N_8746,N_8493,N_8527);
and U8747 (N_8747,N_8531,N_8497);
nor U8748 (N_8748,N_8591,N_8543);
nor U8749 (N_8749,N_8429,N_8599);
and U8750 (N_8750,N_8506,N_8468);
nor U8751 (N_8751,N_8486,N_8445);
or U8752 (N_8752,N_8434,N_8468);
nor U8753 (N_8753,N_8552,N_8415);
nand U8754 (N_8754,N_8459,N_8469);
or U8755 (N_8755,N_8448,N_8483);
or U8756 (N_8756,N_8477,N_8443);
or U8757 (N_8757,N_8445,N_8449);
and U8758 (N_8758,N_8495,N_8472);
nand U8759 (N_8759,N_8404,N_8541);
or U8760 (N_8760,N_8524,N_8467);
nand U8761 (N_8761,N_8440,N_8404);
and U8762 (N_8762,N_8447,N_8599);
nor U8763 (N_8763,N_8594,N_8526);
xor U8764 (N_8764,N_8597,N_8488);
nor U8765 (N_8765,N_8476,N_8509);
and U8766 (N_8766,N_8466,N_8480);
and U8767 (N_8767,N_8489,N_8561);
and U8768 (N_8768,N_8574,N_8567);
nor U8769 (N_8769,N_8436,N_8479);
and U8770 (N_8770,N_8531,N_8412);
or U8771 (N_8771,N_8455,N_8490);
xor U8772 (N_8772,N_8483,N_8562);
and U8773 (N_8773,N_8544,N_8469);
nand U8774 (N_8774,N_8488,N_8555);
xor U8775 (N_8775,N_8578,N_8499);
xor U8776 (N_8776,N_8469,N_8458);
and U8777 (N_8777,N_8556,N_8500);
nor U8778 (N_8778,N_8551,N_8460);
nor U8779 (N_8779,N_8428,N_8592);
nand U8780 (N_8780,N_8454,N_8505);
nor U8781 (N_8781,N_8598,N_8590);
xnor U8782 (N_8782,N_8474,N_8517);
and U8783 (N_8783,N_8404,N_8547);
nor U8784 (N_8784,N_8488,N_8539);
xnor U8785 (N_8785,N_8556,N_8580);
or U8786 (N_8786,N_8562,N_8440);
xnor U8787 (N_8787,N_8534,N_8426);
or U8788 (N_8788,N_8552,N_8402);
nor U8789 (N_8789,N_8557,N_8486);
or U8790 (N_8790,N_8536,N_8488);
and U8791 (N_8791,N_8424,N_8568);
xnor U8792 (N_8792,N_8456,N_8574);
or U8793 (N_8793,N_8544,N_8586);
nand U8794 (N_8794,N_8419,N_8420);
or U8795 (N_8795,N_8420,N_8555);
or U8796 (N_8796,N_8584,N_8429);
or U8797 (N_8797,N_8501,N_8484);
nor U8798 (N_8798,N_8516,N_8592);
nand U8799 (N_8799,N_8486,N_8522);
xor U8800 (N_8800,N_8601,N_8714);
nor U8801 (N_8801,N_8639,N_8759);
xnor U8802 (N_8802,N_8700,N_8726);
or U8803 (N_8803,N_8669,N_8785);
nor U8804 (N_8804,N_8768,N_8612);
nor U8805 (N_8805,N_8711,N_8692);
nor U8806 (N_8806,N_8678,N_8771);
and U8807 (N_8807,N_8615,N_8741);
or U8808 (N_8808,N_8790,N_8701);
and U8809 (N_8809,N_8721,N_8655);
nand U8810 (N_8810,N_8732,N_8689);
xor U8811 (N_8811,N_8784,N_8789);
nor U8812 (N_8812,N_8608,N_8611);
and U8813 (N_8813,N_8781,N_8643);
nand U8814 (N_8814,N_8753,N_8691);
and U8815 (N_8815,N_8617,N_8751);
xnor U8816 (N_8816,N_8645,N_8738);
nor U8817 (N_8817,N_8610,N_8776);
nand U8818 (N_8818,N_8736,N_8698);
nand U8819 (N_8819,N_8798,N_8631);
nor U8820 (N_8820,N_8740,N_8687);
xor U8821 (N_8821,N_8635,N_8626);
nor U8822 (N_8822,N_8719,N_8630);
xnor U8823 (N_8823,N_8760,N_8782);
nand U8824 (N_8824,N_8675,N_8683);
nor U8825 (N_8825,N_8793,N_8727);
nor U8826 (N_8826,N_8786,N_8702);
nand U8827 (N_8827,N_8684,N_8797);
nor U8828 (N_8828,N_8642,N_8734);
nor U8829 (N_8829,N_8715,N_8633);
or U8830 (N_8830,N_8706,N_8616);
or U8831 (N_8831,N_8624,N_8755);
and U8832 (N_8832,N_8762,N_8713);
nand U8833 (N_8833,N_8757,N_8622);
or U8834 (N_8834,N_8685,N_8653);
or U8835 (N_8835,N_8688,N_8764);
nor U8836 (N_8836,N_8662,N_8614);
and U8837 (N_8837,N_8660,N_8791);
nor U8838 (N_8838,N_8632,N_8658);
xnor U8839 (N_8839,N_8703,N_8694);
nor U8840 (N_8840,N_8665,N_8603);
nor U8841 (N_8841,N_8609,N_8710);
or U8842 (N_8842,N_8627,N_8628);
nand U8843 (N_8843,N_8750,N_8663);
nand U8844 (N_8844,N_8780,N_8772);
xor U8845 (N_8845,N_8697,N_8657);
or U8846 (N_8846,N_8605,N_8725);
and U8847 (N_8847,N_8641,N_8766);
nor U8848 (N_8848,N_8744,N_8668);
xor U8849 (N_8849,N_8718,N_8625);
or U8850 (N_8850,N_8723,N_8746);
nor U8851 (N_8851,N_8705,N_8737);
or U8852 (N_8852,N_8752,N_8777);
nor U8853 (N_8853,N_8717,N_8681);
nand U8854 (N_8854,N_8739,N_8621);
nor U8855 (N_8855,N_8792,N_8613);
nor U8856 (N_8856,N_8730,N_8620);
or U8857 (N_8857,N_8699,N_8656);
xor U8858 (N_8858,N_8795,N_8619);
and U8859 (N_8859,N_8644,N_8720);
xor U8860 (N_8860,N_8783,N_8646);
xnor U8861 (N_8861,N_8659,N_8788);
or U8862 (N_8862,N_8634,N_8763);
nor U8863 (N_8863,N_8724,N_8667);
nor U8864 (N_8864,N_8629,N_8652);
nor U8865 (N_8865,N_8770,N_8636);
nor U8866 (N_8866,N_8745,N_8649);
nor U8867 (N_8867,N_8775,N_8661);
nand U8868 (N_8868,N_8618,N_8765);
and U8869 (N_8869,N_8742,N_8679);
or U8870 (N_8870,N_8607,N_8693);
nand U8871 (N_8871,N_8637,N_8638);
nor U8872 (N_8872,N_8754,N_8606);
nor U8873 (N_8873,N_8794,N_8704);
nand U8874 (N_8874,N_8749,N_8674);
nor U8875 (N_8875,N_8735,N_8716);
or U8876 (N_8876,N_8767,N_8650);
xor U8877 (N_8877,N_8731,N_8729);
nand U8878 (N_8878,N_8670,N_8696);
and U8879 (N_8879,N_8682,N_8680);
nor U8880 (N_8880,N_8787,N_8651);
and U8881 (N_8881,N_8671,N_8796);
or U8882 (N_8882,N_8602,N_8677);
xnor U8883 (N_8883,N_8623,N_8756);
or U8884 (N_8884,N_8769,N_8712);
nand U8885 (N_8885,N_8640,N_8707);
or U8886 (N_8886,N_8648,N_8690);
nor U8887 (N_8887,N_8778,N_8774);
xor U8888 (N_8888,N_8743,N_8654);
nand U8889 (N_8889,N_8748,N_8779);
and U8890 (N_8890,N_8728,N_8672);
nor U8891 (N_8891,N_8747,N_8722);
nor U8892 (N_8892,N_8758,N_8708);
nor U8893 (N_8893,N_8686,N_8664);
and U8894 (N_8894,N_8600,N_8799);
and U8895 (N_8895,N_8647,N_8773);
or U8896 (N_8896,N_8709,N_8676);
xnor U8897 (N_8897,N_8666,N_8673);
nand U8898 (N_8898,N_8695,N_8761);
nand U8899 (N_8899,N_8733,N_8604);
or U8900 (N_8900,N_8618,N_8650);
nand U8901 (N_8901,N_8700,N_8617);
and U8902 (N_8902,N_8728,N_8723);
nor U8903 (N_8903,N_8781,N_8617);
or U8904 (N_8904,N_8647,N_8702);
nand U8905 (N_8905,N_8609,N_8699);
nand U8906 (N_8906,N_8626,N_8659);
and U8907 (N_8907,N_8645,N_8656);
and U8908 (N_8908,N_8733,N_8765);
or U8909 (N_8909,N_8725,N_8774);
xor U8910 (N_8910,N_8682,N_8746);
xor U8911 (N_8911,N_8670,N_8694);
xor U8912 (N_8912,N_8629,N_8745);
nor U8913 (N_8913,N_8607,N_8653);
nor U8914 (N_8914,N_8667,N_8676);
nor U8915 (N_8915,N_8784,N_8793);
and U8916 (N_8916,N_8606,N_8643);
xnor U8917 (N_8917,N_8707,N_8784);
and U8918 (N_8918,N_8712,N_8683);
xnor U8919 (N_8919,N_8634,N_8721);
nand U8920 (N_8920,N_8734,N_8671);
and U8921 (N_8921,N_8796,N_8734);
xor U8922 (N_8922,N_8777,N_8698);
xor U8923 (N_8923,N_8733,N_8686);
nand U8924 (N_8924,N_8733,N_8739);
nor U8925 (N_8925,N_8604,N_8616);
nand U8926 (N_8926,N_8636,N_8639);
nor U8927 (N_8927,N_8720,N_8658);
and U8928 (N_8928,N_8704,N_8667);
xnor U8929 (N_8929,N_8685,N_8675);
nor U8930 (N_8930,N_8734,N_8602);
nor U8931 (N_8931,N_8631,N_8703);
and U8932 (N_8932,N_8684,N_8641);
nand U8933 (N_8933,N_8625,N_8719);
and U8934 (N_8934,N_8646,N_8762);
xor U8935 (N_8935,N_8724,N_8796);
xnor U8936 (N_8936,N_8700,N_8702);
and U8937 (N_8937,N_8624,N_8738);
nor U8938 (N_8938,N_8799,N_8642);
and U8939 (N_8939,N_8609,N_8633);
or U8940 (N_8940,N_8784,N_8770);
nor U8941 (N_8941,N_8782,N_8751);
and U8942 (N_8942,N_8787,N_8608);
or U8943 (N_8943,N_8602,N_8609);
or U8944 (N_8944,N_8710,N_8628);
and U8945 (N_8945,N_8631,N_8636);
nor U8946 (N_8946,N_8654,N_8622);
nor U8947 (N_8947,N_8701,N_8762);
or U8948 (N_8948,N_8709,N_8758);
and U8949 (N_8949,N_8652,N_8659);
or U8950 (N_8950,N_8691,N_8642);
xnor U8951 (N_8951,N_8705,N_8654);
xor U8952 (N_8952,N_8735,N_8656);
nand U8953 (N_8953,N_8764,N_8778);
or U8954 (N_8954,N_8750,N_8638);
nor U8955 (N_8955,N_8799,N_8743);
or U8956 (N_8956,N_8652,N_8721);
xnor U8957 (N_8957,N_8738,N_8732);
xor U8958 (N_8958,N_8648,N_8643);
and U8959 (N_8959,N_8751,N_8726);
nor U8960 (N_8960,N_8692,N_8687);
and U8961 (N_8961,N_8675,N_8741);
nand U8962 (N_8962,N_8607,N_8708);
nand U8963 (N_8963,N_8705,N_8718);
and U8964 (N_8964,N_8763,N_8622);
or U8965 (N_8965,N_8770,N_8795);
nor U8966 (N_8966,N_8713,N_8644);
and U8967 (N_8967,N_8606,N_8744);
and U8968 (N_8968,N_8770,N_8701);
xor U8969 (N_8969,N_8623,N_8720);
or U8970 (N_8970,N_8783,N_8722);
and U8971 (N_8971,N_8636,N_8763);
or U8972 (N_8972,N_8659,N_8717);
and U8973 (N_8973,N_8777,N_8683);
or U8974 (N_8974,N_8700,N_8788);
nor U8975 (N_8975,N_8689,N_8685);
nand U8976 (N_8976,N_8632,N_8751);
and U8977 (N_8977,N_8743,N_8770);
nand U8978 (N_8978,N_8612,N_8701);
xnor U8979 (N_8979,N_8744,N_8650);
nor U8980 (N_8980,N_8658,N_8654);
or U8981 (N_8981,N_8629,N_8668);
xor U8982 (N_8982,N_8608,N_8676);
nand U8983 (N_8983,N_8783,N_8680);
nand U8984 (N_8984,N_8691,N_8611);
xor U8985 (N_8985,N_8737,N_8651);
or U8986 (N_8986,N_8776,N_8750);
nor U8987 (N_8987,N_8725,N_8690);
and U8988 (N_8988,N_8723,N_8761);
nor U8989 (N_8989,N_8712,N_8789);
and U8990 (N_8990,N_8683,N_8607);
and U8991 (N_8991,N_8752,N_8707);
and U8992 (N_8992,N_8704,N_8651);
xnor U8993 (N_8993,N_8744,N_8769);
nand U8994 (N_8994,N_8607,N_8704);
nand U8995 (N_8995,N_8772,N_8765);
nor U8996 (N_8996,N_8766,N_8767);
or U8997 (N_8997,N_8694,N_8778);
xor U8998 (N_8998,N_8740,N_8630);
nand U8999 (N_8999,N_8727,N_8606);
nor U9000 (N_9000,N_8809,N_8863);
xnor U9001 (N_9001,N_8896,N_8819);
and U9002 (N_9002,N_8879,N_8915);
nor U9003 (N_9003,N_8927,N_8867);
nand U9004 (N_9004,N_8839,N_8900);
nor U9005 (N_9005,N_8903,N_8843);
nor U9006 (N_9006,N_8953,N_8835);
nand U9007 (N_9007,N_8911,N_8984);
xor U9008 (N_9008,N_8945,N_8821);
nand U9009 (N_9009,N_8800,N_8929);
xor U9010 (N_9010,N_8926,N_8967);
nand U9011 (N_9011,N_8972,N_8988);
xor U9012 (N_9012,N_8996,N_8857);
xor U9013 (N_9013,N_8815,N_8957);
or U9014 (N_9014,N_8912,N_8851);
xnor U9015 (N_9015,N_8810,N_8824);
and U9016 (N_9016,N_8891,N_8985);
or U9017 (N_9017,N_8860,N_8889);
or U9018 (N_9018,N_8875,N_8958);
xor U9019 (N_9019,N_8861,N_8812);
xor U9020 (N_9020,N_8979,N_8906);
xnor U9021 (N_9021,N_8924,N_8983);
and U9022 (N_9022,N_8943,N_8878);
or U9023 (N_9023,N_8910,N_8997);
xor U9024 (N_9024,N_8993,N_8807);
nand U9025 (N_9025,N_8873,N_8989);
and U9026 (N_9026,N_8959,N_8806);
and U9027 (N_9027,N_8990,N_8951);
nor U9028 (N_9028,N_8838,N_8874);
xnor U9029 (N_9029,N_8881,N_8830);
nor U9030 (N_9030,N_8955,N_8898);
or U9031 (N_9031,N_8836,N_8871);
xnor U9032 (N_9032,N_8828,N_8947);
xor U9033 (N_9033,N_8919,N_8901);
xnor U9034 (N_9034,N_8849,N_8992);
nand U9035 (N_9035,N_8834,N_8845);
nand U9036 (N_9036,N_8892,N_8952);
nand U9037 (N_9037,N_8963,N_8969);
or U9038 (N_9038,N_8801,N_8888);
nand U9039 (N_9039,N_8877,N_8923);
or U9040 (N_9040,N_8960,N_8935);
and U9041 (N_9041,N_8904,N_8862);
nand U9042 (N_9042,N_8976,N_8991);
nand U9043 (N_9043,N_8855,N_8921);
and U9044 (N_9044,N_8965,N_8980);
or U9045 (N_9045,N_8887,N_8859);
xor U9046 (N_9046,N_8975,N_8995);
xor U9047 (N_9047,N_8981,N_8894);
xor U9048 (N_9048,N_8814,N_8803);
nand U9049 (N_9049,N_8933,N_8864);
nand U9050 (N_9050,N_8987,N_8837);
xnor U9051 (N_9051,N_8964,N_8922);
or U9052 (N_9052,N_8826,N_8968);
nor U9053 (N_9053,N_8832,N_8928);
xor U9054 (N_9054,N_8902,N_8946);
nand U9055 (N_9055,N_8913,N_8982);
nand U9056 (N_9056,N_8872,N_8973);
or U9057 (N_9057,N_8876,N_8936);
nor U9058 (N_9058,N_8827,N_8914);
and U9059 (N_9059,N_8885,N_8941);
or U9060 (N_9060,N_8938,N_8842);
xnor U9061 (N_9061,N_8931,N_8907);
xor U9062 (N_9062,N_8848,N_8934);
xor U9063 (N_9063,N_8970,N_8818);
nand U9064 (N_9064,N_8804,N_8956);
nand U9065 (N_9065,N_8939,N_8829);
or U9066 (N_9066,N_8823,N_8944);
nand U9067 (N_9067,N_8948,N_8978);
nand U9068 (N_9068,N_8866,N_8852);
or U9069 (N_9069,N_8890,N_8940);
nand U9070 (N_9070,N_8820,N_8954);
xnor U9071 (N_9071,N_8908,N_8966);
xnor U9072 (N_9072,N_8974,N_8977);
xnor U9073 (N_9073,N_8816,N_8808);
nand U9074 (N_9074,N_8822,N_8949);
or U9075 (N_9075,N_8942,N_8999);
or U9076 (N_9076,N_8937,N_8998);
nand U9077 (N_9077,N_8895,N_8883);
nor U9078 (N_9078,N_8918,N_8884);
nand U9079 (N_9079,N_8869,N_8920);
nor U9080 (N_9080,N_8950,N_8813);
and U9081 (N_9081,N_8841,N_8805);
and U9082 (N_9082,N_8853,N_8916);
and U9083 (N_9083,N_8986,N_8870);
nor U9084 (N_9084,N_8909,N_8865);
or U9085 (N_9085,N_8854,N_8802);
and U9086 (N_9086,N_8930,N_8850);
and U9087 (N_9087,N_8844,N_8833);
and U9088 (N_9088,N_8846,N_8994);
or U9089 (N_9089,N_8925,N_8893);
or U9090 (N_9090,N_8886,N_8932);
or U9091 (N_9091,N_8962,N_8971);
and U9092 (N_9092,N_8917,N_8847);
nor U9093 (N_9093,N_8825,N_8831);
nor U9094 (N_9094,N_8961,N_8897);
nor U9095 (N_9095,N_8882,N_8899);
or U9096 (N_9096,N_8880,N_8840);
and U9097 (N_9097,N_8811,N_8868);
and U9098 (N_9098,N_8856,N_8858);
and U9099 (N_9099,N_8817,N_8905);
or U9100 (N_9100,N_8947,N_8872);
and U9101 (N_9101,N_8879,N_8903);
or U9102 (N_9102,N_8903,N_8812);
xnor U9103 (N_9103,N_8870,N_8833);
nor U9104 (N_9104,N_8930,N_8811);
and U9105 (N_9105,N_8941,N_8835);
and U9106 (N_9106,N_8977,N_8915);
nor U9107 (N_9107,N_8917,N_8859);
or U9108 (N_9108,N_8815,N_8824);
nor U9109 (N_9109,N_8819,N_8931);
xnor U9110 (N_9110,N_8913,N_8828);
or U9111 (N_9111,N_8813,N_8911);
nand U9112 (N_9112,N_8876,N_8939);
and U9113 (N_9113,N_8912,N_8891);
nor U9114 (N_9114,N_8830,N_8854);
nand U9115 (N_9115,N_8946,N_8833);
or U9116 (N_9116,N_8974,N_8842);
nor U9117 (N_9117,N_8880,N_8904);
and U9118 (N_9118,N_8981,N_8830);
or U9119 (N_9119,N_8808,N_8981);
and U9120 (N_9120,N_8926,N_8826);
nand U9121 (N_9121,N_8900,N_8999);
nor U9122 (N_9122,N_8893,N_8962);
xnor U9123 (N_9123,N_8993,N_8906);
nand U9124 (N_9124,N_8942,N_8937);
nand U9125 (N_9125,N_8862,N_8844);
and U9126 (N_9126,N_8884,N_8916);
nor U9127 (N_9127,N_8874,N_8881);
xor U9128 (N_9128,N_8883,N_8922);
or U9129 (N_9129,N_8884,N_8895);
nor U9130 (N_9130,N_8900,N_8849);
xor U9131 (N_9131,N_8883,N_8806);
or U9132 (N_9132,N_8950,N_8865);
nand U9133 (N_9133,N_8882,N_8848);
nand U9134 (N_9134,N_8939,N_8823);
and U9135 (N_9135,N_8961,N_8866);
nand U9136 (N_9136,N_8890,N_8894);
xor U9137 (N_9137,N_8890,N_8922);
nor U9138 (N_9138,N_8812,N_8809);
nand U9139 (N_9139,N_8998,N_8935);
and U9140 (N_9140,N_8870,N_8856);
xnor U9141 (N_9141,N_8941,N_8905);
nor U9142 (N_9142,N_8992,N_8980);
and U9143 (N_9143,N_8815,N_8950);
and U9144 (N_9144,N_8883,N_8838);
and U9145 (N_9145,N_8808,N_8853);
xnor U9146 (N_9146,N_8895,N_8910);
nor U9147 (N_9147,N_8874,N_8849);
or U9148 (N_9148,N_8843,N_8801);
nand U9149 (N_9149,N_8974,N_8952);
xnor U9150 (N_9150,N_8801,N_8989);
nand U9151 (N_9151,N_8902,N_8872);
or U9152 (N_9152,N_8961,N_8941);
nand U9153 (N_9153,N_8932,N_8804);
xor U9154 (N_9154,N_8823,N_8959);
nor U9155 (N_9155,N_8836,N_8977);
xor U9156 (N_9156,N_8846,N_8804);
xor U9157 (N_9157,N_8856,N_8894);
and U9158 (N_9158,N_8821,N_8856);
nand U9159 (N_9159,N_8808,N_8801);
nor U9160 (N_9160,N_8840,N_8823);
nand U9161 (N_9161,N_8889,N_8825);
nor U9162 (N_9162,N_8889,N_8911);
nand U9163 (N_9163,N_8881,N_8824);
and U9164 (N_9164,N_8883,N_8810);
or U9165 (N_9165,N_8809,N_8885);
xor U9166 (N_9166,N_8845,N_8944);
and U9167 (N_9167,N_8904,N_8853);
or U9168 (N_9168,N_8978,N_8833);
nor U9169 (N_9169,N_8838,N_8900);
and U9170 (N_9170,N_8968,N_8864);
xnor U9171 (N_9171,N_8992,N_8857);
xor U9172 (N_9172,N_8948,N_8985);
xnor U9173 (N_9173,N_8850,N_8805);
nor U9174 (N_9174,N_8914,N_8870);
nor U9175 (N_9175,N_8991,N_8881);
xnor U9176 (N_9176,N_8836,N_8852);
nor U9177 (N_9177,N_8873,N_8825);
nor U9178 (N_9178,N_8830,N_8895);
xor U9179 (N_9179,N_8850,N_8905);
xor U9180 (N_9180,N_8841,N_8815);
nand U9181 (N_9181,N_8998,N_8814);
xor U9182 (N_9182,N_8805,N_8955);
nand U9183 (N_9183,N_8903,N_8934);
or U9184 (N_9184,N_8889,N_8859);
nand U9185 (N_9185,N_8886,N_8979);
or U9186 (N_9186,N_8913,N_8997);
nor U9187 (N_9187,N_8917,N_8967);
nor U9188 (N_9188,N_8923,N_8999);
nand U9189 (N_9189,N_8983,N_8991);
or U9190 (N_9190,N_8928,N_8854);
and U9191 (N_9191,N_8940,N_8938);
or U9192 (N_9192,N_8894,N_8946);
nand U9193 (N_9193,N_8966,N_8910);
nor U9194 (N_9194,N_8939,N_8807);
and U9195 (N_9195,N_8862,N_8926);
nor U9196 (N_9196,N_8915,N_8927);
nand U9197 (N_9197,N_8992,N_8871);
xnor U9198 (N_9198,N_8963,N_8927);
nand U9199 (N_9199,N_8984,N_8986);
nor U9200 (N_9200,N_9158,N_9152);
xnor U9201 (N_9201,N_9086,N_9065);
and U9202 (N_9202,N_9096,N_9002);
nand U9203 (N_9203,N_9131,N_9102);
and U9204 (N_9204,N_9042,N_9198);
or U9205 (N_9205,N_9192,N_9009);
nand U9206 (N_9206,N_9024,N_9100);
nor U9207 (N_9207,N_9146,N_9163);
nor U9208 (N_9208,N_9187,N_9125);
nand U9209 (N_9209,N_9046,N_9080);
and U9210 (N_9210,N_9008,N_9175);
or U9211 (N_9211,N_9129,N_9144);
or U9212 (N_9212,N_9179,N_9030);
nand U9213 (N_9213,N_9185,N_9029);
and U9214 (N_9214,N_9067,N_9013);
nand U9215 (N_9215,N_9075,N_9184);
nand U9216 (N_9216,N_9106,N_9082);
or U9217 (N_9217,N_9091,N_9035);
or U9218 (N_9218,N_9006,N_9156);
and U9219 (N_9219,N_9007,N_9188);
and U9220 (N_9220,N_9182,N_9189);
and U9221 (N_9221,N_9142,N_9137);
nand U9222 (N_9222,N_9059,N_9048);
or U9223 (N_9223,N_9010,N_9181);
and U9224 (N_9224,N_9127,N_9066);
or U9225 (N_9225,N_9001,N_9000);
and U9226 (N_9226,N_9136,N_9151);
nor U9227 (N_9227,N_9094,N_9108);
or U9228 (N_9228,N_9003,N_9078);
or U9229 (N_9229,N_9055,N_9085);
nor U9230 (N_9230,N_9041,N_9018);
nor U9231 (N_9231,N_9093,N_9112);
xnor U9232 (N_9232,N_9022,N_9070);
nor U9233 (N_9233,N_9107,N_9191);
and U9234 (N_9234,N_9045,N_9026);
xnor U9235 (N_9235,N_9101,N_9178);
and U9236 (N_9236,N_9133,N_9072);
nand U9237 (N_9237,N_9060,N_9155);
nor U9238 (N_9238,N_9199,N_9088);
or U9239 (N_9239,N_9143,N_9190);
xnor U9240 (N_9240,N_9173,N_9005);
nand U9241 (N_9241,N_9183,N_9110);
nor U9242 (N_9242,N_9103,N_9165);
nor U9243 (N_9243,N_9063,N_9083);
xnor U9244 (N_9244,N_9126,N_9104);
nor U9245 (N_9245,N_9154,N_9164);
nor U9246 (N_9246,N_9031,N_9161);
or U9247 (N_9247,N_9115,N_9180);
xor U9248 (N_9248,N_9122,N_9134);
xnor U9249 (N_9249,N_9068,N_9186);
or U9250 (N_9250,N_9141,N_9105);
xnor U9251 (N_9251,N_9077,N_9135);
xnor U9252 (N_9252,N_9069,N_9027);
nand U9253 (N_9253,N_9120,N_9049);
nand U9254 (N_9254,N_9034,N_9089);
nor U9255 (N_9255,N_9123,N_9130);
nor U9256 (N_9256,N_9171,N_9021);
nand U9257 (N_9257,N_9124,N_9062);
and U9258 (N_9258,N_9015,N_9074);
and U9259 (N_9259,N_9140,N_9044);
xnor U9260 (N_9260,N_9116,N_9019);
or U9261 (N_9261,N_9043,N_9097);
xnor U9262 (N_9262,N_9177,N_9132);
and U9263 (N_9263,N_9092,N_9016);
nand U9264 (N_9264,N_9157,N_9047);
and U9265 (N_9265,N_9028,N_9017);
and U9266 (N_9266,N_9176,N_9117);
and U9267 (N_9267,N_9118,N_9172);
nand U9268 (N_9268,N_9098,N_9038);
xnor U9269 (N_9269,N_9139,N_9193);
and U9270 (N_9270,N_9169,N_9033);
and U9271 (N_9271,N_9195,N_9087);
or U9272 (N_9272,N_9051,N_9111);
or U9273 (N_9273,N_9159,N_9196);
or U9274 (N_9274,N_9081,N_9197);
and U9275 (N_9275,N_9099,N_9153);
nand U9276 (N_9276,N_9147,N_9079);
nand U9277 (N_9277,N_9052,N_9076);
xor U9278 (N_9278,N_9014,N_9054);
nand U9279 (N_9279,N_9114,N_9121);
nor U9280 (N_9280,N_9145,N_9025);
and U9281 (N_9281,N_9061,N_9050);
nor U9282 (N_9282,N_9039,N_9119);
and U9283 (N_9283,N_9064,N_9058);
and U9284 (N_9284,N_9160,N_9071);
nor U9285 (N_9285,N_9040,N_9012);
nor U9286 (N_9286,N_9194,N_9095);
or U9287 (N_9287,N_9053,N_9056);
and U9288 (N_9288,N_9128,N_9167);
nand U9289 (N_9289,N_9113,N_9020);
and U9290 (N_9290,N_9170,N_9036);
nor U9291 (N_9291,N_9032,N_9138);
xnor U9292 (N_9292,N_9037,N_9023);
nand U9293 (N_9293,N_9073,N_9168);
nor U9294 (N_9294,N_9109,N_9084);
and U9295 (N_9295,N_9148,N_9090);
xnor U9296 (N_9296,N_9150,N_9162);
nand U9297 (N_9297,N_9011,N_9166);
nor U9298 (N_9298,N_9057,N_9004);
xnor U9299 (N_9299,N_9149,N_9174);
and U9300 (N_9300,N_9117,N_9039);
nand U9301 (N_9301,N_9158,N_9113);
xnor U9302 (N_9302,N_9136,N_9027);
or U9303 (N_9303,N_9167,N_9070);
or U9304 (N_9304,N_9152,N_9034);
and U9305 (N_9305,N_9039,N_9147);
nor U9306 (N_9306,N_9031,N_9041);
or U9307 (N_9307,N_9155,N_9011);
nand U9308 (N_9308,N_9028,N_9175);
nand U9309 (N_9309,N_9177,N_9140);
or U9310 (N_9310,N_9089,N_9184);
xnor U9311 (N_9311,N_9009,N_9133);
or U9312 (N_9312,N_9008,N_9194);
and U9313 (N_9313,N_9178,N_9022);
nand U9314 (N_9314,N_9033,N_9004);
nor U9315 (N_9315,N_9041,N_9159);
and U9316 (N_9316,N_9046,N_9011);
xnor U9317 (N_9317,N_9115,N_9055);
nand U9318 (N_9318,N_9004,N_9006);
nor U9319 (N_9319,N_9030,N_9133);
nand U9320 (N_9320,N_9038,N_9076);
xor U9321 (N_9321,N_9147,N_9132);
nor U9322 (N_9322,N_9137,N_9178);
nand U9323 (N_9323,N_9039,N_9141);
or U9324 (N_9324,N_9199,N_9132);
nand U9325 (N_9325,N_9173,N_9040);
xor U9326 (N_9326,N_9120,N_9126);
nand U9327 (N_9327,N_9145,N_9108);
nor U9328 (N_9328,N_9109,N_9126);
xor U9329 (N_9329,N_9038,N_9149);
nor U9330 (N_9330,N_9089,N_9164);
xnor U9331 (N_9331,N_9061,N_9074);
xor U9332 (N_9332,N_9185,N_9105);
nor U9333 (N_9333,N_9025,N_9133);
nor U9334 (N_9334,N_9039,N_9027);
xor U9335 (N_9335,N_9163,N_9154);
nand U9336 (N_9336,N_9000,N_9149);
and U9337 (N_9337,N_9006,N_9098);
or U9338 (N_9338,N_9030,N_9155);
nor U9339 (N_9339,N_9097,N_9164);
xor U9340 (N_9340,N_9051,N_9038);
nand U9341 (N_9341,N_9010,N_9048);
nand U9342 (N_9342,N_9092,N_9181);
or U9343 (N_9343,N_9027,N_9052);
and U9344 (N_9344,N_9019,N_9059);
nand U9345 (N_9345,N_9198,N_9130);
xnor U9346 (N_9346,N_9019,N_9155);
and U9347 (N_9347,N_9166,N_9032);
xor U9348 (N_9348,N_9108,N_9063);
xnor U9349 (N_9349,N_9126,N_9188);
nor U9350 (N_9350,N_9042,N_9033);
and U9351 (N_9351,N_9018,N_9035);
and U9352 (N_9352,N_9184,N_9023);
xnor U9353 (N_9353,N_9073,N_9102);
and U9354 (N_9354,N_9061,N_9187);
and U9355 (N_9355,N_9136,N_9128);
nand U9356 (N_9356,N_9005,N_9143);
xnor U9357 (N_9357,N_9110,N_9106);
nor U9358 (N_9358,N_9158,N_9038);
nand U9359 (N_9359,N_9094,N_9074);
and U9360 (N_9360,N_9193,N_9059);
or U9361 (N_9361,N_9050,N_9055);
nand U9362 (N_9362,N_9098,N_9168);
and U9363 (N_9363,N_9127,N_9104);
or U9364 (N_9364,N_9175,N_9158);
xor U9365 (N_9365,N_9068,N_9161);
and U9366 (N_9366,N_9144,N_9029);
nor U9367 (N_9367,N_9113,N_9024);
and U9368 (N_9368,N_9058,N_9030);
nor U9369 (N_9369,N_9014,N_9053);
nand U9370 (N_9370,N_9163,N_9150);
nand U9371 (N_9371,N_9090,N_9083);
nand U9372 (N_9372,N_9022,N_9139);
or U9373 (N_9373,N_9180,N_9163);
or U9374 (N_9374,N_9192,N_9157);
nor U9375 (N_9375,N_9110,N_9199);
and U9376 (N_9376,N_9142,N_9117);
nor U9377 (N_9377,N_9072,N_9021);
nand U9378 (N_9378,N_9199,N_9085);
and U9379 (N_9379,N_9072,N_9013);
nor U9380 (N_9380,N_9141,N_9116);
or U9381 (N_9381,N_9001,N_9118);
nor U9382 (N_9382,N_9102,N_9097);
or U9383 (N_9383,N_9125,N_9165);
nand U9384 (N_9384,N_9092,N_9152);
or U9385 (N_9385,N_9176,N_9188);
xnor U9386 (N_9386,N_9105,N_9029);
and U9387 (N_9387,N_9195,N_9182);
and U9388 (N_9388,N_9020,N_9039);
and U9389 (N_9389,N_9060,N_9097);
and U9390 (N_9390,N_9074,N_9195);
nor U9391 (N_9391,N_9042,N_9060);
or U9392 (N_9392,N_9099,N_9017);
nor U9393 (N_9393,N_9123,N_9180);
xnor U9394 (N_9394,N_9093,N_9169);
and U9395 (N_9395,N_9169,N_9084);
nor U9396 (N_9396,N_9013,N_9105);
nand U9397 (N_9397,N_9026,N_9037);
nor U9398 (N_9398,N_9139,N_9129);
and U9399 (N_9399,N_9022,N_9056);
xor U9400 (N_9400,N_9386,N_9251);
or U9401 (N_9401,N_9306,N_9276);
nand U9402 (N_9402,N_9269,N_9233);
or U9403 (N_9403,N_9293,N_9289);
xor U9404 (N_9404,N_9372,N_9263);
xnor U9405 (N_9405,N_9349,N_9390);
nand U9406 (N_9406,N_9204,N_9333);
or U9407 (N_9407,N_9353,N_9341);
xor U9408 (N_9408,N_9359,N_9365);
or U9409 (N_9409,N_9312,N_9255);
nor U9410 (N_9410,N_9317,N_9313);
xor U9411 (N_9411,N_9331,N_9260);
or U9412 (N_9412,N_9361,N_9231);
or U9413 (N_9413,N_9393,N_9392);
and U9414 (N_9414,N_9277,N_9261);
and U9415 (N_9415,N_9399,N_9250);
nand U9416 (N_9416,N_9258,N_9213);
nand U9417 (N_9417,N_9253,N_9224);
or U9418 (N_9418,N_9225,N_9323);
or U9419 (N_9419,N_9278,N_9286);
or U9420 (N_9420,N_9389,N_9299);
nor U9421 (N_9421,N_9264,N_9325);
nor U9422 (N_9422,N_9248,N_9375);
nor U9423 (N_9423,N_9214,N_9234);
and U9424 (N_9424,N_9377,N_9284);
xor U9425 (N_9425,N_9266,N_9236);
nand U9426 (N_9426,N_9394,N_9387);
nand U9427 (N_9427,N_9357,N_9380);
xor U9428 (N_9428,N_9209,N_9339);
nand U9429 (N_9429,N_9208,N_9303);
nand U9430 (N_9430,N_9205,N_9379);
nor U9431 (N_9431,N_9279,N_9202);
and U9432 (N_9432,N_9291,N_9369);
or U9433 (N_9433,N_9388,N_9232);
or U9434 (N_9434,N_9322,N_9211);
or U9435 (N_9435,N_9239,N_9241);
xor U9436 (N_9436,N_9366,N_9304);
nor U9437 (N_9437,N_9355,N_9210);
or U9438 (N_9438,N_9282,N_9351);
nor U9439 (N_9439,N_9216,N_9324);
nor U9440 (N_9440,N_9391,N_9384);
xnor U9441 (N_9441,N_9310,N_9271);
or U9442 (N_9442,N_9247,N_9398);
and U9443 (N_9443,N_9226,N_9295);
and U9444 (N_9444,N_9207,N_9337);
or U9445 (N_9445,N_9320,N_9319);
nor U9446 (N_9446,N_9254,N_9382);
or U9447 (N_9447,N_9294,N_9381);
nor U9448 (N_9448,N_9274,N_9334);
xor U9449 (N_9449,N_9246,N_9281);
or U9450 (N_9450,N_9395,N_9302);
nor U9451 (N_9451,N_9376,N_9200);
or U9452 (N_9452,N_9354,N_9308);
nand U9453 (N_9453,N_9328,N_9300);
xnor U9454 (N_9454,N_9307,N_9288);
nand U9455 (N_9455,N_9373,N_9378);
or U9456 (N_9456,N_9356,N_9343);
nand U9457 (N_9457,N_9348,N_9223);
nand U9458 (N_9458,N_9275,N_9252);
xor U9459 (N_9459,N_9221,N_9259);
xnor U9460 (N_9460,N_9330,N_9243);
xnor U9461 (N_9461,N_9273,N_9314);
or U9462 (N_9462,N_9297,N_9374);
or U9463 (N_9463,N_9358,N_9336);
xnor U9464 (N_9464,N_9346,N_9270);
nor U9465 (N_9465,N_9242,N_9283);
nor U9466 (N_9466,N_9338,N_9350);
nand U9467 (N_9467,N_9218,N_9257);
nand U9468 (N_9468,N_9245,N_9332);
or U9469 (N_9469,N_9327,N_9309);
nor U9470 (N_9470,N_9383,N_9256);
nor U9471 (N_9471,N_9206,N_9342);
xnor U9472 (N_9472,N_9315,N_9230);
or U9473 (N_9473,N_9385,N_9235);
and U9474 (N_9474,N_9311,N_9268);
and U9475 (N_9475,N_9396,N_9321);
nor U9476 (N_9476,N_9280,N_9215);
or U9477 (N_9477,N_9362,N_9217);
xnor U9478 (N_9478,N_9237,N_9367);
xor U9479 (N_9479,N_9272,N_9203);
nand U9480 (N_9480,N_9287,N_9371);
or U9481 (N_9481,N_9329,N_9316);
xor U9482 (N_9482,N_9363,N_9326);
and U9483 (N_9483,N_9370,N_9267);
nand U9484 (N_9484,N_9227,N_9285);
and U9485 (N_9485,N_9229,N_9352);
nand U9486 (N_9486,N_9219,N_9222);
nand U9487 (N_9487,N_9262,N_9318);
nor U9488 (N_9488,N_9344,N_9220);
xnor U9489 (N_9489,N_9249,N_9301);
nor U9490 (N_9490,N_9340,N_9360);
xor U9491 (N_9491,N_9345,N_9240);
and U9492 (N_9492,N_9238,N_9305);
xor U9493 (N_9493,N_9298,N_9347);
nand U9494 (N_9494,N_9201,N_9212);
and U9495 (N_9495,N_9244,N_9364);
nor U9496 (N_9496,N_9265,N_9228);
and U9497 (N_9497,N_9296,N_9335);
xnor U9498 (N_9498,N_9397,N_9290);
and U9499 (N_9499,N_9368,N_9292);
or U9500 (N_9500,N_9395,N_9297);
nor U9501 (N_9501,N_9298,N_9334);
nor U9502 (N_9502,N_9297,N_9205);
and U9503 (N_9503,N_9279,N_9271);
nand U9504 (N_9504,N_9390,N_9303);
xnor U9505 (N_9505,N_9301,N_9303);
nor U9506 (N_9506,N_9260,N_9202);
nand U9507 (N_9507,N_9225,N_9333);
or U9508 (N_9508,N_9242,N_9209);
nor U9509 (N_9509,N_9305,N_9246);
nand U9510 (N_9510,N_9331,N_9294);
nor U9511 (N_9511,N_9337,N_9324);
xnor U9512 (N_9512,N_9215,N_9203);
and U9513 (N_9513,N_9325,N_9243);
nor U9514 (N_9514,N_9253,N_9214);
and U9515 (N_9515,N_9375,N_9257);
and U9516 (N_9516,N_9221,N_9267);
nor U9517 (N_9517,N_9208,N_9252);
nand U9518 (N_9518,N_9223,N_9326);
and U9519 (N_9519,N_9299,N_9385);
and U9520 (N_9520,N_9258,N_9231);
xor U9521 (N_9521,N_9247,N_9375);
and U9522 (N_9522,N_9268,N_9343);
nor U9523 (N_9523,N_9226,N_9278);
xnor U9524 (N_9524,N_9290,N_9395);
nand U9525 (N_9525,N_9384,N_9376);
nor U9526 (N_9526,N_9281,N_9215);
or U9527 (N_9527,N_9255,N_9291);
or U9528 (N_9528,N_9214,N_9341);
xor U9529 (N_9529,N_9365,N_9379);
nor U9530 (N_9530,N_9241,N_9333);
nor U9531 (N_9531,N_9332,N_9382);
and U9532 (N_9532,N_9339,N_9314);
nor U9533 (N_9533,N_9235,N_9206);
nor U9534 (N_9534,N_9387,N_9365);
or U9535 (N_9535,N_9367,N_9291);
nor U9536 (N_9536,N_9212,N_9332);
xnor U9537 (N_9537,N_9259,N_9385);
xnor U9538 (N_9538,N_9270,N_9225);
nor U9539 (N_9539,N_9327,N_9373);
and U9540 (N_9540,N_9266,N_9397);
nand U9541 (N_9541,N_9289,N_9315);
and U9542 (N_9542,N_9310,N_9222);
xor U9543 (N_9543,N_9260,N_9318);
xor U9544 (N_9544,N_9363,N_9266);
or U9545 (N_9545,N_9273,N_9310);
or U9546 (N_9546,N_9387,N_9259);
nor U9547 (N_9547,N_9259,N_9205);
nor U9548 (N_9548,N_9337,N_9375);
xnor U9549 (N_9549,N_9324,N_9252);
and U9550 (N_9550,N_9383,N_9254);
nand U9551 (N_9551,N_9313,N_9323);
xor U9552 (N_9552,N_9276,N_9314);
nand U9553 (N_9553,N_9365,N_9207);
nor U9554 (N_9554,N_9392,N_9301);
or U9555 (N_9555,N_9399,N_9311);
or U9556 (N_9556,N_9373,N_9284);
nor U9557 (N_9557,N_9289,N_9235);
nand U9558 (N_9558,N_9269,N_9377);
xor U9559 (N_9559,N_9355,N_9307);
or U9560 (N_9560,N_9341,N_9242);
or U9561 (N_9561,N_9328,N_9215);
or U9562 (N_9562,N_9237,N_9219);
nand U9563 (N_9563,N_9303,N_9331);
nand U9564 (N_9564,N_9363,N_9248);
or U9565 (N_9565,N_9364,N_9291);
nor U9566 (N_9566,N_9226,N_9398);
and U9567 (N_9567,N_9207,N_9321);
or U9568 (N_9568,N_9210,N_9224);
xnor U9569 (N_9569,N_9231,N_9201);
nor U9570 (N_9570,N_9309,N_9266);
xnor U9571 (N_9571,N_9374,N_9222);
nand U9572 (N_9572,N_9296,N_9252);
nor U9573 (N_9573,N_9217,N_9210);
nand U9574 (N_9574,N_9209,N_9358);
or U9575 (N_9575,N_9297,N_9343);
nand U9576 (N_9576,N_9206,N_9297);
or U9577 (N_9577,N_9261,N_9238);
nor U9578 (N_9578,N_9370,N_9204);
or U9579 (N_9579,N_9285,N_9376);
xor U9580 (N_9580,N_9369,N_9230);
xnor U9581 (N_9581,N_9300,N_9269);
and U9582 (N_9582,N_9263,N_9252);
or U9583 (N_9583,N_9306,N_9284);
nor U9584 (N_9584,N_9346,N_9311);
nor U9585 (N_9585,N_9293,N_9213);
or U9586 (N_9586,N_9341,N_9393);
and U9587 (N_9587,N_9287,N_9218);
and U9588 (N_9588,N_9387,N_9236);
nor U9589 (N_9589,N_9326,N_9281);
xnor U9590 (N_9590,N_9227,N_9268);
or U9591 (N_9591,N_9211,N_9304);
xor U9592 (N_9592,N_9267,N_9395);
and U9593 (N_9593,N_9355,N_9376);
or U9594 (N_9594,N_9359,N_9337);
xnor U9595 (N_9595,N_9325,N_9350);
nor U9596 (N_9596,N_9268,N_9248);
nor U9597 (N_9597,N_9275,N_9362);
xnor U9598 (N_9598,N_9399,N_9228);
and U9599 (N_9599,N_9327,N_9259);
and U9600 (N_9600,N_9405,N_9473);
nand U9601 (N_9601,N_9494,N_9551);
xor U9602 (N_9602,N_9592,N_9556);
nand U9603 (N_9603,N_9583,N_9444);
xor U9604 (N_9604,N_9442,N_9531);
nand U9605 (N_9605,N_9543,N_9560);
and U9606 (N_9606,N_9435,N_9414);
or U9607 (N_9607,N_9509,N_9506);
or U9608 (N_9608,N_9468,N_9572);
and U9609 (N_9609,N_9534,N_9581);
nor U9610 (N_9610,N_9485,N_9481);
xor U9611 (N_9611,N_9587,N_9490);
xor U9612 (N_9612,N_9523,N_9458);
and U9613 (N_9613,N_9537,N_9480);
and U9614 (N_9614,N_9507,N_9486);
or U9615 (N_9615,N_9400,N_9451);
or U9616 (N_9616,N_9597,N_9570);
and U9617 (N_9617,N_9558,N_9484);
or U9618 (N_9618,N_9546,N_9589);
xnor U9619 (N_9619,N_9411,N_9561);
nor U9620 (N_9620,N_9544,N_9429);
nor U9621 (N_9621,N_9408,N_9536);
and U9622 (N_9622,N_9584,N_9409);
nand U9623 (N_9623,N_9436,N_9498);
xnor U9624 (N_9624,N_9530,N_9413);
and U9625 (N_9625,N_9547,N_9449);
or U9626 (N_9626,N_9463,N_9475);
nor U9627 (N_9627,N_9428,N_9474);
nor U9628 (N_9628,N_9532,N_9489);
or U9629 (N_9629,N_9576,N_9564);
nand U9630 (N_9630,N_9496,N_9541);
nor U9631 (N_9631,N_9471,N_9441);
and U9632 (N_9632,N_9401,N_9455);
nor U9633 (N_9633,N_9439,N_9520);
nand U9634 (N_9634,N_9412,N_9450);
nand U9635 (N_9635,N_9482,N_9505);
xnor U9636 (N_9636,N_9548,N_9582);
or U9637 (N_9637,N_9568,N_9577);
or U9638 (N_9638,N_9513,N_9407);
xor U9639 (N_9639,N_9479,N_9448);
xor U9640 (N_9640,N_9539,N_9432);
nand U9641 (N_9641,N_9552,N_9476);
and U9642 (N_9642,N_9467,N_9553);
nand U9643 (N_9643,N_9417,N_9457);
or U9644 (N_9644,N_9565,N_9591);
xor U9645 (N_9645,N_9453,N_9477);
nor U9646 (N_9646,N_9529,N_9503);
or U9647 (N_9647,N_9422,N_9420);
and U9648 (N_9648,N_9491,N_9493);
and U9649 (N_9649,N_9497,N_9433);
xnor U9650 (N_9650,N_9542,N_9465);
and U9651 (N_9651,N_9585,N_9586);
xnor U9652 (N_9652,N_9528,N_9598);
nand U9653 (N_9653,N_9593,N_9562);
xnor U9654 (N_9654,N_9440,N_9522);
or U9655 (N_9655,N_9454,N_9424);
or U9656 (N_9656,N_9418,N_9569);
or U9657 (N_9657,N_9423,N_9447);
nor U9658 (N_9658,N_9416,N_9469);
nand U9659 (N_9659,N_9462,N_9580);
or U9660 (N_9660,N_9526,N_9404);
nand U9661 (N_9661,N_9578,N_9554);
nor U9662 (N_9662,N_9535,N_9415);
xnor U9663 (N_9663,N_9403,N_9550);
nand U9664 (N_9664,N_9430,N_9594);
and U9665 (N_9665,N_9563,N_9518);
or U9666 (N_9666,N_9406,N_9516);
and U9667 (N_9667,N_9437,N_9446);
xor U9668 (N_9668,N_9514,N_9527);
and U9669 (N_9669,N_9460,N_9567);
and U9670 (N_9670,N_9555,N_9559);
or U9671 (N_9671,N_9512,N_9574);
nand U9672 (N_9672,N_9557,N_9402);
xor U9673 (N_9673,N_9515,N_9456);
xor U9674 (N_9674,N_9501,N_9434);
nor U9675 (N_9675,N_9508,N_9464);
xor U9676 (N_9676,N_9483,N_9425);
xnor U9677 (N_9677,N_9533,N_9426);
or U9678 (N_9678,N_9410,N_9588);
or U9679 (N_9679,N_9499,N_9511);
nand U9680 (N_9680,N_9495,N_9421);
or U9681 (N_9681,N_9510,N_9461);
nand U9682 (N_9682,N_9478,N_9595);
nand U9683 (N_9683,N_9492,N_9445);
nand U9684 (N_9684,N_9452,N_9525);
xor U9685 (N_9685,N_9596,N_9549);
or U9686 (N_9686,N_9590,N_9427);
or U9687 (N_9687,N_9443,N_9487);
or U9688 (N_9688,N_9472,N_9470);
nor U9689 (N_9689,N_9573,N_9599);
nand U9690 (N_9690,N_9519,N_9504);
or U9691 (N_9691,N_9488,N_9521);
and U9692 (N_9692,N_9502,N_9545);
or U9693 (N_9693,N_9566,N_9540);
xor U9694 (N_9694,N_9431,N_9524);
and U9695 (N_9695,N_9438,N_9500);
nand U9696 (N_9696,N_9538,N_9571);
or U9697 (N_9697,N_9459,N_9419);
and U9698 (N_9698,N_9575,N_9466);
xor U9699 (N_9699,N_9579,N_9517);
or U9700 (N_9700,N_9516,N_9441);
nor U9701 (N_9701,N_9547,N_9433);
and U9702 (N_9702,N_9474,N_9465);
nand U9703 (N_9703,N_9561,N_9496);
nand U9704 (N_9704,N_9581,N_9591);
xor U9705 (N_9705,N_9403,N_9470);
xnor U9706 (N_9706,N_9536,N_9541);
or U9707 (N_9707,N_9502,N_9461);
xnor U9708 (N_9708,N_9437,N_9592);
nand U9709 (N_9709,N_9421,N_9457);
or U9710 (N_9710,N_9415,N_9499);
or U9711 (N_9711,N_9583,N_9441);
nand U9712 (N_9712,N_9528,N_9441);
nor U9713 (N_9713,N_9433,N_9536);
or U9714 (N_9714,N_9460,N_9592);
nand U9715 (N_9715,N_9459,N_9583);
nand U9716 (N_9716,N_9529,N_9587);
xnor U9717 (N_9717,N_9476,N_9413);
nand U9718 (N_9718,N_9539,N_9541);
nand U9719 (N_9719,N_9576,N_9444);
nor U9720 (N_9720,N_9569,N_9505);
nand U9721 (N_9721,N_9595,N_9508);
nor U9722 (N_9722,N_9579,N_9529);
nor U9723 (N_9723,N_9401,N_9446);
or U9724 (N_9724,N_9480,N_9574);
xor U9725 (N_9725,N_9500,N_9596);
and U9726 (N_9726,N_9425,N_9555);
nand U9727 (N_9727,N_9465,N_9583);
nor U9728 (N_9728,N_9520,N_9459);
xor U9729 (N_9729,N_9485,N_9449);
nor U9730 (N_9730,N_9532,N_9457);
or U9731 (N_9731,N_9539,N_9543);
or U9732 (N_9732,N_9496,N_9478);
or U9733 (N_9733,N_9433,N_9590);
xnor U9734 (N_9734,N_9466,N_9599);
nor U9735 (N_9735,N_9520,N_9416);
or U9736 (N_9736,N_9588,N_9475);
nand U9737 (N_9737,N_9407,N_9586);
and U9738 (N_9738,N_9448,N_9456);
nand U9739 (N_9739,N_9589,N_9473);
or U9740 (N_9740,N_9455,N_9497);
nor U9741 (N_9741,N_9469,N_9542);
or U9742 (N_9742,N_9526,N_9585);
and U9743 (N_9743,N_9432,N_9586);
nand U9744 (N_9744,N_9543,N_9460);
xnor U9745 (N_9745,N_9470,N_9552);
xnor U9746 (N_9746,N_9597,N_9439);
nor U9747 (N_9747,N_9530,N_9480);
xnor U9748 (N_9748,N_9559,N_9434);
or U9749 (N_9749,N_9547,N_9441);
or U9750 (N_9750,N_9548,N_9588);
nor U9751 (N_9751,N_9584,N_9406);
xnor U9752 (N_9752,N_9449,N_9593);
xor U9753 (N_9753,N_9544,N_9430);
xnor U9754 (N_9754,N_9555,N_9400);
nand U9755 (N_9755,N_9585,N_9554);
xnor U9756 (N_9756,N_9408,N_9527);
nand U9757 (N_9757,N_9528,N_9544);
nor U9758 (N_9758,N_9465,N_9516);
nand U9759 (N_9759,N_9561,N_9415);
xnor U9760 (N_9760,N_9585,N_9475);
and U9761 (N_9761,N_9529,N_9569);
xor U9762 (N_9762,N_9429,N_9547);
or U9763 (N_9763,N_9596,N_9571);
xnor U9764 (N_9764,N_9597,N_9411);
nand U9765 (N_9765,N_9594,N_9446);
nand U9766 (N_9766,N_9449,N_9483);
or U9767 (N_9767,N_9417,N_9573);
or U9768 (N_9768,N_9442,N_9552);
nor U9769 (N_9769,N_9448,N_9485);
nand U9770 (N_9770,N_9494,N_9536);
and U9771 (N_9771,N_9414,N_9556);
nor U9772 (N_9772,N_9437,N_9503);
nand U9773 (N_9773,N_9515,N_9475);
nand U9774 (N_9774,N_9593,N_9460);
and U9775 (N_9775,N_9522,N_9457);
or U9776 (N_9776,N_9500,N_9499);
nor U9777 (N_9777,N_9434,N_9498);
and U9778 (N_9778,N_9478,N_9548);
and U9779 (N_9779,N_9480,N_9501);
nand U9780 (N_9780,N_9416,N_9444);
nor U9781 (N_9781,N_9439,N_9516);
or U9782 (N_9782,N_9560,N_9424);
nor U9783 (N_9783,N_9498,N_9480);
xor U9784 (N_9784,N_9591,N_9404);
and U9785 (N_9785,N_9513,N_9411);
xor U9786 (N_9786,N_9556,N_9597);
or U9787 (N_9787,N_9575,N_9494);
nor U9788 (N_9788,N_9524,N_9479);
xor U9789 (N_9789,N_9436,N_9482);
nand U9790 (N_9790,N_9495,N_9493);
xor U9791 (N_9791,N_9570,N_9578);
or U9792 (N_9792,N_9446,N_9509);
xnor U9793 (N_9793,N_9474,N_9549);
nor U9794 (N_9794,N_9424,N_9401);
and U9795 (N_9795,N_9584,N_9457);
nand U9796 (N_9796,N_9430,N_9401);
nor U9797 (N_9797,N_9423,N_9498);
nand U9798 (N_9798,N_9503,N_9585);
or U9799 (N_9799,N_9526,N_9533);
or U9800 (N_9800,N_9631,N_9780);
or U9801 (N_9801,N_9776,N_9723);
or U9802 (N_9802,N_9691,N_9601);
or U9803 (N_9803,N_9615,N_9607);
nand U9804 (N_9804,N_9630,N_9725);
nand U9805 (N_9805,N_9623,N_9644);
or U9806 (N_9806,N_9744,N_9711);
nand U9807 (N_9807,N_9665,N_9616);
nand U9808 (N_9808,N_9753,N_9778);
xnor U9809 (N_9809,N_9693,N_9710);
and U9810 (N_9810,N_9699,N_9669);
nand U9811 (N_9811,N_9657,N_9739);
nor U9812 (N_9812,N_9618,N_9673);
or U9813 (N_9813,N_9685,N_9726);
nor U9814 (N_9814,N_9654,N_9767);
nor U9815 (N_9815,N_9795,N_9611);
nand U9816 (N_9816,N_9689,N_9708);
xor U9817 (N_9817,N_9661,N_9770);
or U9818 (N_9818,N_9786,N_9676);
nor U9819 (N_9819,N_9651,N_9758);
nor U9820 (N_9820,N_9677,N_9701);
or U9821 (N_9821,N_9757,N_9694);
or U9822 (N_9822,N_9690,N_9604);
nor U9823 (N_9823,N_9696,N_9687);
or U9824 (N_9824,N_9796,N_9781);
xor U9825 (N_9825,N_9771,N_9692);
or U9826 (N_9826,N_9626,N_9737);
xor U9827 (N_9827,N_9797,N_9750);
xnor U9828 (N_9828,N_9709,N_9613);
or U9829 (N_9829,N_9731,N_9730);
nand U9830 (N_9830,N_9603,N_9674);
or U9831 (N_9831,N_9652,N_9783);
and U9832 (N_9832,N_9791,N_9612);
or U9833 (N_9833,N_9754,N_9799);
xnor U9834 (N_9834,N_9659,N_9794);
nand U9835 (N_9835,N_9798,N_9642);
or U9836 (N_9836,N_9756,N_9614);
nor U9837 (N_9837,N_9742,N_9773);
nand U9838 (N_9838,N_9628,N_9682);
or U9839 (N_9839,N_9672,N_9637);
and U9840 (N_9840,N_9627,N_9624);
xnor U9841 (N_9841,N_9784,N_9740);
nand U9842 (N_9842,N_9734,N_9622);
xnor U9843 (N_9843,N_9675,N_9720);
nor U9844 (N_9844,N_9751,N_9714);
or U9845 (N_9845,N_9688,N_9768);
nand U9846 (N_9846,N_9777,N_9732);
and U9847 (N_9847,N_9666,N_9729);
nor U9848 (N_9848,N_9741,N_9650);
or U9849 (N_9849,N_9761,N_9625);
nand U9850 (N_9850,N_9782,N_9629);
or U9851 (N_9851,N_9721,N_9608);
xor U9852 (N_9852,N_9712,N_9619);
nand U9853 (N_9853,N_9647,N_9620);
or U9854 (N_9854,N_9738,N_9635);
xnor U9855 (N_9855,N_9787,N_9755);
or U9856 (N_9856,N_9762,N_9667);
or U9857 (N_9857,N_9698,N_9736);
and U9858 (N_9858,N_9646,N_9715);
and U9859 (N_9859,N_9681,N_9785);
and U9860 (N_9860,N_9640,N_9719);
nor U9861 (N_9861,N_9705,N_9605);
or U9862 (N_9862,N_9733,N_9609);
nor U9863 (N_9863,N_9632,N_9769);
and U9864 (N_9864,N_9789,N_9790);
or U9865 (N_9865,N_9765,N_9643);
nand U9866 (N_9866,N_9718,N_9636);
nor U9867 (N_9867,N_9748,N_9716);
xnor U9868 (N_9868,N_9658,N_9764);
and U9869 (N_9869,N_9697,N_9772);
or U9870 (N_9870,N_9684,N_9722);
nand U9871 (N_9871,N_9606,N_9700);
nand U9872 (N_9872,N_9671,N_9717);
or U9873 (N_9873,N_9683,N_9713);
or U9874 (N_9874,N_9788,N_9728);
nand U9875 (N_9875,N_9679,N_9775);
xnor U9876 (N_9876,N_9686,N_9747);
nor U9877 (N_9877,N_9617,N_9746);
or U9878 (N_9878,N_9727,N_9678);
nor U9879 (N_9879,N_9707,N_9792);
and U9880 (N_9880,N_9745,N_9653);
and U9881 (N_9881,N_9664,N_9779);
and U9882 (N_9882,N_9662,N_9655);
nand U9883 (N_9883,N_9793,N_9621);
nand U9884 (N_9884,N_9638,N_9668);
and U9885 (N_9885,N_9660,N_9759);
xnor U9886 (N_9886,N_9704,N_9634);
and U9887 (N_9887,N_9760,N_9610);
nor U9888 (N_9888,N_9735,N_9633);
xnor U9889 (N_9889,N_9749,N_9600);
nand U9890 (N_9890,N_9724,N_9766);
or U9891 (N_9891,N_9763,N_9663);
or U9892 (N_9892,N_9649,N_9680);
or U9893 (N_9893,N_9702,N_9706);
nand U9894 (N_9894,N_9602,N_9656);
nand U9895 (N_9895,N_9695,N_9645);
nand U9896 (N_9896,N_9639,N_9670);
xnor U9897 (N_9897,N_9641,N_9743);
or U9898 (N_9898,N_9774,N_9648);
and U9899 (N_9899,N_9752,N_9703);
or U9900 (N_9900,N_9727,N_9706);
xnor U9901 (N_9901,N_9665,N_9762);
nor U9902 (N_9902,N_9754,N_9692);
and U9903 (N_9903,N_9711,N_9664);
nor U9904 (N_9904,N_9622,N_9760);
nand U9905 (N_9905,N_9642,N_9677);
or U9906 (N_9906,N_9638,N_9631);
nor U9907 (N_9907,N_9777,N_9666);
or U9908 (N_9908,N_9679,N_9646);
xor U9909 (N_9909,N_9756,N_9622);
or U9910 (N_9910,N_9745,N_9615);
or U9911 (N_9911,N_9668,N_9660);
or U9912 (N_9912,N_9707,N_9764);
or U9913 (N_9913,N_9628,N_9661);
nor U9914 (N_9914,N_9712,N_9662);
xor U9915 (N_9915,N_9728,N_9631);
or U9916 (N_9916,N_9783,N_9623);
nor U9917 (N_9917,N_9627,N_9796);
or U9918 (N_9918,N_9618,N_9791);
and U9919 (N_9919,N_9761,N_9727);
and U9920 (N_9920,N_9757,N_9674);
xnor U9921 (N_9921,N_9626,N_9673);
xor U9922 (N_9922,N_9772,N_9737);
nor U9923 (N_9923,N_9767,N_9684);
or U9924 (N_9924,N_9609,N_9734);
xor U9925 (N_9925,N_9641,N_9688);
and U9926 (N_9926,N_9680,N_9764);
and U9927 (N_9927,N_9709,N_9638);
xnor U9928 (N_9928,N_9639,N_9734);
xnor U9929 (N_9929,N_9685,N_9617);
nor U9930 (N_9930,N_9691,N_9730);
or U9931 (N_9931,N_9670,N_9724);
nor U9932 (N_9932,N_9751,N_9746);
nor U9933 (N_9933,N_9617,N_9634);
xor U9934 (N_9934,N_9749,N_9677);
nand U9935 (N_9935,N_9637,N_9783);
nand U9936 (N_9936,N_9677,N_9610);
nand U9937 (N_9937,N_9702,N_9742);
nor U9938 (N_9938,N_9794,N_9604);
nor U9939 (N_9939,N_9659,N_9792);
xor U9940 (N_9940,N_9748,N_9650);
or U9941 (N_9941,N_9603,N_9646);
nand U9942 (N_9942,N_9708,N_9686);
nor U9943 (N_9943,N_9713,N_9613);
xnor U9944 (N_9944,N_9645,N_9659);
or U9945 (N_9945,N_9646,N_9798);
and U9946 (N_9946,N_9781,N_9667);
nor U9947 (N_9947,N_9703,N_9795);
nand U9948 (N_9948,N_9637,N_9618);
or U9949 (N_9949,N_9700,N_9789);
or U9950 (N_9950,N_9643,N_9746);
nand U9951 (N_9951,N_9733,N_9796);
nand U9952 (N_9952,N_9659,N_9689);
or U9953 (N_9953,N_9677,N_9768);
xnor U9954 (N_9954,N_9719,N_9618);
nor U9955 (N_9955,N_9708,N_9707);
and U9956 (N_9956,N_9721,N_9772);
xnor U9957 (N_9957,N_9642,N_9710);
or U9958 (N_9958,N_9740,N_9614);
nand U9959 (N_9959,N_9753,N_9704);
or U9960 (N_9960,N_9723,N_9796);
nand U9961 (N_9961,N_9665,N_9744);
nand U9962 (N_9962,N_9607,N_9799);
nor U9963 (N_9963,N_9696,N_9668);
or U9964 (N_9964,N_9782,N_9729);
nand U9965 (N_9965,N_9603,N_9619);
nor U9966 (N_9966,N_9660,N_9622);
xor U9967 (N_9967,N_9732,N_9753);
nor U9968 (N_9968,N_9654,N_9791);
nand U9969 (N_9969,N_9695,N_9615);
xnor U9970 (N_9970,N_9681,N_9779);
xor U9971 (N_9971,N_9751,N_9734);
and U9972 (N_9972,N_9601,N_9610);
nand U9973 (N_9973,N_9719,N_9769);
xnor U9974 (N_9974,N_9606,N_9662);
and U9975 (N_9975,N_9602,N_9674);
and U9976 (N_9976,N_9684,N_9799);
and U9977 (N_9977,N_9749,N_9671);
or U9978 (N_9978,N_9670,N_9757);
nand U9979 (N_9979,N_9689,N_9651);
nor U9980 (N_9980,N_9650,N_9707);
and U9981 (N_9981,N_9747,N_9765);
nor U9982 (N_9982,N_9687,N_9765);
nand U9983 (N_9983,N_9664,N_9635);
xor U9984 (N_9984,N_9632,N_9708);
xnor U9985 (N_9985,N_9755,N_9640);
or U9986 (N_9986,N_9788,N_9689);
and U9987 (N_9987,N_9609,N_9678);
xnor U9988 (N_9988,N_9647,N_9795);
nor U9989 (N_9989,N_9712,N_9737);
nor U9990 (N_9990,N_9762,N_9747);
nand U9991 (N_9991,N_9681,N_9641);
or U9992 (N_9992,N_9721,N_9637);
nor U9993 (N_9993,N_9639,N_9773);
xnor U9994 (N_9994,N_9631,N_9620);
nand U9995 (N_9995,N_9763,N_9616);
and U9996 (N_9996,N_9703,N_9667);
nor U9997 (N_9997,N_9615,N_9692);
and U9998 (N_9998,N_9737,N_9738);
and U9999 (N_9999,N_9615,N_9663);
xnor U10000 (N_10000,N_9918,N_9895);
xor U10001 (N_10001,N_9999,N_9973);
and U10002 (N_10002,N_9938,N_9944);
or U10003 (N_10003,N_9940,N_9836);
and U10004 (N_10004,N_9972,N_9904);
nand U10005 (N_10005,N_9804,N_9923);
or U10006 (N_10006,N_9993,N_9911);
nor U10007 (N_10007,N_9849,N_9996);
or U10008 (N_10008,N_9912,N_9991);
and U10009 (N_10009,N_9974,N_9975);
and U10010 (N_10010,N_9947,N_9983);
nand U10011 (N_10011,N_9984,N_9812);
xor U10012 (N_10012,N_9942,N_9919);
nand U10013 (N_10013,N_9841,N_9946);
xor U10014 (N_10014,N_9985,N_9910);
or U10015 (N_10015,N_9879,N_9847);
nand U10016 (N_10016,N_9901,N_9851);
nor U10017 (N_10017,N_9821,N_9833);
nor U10018 (N_10018,N_9844,N_9933);
and U10019 (N_10019,N_9855,N_9891);
nand U10020 (N_10020,N_9992,N_9835);
and U10021 (N_10021,N_9979,N_9894);
nand U10022 (N_10022,N_9888,N_9810);
nand U10023 (N_10023,N_9956,N_9902);
nand U10024 (N_10024,N_9856,N_9837);
and U10025 (N_10025,N_9830,N_9969);
or U10026 (N_10026,N_9823,N_9858);
nor U10027 (N_10027,N_9866,N_9827);
and U10028 (N_10028,N_9868,N_9890);
nand U10029 (N_10029,N_9854,N_9863);
or U10030 (N_10030,N_9892,N_9882);
and U10031 (N_10031,N_9997,N_9869);
and U10032 (N_10032,N_9801,N_9929);
nand U10033 (N_10033,N_9920,N_9930);
or U10034 (N_10034,N_9907,N_9875);
nand U10035 (N_10035,N_9957,N_9839);
nand U10036 (N_10036,N_9840,N_9814);
and U10037 (N_10037,N_9934,N_9880);
or U10038 (N_10038,N_9909,N_9865);
xor U10039 (N_10039,N_9903,N_9898);
and U10040 (N_10040,N_9932,N_9885);
or U10041 (N_10041,N_9838,N_9926);
nand U10042 (N_10042,N_9873,N_9958);
xnor U10043 (N_10043,N_9915,N_9914);
nand U10044 (N_10044,N_9828,N_9951);
nand U10045 (N_10045,N_9803,N_9809);
and U10046 (N_10046,N_9978,N_9941);
xnor U10047 (N_10047,N_9845,N_9995);
and U10048 (N_10048,N_9964,N_9832);
or U10049 (N_10049,N_9883,N_9927);
nand U10050 (N_10050,N_9916,N_9913);
or U10051 (N_10051,N_9897,N_9900);
or U10052 (N_10052,N_9961,N_9952);
xor U10053 (N_10053,N_9867,N_9936);
nand U10054 (N_10054,N_9943,N_9928);
and U10055 (N_10055,N_9822,N_9989);
and U10056 (N_10056,N_9813,N_9981);
xnor U10057 (N_10057,N_9965,N_9831);
xor U10058 (N_10058,N_9807,N_9870);
and U10059 (N_10059,N_9948,N_9861);
xnor U10060 (N_10060,N_9802,N_9817);
nor U10061 (N_10061,N_9955,N_9800);
nand U10062 (N_10062,N_9889,N_9877);
nor U10063 (N_10063,N_9829,N_9860);
nand U10064 (N_10064,N_9884,N_9846);
xor U10065 (N_10065,N_9917,N_9976);
xor U10066 (N_10066,N_9815,N_9834);
nand U10067 (N_10067,N_9874,N_9811);
nor U10068 (N_10068,N_9954,N_9925);
nand U10069 (N_10069,N_9990,N_9908);
nor U10070 (N_10070,N_9994,N_9806);
nor U10071 (N_10071,N_9864,N_9986);
and U10072 (N_10072,N_9937,N_9805);
nand U10073 (N_10073,N_9843,N_9872);
nand U10074 (N_10074,N_9924,N_9967);
nand U10075 (N_10075,N_9922,N_9905);
and U10076 (N_10076,N_9887,N_9852);
xnor U10077 (N_10077,N_9881,N_9931);
nand U10078 (N_10078,N_9971,N_9853);
nor U10079 (N_10079,N_9871,N_9935);
or U10080 (N_10080,N_9859,N_9819);
nor U10081 (N_10081,N_9818,N_9826);
nor U10082 (N_10082,N_9960,N_9998);
nor U10083 (N_10083,N_9848,N_9824);
and U10084 (N_10084,N_9876,N_9862);
nand U10085 (N_10085,N_9878,N_9825);
nor U10086 (N_10086,N_9982,N_9893);
nor U10087 (N_10087,N_9963,N_9959);
xnor U10088 (N_10088,N_9977,N_9820);
and U10089 (N_10089,N_9968,N_9945);
or U10090 (N_10090,N_9970,N_9939);
nor U10091 (N_10091,N_9850,N_9950);
or U10092 (N_10092,N_9906,N_9896);
or U10093 (N_10093,N_9953,N_9857);
nor U10094 (N_10094,N_9966,N_9980);
nand U10095 (N_10095,N_9899,N_9921);
nor U10096 (N_10096,N_9987,N_9962);
or U10097 (N_10097,N_9886,N_9949);
nand U10098 (N_10098,N_9988,N_9842);
and U10099 (N_10099,N_9808,N_9816);
and U10100 (N_10100,N_9807,N_9958);
nand U10101 (N_10101,N_9952,N_9803);
nand U10102 (N_10102,N_9900,N_9891);
or U10103 (N_10103,N_9802,N_9841);
xor U10104 (N_10104,N_9805,N_9973);
or U10105 (N_10105,N_9942,N_9954);
and U10106 (N_10106,N_9967,N_9932);
xor U10107 (N_10107,N_9898,N_9966);
nand U10108 (N_10108,N_9925,N_9905);
xor U10109 (N_10109,N_9949,N_9847);
nand U10110 (N_10110,N_9868,N_9907);
nor U10111 (N_10111,N_9953,N_9882);
nor U10112 (N_10112,N_9921,N_9877);
nand U10113 (N_10113,N_9937,N_9958);
nand U10114 (N_10114,N_9806,N_9913);
xnor U10115 (N_10115,N_9958,N_9880);
xnor U10116 (N_10116,N_9947,N_9942);
nor U10117 (N_10117,N_9996,N_9986);
nand U10118 (N_10118,N_9833,N_9800);
nand U10119 (N_10119,N_9855,N_9912);
nor U10120 (N_10120,N_9858,N_9977);
nor U10121 (N_10121,N_9939,N_9991);
and U10122 (N_10122,N_9859,N_9972);
nor U10123 (N_10123,N_9836,N_9878);
xnor U10124 (N_10124,N_9968,N_9831);
or U10125 (N_10125,N_9861,N_9923);
nand U10126 (N_10126,N_9847,N_9842);
xor U10127 (N_10127,N_9856,N_9876);
nand U10128 (N_10128,N_9819,N_9908);
and U10129 (N_10129,N_9819,N_9978);
and U10130 (N_10130,N_9906,N_9956);
nor U10131 (N_10131,N_9802,N_9988);
or U10132 (N_10132,N_9872,N_9839);
or U10133 (N_10133,N_9945,N_9801);
or U10134 (N_10134,N_9948,N_9892);
or U10135 (N_10135,N_9953,N_9834);
xor U10136 (N_10136,N_9890,N_9861);
nor U10137 (N_10137,N_9835,N_9971);
and U10138 (N_10138,N_9974,N_9826);
nor U10139 (N_10139,N_9903,N_9883);
nand U10140 (N_10140,N_9912,N_9986);
or U10141 (N_10141,N_9808,N_9863);
xor U10142 (N_10142,N_9988,N_9923);
xor U10143 (N_10143,N_9922,N_9858);
nand U10144 (N_10144,N_9849,N_9883);
nand U10145 (N_10145,N_9830,N_9957);
or U10146 (N_10146,N_9932,N_9854);
nor U10147 (N_10147,N_9998,N_9844);
or U10148 (N_10148,N_9987,N_9831);
or U10149 (N_10149,N_9989,N_9852);
xor U10150 (N_10150,N_9994,N_9859);
and U10151 (N_10151,N_9952,N_9894);
nand U10152 (N_10152,N_9824,N_9928);
and U10153 (N_10153,N_9880,N_9893);
nor U10154 (N_10154,N_9957,N_9977);
or U10155 (N_10155,N_9896,N_9859);
nor U10156 (N_10156,N_9803,N_9898);
nor U10157 (N_10157,N_9927,N_9801);
nand U10158 (N_10158,N_9826,N_9929);
xnor U10159 (N_10159,N_9991,N_9900);
or U10160 (N_10160,N_9992,N_9981);
and U10161 (N_10161,N_9883,N_9934);
xnor U10162 (N_10162,N_9880,N_9913);
and U10163 (N_10163,N_9843,N_9994);
nor U10164 (N_10164,N_9817,N_9896);
xnor U10165 (N_10165,N_9832,N_9955);
nand U10166 (N_10166,N_9981,N_9824);
nand U10167 (N_10167,N_9860,N_9970);
or U10168 (N_10168,N_9874,N_9950);
xnor U10169 (N_10169,N_9868,N_9813);
or U10170 (N_10170,N_9865,N_9941);
nor U10171 (N_10171,N_9924,N_9852);
or U10172 (N_10172,N_9802,N_9924);
xnor U10173 (N_10173,N_9983,N_9846);
or U10174 (N_10174,N_9914,N_9922);
or U10175 (N_10175,N_9860,N_9901);
xnor U10176 (N_10176,N_9945,N_9810);
and U10177 (N_10177,N_9845,N_9806);
nand U10178 (N_10178,N_9898,N_9875);
xnor U10179 (N_10179,N_9896,N_9993);
nand U10180 (N_10180,N_9895,N_9884);
nor U10181 (N_10181,N_9905,N_9973);
or U10182 (N_10182,N_9901,N_9955);
nand U10183 (N_10183,N_9838,N_9993);
nand U10184 (N_10184,N_9958,N_9949);
and U10185 (N_10185,N_9821,N_9870);
nand U10186 (N_10186,N_9873,N_9995);
and U10187 (N_10187,N_9886,N_9899);
and U10188 (N_10188,N_9906,N_9975);
nor U10189 (N_10189,N_9932,N_9904);
nor U10190 (N_10190,N_9969,N_9959);
nor U10191 (N_10191,N_9816,N_9839);
xor U10192 (N_10192,N_9848,N_9816);
and U10193 (N_10193,N_9836,N_9853);
nand U10194 (N_10194,N_9952,N_9874);
nor U10195 (N_10195,N_9853,N_9802);
xor U10196 (N_10196,N_9901,N_9910);
xnor U10197 (N_10197,N_9989,N_9838);
and U10198 (N_10198,N_9863,N_9806);
or U10199 (N_10199,N_9856,N_9946);
nand U10200 (N_10200,N_10109,N_10016);
or U10201 (N_10201,N_10011,N_10147);
nand U10202 (N_10202,N_10086,N_10029);
or U10203 (N_10203,N_10184,N_10192);
nand U10204 (N_10204,N_10144,N_10189);
nor U10205 (N_10205,N_10183,N_10045);
or U10206 (N_10206,N_10176,N_10094);
and U10207 (N_10207,N_10079,N_10167);
xnor U10208 (N_10208,N_10175,N_10073);
or U10209 (N_10209,N_10025,N_10092);
and U10210 (N_10210,N_10165,N_10164);
or U10211 (N_10211,N_10170,N_10133);
and U10212 (N_10212,N_10040,N_10120);
nor U10213 (N_10213,N_10070,N_10131);
nor U10214 (N_10214,N_10121,N_10013);
or U10215 (N_10215,N_10108,N_10077);
and U10216 (N_10216,N_10148,N_10173);
or U10217 (N_10217,N_10015,N_10096);
nand U10218 (N_10218,N_10190,N_10141);
nor U10219 (N_10219,N_10138,N_10123);
or U10220 (N_10220,N_10132,N_10038);
nor U10221 (N_10221,N_10020,N_10156);
and U10222 (N_10222,N_10056,N_10052);
and U10223 (N_10223,N_10057,N_10030);
nand U10224 (N_10224,N_10129,N_10116);
or U10225 (N_10225,N_10027,N_10128);
and U10226 (N_10226,N_10012,N_10095);
or U10227 (N_10227,N_10060,N_10023);
or U10228 (N_10228,N_10160,N_10162);
and U10229 (N_10229,N_10078,N_10181);
or U10230 (N_10230,N_10054,N_10062);
xor U10231 (N_10231,N_10171,N_10082);
or U10232 (N_10232,N_10019,N_10179);
nor U10233 (N_10233,N_10169,N_10196);
or U10234 (N_10234,N_10093,N_10069);
xnor U10235 (N_10235,N_10145,N_10099);
xnor U10236 (N_10236,N_10187,N_10104);
nor U10237 (N_10237,N_10002,N_10199);
or U10238 (N_10238,N_10032,N_10140);
and U10239 (N_10239,N_10009,N_10044);
nand U10240 (N_10240,N_10061,N_10146);
or U10241 (N_10241,N_10010,N_10103);
xnor U10242 (N_10242,N_10067,N_10053);
nor U10243 (N_10243,N_10098,N_10112);
nand U10244 (N_10244,N_10126,N_10188);
and U10245 (N_10245,N_10100,N_10008);
or U10246 (N_10246,N_10193,N_10155);
or U10247 (N_10247,N_10071,N_10075);
nand U10248 (N_10248,N_10127,N_10034);
nor U10249 (N_10249,N_10174,N_10178);
nor U10250 (N_10250,N_10097,N_10042);
nor U10251 (N_10251,N_10033,N_10143);
and U10252 (N_10252,N_10024,N_10035);
xor U10253 (N_10253,N_10087,N_10134);
nor U10254 (N_10254,N_10076,N_10041);
xnor U10255 (N_10255,N_10125,N_10047);
xnor U10256 (N_10256,N_10000,N_10072);
xnor U10257 (N_10257,N_10022,N_10113);
xnor U10258 (N_10258,N_10185,N_10111);
and U10259 (N_10259,N_10177,N_10055);
xnor U10260 (N_10260,N_10115,N_10037);
or U10261 (N_10261,N_10017,N_10194);
nor U10262 (N_10262,N_10110,N_10039);
xor U10263 (N_10263,N_10084,N_10149);
and U10264 (N_10264,N_10139,N_10168);
or U10265 (N_10265,N_10163,N_10137);
nor U10266 (N_10266,N_10068,N_10136);
and U10267 (N_10267,N_10074,N_10048);
and U10268 (N_10268,N_10028,N_10036);
xnor U10269 (N_10269,N_10150,N_10021);
nor U10270 (N_10270,N_10004,N_10089);
or U10271 (N_10271,N_10153,N_10091);
or U10272 (N_10272,N_10158,N_10066);
and U10273 (N_10273,N_10063,N_10114);
or U10274 (N_10274,N_10050,N_10006);
and U10275 (N_10275,N_10101,N_10159);
xor U10276 (N_10276,N_10014,N_10026);
nor U10277 (N_10277,N_10001,N_10106);
nor U10278 (N_10278,N_10180,N_10197);
xnor U10279 (N_10279,N_10105,N_10080);
xnor U10280 (N_10280,N_10058,N_10102);
nor U10281 (N_10281,N_10107,N_10065);
or U10282 (N_10282,N_10051,N_10003);
and U10283 (N_10283,N_10083,N_10088);
and U10284 (N_10284,N_10182,N_10043);
xor U10285 (N_10285,N_10090,N_10081);
xnor U10286 (N_10286,N_10142,N_10118);
xnor U10287 (N_10287,N_10161,N_10154);
nand U10288 (N_10288,N_10130,N_10085);
nand U10289 (N_10289,N_10157,N_10166);
nor U10290 (N_10290,N_10135,N_10046);
or U10291 (N_10291,N_10064,N_10195);
nor U10292 (N_10292,N_10152,N_10186);
xnor U10293 (N_10293,N_10031,N_10191);
nand U10294 (N_10294,N_10005,N_10151);
or U10295 (N_10295,N_10119,N_10007);
xor U10296 (N_10296,N_10049,N_10117);
or U10297 (N_10297,N_10059,N_10198);
and U10298 (N_10298,N_10018,N_10124);
xor U10299 (N_10299,N_10122,N_10172);
and U10300 (N_10300,N_10087,N_10027);
xnor U10301 (N_10301,N_10144,N_10104);
xnor U10302 (N_10302,N_10076,N_10094);
xnor U10303 (N_10303,N_10180,N_10181);
nand U10304 (N_10304,N_10101,N_10199);
nand U10305 (N_10305,N_10157,N_10195);
nor U10306 (N_10306,N_10002,N_10064);
nand U10307 (N_10307,N_10040,N_10157);
or U10308 (N_10308,N_10197,N_10032);
or U10309 (N_10309,N_10123,N_10110);
xor U10310 (N_10310,N_10102,N_10084);
xnor U10311 (N_10311,N_10193,N_10065);
nor U10312 (N_10312,N_10052,N_10130);
or U10313 (N_10313,N_10170,N_10006);
xnor U10314 (N_10314,N_10178,N_10128);
nand U10315 (N_10315,N_10194,N_10187);
xor U10316 (N_10316,N_10152,N_10142);
nor U10317 (N_10317,N_10152,N_10069);
xor U10318 (N_10318,N_10154,N_10081);
or U10319 (N_10319,N_10120,N_10048);
and U10320 (N_10320,N_10165,N_10139);
nor U10321 (N_10321,N_10131,N_10107);
nand U10322 (N_10322,N_10122,N_10072);
xor U10323 (N_10323,N_10087,N_10162);
nand U10324 (N_10324,N_10051,N_10187);
nor U10325 (N_10325,N_10011,N_10030);
nor U10326 (N_10326,N_10082,N_10070);
xor U10327 (N_10327,N_10190,N_10000);
xnor U10328 (N_10328,N_10095,N_10004);
nand U10329 (N_10329,N_10138,N_10083);
nor U10330 (N_10330,N_10044,N_10008);
nor U10331 (N_10331,N_10119,N_10184);
xnor U10332 (N_10332,N_10068,N_10177);
and U10333 (N_10333,N_10112,N_10186);
nor U10334 (N_10334,N_10079,N_10005);
or U10335 (N_10335,N_10102,N_10014);
nor U10336 (N_10336,N_10181,N_10029);
and U10337 (N_10337,N_10132,N_10137);
or U10338 (N_10338,N_10188,N_10017);
nand U10339 (N_10339,N_10157,N_10013);
and U10340 (N_10340,N_10145,N_10170);
nand U10341 (N_10341,N_10065,N_10137);
or U10342 (N_10342,N_10131,N_10139);
xnor U10343 (N_10343,N_10084,N_10152);
xor U10344 (N_10344,N_10121,N_10120);
xor U10345 (N_10345,N_10083,N_10041);
or U10346 (N_10346,N_10149,N_10108);
nor U10347 (N_10347,N_10113,N_10082);
or U10348 (N_10348,N_10061,N_10179);
nor U10349 (N_10349,N_10113,N_10159);
nor U10350 (N_10350,N_10137,N_10036);
xor U10351 (N_10351,N_10037,N_10190);
nor U10352 (N_10352,N_10010,N_10024);
and U10353 (N_10353,N_10148,N_10150);
and U10354 (N_10354,N_10027,N_10176);
and U10355 (N_10355,N_10143,N_10132);
nor U10356 (N_10356,N_10180,N_10063);
and U10357 (N_10357,N_10145,N_10044);
or U10358 (N_10358,N_10039,N_10087);
or U10359 (N_10359,N_10197,N_10017);
or U10360 (N_10360,N_10060,N_10150);
nor U10361 (N_10361,N_10117,N_10142);
xnor U10362 (N_10362,N_10011,N_10094);
nand U10363 (N_10363,N_10032,N_10089);
or U10364 (N_10364,N_10191,N_10081);
xnor U10365 (N_10365,N_10103,N_10078);
nand U10366 (N_10366,N_10083,N_10047);
nor U10367 (N_10367,N_10063,N_10166);
or U10368 (N_10368,N_10160,N_10106);
nand U10369 (N_10369,N_10016,N_10178);
and U10370 (N_10370,N_10048,N_10031);
and U10371 (N_10371,N_10116,N_10151);
nor U10372 (N_10372,N_10151,N_10095);
xnor U10373 (N_10373,N_10081,N_10017);
xnor U10374 (N_10374,N_10172,N_10058);
nor U10375 (N_10375,N_10013,N_10174);
nor U10376 (N_10376,N_10172,N_10188);
nand U10377 (N_10377,N_10087,N_10080);
nor U10378 (N_10378,N_10055,N_10159);
nor U10379 (N_10379,N_10056,N_10105);
or U10380 (N_10380,N_10009,N_10140);
or U10381 (N_10381,N_10026,N_10066);
nor U10382 (N_10382,N_10145,N_10151);
nand U10383 (N_10383,N_10100,N_10170);
nor U10384 (N_10384,N_10094,N_10187);
nand U10385 (N_10385,N_10159,N_10156);
xor U10386 (N_10386,N_10139,N_10092);
nor U10387 (N_10387,N_10127,N_10118);
xnor U10388 (N_10388,N_10051,N_10163);
or U10389 (N_10389,N_10049,N_10036);
nand U10390 (N_10390,N_10001,N_10020);
and U10391 (N_10391,N_10192,N_10073);
nand U10392 (N_10392,N_10042,N_10006);
nor U10393 (N_10393,N_10118,N_10198);
nand U10394 (N_10394,N_10140,N_10046);
and U10395 (N_10395,N_10137,N_10150);
nor U10396 (N_10396,N_10005,N_10086);
nand U10397 (N_10397,N_10058,N_10063);
nor U10398 (N_10398,N_10002,N_10066);
xor U10399 (N_10399,N_10125,N_10045);
nor U10400 (N_10400,N_10264,N_10351);
or U10401 (N_10401,N_10304,N_10397);
or U10402 (N_10402,N_10398,N_10288);
and U10403 (N_10403,N_10231,N_10307);
nor U10404 (N_10404,N_10202,N_10215);
and U10405 (N_10405,N_10333,N_10284);
xor U10406 (N_10406,N_10219,N_10286);
nand U10407 (N_10407,N_10381,N_10263);
and U10408 (N_10408,N_10206,N_10208);
or U10409 (N_10409,N_10212,N_10309);
xor U10410 (N_10410,N_10311,N_10220);
nand U10411 (N_10411,N_10200,N_10294);
and U10412 (N_10412,N_10383,N_10268);
nor U10413 (N_10413,N_10386,N_10385);
nor U10414 (N_10414,N_10322,N_10356);
or U10415 (N_10415,N_10342,N_10295);
nor U10416 (N_10416,N_10378,N_10271);
nor U10417 (N_10417,N_10203,N_10321);
nor U10418 (N_10418,N_10269,N_10282);
and U10419 (N_10419,N_10375,N_10319);
xor U10420 (N_10420,N_10298,N_10204);
nand U10421 (N_10421,N_10227,N_10260);
xor U10422 (N_10422,N_10313,N_10337);
nor U10423 (N_10423,N_10368,N_10306);
and U10424 (N_10424,N_10303,N_10254);
nand U10425 (N_10425,N_10275,N_10350);
and U10426 (N_10426,N_10232,N_10392);
xor U10427 (N_10427,N_10382,N_10222);
nor U10428 (N_10428,N_10218,N_10205);
nor U10429 (N_10429,N_10252,N_10315);
nand U10430 (N_10430,N_10221,N_10334);
and U10431 (N_10431,N_10259,N_10230);
or U10432 (N_10432,N_10236,N_10238);
nor U10433 (N_10433,N_10352,N_10248);
nand U10434 (N_10434,N_10363,N_10323);
or U10435 (N_10435,N_10336,N_10270);
and U10436 (N_10436,N_10296,N_10394);
and U10437 (N_10437,N_10240,N_10354);
or U10438 (N_10438,N_10244,N_10289);
or U10439 (N_10439,N_10267,N_10370);
and U10440 (N_10440,N_10285,N_10250);
and U10441 (N_10441,N_10340,N_10390);
nor U10442 (N_10442,N_10364,N_10343);
and U10443 (N_10443,N_10345,N_10330);
or U10444 (N_10444,N_10339,N_10272);
nand U10445 (N_10445,N_10224,N_10242);
or U10446 (N_10446,N_10277,N_10257);
nor U10447 (N_10447,N_10366,N_10325);
or U10448 (N_10448,N_10251,N_10210);
and U10449 (N_10449,N_10332,N_10360);
xor U10450 (N_10450,N_10256,N_10358);
and U10451 (N_10451,N_10389,N_10226);
or U10452 (N_10452,N_10258,N_10217);
nand U10453 (N_10453,N_10237,N_10367);
and U10454 (N_10454,N_10291,N_10374);
or U10455 (N_10455,N_10239,N_10276);
xnor U10456 (N_10456,N_10326,N_10201);
nor U10457 (N_10457,N_10380,N_10233);
xor U10458 (N_10458,N_10369,N_10207);
or U10459 (N_10459,N_10361,N_10261);
nand U10460 (N_10460,N_10211,N_10355);
and U10461 (N_10461,N_10249,N_10341);
nand U10462 (N_10462,N_10353,N_10225);
nand U10463 (N_10463,N_10229,N_10316);
xnor U10464 (N_10464,N_10287,N_10396);
xor U10465 (N_10465,N_10310,N_10262);
xor U10466 (N_10466,N_10302,N_10388);
nand U10467 (N_10467,N_10348,N_10349);
nand U10468 (N_10468,N_10359,N_10243);
and U10469 (N_10469,N_10328,N_10317);
nor U10470 (N_10470,N_10347,N_10223);
xnor U10471 (N_10471,N_10376,N_10253);
or U10472 (N_10472,N_10228,N_10247);
and U10473 (N_10473,N_10346,N_10235);
or U10474 (N_10474,N_10312,N_10273);
and U10475 (N_10475,N_10314,N_10216);
or U10476 (N_10476,N_10329,N_10384);
or U10477 (N_10477,N_10241,N_10283);
or U10478 (N_10478,N_10209,N_10245);
nor U10479 (N_10479,N_10335,N_10324);
xnor U10480 (N_10480,N_10214,N_10377);
or U10481 (N_10481,N_10246,N_10365);
or U10482 (N_10482,N_10387,N_10213);
xor U10483 (N_10483,N_10357,N_10293);
nand U10484 (N_10484,N_10395,N_10372);
nor U10485 (N_10485,N_10379,N_10344);
nor U10486 (N_10486,N_10299,N_10331);
nor U10487 (N_10487,N_10280,N_10255);
or U10488 (N_10488,N_10281,N_10292);
and U10489 (N_10489,N_10327,N_10297);
and U10490 (N_10490,N_10301,N_10278);
xor U10491 (N_10491,N_10320,N_10362);
and U10492 (N_10492,N_10393,N_10308);
and U10493 (N_10493,N_10338,N_10300);
and U10494 (N_10494,N_10305,N_10265);
xnor U10495 (N_10495,N_10274,N_10391);
nand U10496 (N_10496,N_10373,N_10279);
nor U10497 (N_10497,N_10371,N_10234);
nor U10498 (N_10498,N_10399,N_10266);
or U10499 (N_10499,N_10290,N_10318);
nor U10500 (N_10500,N_10359,N_10212);
or U10501 (N_10501,N_10390,N_10297);
xor U10502 (N_10502,N_10367,N_10376);
or U10503 (N_10503,N_10210,N_10286);
or U10504 (N_10504,N_10319,N_10262);
nand U10505 (N_10505,N_10228,N_10395);
and U10506 (N_10506,N_10298,N_10353);
nand U10507 (N_10507,N_10201,N_10395);
or U10508 (N_10508,N_10360,N_10349);
nor U10509 (N_10509,N_10377,N_10319);
nor U10510 (N_10510,N_10341,N_10270);
nor U10511 (N_10511,N_10309,N_10235);
or U10512 (N_10512,N_10208,N_10237);
xnor U10513 (N_10513,N_10282,N_10356);
and U10514 (N_10514,N_10364,N_10205);
nor U10515 (N_10515,N_10226,N_10244);
or U10516 (N_10516,N_10303,N_10261);
xor U10517 (N_10517,N_10368,N_10246);
or U10518 (N_10518,N_10245,N_10360);
or U10519 (N_10519,N_10210,N_10380);
nor U10520 (N_10520,N_10293,N_10319);
nor U10521 (N_10521,N_10388,N_10348);
and U10522 (N_10522,N_10260,N_10338);
and U10523 (N_10523,N_10207,N_10250);
and U10524 (N_10524,N_10368,N_10337);
or U10525 (N_10525,N_10289,N_10314);
or U10526 (N_10526,N_10341,N_10200);
nor U10527 (N_10527,N_10254,N_10214);
xor U10528 (N_10528,N_10257,N_10235);
or U10529 (N_10529,N_10207,N_10330);
xor U10530 (N_10530,N_10297,N_10343);
or U10531 (N_10531,N_10371,N_10215);
and U10532 (N_10532,N_10256,N_10296);
xor U10533 (N_10533,N_10245,N_10272);
nand U10534 (N_10534,N_10334,N_10377);
nor U10535 (N_10535,N_10214,N_10394);
nor U10536 (N_10536,N_10318,N_10249);
or U10537 (N_10537,N_10281,N_10215);
xor U10538 (N_10538,N_10380,N_10219);
and U10539 (N_10539,N_10396,N_10305);
and U10540 (N_10540,N_10231,N_10237);
nor U10541 (N_10541,N_10247,N_10399);
and U10542 (N_10542,N_10204,N_10365);
and U10543 (N_10543,N_10249,N_10353);
nor U10544 (N_10544,N_10372,N_10290);
nand U10545 (N_10545,N_10250,N_10304);
or U10546 (N_10546,N_10287,N_10205);
nor U10547 (N_10547,N_10212,N_10336);
and U10548 (N_10548,N_10204,N_10219);
or U10549 (N_10549,N_10279,N_10292);
nor U10550 (N_10550,N_10221,N_10385);
nor U10551 (N_10551,N_10374,N_10303);
and U10552 (N_10552,N_10350,N_10345);
nand U10553 (N_10553,N_10383,N_10278);
and U10554 (N_10554,N_10250,N_10237);
or U10555 (N_10555,N_10385,N_10345);
and U10556 (N_10556,N_10353,N_10259);
and U10557 (N_10557,N_10335,N_10206);
xnor U10558 (N_10558,N_10373,N_10317);
nor U10559 (N_10559,N_10253,N_10315);
nor U10560 (N_10560,N_10219,N_10393);
xor U10561 (N_10561,N_10346,N_10250);
nand U10562 (N_10562,N_10262,N_10271);
xnor U10563 (N_10563,N_10302,N_10297);
and U10564 (N_10564,N_10255,N_10213);
nand U10565 (N_10565,N_10241,N_10239);
nor U10566 (N_10566,N_10290,N_10389);
or U10567 (N_10567,N_10273,N_10302);
or U10568 (N_10568,N_10359,N_10235);
nor U10569 (N_10569,N_10251,N_10260);
nand U10570 (N_10570,N_10268,N_10353);
xor U10571 (N_10571,N_10255,N_10273);
xor U10572 (N_10572,N_10323,N_10357);
xor U10573 (N_10573,N_10359,N_10285);
or U10574 (N_10574,N_10378,N_10330);
or U10575 (N_10575,N_10223,N_10318);
and U10576 (N_10576,N_10253,N_10231);
and U10577 (N_10577,N_10337,N_10290);
nand U10578 (N_10578,N_10345,N_10299);
and U10579 (N_10579,N_10237,N_10260);
or U10580 (N_10580,N_10205,N_10393);
and U10581 (N_10581,N_10328,N_10396);
nand U10582 (N_10582,N_10206,N_10364);
and U10583 (N_10583,N_10283,N_10264);
nand U10584 (N_10584,N_10395,N_10396);
xnor U10585 (N_10585,N_10350,N_10274);
or U10586 (N_10586,N_10300,N_10394);
nor U10587 (N_10587,N_10304,N_10281);
nor U10588 (N_10588,N_10207,N_10360);
nor U10589 (N_10589,N_10208,N_10285);
and U10590 (N_10590,N_10217,N_10237);
and U10591 (N_10591,N_10265,N_10289);
or U10592 (N_10592,N_10264,N_10368);
nor U10593 (N_10593,N_10262,N_10274);
nand U10594 (N_10594,N_10200,N_10300);
nor U10595 (N_10595,N_10318,N_10316);
nor U10596 (N_10596,N_10384,N_10354);
and U10597 (N_10597,N_10304,N_10228);
xor U10598 (N_10598,N_10383,N_10382);
nand U10599 (N_10599,N_10214,N_10331);
nand U10600 (N_10600,N_10511,N_10591);
and U10601 (N_10601,N_10432,N_10472);
or U10602 (N_10602,N_10451,N_10575);
nor U10603 (N_10603,N_10436,N_10477);
xor U10604 (N_10604,N_10458,N_10530);
xnor U10605 (N_10605,N_10518,N_10596);
nand U10606 (N_10606,N_10584,N_10479);
nor U10607 (N_10607,N_10510,N_10507);
xnor U10608 (N_10608,N_10455,N_10470);
nor U10609 (N_10609,N_10486,N_10571);
and U10610 (N_10610,N_10504,N_10529);
xor U10611 (N_10611,N_10446,N_10498);
nor U10612 (N_10612,N_10496,N_10559);
or U10613 (N_10613,N_10429,N_10563);
nand U10614 (N_10614,N_10461,N_10422);
or U10615 (N_10615,N_10469,N_10505);
nor U10616 (N_10616,N_10454,N_10536);
xor U10617 (N_10617,N_10524,N_10547);
and U10618 (N_10618,N_10474,N_10439);
nand U10619 (N_10619,N_10573,N_10531);
xnor U10620 (N_10620,N_10583,N_10445);
nand U10621 (N_10621,N_10440,N_10544);
or U10622 (N_10622,N_10406,N_10585);
or U10623 (N_10623,N_10401,N_10516);
nand U10624 (N_10624,N_10599,N_10560);
or U10625 (N_10625,N_10471,N_10586);
nor U10626 (N_10626,N_10542,N_10501);
and U10627 (N_10627,N_10411,N_10499);
nor U10628 (N_10628,N_10490,N_10414);
and U10629 (N_10629,N_10582,N_10551);
nand U10630 (N_10630,N_10519,N_10562);
nand U10631 (N_10631,N_10595,N_10549);
and U10632 (N_10632,N_10447,N_10513);
and U10633 (N_10633,N_10523,N_10478);
nor U10634 (N_10634,N_10423,N_10512);
xor U10635 (N_10635,N_10443,N_10462);
and U10636 (N_10636,N_10533,N_10400);
nand U10637 (N_10637,N_10572,N_10466);
nand U10638 (N_10638,N_10550,N_10494);
nand U10639 (N_10639,N_10412,N_10548);
or U10640 (N_10640,N_10532,N_10488);
nor U10641 (N_10641,N_10558,N_10410);
or U10642 (N_10642,N_10580,N_10569);
xnor U10643 (N_10643,N_10409,N_10565);
and U10644 (N_10644,N_10438,N_10546);
and U10645 (N_10645,N_10444,N_10482);
nor U10646 (N_10646,N_10598,N_10592);
and U10647 (N_10647,N_10537,N_10484);
nand U10648 (N_10648,N_10568,N_10480);
nor U10649 (N_10649,N_10587,N_10538);
xor U10650 (N_10650,N_10473,N_10467);
or U10651 (N_10651,N_10553,N_10434);
nand U10652 (N_10652,N_10402,N_10404);
and U10653 (N_10653,N_10579,N_10424);
and U10654 (N_10654,N_10492,N_10431);
nor U10655 (N_10655,N_10577,N_10416);
nand U10656 (N_10656,N_10552,N_10527);
or U10657 (N_10657,N_10464,N_10426);
nand U10658 (N_10658,N_10500,N_10437);
or U10659 (N_10659,N_10517,N_10475);
and U10660 (N_10660,N_10557,N_10487);
and U10661 (N_10661,N_10556,N_10514);
and U10662 (N_10662,N_10468,N_10459);
nor U10663 (N_10663,N_10522,N_10453);
nand U10664 (N_10664,N_10574,N_10465);
nand U10665 (N_10665,N_10508,N_10457);
and U10666 (N_10666,N_10493,N_10497);
nand U10667 (N_10667,N_10525,N_10427);
and U10668 (N_10668,N_10418,N_10590);
xnor U10669 (N_10669,N_10421,N_10545);
and U10670 (N_10670,N_10506,N_10526);
or U10671 (N_10671,N_10589,N_10528);
xnor U10672 (N_10672,N_10450,N_10435);
xor U10673 (N_10673,N_10489,N_10415);
or U10674 (N_10674,N_10448,N_10555);
nor U10675 (N_10675,N_10534,N_10456);
or U10676 (N_10676,N_10535,N_10594);
and U10677 (N_10677,N_10520,N_10428);
or U10678 (N_10678,N_10515,N_10452);
and U10679 (N_10679,N_10491,N_10483);
xnor U10680 (N_10680,N_10463,N_10539);
nand U10681 (N_10681,N_10460,N_10564);
or U10682 (N_10682,N_10554,N_10570);
and U10683 (N_10683,N_10543,N_10597);
nor U10684 (N_10684,N_10567,N_10581);
nor U10685 (N_10685,N_10405,N_10541);
nand U10686 (N_10686,N_10593,N_10495);
and U10687 (N_10687,N_10420,N_10540);
nor U10688 (N_10688,N_10578,N_10419);
xor U10689 (N_10689,N_10481,N_10408);
nand U10690 (N_10690,N_10561,N_10430);
or U10691 (N_10691,N_10425,N_10441);
nand U10692 (N_10692,N_10566,N_10503);
and U10693 (N_10693,N_10485,N_10449);
and U10694 (N_10694,N_10588,N_10417);
or U10695 (N_10695,N_10502,N_10476);
nand U10696 (N_10696,N_10576,N_10521);
or U10697 (N_10697,N_10403,N_10407);
and U10698 (N_10698,N_10433,N_10509);
nor U10699 (N_10699,N_10413,N_10442);
and U10700 (N_10700,N_10537,N_10400);
nand U10701 (N_10701,N_10579,N_10449);
or U10702 (N_10702,N_10509,N_10568);
and U10703 (N_10703,N_10489,N_10571);
and U10704 (N_10704,N_10460,N_10431);
nor U10705 (N_10705,N_10479,N_10593);
or U10706 (N_10706,N_10405,N_10497);
and U10707 (N_10707,N_10544,N_10475);
or U10708 (N_10708,N_10585,N_10535);
nand U10709 (N_10709,N_10569,N_10572);
nor U10710 (N_10710,N_10414,N_10429);
xor U10711 (N_10711,N_10411,N_10444);
or U10712 (N_10712,N_10546,N_10418);
nor U10713 (N_10713,N_10484,N_10463);
xor U10714 (N_10714,N_10458,N_10435);
nand U10715 (N_10715,N_10530,N_10467);
or U10716 (N_10716,N_10515,N_10517);
nor U10717 (N_10717,N_10523,N_10494);
or U10718 (N_10718,N_10556,N_10493);
and U10719 (N_10719,N_10415,N_10589);
nor U10720 (N_10720,N_10572,N_10530);
xnor U10721 (N_10721,N_10535,N_10442);
nor U10722 (N_10722,N_10540,N_10447);
and U10723 (N_10723,N_10427,N_10516);
xor U10724 (N_10724,N_10459,N_10527);
and U10725 (N_10725,N_10597,N_10477);
or U10726 (N_10726,N_10503,N_10431);
and U10727 (N_10727,N_10535,N_10417);
and U10728 (N_10728,N_10428,N_10570);
xnor U10729 (N_10729,N_10475,N_10469);
or U10730 (N_10730,N_10470,N_10414);
nand U10731 (N_10731,N_10465,N_10454);
and U10732 (N_10732,N_10552,N_10488);
xor U10733 (N_10733,N_10475,N_10535);
and U10734 (N_10734,N_10499,N_10479);
and U10735 (N_10735,N_10501,N_10405);
nand U10736 (N_10736,N_10455,N_10407);
and U10737 (N_10737,N_10469,N_10433);
xor U10738 (N_10738,N_10408,N_10527);
or U10739 (N_10739,N_10414,N_10415);
and U10740 (N_10740,N_10588,N_10400);
and U10741 (N_10741,N_10400,N_10529);
or U10742 (N_10742,N_10480,N_10490);
nand U10743 (N_10743,N_10491,N_10488);
or U10744 (N_10744,N_10424,N_10476);
or U10745 (N_10745,N_10535,N_10555);
and U10746 (N_10746,N_10493,N_10459);
or U10747 (N_10747,N_10408,N_10552);
or U10748 (N_10748,N_10522,N_10574);
nor U10749 (N_10749,N_10470,N_10431);
xor U10750 (N_10750,N_10483,N_10476);
nand U10751 (N_10751,N_10445,N_10427);
xnor U10752 (N_10752,N_10471,N_10493);
nor U10753 (N_10753,N_10530,N_10421);
xor U10754 (N_10754,N_10506,N_10514);
or U10755 (N_10755,N_10598,N_10526);
nand U10756 (N_10756,N_10450,N_10468);
xor U10757 (N_10757,N_10427,N_10467);
xnor U10758 (N_10758,N_10591,N_10449);
nor U10759 (N_10759,N_10500,N_10551);
or U10760 (N_10760,N_10580,N_10471);
nor U10761 (N_10761,N_10500,N_10456);
and U10762 (N_10762,N_10594,N_10415);
nand U10763 (N_10763,N_10552,N_10479);
nor U10764 (N_10764,N_10435,N_10474);
or U10765 (N_10765,N_10542,N_10408);
nand U10766 (N_10766,N_10488,N_10468);
and U10767 (N_10767,N_10568,N_10442);
nand U10768 (N_10768,N_10578,N_10461);
or U10769 (N_10769,N_10432,N_10431);
xor U10770 (N_10770,N_10405,N_10506);
xor U10771 (N_10771,N_10492,N_10475);
xnor U10772 (N_10772,N_10424,N_10410);
xnor U10773 (N_10773,N_10573,N_10452);
xnor U10774 (N_10774,N_10584,N_10532);
and U10775 (N_10775,N_10470,N_10495);
xnor U10776 (N_10776,N_10420,N_10488);
and U10777 (N_10777,N_10447,N_10550);
or U10778 (N_10778,N_10531,N_10422);
and U10779 (N_10779,N_10590,N_10486);
or U10780 (N_10780,N_10575,N_10516);
or U10781 (N_10781,N_10556,N_10508);
or U10782 (N_10782,N_10594,N_10570);
xnor U10783 (N_10783,N_10479,N_10597);
nand U10784 (N_10784,N_10402,N_10482);
and U10785 (N_10785,N_10462,N_10546);
xor U10786 (N_10786,N_10418,N_10560);
and U10787 (N_10787,N_10413,N_10401);
xor U10788 (N_10788,N_10507,N_10433);
and U10789 (N_10789,N_10579,N_10464);
nand U10790 (N_10790,N_10471,N_10491);
or U10791 (N_10791,N_10485,N_10565);
nand U10792 (N_10792,N_10583,N_10547);
xnor U10793 (N_10793,N_10474,N_10481);
nand U10794 (N_10794,N_10483,N_10542);
and U10795 (N_10795,N_10448,N_10554);
xnor U10796 (N_10796,N_10442,N_10510);
xor U10797 (N_10797,N_10462,N_10489);
and U10798 (N_10798,N_10582,N_10509);
and U10799 (N_10799,N_10588,N_10490);
nand U10800 (N_10800,N_10762,N_10691);
nor U10801 (N_10801,N_10673,N_10778);
xor U10802 (N_10802,N_10604,N_10763);
or U10803 (N_10803,N_10771,N_10709);
or U10804 (N_10804,N_10628,N_10662);
nand U10805 (N_10805,N_10623,N_10681);
nor U10806 (N_10806,N_10768,N_10626);
or U10807 (N_10807,N_10666,N_10679);
nor U10808 (N_10808,N_10649,N_10767);
nand U10809 (N_10809,N_10731,N_10601);
nor U10810 (N_10810,N_10715,N_10622);
xor U10811 (N_10811,N_10786,N_10613);
xnor U10812 (N_10812,N_10689,N_10651);
nor U10813 (N_10813,N_10639,N_10722);
nand U10814 (N_10814,N_10738,N_10795);
or U10815 (N_10815,N_10632,N_10706);
nor U10816 (N_10816,N_10744,N_10725);
xnor U10817 (N_10817,N_10707,N_10650);
xnor U10818 (N_10818,N_10684,N_10702);
or U10819 (N_10819,N_10770,N_10774);
xor U10820 (N_10820,N_10605,N_10727);
and U10821 (N_10821,N_10741,N_10678);
nand U10822 (N_10822,N_10796,N_10616);
and U10823 (N_10823,N_10636,N_10618);
and U10824 (N_10824,N_10784,N_10794);
nor U10825 (N_10825,N_10674,N_10728);
nand U10826 (N_10826,N_10782,N_10697);
and U10827 (N_10827,N_10772,N_10756);
xor U10828 (N_10828,N_10627,N_10711);
nor U10829 (N_10829,N_10734,N_10637);
nand U10830 (N_10830,N_10638,N_10695);
and U10831 (N_10831,N_10612,N_10694);
or U10832 (N_10832,N_10781,N_10749);
nor U10833 (N_10833,N_10646,N_10757);
and U10834 (N_10834,N_10773,N_10758);
xor U10835 (N_10835,N_10670,N_10669);
xor U10836 (N_10836,N_10754,N_10745);
xor U10837 (N_10837,N_10641,N_10600);
nor U10838 (N_10838,N_10700,N_10631);
nor U10839 (N_10839,N_10610,N_10617);
nand U10840 (N_10840,N_10789,N_10640);
nor U10841 (N_10841,N_10726,N_10625);
nor U10842 (N_10842,N_10753,N_10765);
xnor U10843 (N_10843,N_10645,N_10696);
and U10844 (N_10844,N_10664,N_10693);
and U10845 (N_10845,N_10732,N_10660);
xnor U10846 (N_10846,N_10698,N_10752);
or U10847 (N_10847,N_10721,N_10634);
and U10848 (N_10848,N_10723,N_10648);
or U10849 (N_10849,N_10740,N_10717);
or U10850 (N_10850,N_10654,N_10718);
nand U10851 (N_10851,N_10611,N_10686);
xor U10852 (N_10852,N_10647,N_10736);
and U10853 (N_10853,N_10792,N_10787);
nand U10854 (N_10854,N_10663,N_10751);
xnor U10855 (N_10855,N_10710,N_10735);
or U10856 (N_10856,N_10682,N_10798);
or U10857 (N_10857,N_10785,N_10750);
xnor U10858 (N_10858,N_10683,N_10733);
or U10859 (N_10859,N_10619,N_10614);
or U10860 (N_10860,N_10661,N_10621);
nor U10861 (N_10861,N_10675,N_10688);
xor U10862 (N_10862,N_10603,N_10720);
nor U10863 (N_10863,N_10642,N_10769);
nand U10864 (N_10864,N_10667,N_10665);
and U10865 (N_10865,N_10635,N_10656);
nor U10866 (N_10866,N_10607,N_10606);
or U10867 (N_10867,N_10685,N_10704);
and U10868 (N_10868,N_10680,N_10692);
nor U10869 (N_10869,N_10668,N_10714);
nand U10870 (N_10870,N_10633,N_10747);
or U10871 (N_10871,N_10615,N_10703);
nor U10872 (N_10872,N_10701,N_10671);
nand U10873 (N_10873,N_10730,N_10797);
xnor U10874 (N_10874,N_10652,N_10659);
or U10875 (N_10875,N_10783,N_10676);
nor U10876 (N_10876,N_10620,N_10759);
xnor U10877 (N_10877,N_10629,N_10776);
or U10878 (N_10878,N_10609,N_10780);
nand U10879 (N_10879,N_10799,N_10653);
or U10880 (N_10880,N_10724,N_10624);
xnor U10881 (N_10881,N_10788,N_10761);
and U10882 (N_10882,N_10657,N_10630);
or U10883 (N_10883,N_10766,N_10705);
xor U10884 (N_10884,N_10742,N_10793);
nand U10885 (N_10885,N_10748,N_10713);
nand U10886 (N_10886,N_10643,N_10716);
nor U10887 (N_10887,N_10719,N_10602);
nor U10888 (N_10888,N_10791,N_10708);
or U10889 (N_10889,N_10690,N_10760);
nand U10890 (N_10890,N_10777,N_10655);
nand U10891 (N_10891,N_10764,N_10746);
xor U10892 (N_10892,N_10677,N_10644);
xnor U10893 (N_10893,N_10699,N_10672);
xor U10894 (N_10894,N_10775,N_10608);
or U10895 (N_10895,N_10687,N_10779);
xor U10896 (N_10896,N_10737,N_10743);
xor U10897 (N_10897,N_10755,N_10658);
nand U10898 (N_10898,N_10739,N_10712);
and U10899 (N_10899,N_10790,N_10729);
and U10900 (N_10900,N_10750,N_10796);
and U10901 (N_10901,N_10656,N_10621);
and U10902 (N_10902,N_10718,N_10662);
xor U10903 (N_10903,N_10656,N_10712);
nor U10904 (N_10904,N_10600,N_10705);
xor U10905 (N_10905,N_10760,N_10700);
and U10906 (N_10906,N_10782,N_10756);
nand U10907 (N_10907,N_10733,N_10663);
nor U10908 (N_10908,N_10710,N_10717);
and U10909 (N_10909,N_10689,N_10782);
or U10910 (N_10910,N_10703,N_10717);
nand U10911 (N_10911,N_10626,N_10688);
nor U10912 (N_10912,N_10668,N_10681);
and U10913 (N_10913,N_10753,N_10797);
xnor U10914 (N_10914,N_10776,N_10782);
and U10915 (N_10915,N_10684,N_10725);
nor U10916 (N_10916,N_10663,N_10637);
nor U10917 (N_10917,N_10788,N_10676);
nand U10918 (N_10918,N_10604,N_10722);
nor U10919 (N_10919,N_10694,N_10628);
nor U10920 (N_10920,N_10759,N_10776);
and U10921 (N_10921,N_10684,N_10745);
nor U10922 (N_10922,N_10634,N_10765);
nand U10923 (N_10923,N_10683,N_10762);
or U10924 (N_10924,N_10749,N_10626);
xor U10925 (N_10925,N_10772,N_10618);
xor U10926 (N_10926,N_10650,N_10651);
and U10927 (N_10927,N_10644,N_10797);
nand U10928 (N_10928,N_10722,N_10719);
or U10929 (N_10929,N_10714,N_10709);
and U10930 (N_10930,N_10621,N_10731);
xnor U10931 (N_10931,N_10600,N_10694);
nor U10932 (N_10932,N_10635,N_10647);
and U10933 (N_10933,N_10759,N_10762);
and U10934 (N_10934,N_10724,N_10603);
or U10935 (N_10935,N_10742,N_10620);
xor U10936 (N_10936,N_10695,N_10628);
or U10937 (N_10937,N_10623,N_10609);
and U10938 (N_10938,N_10717,N_10711);
or U10939 (N_10939,N_10725,N_10658);
and U10940 (N_10940,N_10749,N_10600);
xnor U10941 (N_10941,N_10664,N_10759);
and U10942 (N_10942,N_10782,N_10695);
or U10943 (N_10943,N_10793,N_10717);
and U10944 (N_10944,N_10634,N_10604);
nor U10945 (N_10945,N_10686,N_10625);
nor U10946 (N_10946,N_10752,N_10762);
or U10947 (N_10947,N_10642,N_10604);
xor U10948 (N_10948,N_10753,N_10609);
nor U10949 (N_10949,N_10718,N_10630);
nor U10950 (N_10950,N_10676,N_10747);
and U10951 (N_10951,N_10699,N_10639);
xnor U10952 (N_10952,N_10787,N_10630);
nand U10953 (N_10953,N_10605,N_10615);
nand U10954 (N_10954,N_10769,N_10670);
nor U10955 (N_10955,N_10723,N_10790);
nand U10956 (N_10956,N_10695,N_10657);
nor U10957 (N_10957,N_10784,N_10795);
or U10958 (N_10958,N_10601,N_10662);
nor U10959 (N_10959,N_10628,N_10798);
and U10960 (N_10960,N_10629,N_10689);
nor U10961 (N_10961,N_10737,N_10699);
or U10962 (N_10962,N_10758,N_10658);
or U10963 (N_10963,N_10654,N_10703);
and U10964 (N_10964,N_10732,N_10734);
xor U10965 (N_10965,N_10724,N_10776);
xnor U10966 (N_10966,N_10749,N_10608);
xnor U10967 (N_10967,N_10623,N_10769);
nand U10968 (N_10968,N_10694,N_10705);
or U10969 (N_10969,N_10667,N_10792);
xnor U10970 (N_10970,N_10699,N_10703);
or U10971 (N_10971,N_10739,N_10689);
and U10972 (N_10972,N_10786,N_10620);
or U10973 (N_10973,N_10797,N_10636);
or U10974 (N_10974,N_10756,N_10641);
and U10975 (N_10975,N_10659,N_10727);
xor U10976 (N_10976,N_10780,N_10733);
or U10977 (N_10977,N_10619,N_10732);
nand U10978 (N_10978,N_10729,N_10796);
nand U10979 (N_10979,N_10702,N_10677);
xnor U10980 (N_10980,N_10697,N_10662);
nor U10981 (N_10981,N_10691,N_10733);
or U10982 (N_10982,N_10761,N_10740);
xor U10983 (N_10983,N_10767,N_10773);
nor U10984 (N_10984,N_10603,N_10707);
or U10985 (N_10985,N_10648,N_10699);
nor U10986 (N_10986,N_10713,N_10607);
or U10987 (N_10987,N_10790,N_10689);
nand U10988 (N_10988,N_10661,N_10731);
or U10989 (N_10989,N_10701,N_10670);
nor U10990 (N_10990,N_10711,N_10690);
xnor U10991 (N_10991,N_10772,N_10779);
nand U10992 (N_10992,N_10705,N_10740);
nand U10993 (N_10993,N_10720,N_10731);
nand U10994 (N_10994,N_10659,N_10742);
and U10995 (N_10995,N_10702,N_10690);
nor U10996 (N_10996,N_10743,N_10759);
and U10997 (N_10997,N_10607,N_10700);
and U10998 (N_10998,N_10679,N_10789);
nor U10999 (N_10999,N_10768,N_10639);
nor U11000 (N_11000,N_10878,N_10973);
or U11001 (N_11001,N_10832,N_10987);
xnor U11002 (N_11002,N_10890,N_10808);
or U11003 (N_11003,N_10881,N_10826);
xor U11004 (N_11004,N_10993,N_10846);
xor U11005 (N_11005,N_10932,N_10933);
and U11006 (N_11006,N_10925,N_10817);
nor U11007 (N_11007,N_10838,N_10812);
or U11008 (N_11008,N_10942,N_10822);
and U11009 (N_11009,N_10874,N_10835);
nand U11010 (N_11010,N_10887,N_10888);
xnor U11011 (N_11011,N_10869,N_10810);
nand U11012 (N_11012,N_10891,N_10883);
or U11013 (N_11013,N_10940,N_10899);
nor U11014 (N_11014,N_10928,N_10913);
nor U11015 (N_11015,N_10858,N_10930);
nor U11016 (N_11016,N_10844,N_10984);
or U11017 (N_11017,N_10955,N_10959);
xnor U11018 (N_11018,N_10815,N_10964);
nor U11019 (N_11019,N_10864,N_10911);
or U11020 (N_11020,N_10947,N_10893);
nand U11021 (N_11021,N_10965,N_10985);
xnor U11022 (N_11022,N_10927,N_10840);
nor U11023 (N_11023,N_10936,N_10941);
xnor U11024 (N_11024,N_10845,N_10862);
xor U11025 (N_11025,N_10904,N_10912);
or U11026 (N_11026,N_10863,N_10847);
and U11027 (N_11027,N_10828,N_10995);
nor U11028 (N_11028,N_10829,N_10857);
nor U11029 (N_11029,N_10821,N_10915);
xor U11030 (N_11030,N_10989,N_10850);
and U11031 (N_11031,N_10879,N_10825);
and U11032 (N_11032,N_10951,N_10806);
or U11033 (N_11033,N_10923,N_10990);
nand U11034 (N_11034,N_10991,N_10978);
nand U11035 (N_11035,N_10875,N_10924);
nand U11036 (N_11036,N_10804,N_10900);
xor U11037 (N_11037,N_10931,N_10859);
nor U11038 (N_11038,N_10873,N_10895);
nor U11039 (N_11039,N_10811,N_10839);
or U11040 (N_11040,N_10914,N_10866);
xor U11041 (N_11041,N_10937,N_10999);
and U11042 (N_11042,N_10968,N_10934);
xor U11043 (N_11043,N_10938,N_10865);
xnor U11044 (N_11044,N_10919,N_10953);
nand U11045 (N_11045,N_10824,N_10848);
nand U11046 (N_11046,N_10800,N_10926);
nand U11047 (N_11047,N_10809,N_10983);
or U11048 (N_11048,N_10853,N_10819);
and U11049 (N_11049,N_10974,N_10967);
or U11050 (N_11050,N_10861,N_10842);
and U11051 (N_11051,N_10980,N_10880);
nor U11052 (N_11052,N_10929,N_10961);
nor U11053 (N_11053,N_10957,N_10872);
or U11054 (N_11054,N_10996,N_10907);
and U11055 (N_11055,N_10886,N_10909);
nand U11056 (N_11056,N_10870,N_10803);
and U11057 (N_11057,N_10867,N_10949);
xnor U11058 (N_11058,N_10813,N_10877);
nand U11059 (N_11059,N_10833,N_10966);
and U11060 (N_11060,N_10988,N_10834);
nand U11061 (N_11061,N_10948,N_10836);
nand U11062 (N_11062,N_10816,N_10854);
or U11063 (N_11063,N_10994,N_10963);
and U11064 (N_11064,N_10830,N_10897);
xnor U11065 (N_11065,N_10885,N_10820);
and U11066 (N_11066,N_10837,N_10975);
nor U11067 (N_11067,N_10910,N_10943);
nand U11068 (N_11068,N_10971,N_10969);
or U11069 (N_11069,N_10972,N_10871);
nand U11070 (N_11070,N_10843,N_10831);
nor U11071 (N_11071,N_10906,N_10868);
nor U11072 (N_11072,N_10982,N_10805);
and U11073 (N_11073,N_10855,N_10827);
xnor U11074 (N_11074,N_10976,N_10908);
nand U11075 (N_11075,N_10818,N_10902);
nor U11076 (N_11076,N_10954,N_10889);
or U11077 (N_11077,N_10807,N_10921);
xor U11078 (N_11078,N_10952,N_10841);
xor U11079 (N_11079,N_10884,N_10917);
nand U11080 (N_11080,N_10986,N_10935);
xor U11081 (N_11081,N_10998,N_10823);
and U11082 (N_11082,N_10849,N_10814);
nor U11083 (N_11083,N_10979,N_10901);
and U11084 (N_11084,N_10903,N_10916);
nor U11085 (N_11085,N_10856,N_10950);
nand U11086 (N_11086,N_10946,N_10945);
xor U11087 (N_11087,N_10922,N_10960);
xnor U11088 (N_11088,N_10801,N_10802);
nor U11089 (N_11089,N_10939,N_10956);
nor U11090 (N_11090,N_10860,N_10882);
nor U11091 (N_11091,N_10962,N_10905);
and U11092 (N_11092,N_10997,N_10894);
nor U11093 (N_11093,N_10920,N_10852);
and U11094 (N_11094,N_10944,N_10851);
or U11095 (N_11095,N_10898,N_10992);
nand U11096 (N_11096,N_10918,N_10896);
xor U11097 (N_11097,N_10970,N_10981);
nor U11098 (N_11098,N_10977,N_10958);
xnor U11099 (N_11099,N_10876,N_10892);
or U11100 (N_11100,N_10910,N_10904);
and U11101 (N_11101,N_10819,N_10823);
nor U11102 (N_11102,N_10916,N_10850);
nand U11103 (N_11103,N_10942,N_10876);
nor U11104 (N_11104,N_10914,N_10810);
xor U11105 (N_11105,N_10983,N_10968);
nor U11106 (N_11106,N_10838,N_10969);
or U11107 (N_11107,N_10849,N_10940);
nor U11108 (N_11108,N_10934,N_10908);
or U11109 (N_11109,N_10802,N_10810);
xnor U11110 (N_11110,N_10877,N_10928);
or U11111 (N_11111,N_10817,N_10918);
or U11112 (N_11112,N_10935,N_10984);
nand U11113 (N_11113,N_10984,N_10904);
nor U11114 (N_11114,N_10828,N_10855);
xnor U11115 (N_11115,N_10908,N_10930);
or U11116 (N_11116,N_10817,N_10879);
nor U11117 (N_11117,N_10901,N_10837);
nand U11118 (N_11118,N_10857,N_10812);
nor U11119 (N_11119,N_10952,N_10905);
xnor U11120 (N_11120,N_10854,N_10895);
nand U11121 (N_11121,N_10855,N_10931);
nor U11122 (N_11122,N_10947,N_10943);
and U11123 (N_11123,N_10910,N_10959);
nor U11124 (N_11124,N_10843,N_10973);
or U11125 (N_11125,N_10967,N_10845);
and U11126 (N_11126,N_10850,N_10933);
or U11127 (N_11127,N_10995,N_10936);
or U11128 (N_11128,N_10921,N_10838);
or U11129 (N_11129,N_10843,N_10896);
and U11130 (N_11130,N_10966,N_10804);
nand U11131 (N_11131,N_10947,N_10940);
nor U11132 (N_11132,N_10897,N_10962);
xor U11133 (N_11133,N_10950,N_10975);
nand U11134 (N_11134,N_10838,N_10952);
nand U11135 (N_11135,N_10992,N_10881);
nand U11136 (N_11136,N_10888,N_10899);
nor U11137 (N_11137,N_10891,N_10886);
and U11138 (N_11138,N_10818,N_10834);
or U11139 (N_11139,N_10884,N_10963);
and U11140 (N_11140,N_10934,N_10838);
nand U11141 (N_11141,N_10900,N_10910);
xor U11142 (N_11142,N_10929,N_10815);
or U11143 (N_11143,N_10838,N_10815);
or U11144 (N_11144,N_10844,N_10998);
and U11145 (N_11145,N_10856,N_10948);
nand U11146 (N_11146,N_10985,N_10934);
nor U11147 (N_11147,N_10998,N_10901);
xnor U11148 (N_11148,N_10988,N_10937);
xnor U11149 (N_11149,N_10969,N_10894);
nand U11150 (N_11150,N_10922,N_10923);
nand U11151 (N_11151,N_10933,N_10913);
or U11152 (N_11152,N_10849,N_10832);
nand U11153 (N_11153,N_10931,N_10932);
nand U11154 (N_11154,N_10829,N_10935);
nor U11155 (N_11155,N_10831,N_10963);
xor U11156 (N_11156,N_10958,N_10911);
and U11157 (N_11157,N_10957,N_10905);
nand U11158 (N_11158,N_10895,N_10812);
xnor U11159 (N_11159,N_10811,N_10889);
xor U11160 (N_11160,N_10980,N_10868);
or U11161 (N_11161,N_10958,N_10837);
nand U11162 (N_11162,N_10921,N_10945);
xnor U11163 (N_11163,N_10965,N_10890);
xnor U11164 (N_11164,N_10864,N_10933);
nor U11165 (N_11165,N_10940,N_10955);
or U11166 (N_11166,N_10955,N_10856);
nand U11167 (N_11167,N_10817,N_10928);
nor U11168 (N_11168,N_10835,N_10866);
nand U11169 (N_11169,N_10900,N_10991);
or U11170 (N_11170,N_10995,N_10992);
nor U11171 (N_11171,N_10835,N_10939);
and U11172 (N_11172,N_10862,N_10906);
and U11173 (N_11173,N_10864,N_10932);
nand U11174 (N_11174,N_10918,N_10910);
nor U11175 (N_11175,N_10863,N_10946);
xor U11176 (N_11176,N_10999,N_10983);
and U11177 (N_11177,N_10912,N_10945);
or U11178 (N_11178,N_10853,N_10804);
nor U11179 (N_11179,N_10842,N_10973);
and U11180 (N_11180,N_10948,N_10915);
or U11181 (N_11181,N_10811,N_10885);
and U11182 (N_11182,N_10879,N_10993);
and U11183 (N_11183,N_10829,N_10999);
xnor U11184 (N_11184,N_10904,N_10877);
or U11185 (N_11185,N_10825,N_10999);
or U11186 (N_11186,N_10997,N_10942);
nand U11187 (N_11187,N_10976,N_10913);
xor U11188 (N_11188,N_10865,N_10987);
xnor U11189 (N_11189,N_10971,N_10894);
and U11190 (N_11190,N_10807,N_10852);
xor U11191 (N_11191,N_10872,N_10955);
xor U11192 (N_11192,N_10864,N_10958);
and U11193 (N_11193,N_10844,N_10833);
nor U11194 (N_11194,N_10992,N_10884);
nand U11195 (N_11195,N_10848,N_10990);
nor U11196 (N_11196,N_10993,N_10962);
nor U11197 (N_11197,N_10947,N_10802);
and U11198 (N_11198,N_10978,N_10800);
xnor U11199 (N_11199,N_10885,N_10964);
nor U11200 (N_11200,N_11057,N_11159);
and U11201 (N_11201,N_11016,N_11158);
nand U11202 (N_11202,N_11181,N_11185);
xnor U11203 (N_11203,N_11108,N_11167);
nand U11204 (N_11204,N_11135,N_11093);
nand U11205 (N_11205,N_11022,N_11109);
nor U11206 (N_11206,N_11037,N_11126);
xor U11207 (N_11207,N_11089,N_11060);
nand U11208 (N_11208,N_11059,N_11171);
nor U11209 (N_11209,N_11165,N_11003);
xor U11210 (N_11210,N_11144,N_11192);
xnor U11211 (N_11211,N_11116,N_11096);
nor U11212 (N_11212,N_11005,N_11061);
and U11213 (N_11213,N_11070,N_11163);
xnor U11214 (N_11214,N_11190,N_11098);
or U11215 (N_11215,N_11161,N_11151);
nor U11216 (N_11216,N_11041,N_11048);
and U11217 (N_11217,N_11026,N_11085);
xnor U11218 (N_11218,N_11049,N_11001);
or U11219 (N_11219,N_11047,N_11145);
nor U11220 (N_11220,N_11064,N_11110);
and U11221 (N_11221,N_11076,N_11113);
xor U11222 (N_11222,N_11103,N_11011);
and U11223 (N_11223,N_11078,N_11174);
nor U11224 (N_11224,N_11067,N_11117);
or U11225 (N_11225,N_11183,N_11164);
and U11226 (N_11226,N_11191,N_11000);
and U11227 (N_11227,N_11032,N_11062);
nor U11228 (N_11228,N_11106,N_11019);
and U11229 (N_11229,N_11043,N_11054);
and U11230 (N_11230,N_11199,N_11080);
and U11231 (N_11231,N_11086,N_11141);
nor U11232 (N_11232,N_11176,N_11157);
nor U11233 (N_11233,N_11081,N_11197);
and U11234 (N_11234,N_11036,N_11087);
xnor U11235 (N_11235,N_11138,N_11025);
or U11236 (N_11236,N_11129,N_11133);
nand U11237 (N_11237,N_11046,N_11018);
xnor U11238 (N_11238,N_11173,N_11149);
or U11239 (N_11239,N_11188,N_11039);
and U11240 (N_11240,N_11187,N_11162);
xor U11241 (N_11241,N_11071,N_11132);
nor U11242 (N_11242,N_11056,N_11172);
and U11243 (N_11243,N_11083,N_11128);
xor U11244 (N_11244,N_11051,N_11123);
and U11245 (N_11245,N_11063,N_11186);
and U11246 (N_11246,N_11122,N_11134);
nand U11247 (N_11247,N_11169,N_11177);
xor U11248 (N_11248,N_11102,N_11120);
xnor U11249 (N_11249,N_11013,N_11155);
nand U11250 (N_11250,N_11075,N_11182);
xnor U11251 (N_11251,N_11124,N_11111);
nand U11252 (N_11252,N_11017,N_11184);
nor U11253 (N_11253,N_11107,N_11092);
or U11254 (N_11254,N_11139,N_11007);
nor U11255 (N_11255,N_11195,N_11058);
or U11256 (N_11256,N_11194,N_11130);
nand U11257 (N_11257,N_11112,N_11137);
and U11258 (N_11258,N_11031,N_11028);
xnor U11259 (N_11259,N_11015,N_11038);
xnor U11260 (N_11260,N_11150,N_11077);
or U11261 (N_11261,N_11027,N_11082);
or U11262 (N_11262,N_11091,N_11053);
xor U11263 (N_11263,N_11193,N_11127);
nor U11264 (N_11264,N_11146,N_11050);
or U11265 (N_11265,N_11156,N_11142);
xor U11266 (N_11266,N_11074,N_11180);
or U11267 (N_11267,N_11088,N_11079);
or U11268 (N_11268,N_11196,N_11002);
xnor U11269 (N_11269,N_11065,N_11147);
nor U11270 (N_11270,N_11040,N_11198);
and U11271 (N_11271,N_11168,N_11009);
xor U11272 (N_11272,N_11024,N_11066);
and U11273 (N_11273,N_11068,N_11189);
nand U11274 (N_11274,N_11069,N_11136);
nand U11275 (N_11275,N_11104,N_11119);
or U11276 (N_11276,N_11006,N_11125);
nor U11277 (N_11277,N_11115,N_11095);
and U11278 (N_11278,N_11148,N_11178);
nand U11279 (N_11279,N_11105,N_11045);
nand U11280 (N_11280,N_11023,N_11030);
or U11281 (N_11281,N_11084,N_11021);
and U11282 (N_11282,N_11153,N_11099);
and U11283 (N_11283,N_11175,N_11140);
and U11284 (N_11284,N_11029,N_11166);
or U11285 (N_11285,N_11143,N_11012);
or U11286 (N_11286,N_11114,N_11094);
nand U11287 (N_11287,N_11170,N_11044);
nor U11288 (N_11288,N_11118,N_11055);
xor U11289 (N_11289,N_11160,N_11034);
nor U11290 (N_11290,N_11090,N_11073);
nor U11291 (N_11291,N_11008,N_11052);
and U11292 (N_11292,N_11004,N_11152);
nand U11293 (N_11293,N_11100,N_11035);
nand U11294 (N_11294,N_11121,N_11014);
or U11295 (N_11295,N_11097,N_11072);
xnor U11296 (N_11296,N_11154,N_11010);
nor U11297 (N_11297,N_11179,N_11020);
and U11298 (N_11298,N_11042,N_11131);
nor U11299 (N_11299,N_11101,N_11033);
and U11300 (N_11300,N_11115,N_11165);
or U11301 (N_11301,N_11038,N_11073);
nand U11302 (N_11302,N_11080,N_11053);
or U11303 (N_11303,N_11049,N_11026);
nand U11304 (N_11304,N_11023,N_11050);
or U11305 (N_11305,N_11123,N_11187);
xor U11306 (N_11306,N_11069,N_11017);
xor U11307 (N_11307,N_11084,N_11199);
nor U11308 (N_11308,N_11171,N_11049);
xor U11309 (N_11309,N_11008,N_11127);
or U11310 (N_11310,N_11010,N_11166);
and U11311 (N_11311,N_11162,N_11191);
and U11312 (N_11312,N_11139,N_11197);
nor U11313 (N_11313,N_11036,N_11122);
or U11314 (N_11314,N_11046,N_11004);
and U11315 (N_11315,N_11180,N_11059);
or U11316 (N_11316,N_11194,N_11009);
nor U11317 (N_11317,N_11053,N_11128);
nand U11318 (N_11318,N_11009,N_11054);
or U11319 (N_11319,N_11142,N_11096);
nand U11320 (N_11320,N_11007,N_11164);
nor U11321 (N_11321,N_11131,N_11098);
nand U11322 (N_11322,N_11054,N_11104);
nor U11323 (N_11323,N_11139,N_11120);
nand U11324 (N_11324,N_11175,N_11078);
nand U11325 (N_11325,N_11118,N_11158);
and U11326 (N_11326,N_11173,N_11181);
xnor U11327 (N_11327,N_11156,N_11182);
and U11328 (N_11328,N_11126,N_11143);
nand U11329 (N_11329,N_11182,N_11084);
xor U11330 (N_11330,N_11043,N_11040);
nor U11331 (N_11331,N_11064,N_11157);
nand U11332 (N_11332,N_11052,N_11083);
and U11333 (N_11333,N_11132,N_11122);
nand U11334 (N_11334,N_11109,N_11088);
nor U11335 (N_11335,N_11015,N_11086);
nor U11336 (N_11336,N_11144,N_11035);
and U11337 (N_11337,N_11180,N_11184);
or U11338 (N_11338,N_11036,N_11196);
nand U11339 (N_11339,N_11004,N_11151);
nand U11340 (N_11340,N_11090,N_11166);
xnor U11341 (N_11341,N_11051,N_11031);
or U11342 (N_11342,N_11174,N_11125);
nand U11343 (N_11343,N_11088,N_11137);
nor U11344 (N_11344,N_11166,N_11092);
and U11345 (N_11345,N_11086,N_11135);
xnor U11346 (N_11346,N_11140,N_11195);
or U11347 (N_11347,N_11078,N_11145);
nor U11348 (N_11348,N_11123,N_11179);
nor U11349 (N_11349,N_11091,N_11004);
nand U11350 (N_11350,N_11135,N_11168);
or U11351 (N_11351,N_11118,N_11024);
xnor U11352 (N_11352,N_11160,N_11079);
or U11353 (N_11353,N_11098,N_11068);
or U11354 (N_11354,N_11042,N_11097);
and U11355 (N_11355,N_11102,N_11032);
nor U11356 (N_11356,N_11120,N_11090);
xnor U11357 (N_11357,N_11085,N_11112);
nand U11358 (N_11358,N_11008,N_11034);
and U11359 (N_11359,N_11056,N_11015);
xnor U11360 (N_11360,N_11021,N_11191);
or U11361 (N_11361,N_11064,N_11173);
or U11362 (N_11362,N_11178,N_11146);
and U11363 (N_11363,N_11189,N_11199);
nand U11364 (N_11364,N_11154,N_11035);
or U11365 (N_11365,N_11163,N_11076);
nor U11366 (N_11366,N_11171,N_11187);
nor U11367 (N_11367,N_11045,N_11140);
xor U11368 (N_11368,N_11144,N_11148);
or U11369 (N_11369,N_11090,N_11151);
nand U11370 (N_11370,N_11030,N_11088);
xnor U11371 (N_11371,N_11071,N_11027);
nor U11372 (N_11372,N_11036,N_11003);
or U11373 (N_11373,N_11159,N_11146);
xor U11374 (N_11374,N_11001,N_11123);
and U11375 (N_11375,N_11113,N_11170);
nor U11376 (N_11376,N_11046,N_11073);
nand U11377 (N_11377,N_11180,N_11131);
and U11378 (N_11378,N_11039,N_11058);
and U11379 (N_11379,N_11048,N_11121);
nor U11380 (N_11380,N_11192,N_11089);
and U11381 (N_11381,N_11040,N_11176);
nand U11382 (N_11382,N_11052,N_11175);
xor U11383 (N_11383,N_11178,N_11021);
nand U11384 (N_11384,N_11169,N_11172);
and U11385 (N_11385,N_11189,N_11105);
and U11386 (N_11386,N_11004,N_11020);
or U11387 (N_11387,N_11019,N_11077);
nand U11388 (N_11388,N_11153,N_11137);
or U11389 (N_11389,N_11066,N_11109);
nor U11390 (N_11390,N_11016,N_11147);
nor U11391 (N_11391,N_11171,N_11089);
and U11392 (N_11392,N_11040,N_11077);
xor U11393 (N_11393,N_11092,N_11181);
or U11394 (N_11394,N_11026,N_11198);
or U11395 (N_11395,N_11128,N_11119);
or U11396 (N_11396,N_11058,N_11109);
nand U11397 (N_11397,N_11191,N_11093);
nand U11398 (N_11398,N_11099,N_11086);
and U11399 (N_11399,N_11109,N_11070);
nor U11400 (N_11400,N_11245,N_11262);
nor U11401 (N_11401,N_11382,N_11250);
nand U11402 (N_11402,N_11213,N_11383);
and U11403 (N_11403,N_11352,N_11323);
and U11404 (N_11404,N_11210,N_11324);
nor U11405 (N_11405,N_11274,N_11248);
and U11406 (N_11406,N_11345,N_11273);
nor U11407 (N_11407,N_11295,N_11353);
and U11408 (N_11408,N_11346,N_11389);
or U11409 (N_11409,N_11219,N_11293);
and U11410 (N_11410,N_11317,N_11364);
nand U11411 (N_11411,N_11269,N_11392);
and U11412 (N_11412,N_11211,N_11270);
and U11413 (N_11413,N_11291,N_11350);
and U11414 (N_11414,N_11339,N_11377);
nor U11415 (N_11415,N_11331,N_11303);
or U11416 (N_11416,N_11257,N_11218);
and U11417 (N_11417,N_11276,N_11216);
nor U11418 (N_11418,N_11393,N_11264);
and U11419 (N_11419,N_11252,N_11385);
or U11420 (N_11420,N_11343,N_11222);
or U11421 (N_11421,N_11304,N_11285);
and U11422 (N_11422,N_11230,N_11200);
xor U11423 (N_11423,N_11326,N_11306);
nor U11424 (N_11424,N_11292,N_11333);
or U11425 (N_11425,N_11309,N_11358);
xnor U11426 (N_11426,N_11225,N_11281);
nor U11427 (N_11427,N_11277,N_11266);
nand U11428 (N_11428,N_11207,N_11267);
nor U11429 (N_11429,N_11336,N_11361);
xnor U11430 (N_11430,N_11286,N_11357);
and U11431 (N_11431,N_11391,N_11373);
xor U11432 (N_11432,N_11355,N_11302);
and U11433 (N_11433,N_11397,N_11201);
and U11434 (N_11434,N_11351,N_11314);
or U11435 (N_11435,N_11371,N_11388);
and U11436 (N_11436,N_11279,N_11372);
nor U11437 (N_11437,N_11249,N_11239);
nor U11438 (N_11438,N_11254,N_11311);
or U11439 (N_11439,N_11214,N_11294);
xor U11440 (N_11440,N_11272,N_11227);
and U11441 (N_11441,N_11212,N_11318);
xnor U11442 (N_11442,N_11356,N_11390);
nor U11443 (N_11443,N_11365,N_11289);
nand U11444 (N_11444,N_11229,N_11315);
nor U11445 (N_11445,N_11299,N_11244);
and U11446 (N_11446,N_11321,N_11246);
nor U11447 (N_11447,N_11387,N_11320);
and U11448 (N_11448,N_11235,N_11398);
nor U11449 (N_11449,N_11379,N_11241);
nor U11450 (N_11450,N_11381,N_11236);
xor U11451 (N_11451,N_11375,N_11349);
xnor U11452 (N_11452,N_11386,N_11367);
nor U11453 (N_11453,N_11283,N_11237);
nand U11454 (N_11454,N_11275,N_11362);
or U11455 (N_11455,N_11203,N_11298);
or U11456 (N_11456,N_11243,N_11327);
nor U11457 (N_11457,N_11310,N_11209);
xnor U11458 (N_11458,N_11217,N_11215);
and U11459 (N_11459,N_11278,N_11232);
xor U11460 (N_11460,N_11208,N_11226);
and U11461 (N_11461,N_11337,N_11322);
nand U11462 (N_11462,N_11259,N_11247);
or U11463 (N_11463,N_11300,N_11376);
and U11464 (N_11464,N_11338,N_11296);
and U11465 (N_11465,N_11335,N_11368);
nor U11466 (N_11466,N_11370,N_11301);
or U11467 (N_11467,N_11284,N_11265);
nand U11468 (N_11468,N_11233,N_11251);
nor U11469 (N_11469,N_11205,N_11334);
and U11470 (N_11470,N_11328,N_11255);
nor U11471 (N_11471,N_11384,N_11261);
nand U11472 (N_11472,N_11378,N_11268);
and U11473 (N_11473,N_11258,N_11342);
nor U11474 (N_11474,N_11360,N_11374);
and U11475 (N_11475,N_11260,N_11231);
xor U11476 (N_11476,N_11341,N_11271);
nor U11477 (N_11477,N_11263,N_11223);
or U11478 (N_11478,N_11308,N_11240);
and U11479 (N_11479,N_11344,N_11290);
nand U11480 (N_11480,N_11363,N_11394);
xor U11481 (N_11481,N_11202,N_11380);
and U11482 (N_11482,N_11340,N_11220);
xnor U11483 (N_11483,N_11282,N_11238);
nand U11484 (N_11484,N_11313,N_11359);
and U11485 (N_11485,N_11329,N_11297);
xnor U11486 (N_11486,N_11399,N_11288);
nor U11487 (N_11487,N_11395,N_11253);
nor U11488 (N_11488,N_11319,N_11221);
or U11489 (N_11489,N_11287,N_11234);
nand U11490 (N_11490,N_11347,N_11312);
and U11491 (N_11491,N_11228,N_11396);
nand U11492 (N_11492,N_11256,N_11224);
nand U11493 (N_11493,N_11354,N_11242);
xor U11494 (N_11494,N_11325,N_11316);
nor U11495 (N_11495,N_11280,N_11204);
or U11496 (N_11496,N_11307,N_11206);
nand U11497 (N_11497,N_11366,N_11305);
nand U11498 (N_11498,N_11332,N_11330);
nand U11499 (N_11499,N_11369,N_11348);
and U11500 (N_11500,N_11272,N_11260);
xnor U11501 (N_11501,N_11388,N_11270);
nor U11502 (N_11502,N_11399,N_11225);
nand U11503 (N_11503,N_11380,N_11368);
nor U11504 (N_11504,N_11272,N_11282);
nor U11505 (N_11505,N_11251,N_11203);
or U11506 (N_11506,N_11376,N_11358);
or U11507 (N_11507,N_11368,N_11325);
nand U11508 (N_11508,N_11387,N_11229);
nand U11509 (N_11509,N_11247,N_11361);
nor U11510 (N_11510,N_11262,N_11381);
nor U11511 (N_11511,N_11305,N_11331);
xnor U11512 (N_11512,N_11288,N_11290);
and U11513 (N_11513,N_11304,N_11324);
nand U11514 (N_11514,N_11318,N_11366);
nor U11515 (N_11515,N_11324,N_11214);
xor U11516 (N_11516,N_11365,N_11376);
nor U11517 (N_11517,N_11354,N_11248);
and U11518 (N_11518,N_11332,N_11320);
or U11519 (N_11519,N_11308,N_11336);
and U11520 (N_11520,N_11396,N_11314);
or U11521 (N_11521,N_11313,N_11325);
nand U11522 (N_11522,N_11377,N_11200);
nand U11523 (N_11523,N_11245,N_11207);
xor U11524 (N_11524,N_11249,N_11247);
or U11525 (N_11525,N_11398,N_11239);
or U11526 (N_11526,N_11280,N_11346);
xnor U11527 (N_11527,N_11311,N_11201);
xor U11528 (N_11528,N_11366,N_11205);
nor U11529 (N_11529,N_11227,N_11305);
and U11530 (N_11530,N_11377,N_11225);
xnor U11531 (N_11531,N_11250,N_11237);
or U11532 (N_11532,N_11297,N_11305);
xnor U11533 (N_11533,N_11381,N_11394);
nand U11534 (N_11534,N_11286,N_11205);
or U11535 (N_11535,N_11379,N_11355);
and U11536 (N_11536,N_11276,N_11275);
nand U11537 (N_11537,N_11360,N_11352);
and U11538 (N_11538,N_11224,N_11268);
xor U11539 (N_11539,N_11232,N_11339);
nand U11540 (N_11540,N_11287,N_11231);
nor U11541 (N_11541,N_11292,N_11237);
and U11542 (N_11542,N_11277,N_11242);
xnor U11543 (N_11543,N_11367,N_11321);
and U11544 (N_11544,N_11260,N_11258);
or U11545 (N_11545,N_11236,N_11345);
or U11546 (N_11546,N_11355,N_11350);
or U11547 (N_11547,N_11385,N_11249);
nand U11548 (N_11548,N_11300,N_11219);
nor U11549 (N_11549,N_11256,N_11316);
nor U11550 (N_11550,N_11388,N_11329);
nor U11551 (N_11551,N_11302,N_11337);
and U11552 (N_11552,N_11294,N_11324);
and U11553 (N_11553,N_11211,N_11294);
xor U11554 (N_11554,N_11370,N_11244);
and U11555 (N_11555,N_11247,N_11236);
nand U11556 (N_11556,N_11219,N_11308);
nand U11557 (N_11557,N_11295,N_11361);
nand U11558 (N_11558,N_11247,N_11337);
and U11559 (N_11559,N_11324,N_11285);
nand U11560 (N_11560,N_11362,N_11322);
and U11561 (N_11561,N_11241,N_11321);
or U11562 (N_11562,N_11337,N_11271);
nand U11563 (N_11563,N_11302,N_11267);
nand U11564 (N_11564,N_11296,N_11247);
xor U11565 (N_11565,N_11216,N_11377);
xnor U11566 (N_11566,N_11327,N_11218);
nor U11567 (N_11567,N_11244,N_11366);
nand U11568 (N_11568,N_11322,N_11304);
or U11569 (N_11569,N_11362,N_11223);
nor U11570 (N_11570,N_11279,N_11334);
and U11571 (N_11571,N_11214,N_11391);
nor U11572 (N_11572,N_11356,N_11261);
nor U11573 (N_11573,N_11227,N_11292);
and U11574 (N_11574,N_11268,N_11267);
nand U11575 (N_11575,N_11274,N_11205);
nand U11576 (N_11576,N_11314,N_11326);
nand U11577 (N_11577,N_11390,N_11351);
and U11578 (N_11578,N_11353,N_11345);
or U11579 (N_11579,N_11372,N_11258);
or U11580 (N_11580,N_11296,N_11268);
nand U11581 (N_11581,N_11387,N_11240);
xnor U11582 (N_11582,N_11279,N_11338);
nand U11583 (N_11583,N_11209,N_11268);
nor U11584 (N_11584,N_11238,N_11358);
and U11585 (N_11585,N_11256,N_11219);
nand U11586 (N_11586,N_11294,N_11302);
nand U11587 (N_11587,N_11328,N_11369);
nand U11588 (N_11588,N_11384,N_11250);
nand U11589 (N_11589,N_11302,N_11218);
and U11590 (N_11590,N_11276,N_11332);
and U11591 (N_11591,N_11359,N_11208);
or U11592 (N_11592,N_11242,N_11373);
and U11593 (N_11593,N_11205,N_11288);
and U11594 (N_11594,N_11236,N_11302);
nor U11595 (N_11595,N_11378,N_11204);
xnor U11596 (N_11596,N_11336,N_11293);
or U11597 (N_11597,N_11290,N_11260);
or U11598 (N_11598,N_11261,N_11218);
or U11599 (N_11599,N_11223,N_11374);
nand U11600 (N_11600,N_11514,N_11518);
or U11601 (N_11601,N_11563,N_11419);
nand U11602 (N_11602,N_11589,N_11431);
nand U11603 (N_11603,N_11460,N_11410);
xnor U11604 (N_11604,N_11425,N_11528);
nor U11605 (N_11605,N_11465,N_11498);
or U11606 (N_11606,N_11547,N_11501);
xnor U11607 (N_11607,N_11457,N_11594);
nor U11608 (N_11608,N_11577,N_11511);
nand U11609 (N_11609,N_11546,N_11529);
and U11610 (N_11610,N_11404,N_11500);
xnor U11611 (N_11611,N_11539,N_11573);
and U11612 (N_11612,N_11400,N_11520);
or U11613 (N_11613,N_11469,N_11434);
xor U11614 (N_11614,N_11543,N_11536);
nand U11615 (N_11615,N_11538,N_11494);
nor U11616 (N_11616,N_11452,N_11456);
and U11617 (N_11617,N_11522,N_11476);
nand U11618 (N_11618,N_11424,N_11593);
nor U11619 (N_11619,N_11565,N_11423);
nor U11620 (N_11620,N_11578,N_11559);
nor U11621 (N_11621,N_11478,N_11416);
xnor U11622 (N_11622,N_11403,N_11549);
nand U11623 (N_11623,N_11422,N_11568);
nor U11624 (N_11624,N_11463,N_11483);
nor U11625 (N_11625,N_11405,N_11412);
nand U11626 (N_11626,N_11592,N_11458);
xor U11627 (N_11627,N_11509,N_11535);
nor U11628 (N_11628,N_11557,N_11414);
xor U11629 (N_11629,N_11502,N_11558);
and U11630 (N_11630,N_11598,N_11560);
and U11631 (N_11631,N_11508,N_11562);
nor U11632 (N_11632,N_11435,N_11490);
or U11633 (N_11633,N_11507,N_11551);
or U11634 (N_11634,N_11503,N_11567);
nand U11635 (N_11635,N_11570,N_11421);
xnor U11636 (N_11636,N_11496,N_11420);
nor U11637 (N_11637,N_11597,N_11527);
nand U11638 (N_11638,N_11532,N_11556);
or U11639 (N_11639,N_11439,N_11588);
or U11640 (N_11640,N_11525,N_11438);
nand U11641 (N_11641,N_11583,N_11409);
or U11642 (N_11642,N_11542,N_11406);
nor U11643 (N_11643,N_11515,N_11459);
nand U11644 (N_11644,N_11487,N_11467);
xor U11645 (N_11645,N_11446,N_11582);
nand U11646 (N_11646,N_11519,N_11426);
nand U11647 (N_11647,N_11440,N_11545);
nor U11648 (N_11648,N_11453,N_11531);
xor U11649 (N_11649,N_11584,N_11462);
nand U11650 (N_11650,N_11552,N_11553);
xor U11651 (N_11651,N_11402,N_11561);
nor U11652 (N_11652,N_11526,N_11464);
nor U11653 (N_11653,N_11447,N_11590);
or U11654 (N_11654,N_11569,N_11571);
nor U11655 (N_11655,N_11566,N_11510);
or U11656 (N_11656,N_11541,N_11432);
and U11657 (N_11657,N_11581,N_11475);
or U11658 (N_11658,N_11479,N_11492);
or U11659 (N_11659,N_11586,N_11437);
xor U11660 (N_11660,N_11513,N_11595);
and U11661 (N_11661,N_11441,N_11599);
or U11662 (N_11662,N_11537,N_11471);
nand U11663 (N_11663,N_11473,N_11488);
nand U11664 (N_11664,N_11524,N_11504);
xnor U11665 (N_11665,N_11444,N_11407);
xnor U11666 (N_11666,N_11481,N_11443);
and U11667 (N_11667,N_11534,N_11575);
nand U11668 (N_11668,N_11485,N_11417);
and U11669 (N_11669,N_11591,N_11480);
or U11670 (N_11670,N_11466,N_11449);
nor U11671 (N_11671,N_11499,N_11516);
xor U11672 (N_11672,N_11484,N_11428);
xnor U11673 (N_11673,N_11486,N_11408);
and U11674 (N_11674,N_11596,N_11530);
and U11675 (N_11675,N_11564,N_11433);
xnor U11676 (N_11676,N_11415,N_11470);
or U11677 (N_11677,N_11482,N_11548);
or U11678 (N_11678,N_11461,N_11451);
xor U11679 (N_11679,N_11495,N_11401);
and U11680 (N_11680,N_11472,N_11512);
nor U11681 (N_11681,N_11429,N_11430);
or U11682 (N_11682,N_11411,N_11576);
nor U11683 (N_11683,N_11442,N_11544);
xor U11684 (N_11684,N_11574,N_11493);
nand U11685 (N_11685,N_11454,N_11436);
xnor U11686 (N_11686,N_11517,N_11585);
or U11687 (N_11687,N_11468,N_11491);
nand U11688 (N_11688,N_11474,N_11506);
nand U11689 (N_11689,N_11427,N_11448);
or U11690 (N_11690,N_11450,N_11540);
nand U11691 (N_11691,N_11505,N_11523);
or U11692 (N_11692,N_11554,N_11550);
nand U11693 (N_11693,N_11580,N_11445);
xor U11694 (N_11694,N_11477,N_11533);
xnor U11695 (N_11695,N_11579,N_11587);
nor U11696 (N_11696,N_11489,N_11572);
or U11697 (N_11697,N_11555,N_11413);
or U11698 (N_11698,N_11497,N_11455);
and U11699 (N_11699,N_11418,N_11521);
and U11700 (N_11700,N_11408,N_11424);
and U11701 (N_11701,N_11404,N_11418);
or U11702 (N_11702,N_11448,N_11439);
xor U11703 (N_11703,N_11435,N_11424);
nand U11704 (N_11704,N_11553,N_11591);
nand U11705 (N_11705,N_11565,N_11589);
and U11706 (N_11706,N_11538,N_11408);
xor U11707 (N_11707,N_11530,N_11584);
xnor U11708 (N_11708,N_11553,N_11459);
nor U11709 (N_11709,N_11404,N_11469);
nor U11710 (N_11710,N_11419,N_11420);
nand U11711 (N_11711,N_11583,N_11422);
nand U11712 (N_11712,N_11550,N_11570);
nand U11713 (N_11713,N_11468,N_11581);
nand U11714 (N_11714,N_11499,N_11472);
nor U11715 (N_11715,N_11550,N_11470);
nor U11716 (N_11716,N_11485,N_11553);
and U11717 (N_11717,N_11500,N_11572);
xnor U11718 (N_11718,N_11400,N_11456);
xor U11719 (N_11719,N_11561,N_11443);
nand U11720 (N_11720,N_11443,N_11510);
xor U11721 (N_11721,N_11540,N_11458);
nor U11722 (N_11722,N_11500,N_11478);
xnor U11723 (N_11723,N_11465,N_11408);
xnor U11724 (N_11724,N_11507,N_11461);
nor U11725 (N_11725,N_11495,N_11444);
and U11726 (N_11726,N_11582,N_11578);
or U11727 (N_11727,N_11566,N_11538);
and U11728 (N_11728,N_11563,N_11538);
xor U11729 (N_11729,N_11575,N_11452);
nor U11730 (N_11730,N_11433,N_11495);
or U11731 (N_11731,N_11538,N_11507);
nand U11732 (N_11732,N_11520,N_11495);
nor U11733 (N_11733,N_11532,N_11540);
xnor U11734 (N_11734,N_11444,N_11468);
nor U11735 (N_11735,N_11556,N_11597);
nor U11736 (N_11736,N_11515,N_11468);
or U11737 (N_11737,N_11525,N_11513);
and U11738 (N_11738,N_11442,N_11514);
nor U11739 (N_11739,N_11569,N_11469);
xor U11740 (N_11740,N_11478,N_11523);
and U11741 (N_11741,N_11561,N_11455);
and U11742 (N_11742,N_11528,N_11468);
nor U11743 (N_11743,N_11426,N_11524);
nor U11744 (N_11744,N_11544,N_11440);
or U11745 (N_11745,N_11545,N_11455);
or U11746 (N_11746,N_11439,N_11473);
xor U11747 (N_11747,N_11495,N_11585);
nand U11748 (N_11748,N_11498,N_11533);
nand U11749 (N_11749,N_11528,N_11489);
nor U11750 (N_11750,N_11525,N_11566);
nor U11751 (N_11751,N_11475,N_11440);
or U11752 (N_11752,N_11531,N_11569);
xor U11753 (N_11753,N_11589,N_11519);
and U11754 (N_11754,N_11480,N_11538);
nand U11755 (N_11755,N_11462,N_11519);
or U11756 (N_11756,N_11427,N_11520);
and U11757 (N_11757,N_11415,N_11468);
or U11758 (N_11758,N_11489,N_11596);
or U11759 (N_11759,N_11574,N_11486);
and U11760 (N_11760,N_11584,N_11411);
nor U11761 (N_11761,N_11405,N_11486);
and U11762 (N_11762,N_11592,N_11531);
nand U11763 (N_11763,N_11499,N_11481);
nand U11764 (N_11764,N_11444,N_11545);
and U11765 (N_11765,N_11418,N_11477);
xnor U11766 (N_11766,N_11525,N_11401);
xor U11767 (N_11767,N_11575,N_11431);
and U11768 (N_11768,N_11567,N_11484);
nor U11769 (N_11769,N_11508,N_11409);
nand U11770 (N_11770,N_11509,N_11485);
or U11771 (N_11771,N_11556,N_11541);
nand U11772 (N_11772,N_11465,N_11512);
and U11773 (N_11773,N_11474,N_11528);
and U11774 (N_11774,N_11442,N_11552);
and U11775 (N_11775,N_11590,N_11551);
nand U11776 (N_11776,N_11469,N_11573);
and U11777 (N_11777,N_11507,N_11416);
and U11778 (N_11778,N_11564,N_11548);
xnor U11779 (N_11779,N_11445,N_11433);
or U11780 (N_11780,N_11593,N_11432);
and U11781 (N_11781,N_11467,N_11573);
nand U11782 (N_11782,N_11427,N_11414);
nand U11783 (N_11783,N_11545,N_11588);
nand U11784 (N_11784,N_11596,N_11515);
or U11785 (N_11785,N_11429,N_11575);
xnor U11786 (N_11786,N_11552,N_11502);
nand U11787 (N_11787,N_11547,N_11584);
xnor U11788 (N_11788,N_11423,N_11480);
nor U11789 (N_11789,N_11575,N_11503);
xnor U11790 (N_11790,N_11402,N_11560);
nand U11791 (N_11791,N_11546,N_11480);
or U11792 (N_11792,N_11535,N_11481);
nand U11793 (N_11793,N_11599,N_11474);
or U11794 (N_11794,N_11574,N_11538);
or U11795 (N_11795,N_11404,N_11587);
nand U11796 (N_11796,N_11467,N_11558);
nor U11797 (N_11797,N_11582,N_11525);
xnor U11798 (N_11798,N_11564,N_11423);
nand U11799 (N_11799,N_11563,N_11468);
nand U11800 (N_11800,N_11744,N_11687);
xnor U11801 (N_11801,N_11696,N_11665);
xnor U11802 (N_11802,N_11742,N_11791);
xnor U11803 (N_11803,N_11761,N_11716);
xnor U11804 (N_11804,N_11783,N_11652);
xnor U11805 (N_11805,N_11616,N_11644);
xor U11806 (N_11806,N_11606,N_11715);
nand U11807 (N_11807,N_11718,N_11629);
nor U11808 (N_11808,N_11610,N_11774);
or U11809 (N_11809,N_11760,N_11755);
or U11810 (N_11810,N_11631,N_11739);
or U11811 (N_11811,N_11793,N_11788);
xnor U11812 (N_11812,N_11766,N_11784);
and U11813 (N_11813,N_11614,N_11638);
or U11814 (N_11814,N_11706,N_11630);
nor U11815 (N_11815,N_11680,N_11640);
xnor U11816 (N_11816,N_11688,N_11769);
xnor U11817 (N_11817,N_11771,N_11778);
or U11818 (N_11818,N_11779,N_11655);
nand U11819 (N_11819,N_11651,N_11679);
xor U11820 (N_11820,N_11666,N_11762);
nand U11821 (N_11821,N_11633,N_11741);
nand U11822 (N_11822,N_11648,N_11722);
or U11823 (N_11823,N_11796,N_11726);
and U11824 (N_11824,N_11734,N_11738);
or U11825 (N_11825,N_11621,N_11709);
or U11826 (N_11826,N_11605,N_11695);
or U11827 (N_11827,N_11659,N_11618);
nor U11828 (N_11828,N_11669,N_11745);
or U11829 (N_11829,N_11748,N_11691);
nand U11830 (N_11830,N_11780,N_11637);
nand U11831 (N_11831,N_11728,N_11746);
nand U11832 (N_11832,N_11699,N_11601);
nand U11833 (N_11833,N_11775,N_11694);
nor U11834 (N_11834,N_11609,N_11649);
or U11835 (N_11835,N_11647,N_11757);
nand U11836 (N_11836,N_11686,N_11681);
or U11837 (N_11837,N_11677,N_11619);
nor U11838 (N_11838,N_11643,N_11704);
or U11839 (N_11839,N_11765,N_11708);
nor U11840 (N_11840,N_11740,N_11636);
nor U11841 (N_11841,N_11710,N_11667);
nor U11842 (N_11842,N_11625,N_11713);
or U11843 (N_11843,N_11627,N_11763);
or U11844 (N_11844,N_11703,N_11712);
nor U11845 (N_11845,N_11777,N_11725);
and U11846 (N_11846,N_11753,N_11639);
or U11847 (N_11847,N_11721,N_11773);
xnor U11848 (N_11848,N_11797,N_11662);
nor U11849 (N_11849,N_11675,N_11671);
xor U11850 (N_11850,N_11600,N_11635);
or U11851 (N_11851,N_11611,N_11617);
nand U11852 (N_11852,N_11727,N_11795);
or U11853 (N_11853,N_11711,N_11705);
nand U11854 (N_11854,N_11731,N_11736);
and U11855 (N_11855,N_11684,N_11717);
or U11856 (N_11856,N_11789,N_11689);
xnor U11857 (N_11857,N_11624,N_11668);
or U11858 (N_11858,N_11607,N_11772);
nand U11859 (N_11859,N_11620,N_11685);
nand U11860 (N_11860,N_11690,N_11794);
nand U11861 (N_11861,N_11626,N_11692);
nand U11862 (N_11862,N_11660,N_11785);
xnor U11863 (N_11863,N_11698,N_11724);
nand U11864 (N_11864,N_11674,N_11656);
nand U11865 (N_11865,N_11653,N_11730);
nor U11866 (N_11866,N_11759,N_11747);
xor U11867 (N_11867,N_11782,N_11768);
nor U11868 (N_11868,N_11786,N_11658);
or U11869 (N_11869,N_11719,N_11714);
or U11870 (N_11870,N_11733,N_11693);
and U11871 (N_11871,N_11664,N_11654);
nand U11872 (N_11872,N_11700,N_11622);
or U11873 (N_11873,N_11781,N_11702);
nor U11874 (N_11874,N_11701,N_11729);
nor U11875 (N_11875,N_11767,N_11672);
nand U11876 (N_11876,N_11770,N_11732);
nand U11877 (N_11877,N_11628,N_11645);
or U11878 (N_11878,N_11799,N_11787);
and U11879 (N_11879,N_11683,N_11790);
and U11880 (N_11880,N_11758,N_11663);
and U11881 (N_11881,N_11678,N_11670);
nor U11882 (N_11882,N_11608,N_11661);
nand U11883 (N_11883,N_11612,N_11615);
nor U11884 (N_11884,N_11735,N_11697);
nor U11885 (N_11885,N_11602,N_11752);
xor U11886 (N_11886,N_11743,N_11754);
and U11887 (N_11887,N_11634,N_11720);
xor U11888 (N_11888,N_11764,N_11632);
and U11889 (N_11889,N_11792,N_11750);
nor U11890 (N_11890,N_11604,N_11613);
xor U11891 (N_11891,N_11603,N_11756);
xor U11892 (N_11892,N_11642,N_11673);
xnor U11893 (N_11893,N_11776,N_11737);
nor U11894 (N_11894,N_11650,N_11723);
and U11895 (N_11895,N_11676,N_11682);
or U11896 (N_11896,N_11749,N_11623);
and U11897 (N_11897,N_11641,N_11707);
nor U11898 (N_11898,N_11646,N_11751);
and U11899 (N_11899,N_11657,N_11798);
xnor U11900 (N_11900,N_11690,N_11621);
xnor U11901 (N_11901,N_11670,N_11701);
or U11902 (N_11902,N_11727,N_11737);
or U11903 (N_11903,N_11724,N_11779);
nand U11904 (N_11904,N_11750,N_11627);
nor U11905 (N_11905,N_11780,N_11766);
and U11906 (N_11906,N_11753,N_11720);
nand U11907 (N_11907,N_11794,N_11613);
or U11908 (N_11908,N_11704,N_11705);
and U11909 (N_11909,N_11784,N_11664);
or U11910 (N_11910,N_11768,N_11740);
and U11911 (N_11911,N_11600,N_11716);
nand U11912 (N_11912,N_11623,N_11713);
and U11913 (N_11913,N_11731,N_11682);
or U11914 (N_11914,N_11723,N_11607);
nor U11915 (N_11915,N_11706,N_11776);
nand U11916 (N_11916,N_11785,N_11762);
xnor U11917 (N_11917,N_11717,N_11700);
nor U11918 (N_11918,N_11730,N_11711);
or U11919 (N_11919,N_11605,N_11685);
xnor U11920 (N_11920,N_11641,N_11621);
or U11921 (N_11921,N_11736,N_11661);
xnor U11922 (N_11922,N_11713,N_11751);
and U11923 (N_11923,N_11731,N_11764);
xnor U11924 (N_11924,N_11657,N_11721);
nor U11925 (N_11925,N_11632,N_11787);
and U11926 (N_11926,N_11746,N_11743);
nand U11927 (N_11927,N_11797,N_11795);
nand U11928 (N_11928,N_11616,N_11714);
xnor U11929 (N_11929,N_11753,N_11647);
nor U11930 (N_11930,N_11641,N_11603);
nand U11931 (N_11931,N_11622,N_11797);
nand U11932 (N_11932,N_11617,N_11680);
nand U11933 (N_11933,N_11647,N_11770);
xor U11934 (N_11934,N_11687,N_11684);
and U11935 (N_11935,N_11752,N_11632);
nand U11936 (N_11936,N_11716,N_11651);
or U11937 (N_11937,N_11751,N_11785);
nand U11938 (N_11938,N_11682,N_11610);
xnor U11939 (N_11939,N_11793,N_11680);
nand U11940 (N_11940,N_11600,N_11740);
nor U11941 (N_11941,N_11613,N_11682);
nor U11942 (N_11942,N_11798,N_11754);
nor U11943 (N_11943,N_11640,N_11695);
or U11944 (N_11944,N_11640,N_11741);
nand U11945 (N_11945,N_11763,N_11692);
nand U11946 (N_11946,N_11729,N_11772);
or U11947 (N_11947,N_11713,N_11756);
xor U11948 (N_11948,N_11756,N_11693);
and U11949 (N_11949,N_11713,N_11604);
or U11950 (N_11950,N_11616,N_11703);
and U11951 (N_11951,N_11746,N_11705);
nand U11952 (N_11952,N_11633,N_11687);
or U11953 (N_11953,N_11651,N_11795);
xnor U11954 (N_11954,N_11627,N_11604);
nor U11955 (N_11955,N_11759,N_11775);
nor U11956 (N_11956,N_11746,N_11780);
and U11957 (N_11957,N_11645,N_11745);
or U11958 (N_11958,N_11606,N_11787);
and U11959 (N_11959,N_11725,N_11740);
xor U11960 (N_11960,N_11648,N_11746);
nor U11961 (N_11961,N_11794,N_11631);
xnor U11962 (N_11962,N_11636,N_11767);
nand U11963 (N_11963,N_11637,N_11734);
and U11964 (N_11964,N_11615,N_11744);
and U11965 (N_11965,N_11779,N_11621);
nand U11966 (N_11966,N_11658,N_11766);
xnor U11967 (N_11967,N_11613,N_11789);
xor U11968 (N_11968,N_11674,N_11651);
nor U11969 (N_11969,N_11603,N_11651);
and U11970 (N_11970,N_11616,N_11645);
xnor U11971 (N_11971,N_11750,N_11774);
nand U11972 (N_11972,N_11676,N_11778);
nor U11973 (N_11973,N_11671,N_11689);
nor U11974 (N_11974,N_11624,N_11686);
or U11975 (N_11975,N_11635,N_11708);
nand U11976 (N_11976,N_11774,N_11671);
nor U11977 (N_11977,N_11619,N_11610);
or U11978 (N_11978,N_11644,N_11618);
nand U11979 (N_11979,N_11621,N_11752);
nor U11980 (N_11980,N_11607,N_11692);
nand U11981 (N_11981,N_11649,N_11677);
nor U11982 (N_11982,N_11661,N_11703);
and U11983 (N_11983,N_11635,N_11741);
nor U11984 (N_11984,N_11770,N_11688);
and U11985 (N_11985,N_11758,N_11625);
nor U11986 (N_11986,N_11604,N_11694);
nand U11987 (N_11987,N_11620,N_11656);
xor U11988 (N_11988,N_11603,N_11722);
and U11989 (N_11989,N_11656,N_11624);
nor U11990 (N_11990,N_11752,N_11747);
nand U11991 (N_11991,N_11722,N_11724);
nor U11992 (N_11992,N_11644,N_11702);
nor U11993 (N_11993,N_11603,N_11749);
or U11994 (N_11994,N_11779,N_11745);
xnor U11995 (N_11995,N_11687,N_11724);
or U11996 (N_11996,N_11696,N_11774);
nor U11997 (N_11997,N_11777,N_11715);
nand U11998 (N_11998,N_11799,N_11771);
nand U11999 (N_11999,N_11710,N_11642);
nand U12000 (N_12000,N_11802,N_11814);
and U12001 (N_12001,N_11945,N_11840);
or U12002 (N_12002,N_11967,N_11807);
nor U12003 (N_12003,N_11920,N_11961);
nor U12004 (N_12004,N_11912,N_11824);
xnor U12005 (N_12005,N_11919,N_11959);
and U12006 (N_12006,N_11991,N_11935);
or U12007 (N_12007,N_11952,N_11985);
or U12008 (N_12008,N_11940,N_11877);
and U12009 (N_12009,N_11960,N_11887);
or U12010 (N_12010,N_11915,N_11990);
and U12011 (N_12011,N_11917,N_11804);
or U12012 (N_12012,N_11871,N_11843);
nor U12013 (N_12013,N_11803,N_11966);
nor U12014 (N_12014,N_11925,N_11949);
xnor U12015 (N_12015,N_11809,N_11812);
or U12016 (N_12016,N_11928,N_11813);
nor U12017 (N_12017,N_11805,N_11930);
nand U12018 (N_12018,N_11980,N_11904);
and U12019 (N_12019,N_11996,N_11842);
and U12020 (N_12020,N_11884,N_11913);
or U12021 (N_12021,N_11823,N_11878);
nand U12022 (N_12022,N_11860,N_11822);
or U12023 (N_12023,N_11825,N_11922);
nor U12024 (N_12024,N_11899,N_11908);
nand U12025 (N_12025,N_11858,N_11821);
nand U12026 (N_12026,N_11881,N_11830);
nand U12027 (N_12027,N_11886,N_11962);
nand U12028 (N_12028,N_11855,N_11907);
or U12029 (N_12029,N_11998,N_11994);
nor U12030 (N_12030,N_11834,N_11890);
and U12031 (N_12031,N_11983,N_11874);
and U12032 (N_12032,N_11995,N_11984);
xnor U12033 (N_12033,N_11936,N_11859);
nor U12034 (N_12034,N_11875,N_11948);
or U12035 (N_12035,N_11851,N_11981);
nor U12036 (N_12036,N_11808,N_11963);
and U12037 (N_12037,N_11927,N_11997);
nand U12038 (N_12038,N_11864,N_11868);
or U12039 (N_12039,N_11934,N_11872);
nand U12040 (N_12040,N_11865,N_11918);
nor U12041 (N_12041,N_11818,N_11979);
or U12042 (N_12042,N_11838,N_11953);
xnor U12043 (N_12043,N_11982,N_11911);
or U12044 (N_12044,N_11801,N_11942);
nand U12045 (N_12045,N_11856,N_11971);
or U12046 (N_12046,N_11883,N_11891);
xnor U12047 (N_12047,N_11900,N_11906);
nor U12048 (N_12048,N_11950,N_11944);
xor U12049 (N_12049,N_11810,N_11895);
and U12050 (N_12050,N_11894,N_11847);
and U12051 (N_12051,N_11866,N_11815);
nor U12052 (N_12052,N_11846,N_11880);
xor U12053 (N_12053,N_11863,N_11977);
and U12054 (N_12054,N_11987,N_11951);
nand U12055 (N_12055,N_11896,N_11969);
nand U12056 (N_12056,N_11921,N_11903);
xor U12057 (N_12057,N_11819,N_11836);
nor U12058 (N_12058,N_11811,N_11873);
xor U12059 (N_12059,N_11964,N_11816);
nor U12060 (N_12060,N_11939,N_11909);
nor U12061 (N_12061,N_11926,N_11937);
xnor U12062 (N_12062,N_11905,N_11817);
nor U12063 (N_12063,N_11888,N_11898);
and U12064 (N_12064,N_11892,N_11955);
nor U12065 (N_12065,N_11941,N_11829);
or U12066 (N_12066,N_11968,N_11889);
xor U12067 (N_12067,N_11993,N_11869);
xnor U12068 (N_12068,N_11879,N_11897);
nand U12069 (N_12069,N_11943,N_11885);
nor U12070 (N_12070,N_11999,N_11835);
nand U12071 (N_12071,N_11849,N_11931);
or U12072 (N_12072,N_11832,N_11957);
nand U12073 (N_12073,N_11970,N_11965);
and U12074 (N_12074,N_11956,N_11972);
nor U12075 (N_12075,N_11848,N_11854);
and U12076 (N_12076,N_11853,N_11841);
and U12077 (N_12077,N_11827,N_11833);
nor U12078 (N_12078,N_11916,N_11844);
nor U12079 (N_12079,N_11933,N_11958);
nor U12080 (N_12080,N_11992,N_11882);
xor U12081 (N_12081,N_11852,N_11978);
nand U12082 (N_12082,N_11861,N_11870);
nand U12083 (N_12083,N_11826,N_11932);
nand U12084 (N_12084,N_11914,N_11893);
xnor U12085 (N_12085,N_11929,N_11862);
nor U12086 (N_12086,N_11923,N_11946);
or U12087 (N_12087,N_11947,N_11901);
nor U12088 (N_12088,N_11831,N_11839);
xor U12089 (N_12089,N_11976,N_11857);
and U12090 (N_12090,N_11988,N_11845);
or U12091 (N_12091,N_11989,N_11938);
xnor U12092 (N_12092,N_11837,N_11806);
xnor U12093 (N_12093,N_11975,N_11954);
xnor U12094 (N_12094,N_11924,N_11820);
xor U12095 (N_12095,N_11974,N_11986);
xor U12096 (N_12096,N_11973,N_11910);
or U12097 (N_12097,N_11867,N_11902);
and U12098 (N_12098,N_11800,N_11828);
and U12099 (N_12099,N_11876,N_11850);
xnor U12100 (N_12100,N_11932,N_11966);
and U12101 (N_12101,N_11991,N_11898);
and U12102 (N_12102,N_11925,N_11940);
xnor U12103 (N_12103,N_11906,N_11922);
and U12104 (N_12104,N_11928,N_11973);
and U12105 (N_12105,N_11921,N_11824);
and U12106 (N_12106,N_11870,N_11805);
nand U12107 (N_12107,N_11944,N_11826);
xnor U12108 (N_12108,N_11834,N_11886);
xnor U12109 (N_12109,N_11996,N_11837);
nand U12110 (N_12110,N_11888,N_11918);
and U12111 (N_12111,N_11975,N_11842);
nand U12112 (N_12112,N_11873,N_11902);
nor U12113 (N_12113,N_11981,N_11856);
xor U12114 (N_12114,N_11991,N_11932);
nand U12115 (N_12115,N_11914,N_11860);
or U12116 (N_12116,N_11978,N_11880);
or U12117 (N_12117,N_11842,N_11845);
xor U12118 (N_12118,N_11870,N_11882);
or U12119 (N_12119,N_11866,N_11991);
or U12120 (N_12120,N_11836,N_11840);
or U12121 (N_12121,N_11955,N_11939);
nor U12122 (N_12122,N_11975,N_11895);
nand U12123 (N_12123,N_11824,N_11821);
nor U12124 (N_12124,N_11976,N_11905);
nand U12125 (N_12125,N_11993,N_11985);
and U12126 (N_12126,N_11973,N_11879);
xor U12127 (N_12127,N_11847,N_11933);
nor U12128 (N_12128,N_11890,N_11928);
or U12129 (N_12129,N_11933,N_11974);
nor U12130 (N_12130,N_11970,N_11913);
xor U12131 (N_12131,N_11827,N_11841);
nand U12132 (N_12132,N_11970,N_11860);
or U12133 (N_12133,N_11886,N_11930);
or U12134 (N_12134,N_11927,N_11943);
xnor U12135 (N_12135,N_11800,N_11947);
xor U12136 (N_12136,N_11962,N_11891);
or U12137 (N_12137,N_11981,N_11960);
or U12138 (N_12138,N_11940,N_11927);
and U12139 (N_12139,N_11985,N_11983);
nor U12140 (N_12140,N_11800,N_11897);
or U12141 (N_12141,N_11965,N_11878);
and U12142 (N_12142,N_11976,N_11950);
nand U12143 (N_12143,N_11931,N_11934);
or U12144 (N_12144,N_11848,N_11859);
and U12145 (N_12145,N_11895,N_11920);
nor U12146 (N_12146,N_11948,N_11822);
nand U12147 (N_12147,N_11887,N_11946);
or U12148 (N_12148,N_11921,N_11863);
nor U12149 (N_12149,N_11899,N_11952);
nor U12150 (N_12150,N_11899,N_11819);
nor U12151 (N_12151,N_11983,N_11865);
and U12152 (N_12152,N_11949,N_11939);
nor U12153 (N_12153,N_11823,N_11972);
or U12154 (N_12154,N_11872,N_11939);
nand U12155 (N_12155,N_11867,N_11963);
or U12156 (N_12156,N_11998,N_11846);
nand U12157 (N_12157,N_11980,N_11813);
nand U12158 (N_12158,N_11986,N_11938);
nor U12159 (N_12159,N_11937,N_11910);
nor U12160 (N_12160,N_11904,N_11868);
or U12161 (N_12161,N_11885,N_11989);
xnor U12162 (N_12162,N_11805,N_11983);
nand U12163 (N_12163,N_11957,N_11897);
nor U12164 (N_12164,N_11993,N_11927);
and U12165 (N_12165,N_11834,N_11845);
nand U12166 (N_12166,N_11833,N_11817);
or U12167 (N_12167,N_11865,N_11913);
nor U12168 (N_12168,N_11865,N_11907);
nand U12169 (N_12169,N_11835,N_11889);
nand U12170 (N_12170,N_11828,N_11864);
xnor U12171 (N_12171,N_11891,N_11966);
or U12172 (N_12172,N_11892,N_11872);
and U12173 (N_12173,N_11862,N_11959);
nor U12174 (N_12174,N_11895,N_11939);
nand U12175 (N_12175,N_11947,N_11923);
xnor U12176 (N_12176,N_11884,N_11964);
or U12177 (N_12177,N_11848,N_11862);
nand U12178 (N_12178,N_11832,N_11936);
and U12179 (N_12179,N_11867,N_11901);
nand U12180 (N_12180,N_11956,N_11803);
or U12181 (N_12181,N_11917,N_11926);
xnor U12182 (N_12182,N_11968,N_11912);
or U12183 (N_12183,N_11845,N_11874);
or U12184 (N_12184,N_11820,N_11909);
and U12185 (N_12185,N_11908,N_11809);
and U12186 (N_12186,N_11835,N_11848);
or U12187 (N_12187,N_11875,N_11917);
nor U12188 (N_12188,N_11897,N_11969);
and U12189 (N_12189,N_11942,N_11805);
xnor U12190 (N_12190,N_11848,N_11920);
xor U12191 (N_12191,N_11881,N_11889);
nand U12192 (N_12192,N_11932,N_11862);
nor U12193 (N_12193,N_11810,N_11803);
nand U12194 (N_12194,N_11845,N_11865);
xor U12195 (N_12195,N_11878,N_11867);
xor U12196 (N_12196,N_11923,N_11970);
nand U12197 (N_12197,N_11958,N_11904);
nand U12198 (N_12198,N_11857,N_11807);
and U12199 (N_12199,N_11805,N_11838);
nor U12200 (N_12200,N_12064,N_12197);
nand U12201 (N_12201,N_12167,N_12121);
nand U12202 (N_12202,N_12020,N_12126);
nor U12203 (N_12203,N_12039,N_12159);
nor U12204 (N_12204,N_12022,N_12080);
or U12205 (N_12205,N_12004,N_12062);
or U12206 (N_12206,N_12051,N_12086);
or U12207 (N_12207,N_12036,N_12001);
and U12208 (N_12208,N_12028,N_12161);
nor U12209 (N_12209,N_12168,N_12011);
or U12210 (N_12210,N_12130,N_12122);
nor U12211 (N_12211,N_12015,N_12094);
nor U12212 (N_12212,N_12025,N_12138);
nand U12213 (N_12213,N_12116,N_12089);
nand U12214 (N_12214,N_12145,N_12065);
xnor U12215 (N_12215,N_12131,N_12095);
or U12216 (N_12216,N_12069,N_12074);
or U12217 (N_12217,N_12026,N_12146);
and U12218 (N_12218,N_12085,N_12152);
xnor U12219 (N_12219,N_12093,N_12023);
xnor U12220 (N_12220,N_12190,N_12123);
and U12221 (N_12221,N_12083,N_12115);
nand U12222 (N_12222,N_12073,N_12182);
xnor U12223 (N_12223,N_12029,N_12149);
nor U12224 (N_12224,N_12195,N_12185);
nor U12225 (N_12225,N_12056,N_12194);
xor U12226 (N_12226,N_12114,N_12136);
xor U12227 (N_12227,N_12046,N_12142);
nand U12228 (N_12228,N_12158,N_12128);
and U12229 (N_12229,N_12054,N_12099);
and U12230 (N_12230,N_12030,N_12005);
and U12231 (N_12231,N_12104,N_12079);
xnor U12232 (N_12232,N_12174,N_12192);
nor U12233 (N_12233,N_12016,N_12163);
nand U12234 (N_12234,N_12012,N_12162);
or U12235 (N_12235,N_12171,N_12191);
or U12236 (N_12236,N_12187,N_12118);
xnor U12237 (N_12237,N_12019,N_12150);
nand U12238 (N_12238,N_12105,N_12018);
and U12239 (N_12239,N_12003,N_12166);
nor U12240 (N_12240,N_12169,N_12120);
nor U12241 (N_12241,N_12193,N_12063);
and U12242 (N_12242,N_12188,N_12076);
and U12243 (N_12243,N_12112,N_12058);
or U12244 (N_12244,N_12113,N_12008);
or U12245 (N_12245,N_12091,N_12100);
nand U12246 (N_12246,N_12024,N_12067);
nand U12247 (N_12247,N_12129,N_12071);
or U12248 (N_12248,N_12082,N_12108);
nand U12249 (N_12249,N_12172,N_12178);
nor U12250 (N_12250,N_12135,N_12179);
and U12251 (N_12251,N_12098,N_12141);
or U12252 (N_12252,N_12110,N_12151);
or U12253 (N_12253,N_12137,N_12035);
xnor U12254 (N_12254,N_12045,N_12006);
or U12255 (N_12255,N_12155,N_12119);
and U12256 (N_12256,N_12189,N_12014);
xnor U12257 (N_12257,N_12140,N_12077);
nor U12258 (N_12258,N_12084,N_12009);
and U12259 (N_12259,N_12081,N_12000);
or U12260 (N_12260,N_12052,N_12144);
and U12261 (N_12261,N_12165,N_12090);
xor U12262 (N_12262,N_12041,N_12139);
and U12263 (N_12263,N_12007,N_12038);
and U12264 (N_12264,N_12042,N_12132);
or U12265 (N_12265,N_12047,N_12066);
nor U12266 (N_12266,N_12124,N_12186);
nand U12267 (N_12267,N_12117,N_12002);
and U12268 (N_12268,N_12037,N_12061);
and U12269 (N_12269,N_12176,N_12075);
nor U12270 (N_12270,N_12154,N_12053);
xor U12271 (N_12271,N_12049,N_12183);
and U12272 (N_12272,N_12044,N_12050);
nor U12273 (N_12273,N_12072,N_12102);
or U12274 (N_12274,N_12088,N_12043);
nand U12275 (N_12275,N_12031,N_12157);
nand U12276 (N_12276,N_12107,N_12153);
nand U12277 (N_12277,N_12097,N_12032);
and U12278 (N_12278,N_12101,N_12106);
or U12279 (N_12279,N_12125,N_12111);
nor U12280 (N_12280,N_12060,N_12134);
and U12281 (N_12281,N_12034,N_12196);
or U12282 (N_12282,N_12164,N_12027);
nor U12283 (N_12283,N_12180,N_12070);
xor U12284 (N_12284,N_12127,N_12170);
xnor U12285 (N_12285,N_12175,N_12109);
xnor U12286 (N_12286,N_12013,N_12173);
xnor U12287 (N_12287,N_12148,N_12068);
xnor U12288 (N_12288,N_12087,N_12147);
nor U12289 (N_12289,N_12199,N_12198);
or U12290 (N_12290,N_12143,N_12181);
or U12291 (N_12291,N_12033,N_12078);
nor U12292 (N_12292,N_12177,N_12096);
and U12293 (N_12293,N_12103,N_12040);
nor U12294 (N_12294,N_12184,N_12059);
nand U12295 (N_12295,N_12156,N_12160);
nor U12296 (N_12296,N_12017,N_12133);
or U12297 (N_12297,N_12092,N_12048);
or U12298 (N_12298,N_12010,N_12021);
or U12299 (N_12299,N_12057,N_12055);
xnor U12300 (N_12300,N_12174,N_12078);
xnor U12301 (N_12301,N_12072,N_12168);
or U12302 (N_12302,N_12091,N_12138);
or U12303 (N_12303,N_12081,N_12010);
nand U12304 (N_12304,N_12195,N_12054);
xnor U12305 (N_12305,N_12120,N_12163);
nand U12306 (N_12306,N_12081,N_12119);
nor U12307 (N_12307,N_12000,N_12155);
nor U12308 (N_12308,N_12019,N_12097);
or U12309 (N_12309,N_12164,N_12016);
or U12310 (N_12310,N_12048,N_12132);
and U12311 (N_12311,N_12116,N_12182);
and U12312 (N_12312,N_12148,N_12002);
or U12313 (N_12313,N_12091,N_12196);
or U12314 (N_12314,N_12006,N_12013);
nor U12315 (N_12315,N_12197,N_12089);
and U12316 (N_12316,N_12178,N_12156);
nor U12317 (N_12317,N_12169,N_12111);
and U12318 (N_12318,N_12185,N_12091);
nand U12319 (N_12319,N_12088,N_12037);
xnor U12320 (N_12320,N_12051,N_12183);
or U12321 (N_12321,N_12001,N_12097);
or U12322 (N_12322,N_12095,N_12183);
or U12323 (N_12323,N_12105,N_12024);
and U12324 (N_12324,N_12092,N_12166);
xor U12325 (N_12325,N_12084,N_12143);
nand U12326 (N_12326,N_12140,N_12051);
and U12327 (N_12327,N_12132,N_12157);
and U12328 (N_12328,N_12133,N_12134);
or U12329 (N_12329,N_12014,N_12122);
and U12330 (N_12330,N_12186,N_12104);
and U12331 (N_12331,N_12178,N_12186);
nand U12332 (N_12332,N_12113,N_12060);
and U12333 (N_12333,N_12148,N_12174);
xor U12334 (N_12334,N_12193,N_12118);
or U12335 (N_12335,N_12157,N_12058);
and U12336 (N_12336,N_12028,N_12179);
nand U12337 (N_12337,N_12111,N_12023);
and U12338 (N_12338,N_12035,N_12083);
or U12339 (N_12339,N_12184,N_12077);
and U12340 (N_12340,N_12162,N_12164);
nor U12341 (N_12341,N_12179,N_12062);
or U12342 (N_12342,N_12176,N_12141);
or U12343 (N_12343,N_12173,N_12109);
nor U12344 (N_12344,N_12180,N_12194);
nand U12345 (N_12345,N_12118,N_12042);
xnor U12346 (N_12346,N_12009,N_12024);
or U12347 (N_12347,N_12164,N_12052);
or U12348 (N_12348,N_12049,N_12077);
and U12349 (N_12349,N_12124,N_12037);
and U12350 (N_12350,N_12037,N_12152);
nor U12351 (N_12351,N_12151,N_12085);
nand U12352 (N_12352,N_12019,N_12057);
or U12353 (N_12353,N_12003,N_12066);
nor U12354 (N_12354,N_12061,N_12064);
and U12355 (N_12355,N_12119,N_12061);
nand U12356 (N_12356,N_12006,N_12030);
and U12357 (N_12357,N_12198,N_12137);
nand U12358 (N_12358,N_12160,N_12180);
xnor U12359 (N_12359,N_12060,N_12080);
or U12360 (N_12360,N_12084,N_12023);
nor U12361 (N_12361,N_12137,N_12020);
or U12362 (N_12362,N_12127,N_12019);
and U12363 (N_12363,N_12011,N_12098);
nand U12364 (N_12364,N_12090,N_12048);
or U12365 (N_12365,N_12153,N_12060);
nand U12366 (N_12366,N_12074,N_12031);
or U12367 (N_12367,N_12073,N_12038);
nand U12368 (N_12368,N_12154,N_12116);
nor U12369 (N_12369,N_12161,N_12187);
and U12370 (N_12370,N_12038,N_12099);
nand U12371 (N_12371,N_12030,N_12019);
or U12372 (N_12372,N_12125,N_12142);
xor U12373 (N_12373,N_12149,N_12069);
nand U12374 (N_12374,N_12159,N_12100);
xor U12375 (N_12375,N_12012,N_12027);
xor U12376 (N_12376,N_12029,N_12044);
or U12377 (N_12377,N_12188,N_12145);
and U12378 (N_12378,N_12132,N_12125);
or U12379 (N_12379,N_12149,N_12138);
nand U12380 (N_12380,N_12101,N_12063);
xor U12381 (N_12381,N_12050,N_12074);
nor U12382 (N_12382,N_12049,N_12148);
xor U12383 (N_12383,N_12171,N_12160);
nand U12384 (N_12384,N_12126,N_12196);
and U12385 (N_12385,N_12048,N_12072);
xnor U12386 (N_12386,N_12041,N_12040);
or U12387 (N_12387,N_12182,N_12040);
xnor U12388 (N_12388,N_12117,N_12053);
nor U12389 (N_12389,N_12160,N_12074);
nand U12390 (N_12390,N_12074,N_12044);
nor U12391 (N_12391,N_12097,N_12014);
and U12392 (N_12392,N_12037,N_12057);
and U12393 (N_12393,N_12017,N_12172);
nor U12394 (N_12394,N_12117,N_12124);
xnor U12395 (N_12395,N_12089,N_12168);
nor U12396 (N_12396,N_12076,N_12164);
and U12397 (N_12397,N_12060,N_12103);
nor U12398 (N_12398,N_12052,N_12118);
nand U12399 (N_12399,N_12163,N_12058);
nand U12400 (N_12400,N_12289,N_12270);
and U12401 (N_12401,N_12333,N_12348);
nand U12402 (N_12402,N_12243,N_12278);
nor U12403 (N_12403,N_12203,N_12232);
nand U12404 (N_12404,N_12241,N_12363);
or U12405 (N_12405,N_12223,N_12207);
xnor U12406 (N_12406,N_12376,N_12386);
or U12407 (N_12407,N_12246,N_12364);
or U12408 (N_12408,N_12209,N_12344);
nor U12409 (N_12409,N_12225,N_12211);
xor U12410 (N_12410,N_12313,N_12339);
nor U12411 (N_12411,N_12327,N_12325);
xor U12412 (N_12412,N_12321,N_12240);
nor U12413 (N_12413,N_12249,N_12276);
or U12414 (N_12414,N_12286,N_12271);
nand U12415 (N_12415,N_12347,N_12396);
nor U12416 (N_12416,N_12268,N_12326);
or U12417 (N_12417,N_12329,N_12288);
nor U12418 (N_12418,N_12301,N_12389);
xor U12419 (N_12419,N_12366,N_12295);
nor U12420 (N_12420,N_12315,N_12282);
or U12421 (N_12421,N_12338,N_12201);
or U12422 (N_12422,N_12334,N_12245);
nand U12423 (N_12423,N_12350,N_12222);
xnor U12424 (N_12424,N_12262,N_12320);
nor U12425 (N_12425,N_12224,N_12265);
nor U12426 (N_12426,N_12229,N_12285);
or U12427 (N_12427,N_12216,N_12210);
and U12428 (N_12428,N_12208,N_12252);
nand U12429 (N_12429,N_12353,N_12258);
and U12430 (N_12430,N_12324,N_12269);
xnor U12431 (N_12431,N_12332,N_12390);
and U12432 (N_12432,N_12302,N_12316);
and U12433 (N_12433,N_12261,N_12365);
nor U12434 (N_12434,N_12238,N_12360);
xnor U12435 (N_12435,N_12399,N_12349);
or U12436 (N_12436,N_12356,N_12293);
nand U12437 (N_12437,N_12234,N_12263);
nand U12438 (N_12438,N_12358,N_12228);
xnor U12439 (N_12439,N_12212,N_12250);
and U12440 (N_12440,N_12314,N_12242);
nor U12441 (N_12441,N_12235,N_12279);
or U12442 (N_12442,N_12287,N_12274);
nand U12443 (N_12443,N_12323,N_12373);
and U12444 (N_12444,N_12200,N_12305);
xnor U12445 (N_12445,N_12273,N_12281);
xnor U12446 (N_12446,N_12237,N_12283);
nor U12447 (N_12447,N_12395,N_12371);
nand U12448 (N_12448,N_12205,N_12384);
or U12449 (N_12449,N_12236,N_12379);
nand U12450 (N_12450,N_12394,N_12215);
nand U12451 (N_12451,N_12361,N_12369);
xor U12452 (N_12452,N_12259,N_12256);
and U12453 (N_12453,N_12367,N_12398);
xor U12454 (N_12454,N_12351,N_12254);
and U12455 (N_12455,N_12217,N_12202);
xor U12456 (N_12456,N_12296,N_12392);
nand U12457 (N_12457,N_12357,N_12312);
xnor U12458 (N_12458,N_12337,N_12267);
nand U12459 (N_12459,N_12214,N_12255);
or U12460 (N_12460,N_12391,N_12290);
xor U12461 (N_12461,N_12294,N_12204);
nand U12462 (N_12462,N_12385,N_12382);
nand U12463 (N_12463,N_12219,N_12297);
or U12464 (N_12464,N_12298,N_12330);
and U12465 (N_12465,N_12355,N_12335);
or U12466 (N_12466,N_12336,N_12253);
xor U12467 (N_12467,N_12372,N_12368);
xor U12468 (N_12468,N_12352,N_12277);
xor U12469 (N_12469,N_12393,N_12317);
and U12470 (N_12470,N_12310,N_12354);
or U12471 (N_12471,N_12244,N_12304);
nand U12472 (N_12472,N_12387,N_12362);
or U12473 (N_12473,N_12218,N_12342);
and U12474 (N_12474,N_12343,N_12397);
and U12475 (N_12475,N_12300,N_12233);
xor U12476 (N_12476,N_12378,N_12380);
or U12477 (N_12477,N_12307,N_12275);
or U12478 (N_12478,N_12206,N_12306);
nand U12479 (N_12479,N_12213,N_12309);
nand U12480 (N_12480,N_12341,N_12308);
or U12481 (N_12481,N_12377,N_12299);
xnor U12482 (N_12482,N_12266,N_12221);
xnor U12483 (N_12483,N_12292,N_12247);
and U12484 (N_12484,N_12251,N_12375);
xnor U12485 (N_12485,N_12322,N_12291);
nand U12486 (N_12486,N_12272,N_12359);
or U12487 (N_12487,N_12374,N_12284);
xor U12488 (N_12488,N_12230,N_12340);
nor U12489 (N_12489,N_12319,N_12220);
or U12490 (N_12490,N_12257,N_12331);
and U12491 (N_12491,N_12383,N_12248);
nor U12492 (N_12492,N_12311,N_12231);
nor U12493 (N_12493,N_12280,N_12303);
xnor U12494 (N_12494,N_12227,N_12318);
or U12495 (N_12495,N_12345,N_12264);
nor U12496 (N_12496,N_12226,N_12260);
nor U12497 (N_12497,N_12239,N_12346);
nor U12498 (N_12498,N_12381,N_12328);
and U12499 (N_12499,N_12388,N_12370);
nor U12500 (N_12500,N_12377,N_12388);
or U12501 (N_12501,N_12247,N_12272);
nand U12502 (N_12502,N_12330,N_12366);
xnor U12503 (N_12503,N_12269,N_12288);
nand U12504 (N_12504,N_12378,N_12333);
and U12505 (N_12505,N_12253,N_12331);
xor U12506 (N_12506,N_12260,N_12333);
xnor U12507 (N_12507,N_12388,N_12336);
nand U12508 (N_12508,N_12301,N_12246);
nor U12509 (N_12509,N_12272,N_12350);
xor U12510 (N_12510,N_12245,N_12264);
nor U12511 (N_12511,N_12209,N_12387);
nand U12512 (N_12512,N_12250,N_12200);
or U12513 (N_12513,N_12339,N_12257);
nand U12514 (N_12514,N_12218,N_12203);
nand U12515 (N_12515,N_12272,N_12274);
nand U12516 (N_12516,N_12319,N_12257);
nand U12517 (N_12517,N_12279,N_12332);
nor U12518 (N_12518,N_12338,N_12224);
or U12519 (N_12519,N_12340,N_12310);
or U12520 (N_12520,N_12340,N_12293);
xnor U12521 (N_12521,N_12225,N_12347);
or U12522 (N_12522,N_12398,N_12309);
nand U12523 (N_12523,N_12222,N_12203);
xor U12524 (N_12524,N_12314,N_12210);
or U12525 (N_12525,N_12302,N_12360);
or U12526 (N_12526,N_12332,N_12218);
and U12527 (N_12527,N_12234,N_12334);
and U12528 (N_12528,N_12231,N_12331);
and U12529 (N_12529,N_12321,N_12341);
xnor U12530 (N_12530,N_12374,N_12211);
or U12531 (N_12531,N_12351,N_12285);
and U12532 (N_12532,N_12253,N_12381);
nor U12533 (N_12533,N_12354,N_12387);
xnor U12534 (N_12534,N_12206,N_12392);
nor U12535 (N_12535,N_12249,N_12202);
xnor U12536 (N_12536,N_12372,N_12226);
nand U12537 (N_12537,N_12214,N_12212);
and U12538 (N_12538,N_12288,N_12383);
or U12539 (N_12539,N_12309,N_12320);
xor U12540 (N_12540,N_12324,N_12283);
nand U12541 (N_12541,N_12234,N_12357);
nor U12542 (N_12542,N_12367,N_12210);
or U12543 (N_12543,N_12289,N_12332);
and U12544 (N_12544,N_12235,N_12239);
or U12545 (N_12545,N_12391,N_12229);
or U12546 (N_12546,N_12363,N_12224);
xnor U12547 (N_12547,N_12292,N_12353);
nor U12548 (N_12548,N_12344,N_12399);
and U12549 (N_12549,N_12262,N_12342);
nand U12550 (N_12550,N_12330,N_12329);
or U12551 (N_12551,N_12211,N_12368);
or U12552 (N_12552,N_12288,N_12354);
or U12553 (N_12553,N_12293,N_12305);
and U12554 (N_12554,N_12278,N_12371);
nor U12555 (N_12555,N_12362,N_12342);
nand U12556 (N_12556,N_12237,N_12208);
xnor U12557 (N_12557,N_12326,N_12309);
and U12558 (N_12558,N_12369,N_12201);
and U12559 (N_12559,N_12292,N_12387);
nand U12560 (N_12560,N_12395,N_12321);
and U12561 (N_12561,N_12314,N_12268);
or U12562 (N_12562,N_12308,N_12260);
nor U12563 (N_12563,N_12368,N_12290);
nor U12564 (N_12564,N_12219,N_12339);
nand U12565 (N_12565,N_12368,N_12244);
nand U12566 (N_12566,N_12326,N_12233);
nand U12567 (N_12567,N_12349,N_12343);
xnor U12568 (N_12568,N_12352,N_12371);
and U12569 (N_12569,N_12243,N_12296);
nand U12570 (N_12570,N_12228,N_12373);
nor U12571 (N_12571,N_12394,N_12295);
nand U12572 (N_12572,N_12239,N_12210);
or U12573 (N_12573,N_12386,N_12275);
nand U12574 (N_12574,N_12293,N_12372);
and U12575 (N_12575,N_12356,N_12221);
nor U12576 (N_12576,N_12389,N_12208);
nor U12577 (N_12577,N_12265,N_12234);
and U12578 (N_12578,N_12390,N_12209);
xnor U12579 (N_12579,N_12239,N_12340);
and U12580 (N_12580,N_12271,N_12383);
and U12581 (N_12581,N_12287,N_12236);
nor U12582 (N_12582,N_12316,N_12397);
nand U12583 (N_12583,N_12294,N_12200);
and U12584 (N_12584,N_12212,N_12398);
xor U12585 (N_12585,N_12362,N_12252);
xor U12586 (N_12586,N_12283,N_12320);
and U12587 (N_12587,N_12232,N_12245);
nand U12588 (N_12588,N_12201,N_12266);
nand U12589 (N_12589,N_12325,N_12388);
and U12590 (N_12590,N_12234,N_12209);
and U12591 (N_12591,N_12212,N_12360);
nor U12592 (N_12592,N_12369,N_12373);
nor U12593 (N_12593,N_12393,N_12303);
nor U12594 (N_12594,N_12353,N_12237);
and U12595 (N_12595,N_12207,N_12371);
nor U12596 (N_12596,N_12279,N_12253);
nand U12597 (N_12597,N_12397,N_12322);
xnor U12598 (N_12598,N_12205,N_12278);
and U12599 (N_12599,N_12324,N_12285);
and U12600 (N_12600,N_12439,N_12472);
nand U12601 (N_12601,N_12547,N_12554);
and U12602 (N_12602,N_12443,N_12591);
nand U12603 (N_12603,N_12454,N_12568);
or U12604 (N_12604,N_12465,N_12423);
xor U12605 (N_12605,N_12553,N_12408);
or U12606 (N_12606,N_12557,N_12461);
xnor U12607 (N_12607,N_12415,N_12511);
nand U12608 (N_12608,N_12561,N_12556);
nand U12609 (N_12609,N_12407,N_12411);
and U12610 (N_12610,N_12512,N_12530);
xnor U12611 (N_12611,N_12508,N_12542);
or U12612 (N_12612,N_12495,N_12570);
xor U12613 (N_12613,N_12533,N_12464);
or U12614 (N_12614,N_12589,N_12573);
or U12615 (N_12615,N_12513,N_12492);
nor U12616 (N_12616,N_12565,N_12425);
and U12617 (N_12617,N_12414,N_12469);
and U12618 (N_12618,N_12522,N_12489);
xor U12619 (N_12619,N_12478,N_12456);
nand U12620 (N_12620,N_12545,N_12501);
or U12621 (N_12621,N_12479,N_12577);
or U12622 (N_12622,N_12452,N_12598);
xnor U12623 (N_12623,N_12567,N_12482);
and U12624 (N_12624,N_12449,N_12535);
or U12625 (N_12625,N_12437,N_12442);
nand U12626 (N_12626,N_12592,N_12420);
or U12627 (N_12627,N_12585,N_12559);
and U12628 (N_12628,N_12524,N_12509);
xor U12629 (N_12629,N_12529,N_12597);
or U12630 (N_12630,N_12517,N_12537);
nor U12631 (N_12631,N_12502,N_12453);
nand U12632 (N_12632,N_12587,N_12519);
or U12633 (N_12633,N_12562,N_12419);
or U12634 (N_12634,N_12434,N_12458);
and U12635 (N_12635,N_12560,N_12536);
nor U12636 (N_12636,N_12487,N_12520);
xnor U12637 (N_12637,N_12447,N_12582);
or U12638 (N_12638,N_12563,N_12468);
nor U12639 (N_12639,N_12483,N_12595);
nand U12640 (N_12640,N_12444,N_12599);
nand U12641 (N_12641,N_12543,N_12481);
xor U12642 (N_12642,N_12485,N_12438);
nor U12643 (N_12643,N_12402,N_12540);
and U12644 (N_12644,N_12590,N_12571);
and U12645 (N_12645,N_12475,N_12410);
or U12646 (N_12646,N_12583,N_12596);
or U12647 (N_12647,N_12578,N_12588);
nand U12648 (N_12648,N_12523,N_12499);
or U12649 (N_12649,N_12538,N_12579);
xor U12650 (N_12650,N_12586,N_12555);
and U12651 (N_12651,N_12466,N_12418);
nor U12652 (N_12652,N_12433,N_12566);
nand U12653 (N_12653,N_12500,N_12572);
nor U12654 (N_12654,N_12440,N_12431);
xnor U12655 (N_12655,N_12470,N_12525);
nand U12656 (N_12656,N_12436,N_12497);
nand U12657 (N_12657,N_12409,N_12455);
nand U12658 (N_12658,N_12416,N_12460);
nor U12659 (N_12659,N_12548,N_12575);
and U12660 (N_12660,N_12518,N_12514);
nand U12661 (N_12661,N_12550,N_12480);
and U12662 (N_12662,N_12510,N_12457);
or U12663 (N_12663,N_12463,N_12450);
and U12664 (N_12664,N_12569,N_12486);
xnor U12665 (N_12665,N_12403,N_12441);
nor U12666 (N_12666,N_12526,N_12491);
nand U12667 (N_12667,N_12534,N_12506);
and U12668 (N_12668,N_12421,N_12488);
and U12669 (N_12669,N_12435,N_12504);
nand U12670 (N_12670,N_12404,N_12459);
and U12671 (N_12671,N_12432,N_12594);
xor U12672 (N_12672,N_12412,N_12576);
nor U12673 (N_12673,N_12494,N_12544);
nor U12674 (N_12674,N_12428,N_12498);
nor U12675 (N_12675,N_12552,N_12516);
nor U12676 (N_12676,N_12527,N_12564);
xor U12677 (N_12677,N_12471,N_12473);
or U12678 (N_12678,N_12515,N_12462);
or U12679 (N_12679,N_12406,N_12445);
xor U12680 (N_12680,N_12476,N_12580);
nand U12681 (N_12681,N_12546,N_12474);
or U12682 (N_12682,N_12574,N_12581);
nand U12683 (N_12683,N_12490,N_12401);
nor U12684 (N_12684,N_12427,N_12417);
nor U12685 (N_12685,N_12539,N_12413);
xor U12686 (N_12686,N_12496,N_12551);
nor U12687 (N_12687,N_12451,N_12532);
and U12688 (N_12688,N_12422,N_12521);
nand U12689 (N_12689,N_12584,N_12446);
nor U12690 (N_12690,N_12405,N_12503);
or U12691 (N_12691,N_12507,N_12429);
nand U12692 (N_12692,N_12477,N_12426);
and U12693 (N_12693,N_12541,N_12424);
nor U12694 (N_12694,N_12400,N_12484);
or U12695 (N_12695,N_12448,N_12528);
xnor U12696 (N_12696,N_12430,N_12593);
xor U12697 (N_12697,N_12549,N_12467);
or U12698 (N_12698,N_12505,N_12493);
nor U12699 (N_12699,N_12531,N_12558);
nor U12700 (N_12700,N_12513,N_12490);
nor U12701 (N_12701,N_12585,N_12501);
nor U12702 (N_12702,N_12492,N_12447);
nor U12703 (N_12703,N_12420,N_12459);
xnor U12704 (N_12704,N_12464,N_12525);
xor U12705 (N_12705,N_12482,N_12450);
nor U12706 (N_12706,N_12497,N_12496);
xnor U12707 (N_12707,N_12480,N_12534);
nor U12708 (N_12708,N_12419,N_12475);
xnor U12709 (N_12709,N_12487,N_12562);
nor U12710 (N_12710,N_12400,N_12556);
nand U12711 (N_12711,N_12416,N_12488);
and U12712 (N_12712,N_12462,N_12465);
or U12713 (N_12713,N_12561,N_12477);
or U12714 (N_12714,N_12540,N_12408);
nand U12715 (N_12715,N_12532,N_12431);
nor U12716 (N_12716,N_12527,N_12594);
and U12717 (N_12717,N_12433,N_12435);
or U12718 (N_12718,N_12593,N_12409);
or U12719 (N_12719,N_12422,N_12554);
xnor U12720 (N_12720,N_12421,N_12555);
and U12721 (N_12721,N_12536,N_12507);
xnor U12722 (N_12722,N_12416,N_12477);
nor U12723 (N_12723,N_12541,N_12520);
and U12724 (N_12724,N_12400,N_12568);
nand U12725 (N_12725,N_12568,N_12590);
and U12726 (N_12726,N_12422,N_12549);
nand U12727 (N_12727,N_12505,N_12424);
or U12728 (N_12728,N_12553,N_12561);
and U12729 (N_12729,N_12482,N_12466);
or U12730 (N_12730,N_12446,N_12464);
nand U12731 (N_12731,N_12526,N_12442);
and U12732 (N_12732,N_12549,N_12455);
nor U12733 (N_12733,N_12539,N_12548);
nor U12734 (N_12734,N_12536,N_12584);
or U12735 (N_12735,N_12410,N_12452);
and U12736 (N_12736,N_12518,N_12536);
and U12737 (N_12737,N_12565,N_12400);
xor U12738 (N_12738,N_12593,N_12408);
nand U12739 (N_12739,N_12587,N_12481);
nor U12740 (N_12740,N_12595,N_12480);
nor U12741 (N_12741,N_12501,N_12464);
nand U12742 (N_12742,N_12410,N_12555);
nor U12743 (N_12743,N_12411,N_12466);
xor U12744 (N_12744,N_12404,N_12457);
or U12745 (N_12745,N_12547,N_12524);
nor U12746 (N_12746,N_12483,N_12408);
nor U12747 (N_12747,N_12497,N_12595);
and U12748 (N_12748,N_12546,N_12563);
nand U12749 (N_12749,N_12424,N_12590);
nand U12750 (N_12750,N_12439,N_12404);
and U12751 (N_12751,N_12431,N_12402);
nor U12752 (N_12752,N_12543,N_12506);
or U12753 (N_12753,N_12414,N_12480);
and U12754 (N_12754,N_12500,N_12531);
nand U12755 (N_12755,N_12551,N_12589);
and U12756 (N_12756,N_12535,N_12411);
xnor U12757 (N_12757,N_12573,N_12525);
xor U12758 (N_12758,N_12514,N_12554);
or U12759 (N_12759,N_12553,N_12490);
nand U12760 (N_12760,N_12565,N_12470);
or U12761 (N_12761,N_12552,N_12522);
and U12762 (N_12762,N_12565,N_12547);
nor U12763 (N_12763,N_12533,N_12590);
or U12764 (N_12764,N_12536,N_12410);
and U12765 (N_12765,N_12550,N_12531);
nor U12766 (N_12766,N_12577,N_12483);
nand U12767 (N_12767,N_12566,N_12518);
nand U12768 (N_12768,N_12507,N_12505);
nand U12769 (N_12769,N_12480,N_12540);
and U12770 (N_12770,N_12454,N_12584);
nand U12771 (N_12771,N_12497,N_12486);
nor U12772 (N_12772,N_12419,N_12425);
or U12773 (N_12773,N_12555,N_12546);
xnor U12774 (N_12774,N_12575,N_12436);
and U12775 (N_12775,N_12542,N_12519);
and U12776 (N_12776,N_12464,N_12594);
nor U12777 (N_12777,N_12486,N_12457);
nand U12778 (N_12778,N_12410,N_12561);
or U12779 (N_12779,N_12430,N_12541);
nand U12780 (N_12780,N_12523,N_12459);
nand U12781 (N_12781,N_12422,N_12568);
xor U12782 (N_12782,N_12549,N_12505);
and U12783 (N_12783,N_12486,N_12426);
and U12784 (N_12784,N_12444,N_12567);
and U12785 (N_12785,N_12546,N_12473);
xor U12786 (N_12786,N_12571,N_12505);
and U12787 (N_12787,N_12524,N_12430);
and U12788 (N_12788,N_12504,N_12558);
or U12789 (N_12789,N_12565,N_12592);
nand U12790 (N_12790,N_12439,N_12465);
xnor U12791 (N_12791,N_12433,N_12525);
or U12792 (N_12792,N_12433,N_12462);
or U12793 (N_12793,N_12534,N_12431);
nand U12794 (N_12794,N_12525,N_12561);
nand U12795 (N_12795,N_12553,N_12547);
or U12796 (N_12796,N_12561,N_12489);
nand U12797 (N_12797,N_12468,N_12437);
nor U12798 (N_12798,N_12594,N_12563);
or U12799 (N_12799,N_12459,N_12519);
or U12800 (N_12800,N_12632,N_12753);
xnor U12801 (N_12801,N_12774,N_12718);
and U12802 (N_12802,N_12710,N_12713);
nor U12803 (N_12803,N_12676,N_12734);
xor U12804 (N_12804,N_12649,N_12697);
or U12805 (N_12805,N_12617,N_12664);
or U12806 (N_12806,N_12669,N_12764);
or U12807 (N_12807,N_12742,N_12767);
or U12808 (N_12808,N_12610,N_12611);
or U12809 (N_12809,N_12749,N_12620);
and U12810 (N_12810,N_12738,N_12691);
or U12811 (N_12811,N_12715,N_12681);
or U12812 (N_12812,N_12793,N_12714);
nor U12813 (N_12813,N_12772,N_12607);
xor U12814 (N_12814,N_12616,N_12651);
or U12815 (N_12815,N_12799,N_12618);
xnor U12816 (N_12816,N_12601,N_12604);
nor U12817 (N_12817,N_12762,N_12790);
and U12818 (N_12818,N_12795,N_12638);
nand U12819 (N_12819,N_12686,N_12673);
or U12820 (N_12820,N_12606,N_12675);
nand U12821 (N_12821,N_12736,N_12631);
nor U12822 (N_12822,N_12609,N_12771);
or U12823 (N_12823,N_12747,N_12667);
xnor U12824 (N_12824,N_12706,N_12693);
xor U12825 (N_12825,N_12782,N_12692);
or U12826 (N_12826,N_12623,N_12643);
xnor U12827 (N_12827,N_12724,N_12694);
and U12828 (N_12828,N_12626,N_12754);
or U12829 (N_12829,N_12777,N_12615);
or U12830 (N_12830,N_12683,N_12725);
nand U12831 (N_12831,N_12674,N_12612);
or U12832 (N_12832,N_12729,N_12644);
nor U12833 (N_12833,N_12658,N_12746);
and U12834 (N_12834,N_12639,N_12761);
xor U12835 (N_12835,N_12688,N_12752);
or U12836 (N_12836,N_12656,N_12717);
nand U12837 (N_12837,N_12755,N_12640);
or U12838 (N_12838,N_12744,N_12627);
or U12839 (N_12839,N_12766,N_12657);
nor U12840 (N_12840,N_12653,N_12698);
nor U12841 (N_12841,N_12659,N_12671);
nor U12842 (N_12842,N_12797,N_12655);
nand U12843 (N_12843,N_12677,N_12721);
nor U12844 (N_12844,N_12779,N_12679);
nor U12845 (N_12845,N_12647,N_12719);
or U12846 (N_12846,N_12625,N_12757);
or U12847 (N_12847,N_12684,N_12728);
and U12848 (N_12848,N_12605,N_12743);
nor U12849 (N_12849,N_12758,N_12701);
nor U12850 (N_12850,N_12751,N_12796);
nand U12851 (N_12851,N_12603,N_12662);
nor U12852 (N_12852,N_12711,N_12629);
nor U12853 (N_12853,N_12776,N_12763);
or U12854 (N_12854,N_12712,N_12622);
or U12855 (N_12855,N_12773,N_12784);
nand U12856 (N_12856,N_12633,N_12720);
and U12857 (N_12857,N_12702,N_12678);
or U12858 (N_12858,N_12727,N_12786);
xnor U12859 (N_12859,N_12789,N_12608);
and U12860 (N_12860,N_12652,N_12646);
or U12861 (N_12861,N_12785,N_12630);
xnor U12862 (N_12862,N_12741,N_12672);
and U12863 (N_12863,N_12619,N_12648);
xor U12864 (N_12864,N_12654,N_12794);
xnor U12865 (N_12865,N_12716,N_12775);
or U12866 (N_12866,N_12791,N_12624);
nand U12867 (N_12867,N_12663,N_12628);
xor U12868 (N_12868,N_12769,N_12745);
xor U12869 (N_12869,N_12768,N_12634);
nand U12870 (N_12870,N_12735,N_12726);
xnor U12871 (N_12871,N_12642,N_12740);
and U12872 (N_12872,N_12707,N_12670);
xor U12873 (N_12873,N_12703,N_12760);
and U12874 (N_12874,N_12783,N_12732);
and U12875 (N_12875,N_12690,N_12636);
xor U12876 (N_12876,N_12787,N_12699);
xor U12877 (N_12877,N_12687,N_12668);
nor U12878 (N_12878,N_12650,N_12750);
xor U12879 (N_12879,N_12635,N_12781);
or U12880 (N_12880,N_12723,N_12759);
and U12881 (N_12881,N_12770,N_12733);
nor U12882 (N_12882,N_12685,N_12704);
nor U12883 (N_12883,N_12700,N_12621);
nand U12884 (N_12884,N_12730,N_12765);
and U12885 (N_12885,N_12665,N_12731);
nand U12886 (N_12886,N_12645,N_12689);
or U12887 (N_12887,N_12788,N_12737);
and U12888 (N_12888,N_12722,N_12748);
and U12889 (N_12889,N_12798,N_12780);
xnor U12890 (N_12890,N_12695,N_12602);
nor U12891 (N_12891,N_12708,N_12778);
nand U12892 (N_12892,N_12600,N_12637);
and U12893 (N_12893,N_12756,N_12666);
nand U12894 (N_12894,N_12613,N_12696);
and U12895 (N_12895,N_12709,N_12661);
xnor U12896 (N_12896,N_12739,N_12705);
or U12897 (N_12897,N_12792,N_12641);
and U12898 (N_12898,N_12660,N_12682);
and U12899 (N_12899,N_12680,N_12614);
and U12900 (N_12900,N_12748,N_12694);
xnor U12901 (N_12901,N_12702,N_12760);
and U12902 (N_12902,N_12740,N_12622);
and U12903 (N_12903,N_12656,N_12755);
and U12904 (N_12904,N_12731,N_12695);
xor U12905 (N_12905,N_12606,N_12755);
xor U12906 (N_12906,N_12762,N_12611);
or U12907 (N_12907,N_12621,N_12605);
and U12908 (N_12908,N_12705,N_12734);
and U12909 (N_12909,N_12673,N_12637);
or U12910 (N_12910,N_12795,N_12617);
nor U12911 (N_12911,N_12741,N_12738);
xnor U12912 (N_12912,N_12636,N_12664);
or U12913 (N_12913,N_12676,N_12742);
and U12914 (N_12914,N_12705,N_12770);
xnor U12915 (N_12915,N_12603,N_12613);
nor U12916 (N_12916,N_12657,N_12636);
xor U12917 (N_12917,N_12744,N_12798);
nor U12918 (N_12918,N_12794,N_12715);
or U12919 (N_12919,N_12756,N_12681);
nand U12920 (N_12920,N_12634,N_12641);
nand U12921 (N_12921,N_12677,N_12664);
and U12922 (N_12922,N_12611,N_12785);
or U12923 (N_12923,N_12671,N_12756);
xnor U12924 (N_12924,N_12679,N_12790);
or U12925 (N_12925,N_12684,N_12783);
and U12926 (N_12926,N_12660,N_12653);
xnor U12927 (N_12927,N_12743,N_12685);
nor U12928 (N_12928,N_12666,N_12650);
xor U12929 (N_12929,N_12760,N_12602);
nand U12930 (N_12930,N_12639,N_12622);
nor U12931 (N_12931,N_12695,N_12748);
or U12932 (N_12932,N_12614,N_12609);
or U12933 (N_12933,N_12638,N_12791);
nand U12934 (N_12934,N_12650,N_12609);
nor U12935 (N_12935,N_12643,N_12619);
or U12936 (N_12936,N_12765,N_12767);
xor U12937 (N_12937,N_12660,N_12626);
nor U12938 (N_12938,N_12756,N_12753);
nand U12939 (N_12939,N_12627,N_12758);
or U12940 (N_12940,N_12769,N_12770);
and U12941 (N_12941,N_12730,N_12775);
xnor U12942 (N_12942,N_12621,N_12684);
nand U12943 (N_12943,N_12607,N_12789);
nand U12944 (N_12944,N_12618,N_12677);
or U12945 (N_12945,N_12751,N_12655);
or U12946 (N_12946,N_12734,N_12746);
nand U12947 (N_12947,N_12656,N_12781);
nand U12948 (N_12948,N_12736,N_12641);
xor U12949 (N_12949,N_12691,N_12741);
or U12950 (N_12950,N_12751,N_12604);
xor U12951 (N_12951,N_12605,N_12644);
xnor U12952 (N_12952,N_12635,N_12733);
or U12953 (N_12953,N_12785,N_12793);
or U12954 (N_12954,N_12774,N_12695);
xor U12955 (N_12955,N_12659,N_12607);
nand U12956 (N_12956,N_12746,N_12695);
xor U12957 (N_12957,N_12668,N_12605);
xnor U12958 (N_12958,N_12602,N_12711);
or U12959 (N_12959,N_12771,N_12688);
and U12960 (N_12960,N_12720,N_12617);
and U12961 (N_12961,N_12641,N_12698);
and U12962 (N_12962,N_12774,N_12777);
nor U12963 (N_12963,N_12686,N_12609);
or U12964 (N_12964,N_12716,N_12643);
nor U12965 (N_12965,N_12711,N_12609);
or U12966 (N_12966,N_12626,N_12797);
nor U12967 (N_12967,N_12682,N_12728);
and U12968 (N_12968,N_12633,N_12724);
xnor U12969 (N_12969,N_12684,N_12790);
or U12970 (N_12970,N_12683,N_12792);
nor U12971 (N_12971,N_12743,N_12769);
nand U12972 (N_12972,N_12684,N_12741);
nor U12973 (N_12973,N_12612,N_12753);
or U12974 (N_12974,N_12635,N_12628);
nor U12975 (N_12975,N_12699,N_12739);
nor U12976 (N_12976,N_12647,N_12720);
or U12977 (N_12977,N_12600,N_12733);
or U12978 (N_12978,N_12642,N_12731);
xor U12979 (N_12979,N_12764,N_12619);
and U12980 (N_12980,N_12642,N_12646);
or U12981 (N_12981,N_12648,N_12772);
and U12982 (N_12982,N_12709,N_12663);
nand U12983 (N_12983,N_12791,N_12696);
or U12984 (N_12984,N_12795,N_12690);
and U12985 (N_12985,N_12618,N_12743);
nand U12986 (N_12986,N_12682,N_12625);
nand U12987 (N_12987,N_12737,N_12693);
and U12988 (N_12988,N_12747,N_12788);
and U12989 (N_12989,N_12653,N_12745);
nand U12990 (N_12990,N_12643,N_12729);
nand U12991 (N_12991,N_12634,N_12798);
and U12992 (N_12992,N_12789,N_12601);
and U12993 (N_12993,N_12695,N_12762);
and U12994 (N_12994,N_12683,N_12743);
xnor U12995 (N_12995,N_12674,N_12606);
and U12996 (N_12996,N_12763,N_12701);
and U12997 (N_12997,N_12646,N_12602);
xnor U12998 (N_12998,N_12703,N_12783);
and U12999 (N_12999,N_12656,N_12771);
nor U13000 (N_13000,N_12996,N_12979);
nand U13001 (N_13001,N_12973,N_12892);
nand U13002 (N_13002,N_12843,N_12874);
and U13003 (N_13003,N_12806,N_12923);
nand U13004 (N_13004,N_12981,N_12903);
nor U13005 (N_13005,N_12814,N_12894);
xnor U13006 (N_13006,N_12830,N_12891);
and U13007 (N_13007,N_12847,N_12882);
nand U13008 (N_13008,N_12873,N_12944);
nand U13009 (N_13009,N_12869,N_12964);
nand U13010 (N_13010,N_12933,N_12952);
nand U13011 (N_13011,N_12857,N_12934);
xor U13012 (N_13012,N_12957,N_12966);
xor U13013 (N_13013,N_12938,N_12921);
xnor U13014 (N_13014,N_12901,N_12904);
or U13015 (N_13015,N_12831,N_12883);
and U13016 (N_13016,N_12899,N_12852);
or U13017 (N_13017,N_12870,N_12970);
nor U13018 (N_13018,N_12809,N_12963);
or U13019 (N_13019,N_12922,N_12821);
nand U13020 (N_13020,N_12936,N_12817);
or U13021 (N_13021,N_12910,N_12994);
or U13022 (N_13022,N_12884,N_12879);
nor U13023 (N_13023,N_12807,N_12856);
xnor U13024 (N_13024,N_12916,N_12895);
and U13025 (N_13025,N_12976,N_12949);
nand U13026 (N_13026,N_12876,N_12991);
nor U13027 (N_13027,N_12829,N_12977);
and U13028 (N_13028,N_12826,N_12907);
nor U13029 (N_13029,N_12917,N_12858);
or U13030 (N_13030,N_12862,N_12837);
nand U13031 (N_13031,N_12941,N_12940);
nor U13032 (N_13032,N_12925,N_12812);
and U13033 (N_13033,N_12834,N_12805);
xor U13034 (N_13034,N_12833,N_12965);
nand U13035 (N_13035,N_12943,N_12848);
nor U13036 (N_13036,N_12959,N_12912);
and U13037 (N_13037,N_12924,N_12804);
nand U13038 (N_13038,N_12971,N_12958);
xnor U13039 (N_13039,N_12995,N_12803);
and U13040 (N_13040,N_12983,N_12926);
or U13041 (N_13041,N_12861,N_12824);
xor U13042 (N_13042,N_12802,N_12900);
nand U13043 (N_13043,N_12859,N_12886);
and U13044 (N_13044,N_12911,N_12986);
nand U13045 (N_13045,N_12931,N_12868);
nor U13046 (N_13046,N_12980,N_12816);
nand U13047 (N_13047,N_12937,N_12819);
nor U13048 (N_13048,N_12953,N_12871);
and U13049 (N_13049,N_12942,N_12841);
nand U13050 (N_13050,N_12881,N_12975);
and U13051 (N_13051,N_12918,N_12999);
nor U13052 (N_13052,N_12855,N_12820);
or U13053 (N_13053,N_12984,N_12989);
nor U13054 (N_13054,N_12932,N_12982);
xor U13055 (N_13055,N_12877,N_12908);
nor U13056 (N_13056,N_12962,N_12838);
or U13057 (N_13057,N_12930,N_12955);
and U13058 (N_13058,N_12846,N_12939);
or U13059 (N_13059,N_12815,N_12961);
or U13060 (N_13060,N_12968,N_12887);
nand U13061 (N_13061,N_12993,N_12823);
nor U13062 (N_13062,N_12990,N_12800);
nand U13063 (N_13063,N_12978,N_12872);
nand U13064 (N_13064,N_12997,N_12951);
nor U13065 (N_13065,N_12842,N_12927);
nor U13066 (N_13066,N_12880,N_12935);
and U13067 (N_13067,N_12810,N_12845);
and U13068 (N_13068,N_12905,N_12913);
nor U13069 (N_13069,N_12888,N_12896);
and U13070 (N_13070,N_12836,N_12818);
and U13071 (N_13071,N_12906,N_12956);
xnor U13072 (N_13072,N_12853,N_12960);
nand U13073 (N_13073,N_12844,N_12969);
xor U13074 (N_13074,N_12813,N_12985);
nor U13075 (N_13075,N_12919,N_12864);
xnor U13076 (N_13076,N_12849,N_12992);
and U13077 (N_13077,N_12839,N_12875);
or U13078 (N_13078,N_12878,N_12832);
xnor U13079 (N_13079,N_12885,N_12974);
or U13080 (N_13080,N_12835,N_12801);
and U13081 (N_13081,N_12929,N_12948);
and U13082 (N_13082,N_12988,N_12822);
nand U13083 (N_13083,N_12998,N_12914);
nand U13084 (N_13084,N_12850,N_12897);
and U13085 (N_13085,N_12854,N_12946);
nor U13086 (N_13086,N_12928,N_12860);
nor U13087 (N_13087,N_12828,N_12865);
nand U13088 (N_13088,N_12954,N_12890);
and U13089 (N_13089,N_12863,N_12967);
and U13090 (N_13090,N_12866,N_12827);
or U13091 (N_13091,N_12898,N_12972);
or U13092 (N_13092,N_12893,N_12915);
or U13093 (N_13093,N_12811,N_12867);
or U13094 (N_13094,N_12909,N_12851);
nand U13095 (N_13095,N_12825,N_12920);
nand U13096 (N_13096,N_12947,N_12808);
nand U13097 (N_13097,N_12945,N_12902);
and U13098 (N_13098,N_12950,N_12987);
xor U13099 (N_13099,N_12889,N_12840);
nor U13100 (N_13100,N_12806,N_12839);
and U13101 (N_13101,N_12948,N_12981);
or U13102 (N_13102,N_12878,N_12884);
nand U13103 (N_13103,N_12914,N_12835);
or U13104 (N_13104,N_12912,N_12824);
nor U13105 (N_13105,N_12897,N_12843);
or U13106 (N_13106,N_12937,N_12924);
or U13107 (N_13107,N_12976,N_12943);
or U13108 (N_13108,N_12904,N_12849);
nand U13109 (N_13109,N_12932,N_12827);
nor U13110 (N_13110,N_12824,N_12886);
and U13111 (N_13111,N_12831,N_12904);
or U13112 (N_13112,N_12907,N_12878);
nand U13113 (N_13113,N_12993,N_12982);
or U13114 (N_13114,N_12804,N_12906);
and U13115 (N_13115,N_12889,N_12957);
nor U13116 (N_13116,N_12926,N_12978);
xnor U13117 (N_13117,N_12879,N_12926);
nand U13118 (N_13118,N_12878,N_12929);
and U13119 (N_13119,N_12894,N_12979);
xor U13120 (N_13120,N_12926,N_12959);
nor U13121 (N_13121,N_12974,N_12957);
and U13122 (N_13122,N_12866,N_12962);
and U13123 (N_13123,N_12998,N_12848);
and U13124 (N_13124,N_12841,N_12886);
and U13125 (N_13125,N_12999,N_12899);
xnor U13126 (N_13126,N_12809,N_12824);
nor U13127 (N_13127,N_12957,N_12824);
xor U13128 (N_13128,N_12935,N_12825);
nor U13129 (N_13129,N_12891,N_12922);
nor U13130 (N_13130,N_12914,N_12905);
xnor U13131 (N_13131,N_12833,N_12852);
nand U13132 (N_13132,N_12946,N_12990);
xor U13133 (N_13133,N_12904,N_12994);
or U13134 (N_13134,N_12911,N_12976);
or U13135 (N_13135,N_12804,N_12999);
or U13136 (N_13136,N_12935,N_12955);
xor U13137 (N_13137,N_12868,N_12946);
and U13138 (N_13138,N_12858,N_12971);
or U13139 (N_13139,N_12982,N_12943);
nor U13140 (N_13140,N_12915,N_12897);
xnor U13141 (N_13141,N_12827,N_12876);
xor U13142 (N_13142,N_12833,N_12988);
nor U13143 (N_13143,N_12838,N_12970);
xnor U13144 (N_13144,N_12910,N_12871);
or U13145 (N_13145,N_12982,N_12969);
xnor U13146 (N_13146,N_12914,N_12869);
xnor U13147 (N_13147,N_12899,N_12878);
or U13148 (N_13148,N_12824,N_12999);
nand U13149 (N_13149,N_12837,N_12989);
and U13150 (N_13150,N_12810,N_12963);
xor U13151 (N_13151,N_12870,N_12899);
xnor U13152 (N_13152,N_12953,N_12885);
nand U13153 (N_13153,N_12817,N_12861);
xnor U13154 (N_13154,N_12930,N_12934);
xor U13155 (N_13155,N_12954,N_12869);
and U13156 (N_13156,N_12974,N_12855);
and U13157 (N_13157,N_12889,N_12973);
xnor U13158 (N_13158,N_12999,N_12965);
nor U13159 (N_13159,N_12856,N_12936);
nor U13160 (N_13160,N_12827,N_12893);
or U13161 (N_13161,N_12833,N_12944);
and U13162 (N_13162,N_12957,N_12953);
nand U13163 (N_13163,N_12925,N_12900);
and U13164 (N_13164,N_12941,N_12890);
or U13165 (N_13165,N_12967,N_12893);
nor U13166 (N_13166,N_12976,N_12895);
or U13167 (N_13167,N_12988,N_12831);
xnor U13168 (N_13168,N_12941,N_12959);
or U13169 (N_13169,N_12983,N_12930);
and U13170 (N_13170,N_12832,N_12870);
and U13171 (N_13171,N_12808,N_12869);
nor U13172 (N_13172,N_12830,N_12842);
and U13173 (N_13173,N_12939,N_12809);
xor U13174 (N_13174,N_12835,N_12880);
nor U13175 (N_13175,N_12949,N_12900);
and U13176 (N_13176,N_12853,N_12983);
nor U13177 (N_13177,N_12931,N_12839);
nand U13178 (N_13178,N_12980,N_12943);
and U13179 (N_13179,N_12840,N_12843);
xnor U13180 (N_13180,N_12984,N_12950);
nor U13181 (N_13181,N_12986,N_12834);
xnor U13182 (N_13182,N_12808,N_12816);
nand U13183 (N_13183,N_12827,N_12879);
nand U13184 (N_13184,N_12846,N_12956);
xnor U13185 (N_13185,N_12837,N_12971);
xor U13186 (N_13186,N_12913,N_12898);
nor U13187 (N_13187,N_12964,N_12971);
nand U13188 (N_13188,N_12993,N_12950);
xor U13189 (N_13189,N_12811,N_12923);
xor U13190 (N_13190,N_12893,N_12985);
nor U13191 (N_13191,N_12958,N_12936);
or U13192 (N_13192,N_12907,N_12917);
nand U13193 (N_13193,N_12938,N_12959);
and U13194 (N_13194,N_12904,N_12814);
nor U13195 (N_13195,N_12857,N_12973);
and U13196 (N_13196,N_12860,N_12986);
and U13197 (N_13197,N_12993,N_12807);
or U13198 (N_13198,N_12909,N_12913);
and U13199 (N_13199,N_12937,N_12958);
xnor U13200 (N_13200,N_13128,N_13056);
or U13201 (N_13201,N_13002,N_13024);
xor U13202 (N_13202,N_13155,N_13110);
nand U13203 (N_13203,N_13034,N_13019);
xnor U13204 (N_13204,N_13158,N_13187);
xor U13205 (N_13205,N_13008,N_13177);
xor U13206 (N_13206,N_13072,N_13058);
and U13207 (N_13207,N_13188,N_13036);
nand U13208 (N_13208,N_13140,N_13012);
nor U13209 (N_13209,N_13091,N_13075);
nand U13210 (N_13210,N_13020,N_13013);
xor U13211 (N_13211,N_13004,N_13147);
or U13212 (N_13212,N_13193,N_13044);
or U13213 (N_13213,N_13164,N_13195);
xor U13214 (N_13214,N_13030,N_13102);
xnor U13215 (N_13215,N_13171,N_13098);
and U13216 (N_13216,N_13074,N_13080);
xor U13217 (N_13217,N_13194,N_13041);
nor U13218 (N_13218,N_13060,N_13111);
xor U13219 (N_13219,N_13197,N_13000);
nand U13220 (N_13220,N_13124,N_13154);
nor U13221 (N_13221,N_13067,N_13149);
nor U13222 (N_13222,N_13152,N_13189);
xnor U13223 (N_13223,N_13133,N_13170);
xnor U13224 (N_13224,N_13048,N_13150);
xnor U13225 (N_13225,N_13011,N_13105);
xor U13226 (N_13226,N_13025,N_13139);
and U13227 (N_13227,N_13120,N_13001);
or U13228 (N_13228,N_13179,N_13096);
and U13229 (N_13229,N_13010,N_13039);
and U13230 (N_13230,N_13038,N_13161);
xor U13231 (N_13231,N_13190,N_13042);
and U13232 (N_13232,N_13089,N_13163);
xor U13233 (N_13233,N_13172,N_13126);
or U13234 (N_13234,N_13085,N_13132);
xor U13235 (N_13235,N_13148,N_13095);
nand U13236 (N_13236,N_13077,N_13043);
nand U13237 (N_13237,N_13135,N_13178);
and U13238 (N_13238,N_13099,N_13127);
or U13239 (N_13239,N_13090,N_13183);
nand U13240 (N_13240,N_13159,N_13017);
nor U13241 (N_13241,N_13081,N_13097);
nor U13242 (N_13242,N_13104,N_13108);
xnor U13243 (N_13243,N_13100,N_13141);
nand U13244 (N_13244,N_13144,N_13125);
xor U13245 (N_13245,N_13173,N_13066);
nor U13246 (N_13246,N_13070,N_13050);
nand U13247 (N_13247,N_13079,N_13006);
or U13248 (N_13248,N_13143,N_13018);
or U13249 (N_13249,N_13026,N_13063);
or U13250 (N_13250,N_13047,N_13109);
or U13251 (N_13251,N_13113,N_13134);
nand U13252 (N_13252,N_13093,N_13055);
xnor U13253 (N_13253,N_13033,N_13022);
xor U13254 (N_13254,N_13137,N_13051);
or U13255 (N_13255,N_13136,N_13029);
and U13256 (N_13256,N_13116,N_13174);
nand U13257 (N_13257,N_13054,N_13015);
nor U13258 (N_13258,N_13009,N_13088);
nand U13259 (N_13259,N_13035,N_13166);
nor U13260 (N_13260,N_13073,N_13086);
nand U13261 (N_13261,N_13068,N_13049);
nor U13262 (N_13262,N_13057,N_13021);
or U13263 (N_13263,N_13061,N_13181);
xor U13264 (N_13264,N_13146,N_13175);
or U13265 (N_13265,N_13032,N_13052);
nand U13266 (N_13266,N_13167,N_13145);
nor U13267 (N_13267,N_13083,N_13092);
nor U13268 (N_13268,N_13185,N_13082);
or U13269 (N_13269,N_13084,N_13053);
nand U13270 (N_13270,N_13037,N_13059);
nand U13271 (N_13271,N_13115,N_13065);
or U13272 (N_13272,N_13003,N_13028);
nor U13273 (N_13273,N_13005,N_13192);
nor U13274 (N_13274,N_13101,N_13112);
nand U13275 (N_13275,N_13165,N_13156);
xnor U13276 (N_13276,N_13023,N_13117);
and U13277 (N_13277,N_13076,N_13196);
xor U13278 (N_13278,N_13031,N_13180);
nand U13279 (N_13279,N_13176,N_13198);
and U13280 (N_13280,N_13118,N_13062);
nand U13281 (N_13281,N_13071,N_13182);
xor U13282 (N_13282,N_13186,N_13119);
nor U13283 (N_13283,N_13040,N_13069);
xor U13284 (N_13284,N_13016,N_13064);
and U13285 (N_13285,N_13138,N_13087);
and U13286 (N_13286,N_13162,N_13131);
nor U13287 (N_13287,N_13122,N_13151);
or U13288 (N_13288,N_13107,N_13106);
xor U13289 (N_13289,N_13129,N_13094);
or U13290 (N_13290,N_13160,N_13123);
and U13291 (N_13291,N_13121,N_13157);
or U13292 (N_13292,N_13130,N_13169);
or U13293 (N_13293,N_13103,N_13007);
nand U13294 (N_13294,N_13184,N_13142);
nor U13295 (N_13295,N_13014,N_13045);
and U13296 (N_13296,N_13027,N_13078);
and U13297 (N_13297,N_13168,N_13199);
nand U13298 (N_13298,N_13046,N_13153);
or U13299 (N_13299,N_13191,N_13114);
or U13300 (N_13300,N_13047,N_13086);
nor U13301 (N_13301,N_13050,N_13030);
xnor U13302 (N_13302,N_13078,N_13050);
xor U13303 (N_13303,N_13122,N_13148);
and U13304 (N_13304,N_13177,N_13187);
or U13305 (N_13305,N_13175,N_13163);
nor U13306 (N_13306,N_13131,N_13028);
nand U13307 (N_13307,N_13079,N_13014);
or U13308 (N_13308,N_13186,N_13098);
xnor U13309 (N_13309,N_13109,N_13092);
or U13310 (N_13310,N_13009,N_13044);
nand U13311 (N_13311,N_13036,N_13068);
or U13312 (N_13312,N_13145,N_13009);
and U13313 (N_13313,N_13003,N_13125);
or U13314 (N_13314,N_13030,N_13046);
nor U13315 (N_13315,N_13067,N_13161);
or U13316 (N_13316,N_13186,N_13061);
xnor U13317 (N_13317,N_13067,N_13052);
nor U13318 (N_13318,N_13166,N_13125);
nand U13319 (N_13319,N_13005,N_13140);
and U13320 (N_13320,N_13085,N_13028);
or U13321 (N_13321,N_13046,N_13112);
and U13322 (N_13322,N_13174,N_13123);
nor U13323 (N_13323,N_13087,N_13102);
or U13324 (N_13324,N_13015,N_13138);
nor U13325 (N_13325,N_13125,N_13088);
xnor U13326 (N_13326,N_13141,N_13103);
nand U13327 (N_13327,N_13070,N_13037);
xnor U13328 (N_13328,N_13059,N_13018);
or U13329 (N_13329,N_13066,N_13135);
nand U13330 (N_13330,N_13180,N_13046);
nor U13331 (N_13331,N_13035,N_13061);
xnor U13332 (N_13332,N_13060,N_13183);
nor U13333 (N_13333,N_13121,N_13112);
nand U13334 (N_13334,N_13111,N_13044);
nand U13335 (N_13335,N_13100,N_13073);
nor U13336 (N_13336,N_13017,N_13054);
xnor U13337 (N_13337,N_13071,N_13198);
nor U13338 (N_13338,N_13100,N_13024);
or U13339 (N_13339,N_13127,N_13110);
xnor U13340 (N_13340,N_13124,N_13032);
xnor U13341 (N_13341,N_13021,N_13138);
nand U13342 (N_13342,N_13140,N_13162);
or U13343 (N_13343,N_13188,N_13199);
nor U13344 (N_13344,N_13175,N_13176);
xor U13345 (N_13345,N_13028,N_13053);
and U13346 (N_13346,N_13054,N_13072);
nor U13347 (N_13347,N_13118,N_13056);
xor U13348 (N_13348,N_13005,N_13048);
nand U13349 (N_13349,N_13167,N_13184);
xor U13350 (N_13350,N_13092,N_13015);
or U13351 (N_13351,N_13171,N_13032);
nand U13352 (N_13352,N_13056,N_13187);
and U13353 (N_13353,N_13000,N_13164);
nand U13354 (N_13354,N_13122,N_13104);
or U13355 (N_13355,N_13012,N_13113);
nor U13356 (N_13356,N_13029,N_13160);
and U13357 (N_13357,N_13003,N_13032);
and U13358 (N_13358,N_13084,N_13021);
xnor U13359 (N_13359,N_13173,N_13197);
nand U13360 (N_13360,N_13055,N_13104);
nor U13361 (N_13361,N_13149,N_13090);
or U13362 (N_13362,N_13037,N_13092);
nand U13363 (N_13363,N_13158,N_13020);
nor U13364 (N_13364,N_13028,N_13038);
xor U13365 (N_13365,N_13003,N_13167);
and U13366 (N_13366,N_13185,N_13085);
xnor U13367 (N_13367,N_13074,N_13156);
xnor U13368 (N_13368,N_13063,N_13199);
and U13369 (N_13369,N_13027,N_13116);
and U13370 (N_13370,N_13141,N_13073);
nor U13371 (N_13371,N_13098,N_13044);
nor U13372 (N_13372,N_13198,N_13078);
and U13373 (N_13373,N_13017,N_13021);
nor U13374 (N_13374,N_13172,N_13041);
nand U13375 (N_13375,N_13051,N_13036);
or U13376 (N_13376,N_13142,N_13124);
xor U13377 (N_13377,N_13096,N_13178);
or U13378 (N_13378,N_13052,N_13114);
or U13379 (N_13379,N_13127,N_13010);
nand U13380 (N_13380,N_13008,N_13084);
or U13381 (N_13381,N_13058,N_13029);
nand U13382 (N_13382,N_13154,N_13046);
nand U13383 (N_13383,N_13186,N_13165);
or U13384 (N_13384,N_13158,N_13176);
nand U13385 (N_13385,N_13124,N_13049);
xnor U13386 (N_13386,N_13050,N_13003);
nand U13387 (N_13387,N_13127,N_13138);
and U13388 (N_13388,N_13112,N_13162);
xnor U13389 (N_13389,N_13115,N_13035);
nor U13390 (N_13390,N_13192,N_13178);
xnor U13391 (N_13391,N_13063,N_13183);
xnor U13392 (N_13392,N_13054,N_13074);
nor U13393 (N_13393,N_13019,N_13063);
nor U13394 (N_13394,N_13151,N_13038);
or U13395 (N_13395,N_13090,N_13085);
or U13396 (N_13396,N_13001,N_13040);
and U13397 (N_13397,N_13159,N_13092);
nor U13398 (N_13398,N_13172,N_13076);
and U13399 (N_13399,N_13088,N_13117);
xnor U13400 (N_13400,N_13213,N_13303);
nor U13401 (N_13401,N_13211,N_13339);
and U13402 (N_13402,N_13289,N_13228);
nor U13403 (N_13403,N_13369,N_13234);
or U13404 (N_13404,N_13370,N_13373);
nor U13405 (N_13405,N_13313,N_13237);
nor U13406 (N_13406,N_13280,N_13361);
xnor U13407 (N_13407,N_13271,N_13322);
nand U13408 (N_13408,N_13372,N_13267);
nand U13409 (N_13409,N_13225,N_13387);
and U13410 (N_13410,N_13226,N_13341);
xor U13411 (N_13411,N_13252,N_13342);
nand U13412 (N_13412,N_13246,N_13319);
or U13413 (N_13413,N_13284,N_13354);
or U13414 (N_13414,N_13308,N_13345);
or U13415 (N_13415,N_13212,N_13388);
xor U13416 (N_13416,N_13269,N_13318);
nor U13417 (N_13417,N_13328,N_13258);
nand U13418 (N_13418,N_13360,N_13310);
xor U13419 (N_13419,N_13382,N_13241);
nand U13420 (N_13420,N_13242,N_13386);
xor U13421 (N_13421,N_13222,N_13392);
or U13422 (N_13422,N_13371,N_13279);
xor U13423 (N_13423,N_13300,N_13298);
and U13424 (N_13424,N_13223,N_13283);
and U13425 (N_13425,N_13330,N_13287);
and U13426 (N_13426,N_13274,N_13380);
nand U13427 (N_13427,N_13314,N_13262);
or U13428 (N_13428,N_13253,N_13260);
xor U13429 (N_13429,N_13264,N_13357);
or U13430 (N_13430,N_13320,N_13288);
or U13431 (N_13431,N_13209,N_13385);
and U13432 (N_13432,N_13323,N_13396);
nor U13433 (N_13433,N_13272,N_13340);
and U13434 (N_13434,N_13285,N_13315);
nand U13435 (N_13435,N_13239,N_13210);
nand U13436 (N_13436,N_13335,N_13363);
nand U13437 (N_13437,N_13362,N_13333);
and U13438 (N_13438,N_13336,N_13214);
xnor U13439 (N_13439,N_13378,N_13230);
xor U13440 (N_13440,N_13312,N_13374);
or U13441 (N_13441,N_13397,N_13309);
nand U13442 (N_13442,N_13364,N_13376);
xor U13443 (N_13443,N_13233,N_13200);
xnor U13444 (N_13444,N_13275,N_13299);
xnor U13445 (N_13445,N_13276,N_13250);
nand U13446 (N_13446,N_13384,N_13297);
nor U13447 (N_13447,N_13270,N_13296);
nor U13448 (N_13448,N_13295,N_13366);
or U13449 (N_13449,N_13316,N_13311);
nor U13450 (N_13450,N_13394,N_13218);
nor U13451 (N_13451,N_13367,N_13398);
and U13452 (N_13452,N_13329,N_13273);
or U13453 (N_13453,N_13326,N_13265);
nand U13454 (N_13454,N_13334,N_13205);
xnor U13455 (N_13455,N_13352,N_13263);
nor U13456 (N_13456,N_13338,N_13245);
or U13457 (N_13457,N_13231,N_13207);
or U13458 (N_13458,N_13247,N_13224);
nor U13459 (N_13459,N_13324,N_13390);
nor U13460 (N_13460,N_13327,N_13236);
nor U13461 (N_13461,N_13266,N_13305);
nand U13462 (N_13462,N_13220,N_13393);
xnor U13463 (N_13463,N_13377,N_13355);
or U13464 (N_13464,N_13348,N_13346);
and U13465 (N_13465,N_13259,N_13255);
or U13466 (N_13466,N_13399,N_13395);
xnor U13467 (N_13467,N_13302,N_13290);
or U13468 (N_13468,N_13240,N_13347);
xor U13469 (N_13469,N_13249,N_13317);
xnor U13470 (N_13470,N_13381,N_13254);
or U13471 (N_13471,N_13344,N_13203);
nor U13472 (N_13472,N_13359,N_13391);
or U13473 (N_13473,N_13217,N_13221);
or U13474 (N_13474,N_13286,N_13235);
xnor U13475 (N_13475,N_13208,N_13204);
xor U13476 (N_13476,N_13292,N_13215);
nand U13477 (N_13477,N_13257,N_13202);
nor U13478 (N_13478,N_13293,N_13229);
or U13479 (N_13479,N_13201,N_13206);
and U13480 (N_13480,N_13278,N_13268);
or U13481 (N_13481,N_13389,N_13227);
nand U13482 (N_13482,N_13349,N_13243);
and U13483 (N_13483,N_13219,N_13251);
nand U13484 (N_13484,N_13281,N_13238);
or U13485 (N_13485,N_13232,N_13256);
xnor U13486 (N_13486,N_13248,N_13216);
and U13487 (N_13487,N_13307,N_13301);
or U13488 (N_13488,N_13337,N_13379);
nor U13489 (N_13489,N_13351,N_13294);
nor U13490 (N_13490,N_13277,N_13282);
nand U13491 (N_13491,N_13306,N_13356);
nor U13492 (N_13492,N_13331,N_13343);
or U13493 (N_13493,N_13304,N_13375);
nor U13494 (N_13494,N_13321,N_13358);
and U13495 (N_13495,N_13350,N_13291);
xnor U13496 (N_13496,N_13365,N_13332);
or U13497 (N_13497,N_13261,N_13325);
and U13498 (N_13498,N_13353,N_13244);
or U13499 (N_13499,N_13368,N_13383);
nor U13500 (N_13500,N_13365,N_13366);
xnor U13501 (N_13501,N_13309,N_13349);
nand U13502 (N_13502,N_13340,N_13269);
or U13503 (N_13503,N_13232,N_13322);
and U13504 (N_13504,N_13322,N_13233);
nand U13505 (N_13505,N_13258,N_13214);
nand U13506 (N_13506,N_13354,N_13235);
and U13507 (N_13507,N_13222,N_13325);
and U13508 (N_13508,N_13389,N_13226);
nor U13509 (N_13509,N_13325,N_13233);
nand U13510 (N_13510,N_13337,N_13345);
nor U13511 (N_13511,N_13357,N_13247);
nand U13512 (N_13512,N_13236,N_13349);
nand U13513 (N_13513,N_13279,N_13392);
xor U13514 (N_13514,N_13376,N_13359);
xor U13515 (N_13515,N_13272,N_13223);
and U13516 (N_13516,N_13388,N_13286);
and U13517 (N_13517,N_13356,N_13277);
nand U13518 (N_13518,N_13346,N_13354);
or U13519 (N_13519,N_13227,N_13249);
and U13520 (N_13520,N_13329,N_13353);
and U13521 (N_13521,N_13326,N_13313);
xor U13522 (N_13522,N_13328,N_13206);
or U13523 (N_13523,N_13257,N_13208);
xnor U13524 (N_13524,N_13393,N_13353);
and U13525 (N_13525,N_13249,N_13292);
nor U13526 (N_13526,N_13222,N_13358);
xor U13527 (N_13527,N_13239,N_13217);
or U13528 (N_13528,N_13330,N_13260);
nor U13529 (N_13529,N_13217,N_13399);
nor U13530 (N_13530,N_13270,N_13223);
or U13531 (N_13531,N_13384,N_13201);
or U13532 (N_13532,N_13314,N_13382);
or U13533 (N_13533,N_13230,N_13306);
nor U13534 (N_13534,N_13303,N_13306);
or U13535 (N_13535,N_13312,N_13321);
or U13536 (N_13536,N_13225,N_13314);
nor U13537 (N_13537,N_13213,N_13334);
nor U13538 (N_13538,N_13346,N_13356);
nor U13539 (N_13539,N_13281,N_13262);
nand U13540 (N_13540,N_13211,N_13363);
or U13541 (N_13541,N_13359,N_13369);
nand U13542 (N_13542,N_13261,N_13368);
xnor U13543 (N_13543,N_13231,N_13339);
and U13544 (N_13544,N_13331,N_13235);
nor U13545 (N_13545,N_13386,N_13230);
xnor U13546 (N_13546,N_13300,N_13295);
xnor U13547 (N_13547,N_13308,N_13279);
and U13548 (N_13548,N_13384,N_13320);
xnor U13549 (N_13549,N_13256,N_13226);
or U13550 (N_13550,N_13278,N_13293);
nand U13551 (N_13551,N_13360,N_13227);
nor U13552 (N_13552,N_13221,N_13375);
nand U13553 (N_13553,N_13342,N_13273);
xor U13554 (N_13554,N_13381,N_13253);
nand U13555 (N_13555,N_13342,N_13264);
xor U13556 (N_13556,N_13252,N_13367);
and U13557 (N_13557,N_13349,N_13328);
nand U13558 (N_13558,N_13343,N_13202);
and U13559 (N_13559,N_13346,N_13255);
nand U13560 (N_13560,N_13217,N_13259);
or U13561 (N_13561,N_13252,N_13388);
or U13562 (N_13562,N_13319,N_13320);
or U13563 (N_13563,N_13299,N_13220);
xor U13564 (N_13564,N_13215,N_13350);
or U13565 (N_13565,N_13371,N_13331);
xor U13566 (N_13566,N_13213,N_13263);
nor U13567 (N_13567,N_13201,N_13276);
or U13568 (N_13568,N_13238,N_13245);
and U13569 (N_13569,N_13269,N_13293);
or U13570 (N_13570,N_13293,N_13366);
or U13571 (N_13571,N_13381,N_13284);
and U13572 (N_13572,N_13374,N_13392);
xnor U13573 (N_13573,N_13258,N_13329);
and U13574 (N_13574,N_13378,N_13329);
nand U13575 (N_13575,N_13259,N_13278);
or U13576 (N_13576,N_13399,N_13226);
and U13577 (N_13577,N_13237,N_13371);
or U13578 (N_13578,N_13391,N_13216);
and U13579 (N_13579,N_13290,N_13353);
nor U13580 (N_13580,N_13304,N_13201);
nor U13581 (N_13581,N_13269,N_13317);
or U13582 (N_13582,N_13331,N_13261);
xnor U13583 (N_13583,N_13297,N_13332);
and U13584 (N_13584,N_13373,N_13302);
nand U13585 (N_13585,N_13275,N_13399);
and U13586 (N_13586,N_13230,N_13215);
xor U13587 (N_13587,N_13398,N_13255);
xnor U13588 (N_13588,N_13399,N_13381);
and U13589 (N_13589,N_13383,N_13239);
and U13590 (N_13590,N_13284,N_13261);
and U13591 (N_13591,N_13267,N_13310);
nand U13592 (N_13592,N_13242,N_13306);
nand U13593 (N_13593,N_13241,N_13340);
nand U13594 (N_13594,N_13265,N_13267);
or U13595 (N_13595,N_13395,N_13267);
nor U13596 (N_13596,N_13383,N_13212);
nand U13597 (N_13597,N_13269,N_13368);
and U13598 (N_13598,N_13326,N_13271);
nor U13599 (N_13599,N_13389,N_13222);
and U13600 (N_13600,N_13490,N_13568);
or U13601 (N_13601,N_13412,N_13459);
or U13602 (N_13602,N_13580,N_13483);
or U13603 (N_13603,N_13509,N_13588);
xor U13604 (N_13604,N_13403,N_13503);
xnor U13605 (N_13605,N_13501,N_13504);
nor U13606 (N_13606,N_13423,N_13482);
and U13607 (N_13607,N_13564,N_13439);
or U13608 (N_13608,N_13582,N_13426);
or U13609 (N_13609,N_13430,N_13530);
and U13610 (N_13610,N_13484,N_13432);
xnor U13611 (N_13611,N_13425,N_13409);
xor U13612 (N_13612,N_13587,N_13595);
nor U13613 (N_13613,N_13452,N_13579);
nor U13614 (N_13614,N_13488,N_13494);
and U13615 (N_13615,N_13524,N_13446);
nand U13616 (N_13616,N_13523,N_13518);
xnor U13617 (N_13617,N_13447,N_13497);
nor U13618 (N_13618,N_13450,N_13596);
xnor U13619 (N_13619,N_13591,N_13529);
xnor U13620 (N_13620,N_13462,N_13475);
and U13621 (N_13621,N_13406,N_13440);
nor U13622 (N_13622,N_13480,N_13542);
xor U13623 (N_13623,N_13516,N_13577);
or U13624 (N_13624,N_13508,N_13521);
and U13625 (N_13625,N_13525,N_13566);
xor U13626 (N_13626,N_13526,N_13572);
or U13627 (N_13627,N_13513,N_13506);
or U13628 (N_13628,N_13431,N_13578);
or U13629 (N_13629,N_13520,N_13517);
and U13630 (N_13630,N_13505,N_13556);
or U13631 (N_13631,N_13586,N_13411);
or U13632 (N_13632,N_13463,N_13427);
nand U13633 (N_13633,N_13408,N_13472);
nand U13634 (N_13634,N_13454,N_13569);
and U13635 (N_13635,N_13522,N_13418);
or U13636 (N_13636,N_13428,N_13435);
nor U13637 (N_13637,N_13548,N_13553);
or U13638 (N_13638,N_13543,N_13419);
nor U13639 (N_13639,N_13562,N_13599);
nand U13640 (N_13640,N_13594,N_13443);
nand U13641 (N_13641,N_13555,N_13434);
nand U13642 (N_13642,N_13511,N_13507);
and U13643 (N_13643,N_13550,N_13417);
and U13644 (N_13644,N_13597,N_13545);
and U13645 (N_13645,N_13536,N_13585);
and U13646 (N_13646,N_13534,N_13519);
xnor U13647 (N_13647,N_13539,N_13470);
nor U13648 (N_13648,N_13541,N_13433);
nor U13649 (N_13649,N_13436,N_13478);
or U13650 (N_13650,N_13422,N_13567);
nor U13651 (N_13651,N_13554,N_13481);
or U13652 (N_13652,N_13404,N_13438);
xor U13653 (N_13653,N_13547,N_13400);
xnor U13654 (N_13654,N_13451,N_13474);
nor U13655 (N_13655,N_13448,N_13584);
and U13656 (N_13656,N_13551,N_13535);
and U13657 (N_13657,N_13464,N_13532);
xnor U13658 (N_13658,N_13498,N_13540);
xor U13659 (N_13659,N_13460,N_13544);
and U13660 (N_13660,N_13489,N_13456);
or U13661 (N_13661,N_13495,N_13453);
or U13662 (N_13662,N_13528,N_13563);
nand U13663 (N_13663,N_13473,N_13437);
xor U13664 (N_13664,N_13449,N_13590);
nor U13665 (N_13665,N_13466,N_13560);
or U13666 (N_13666,N_13557,N_13510);
xor U13667 (N_13667,N_13561,N_13429);
and U13668 (N_13668,N_13515,N_13420);
and U13669 (N_13669,N_13598,N_13424);
xor U13670 (N_13670,N_13558,N_13533);
or U13671 (N_13671,N_13575,N_13413);
and U13672 (N_13672,N_13537,N_13538);
or U13673 (N_13673,N_13559,N_13500);
nand U13674 (N_13674,N_13491,N_13589);
nand U13675 (N_13675,N_13476,N_13583);
and U13676 (N_13676,N_13574,N_13461);
nor U13677 (N_13677,N_13487,N_13421);
xor U13678 (N_13678,N_13479,N_13410);
nor U13679 (N_13679,N_13549,N_13405);
xor U13680 (N_13680,N_13416,N_13593);
xor U13681 (N_13681,N_13415,N_13465);
xor U13682 (N_13682,N_13407,N_13546);
xor U13683 (N_13683,N_13441,N_13571);
nand U13684 (N_13684,N_13445,N_13514);
and U13685 (N_13685,N_13502,N_13552);
xor U13686 (N_13686,N_13499,N_13496);
nand U13687 (N_13687,N_13468,N_13565);
nor U13688 (N_13688,N_13486,N_13576);
and U13689 (N_13689,N_13573,N_13471);
or U13690 (N_13690,N_13442,N_13458);
or U13691 (N_13691,N_13414,N_13477);
nor U13692 (N_13692,N_13467,N_13492);
xor U13693 (N_13693,N_13531,N_13444);
or U13694 (N_13694,N_13527,N_13455);
nand U13695 (N_13695,N_13402,N_13581);
nor U13696 (N_13696,N_13457,N_13570);
nor U13697 (N_13697,N_13512,N_13592);
or U13698 (N_13698,N_13485,N_13401);
nor U13699 (N_13699,N_13469,N_13493);
and U13700 (N_13700,N_13517,N_13588);
nand U13701 (N_13701,N_13594,N_13546);
nand U13702 (N_13702,N_13557,N_13465);
xnor U13703 (N_13703,N_13423,N_13428);
and U13704 (N_13704,N_13490,N_13500);
nor U13705 (N_13705,N_13516,N_13502);
and U13706 (N_13706,N_13587,N_13525);
or U13707 (N_13707,N_13508,N_13582);
or U13708 (N_13708,N_13404,N_13502);
xnor U13709 (N_13709,N_13526,N_13433);
xnor U13710 (N_13710,N_13415,N_13414);
xor U13711 (N_13711,N_13428,N_13468);
and U13712 (N_13712,N_13555,N_13512);
nor U13713 (N_13713,N_13530,N_13465);
nor U13714 (N_13714,N_13461,N_13487);
and U13715 (N_13715,N_13502,N_13580);
or U13716 (N_13716,N_13524,N_13476);
nand U13717 (N_13717,N_13557,N_13582);
nand U13718 (N_13718,N_13502,N_13434);
nor U13719 (N_13719,N_13425,N_13548);
xnor U13720 (N_13720,N_13559,N_13435);
nor U13721 (N_13721,N_13419,N_13482);
and U13722 (N_13722,N_13485,N_13503);
nor U13723 (N_13723,N_13583,N_13545);
nand U13724 (N_13724,N_13573,N_13496);
xnor U13725 (N_13725,N_13578,N_13447);
nor U13726 (N_13726,N_13482,N_13518);
and U13727 (N_13727,N_13591,N_13440);
nor U13728 (N_13728,N_13569,N_13490);
nand U13729 (N_13729,N_13500,N_13462);
and U13730 (N_13730,N_13520,N_13400);
or U13731 (N_13731,N_13513,N_13505);
or U13732 (N_13732,N_13530,N_13488);
and U13733 (N_13733,N_13457,N_13436);
xor U13734 (N_13734,N_13571,N_13479);
nor U13735 (N_13735,N_13524,N_13438);
or U13736 (N_13736,N_13519,N_13553);
nor U13737 (N_13737,N_13414,N_13581);
nand U13738 (N_13738,N_13538,N_13474);
nand U13739 (N_13739,N_13415,N_13595);
or U13740 (N_13740,N_13497,N_13502);
nand U13741 (N_13741,N_13500,N_13534);
xnor U13742 (N_13742,N_13406,N_13527);
nor U13743 (N_13743,N_13584,N_13486);
xnor U13744 (N_13744,N_13489,N_13573);
or U13745 (N_13745,N_13488,N_13454);
nand U13746 (N_13746,N_13497,N_13425);
nand U13747 (N_13747,N_13554,N_13556);
or U13748 (N_13748,N_13406,N_13467);
xnor U13749 (N_13749,N_13421,N_13426);
nor U13750 (N_13750,N_13482,N_13407);
and U13751 (N_13751,N_13468,N_13448);
and U13752 (N_13752,N_13492,N_13471);
or U13753 (N_13753,N_13571,N_13492);
nand U13754 (N_13754,N_13459,N_13466);
xor U13755 (N_13755,N_13411,N_13479);
nand U13756 (N_13756,N_13440,N_13472);
xnor U13757 (N_13757,N_13404,N_13537);
nor U13758 (N_13758,N_13552,N_13418);
or U13759 (N_13759,N_13477,N_13568);
nor U13760 (N_13760,N_13586,N_13569);
xnor U13761 (N_13761,N_13511,N_13566);
nand U13762 (N_13762,N_13466,N_13418);
nand U13763 (N_13763,N_13442,N_13559);
nor U13764 (N_13764,N_13592,N_13474);
xnor U13765 (N_13765,N_13438,N_13425);
or U13766 (N_13766,N_13545,N_13487);
xor U13767 (N_13767,N_13487,N_13492);
or U13768 (N_13768,N_13551,N_13566);
nand U13769 (N_13769,N_13430,N_13588);
nor U13770 (N_13770,N_13477,N_13499);
xnor U13771 (N_13771,N_13594,N_13474);
xor U13772 (N_13772,N_13546,N_13571);
nor U13773 (N_13773,N_13516,N_13529);
nand U13774 (N_13774,N_13456,N_13531);
nand U13775 (N_13775,N_13576,N_13521);
or U13776 (N_13776,N_13497,N_13469);
or U13777 (N_13777,N_13446,N_13486);
nand U13778 (N_13778,N_13428,N_13570);
nand U13779 (N_13779,N_13508,N_13437);
or U13780 (N_13780,N_13481,N_13583);
nor U13781 (N_13781,N_13557,N_13596);
xnor U13782 (N_13782,N_13498,N_13595);
or U13783 (N_13783,N_13580,N_13591);
or U13784 (N_13784,N_13422,N_13450);
nand U13785 (N_13785,N_13467,N_13555);
nand U13786 (N_13786,N_13468,N_13576);
nor U13787 (N_13787,N_13528,N_13509);
nor U13788 (N_13788,N_13431,N_13421);
and U13789 (N_13789,N_13418,N_13448);
nand U13790 (N_13790,N_13590,N_13462);
nor U13791 (N_13791,N_13482,N_13562);
or U13792 (N_13792,N_13537,N_13429);
nand U13793 (N_13793,N_13510,N_13453);
or U13794 (N_13794,N_13525,N_13509);
nor U13795 (N_13795,N_13484,N_13508);
xor U13796 (N_13796,N_13543,N_13504);
and U13797 (N_13797,N_13587,N_13428);
and U13798 (N_13798,N_13581,N_13557);
nor U13799 (N_13799,N_13402,N_13444);
or U13800 (N_13800,N_13668,N_13631);
and U13801 (N_13801,N_13669,N_13769);
or U13802 (N_13802,N_13756,N_13762);
or U13803 (N_13803,N_13635,N_13674);
xor U13804 (N_13804,N_13681,N_13745);
xor U13805 (N_13805,N_13725,N_13616);
nand U13806 (N_13806,N_13787,N_13637);
or U13807 (N_13807,N_13751,N_13736);
xor U13808 (N_13808,N_13778,N_13632);
and U13809 (N_13809,N_13663,N_13654);
nor U13810 (N_13810,N_13697,N_13687);
xor U13811 (N_13811,N_13760,N_13780);
or U13812 (N_13812,N_13659,N_13789);
nand U13813 (N_13813,N_13652,N_13673);
xor U13814 (N_13814,N_13757,N_13706);
xor U13815 (N_13815,N_13600,N_13695);
and U13816 (N_13816,N_13624,N_13783);
or U13817 (N_13817,N_13711,N_13726);
and U13818 (N_13818,N_13645,N_13723);
nor U13819 (N_13819,N_13606,N_13660);
and U13820 (N_13820,N_13739,N_13612);
nand U13821 (N_13821,N_13721,N_13773);
and U13822 (N_13822,N_13618,N_13647);
nor U13823 (N_13823,N_13690,N_13639);
and U13824 (N_13824,N_13636,N_13677);
and U13825 (N_13825,N_13771,N_13705);
nor U13826 (N_13826,N_13776,N_13676);
xnor U13827 (N_13827,N_13775,N_13797);
nand U13828 (N_13828,N_13724,N_13621);
nor U13829 (N_13829,N_13692,N_13750);
nor U13830 (N_13830,N_13718,N_13657);
xnor U13831 (N_13831,N_13788,N_13627);
xor U13832 (N_13832,N_13643,N_13719);
xor U13833 (N_13833,N_13613,N_13626);
nor U13834 (N_13834,N_13602,N_13734);
nand U13835 (N_13835,N_13712,N_13717);
nand U13836 (N_13836,N_13671,N_13716);
and U13837 (N_13837,N_13603,N_13672);
nor U13838 (N_13838,N_13714,N_13628);
xnor U13839 (N_13839,N_13753,N_13781);
xor U13840 (N_13840,N_13730,N_13784);
xnor U13841 (N_13841,N_13610,N_13609);
nand U13842 (N_13842,N_13755,N_13766);
nand U13843 (N_13843,N_13633,N_13786);
xnor U13844 (N_13844,N_13664,N_13620);
nor U13845 (N_13845,N_13794,N_13765);
or U13846 (N_13846,N_13683,N_13650);
nand U13847 (N_13847,N_13698,N_13758);
xnor U13848 (N_13848,N_13691,N_13684);
nor U13849 (N_13849,N_13731,N_13715);
and U13850 (N_13850,N_13699,N_13732);
or U13851 (N_13851,N_13763,N_13747);
nor U13852 (N_13852,N_13779,N_13798);
or U13853 (N_13853,N_13707,N_13703);
nand U13854 (N_13854,N_13713,N_13614);
or U13855 (N_13855,N_13764,N_13680);
xnor U13856 (N_13856,N_13770,N_13682);
and U13857 (N_13857,N_13782,N_13611);
nand U13858 (N_13858,N_13744,N_13625);
nor U13859 (N_13859,N_13617,N_13737);
nor U13860 (N_13860,N_13720,N_13641);
nand U13861 (N_13861,N_13607,N_13791);
and U13862 (N_13862,N_13701,N_13665);
and U13863 (N_13863,N_13642,N_13704);
xnor U13864 (N_13864,N_13729,N_13709);
and U13865 (N_13865,N_13678,N_13741);
or U13866 (N_13866,N_13629,N_13666);
nor U13867 (N_13867,N_13601,N_13774);
or U13868 (N_13868,N_13795,N_13749);
nor U13869 (N_13869,N_13777,N_13767);
nand U13870 (N_13870,N_13653,N_13785);
nand U13871 (N_13871,N_13634,N_13793);
and U13872 (N_13872,N_13604,N_13700);
or U13873 (N_13873,N_13623,N_13728);
or U13874 (N_13874,N_13688,N_13615);
xnor U13875 (N_13875,N_13655,N_13649);
and U13876 (N_13876,N_13748,N_13661);
xor U13877 (N_13877,N_13722,N_13796);
and U13878 (N_13878,N_13754,N_13710);
or U13879 (N_13879,N_13662,N_13608);
or U13880 (N_13880,N_13761,N_13759);
or U13881 (N_13881,N_13605,N_13630);
and U13882 (N_13882,N_13708,N_13658);
and U13883 (N_13883,N_13740,N_13656);
or U13884 (N_13884,N_13646,N_13742);
nand U13885 (N_13885,N_13675,N_13640);
and U13886 (N_13886,N_13693,N_13799);
nand U13887 (N_13887,N_13689,N_13670);
or U13888 (N_13888,N_13790,N_13727);
or U13889 (N_13889,N_13685,N_13651);
or U13890 (N_13890,N_13648,N_13772);
xnor U13891 (N_13891,N_13735,N_13752);
xor U13892 (N_13892,N_13768,N_13686);
nor U13893 (N_13893,N_13622,N_13733);
nand U13894 (N_13894,N_13738,N_13792);
and U13895 (N_13895,N_13746,N_13694);
nor U13896 (N_13896,N_13638,N_13743);
xor U13897 (N_13897,N_13696,N_13667);
nand U13898 (N_13898,N_13679,N_13702);
or U13899 (N_13899,N_13619,N_13644);
and U13900 (N_13900,N_13632,N_13731);
or U13901 (N_13901,N_13607,N_13611);
xor U13902 (N_13902,N_13661,N_13716);
and U13903 (N_13903,N_13687,N_13788);
and U13904 (N_13904,N_13775,N_13698);
and U13905 (N_13905,N_13680,N_13719);
and U13906 (N_13906,N_13792,N_13736);
nor U13907 (N_13907,N_13789,N_13795);
xor U13908 (N_13908,N_13719,N_13677);
xnor U13909 (N_13909,N_13743,N_13755);
nor U13910 (N_13910,N_13790,N_13688);
xor U13911 (N_13911,N_13705,N_13752);
nand U13912 (N_13912,N_13675,N_13694);
nor U13913 (N_13913,N_13766,N_13674);
xor U13914 (N_13914,N_13670,N_13664);
nand U13915 (N_13915,N_13784,N_13742);
or U13916 (N_13916,N_13608,N_13723);
nand U13917 (N_13917,N_13794,N_13777);
nand U13918 (N_13918,N_13756,N_13634);
or U13919 (N_13919,N_13634,N_13601);
xor U13920 (N_13920,N_13660,N_13677);
nor U13921 (N_13921,N_13668,N_13681);
xor U13922 (N_13922,N_13788,N_13787);
nor U13923 (N_13923,N_13798,N_13756);
xor U13924 (N_13924,N_13736,N_13644);
and U13925 (N_13925,N_13669,N_13656);
xor U13926 (N_13926,N_13686,N_13653);
xnor U13927 (N_13927,N_13731,N_13779);
xnor U13928 (N_13928,N_13790,N_13757);
nand U13929 (N_13929,N_13744,N_13713);
and U13930 (N_13930,N_13643,N_13660);
or U13931 (N_13931,N_13608,N_13623);
xor U13932 (N_13932,N_13782,N_13682);
and U13933 (N_13933,N_13735,N_13659);
or U13934 (N_13934,N_13651,N_13711);
nor U13935 (N_13935,N_13656,N_13697);
or U13936 (N_13936,N_13789,N_13714);
or U13937 (N_13937,N_13727,N_13753);
xor U13938 (N_13938,N_13650,N_13642);
nand U13939 (N_13939,N_13763,N_13663);
or U13940 (N_13940,N_13665,N_13648);
and U13941 (N_13941,N_13618,N_13667);
xnor U13942 (N_13942,N_13787,N_13735);
and U13943 (N_13943,N_13729,N_13795);
xor U13944 (N_13944,N_13789,N_13759);
or U13945 (N_13945,N_13661,N_13679);
nor U13946 (N_13946,N_13772,N_13797);
nor U13947 (N_13947,N_13797,N_13782);
nor U13948 (N_13948,N_13695,N_13698);
or U13949 (N_13949,N_13758,N_13600);
or U13950 (N_13950,N_13703,N_13662);
and U13951 (N_13951,N_13630,N_13703);
and U13952 (N_13952,N_13622,N_13763);
or U13953 (N_13953,N_13703,N_13658);
and U13954 (N_13954,N_13739,N_13764);
xor U13955 (N_13955,N_13671,N_13696);
or U13956 (N_13956,N_13686,N_13709);
nand U13957 (N_13957,N_13679,N_13726);
nand U13958 (N_13958,N_13670,N_13760);
nand U13959 (N_13959,N_13715,N_13672);
and U13960 (N_13960,N_13719,N_13629);
and U13961 (N_13961,N_13616,N_13688);
nand U13962 (N_13962,N_13739,N_13782);
xor U13963 (N_13963,N_13631,N_13639);
and U13964 (N_13964,N_13613,N_13602);
or U13965 (N_13965,N_13627,N_13601);
or U13966 (N_13966,N_13743,N_13613);
or U13967 (N_13967,N_13728,N_13679);
nand U13968 (N_13968,N_13679,N_13739);
and U13969 (N_13969,N_13732,N_13701);
and U13970 (N_13970,N_13780,N_13721);
nor U13971 (N_13971,N_13650,N_13749);
nand U13972 (N_13972,N_13729,N_13617);
nor U13973 (N_13973,N_13698,N_13652);
nor U13974 (N_13974,N_13780,N_13738);
nor U13975 (N_13975,N_13773,N_13660);
nor U13976 (N_13976,N_13794,N_13636);
or U13977 (N_13977,N_13739,N_13733);
xor U13978 (N_13978,N_13635,N_13792);
nor U13979 (N_13979,N_13737,N_13722);
and U13980 (N_13980,N_13717,N_13678);
xor U13981 (N_13981,N_13715,N_13778);
and U13982 (N_13982,N_13689,N_13602);
nor U13983 (N_13983,N_13799,N_13753);
and U13984 (N_13984,N_13622,N_13792);
nand U13985 (N_13985,N_13625,N_13726);
or U13986 (N_13986,N_13692,N_13679);
xnor U13987 (N_13987,N_13611,N_13622);
xnor U13988 (N_13988,N_13671,N_13719);
or U13989 (N_13989,N_13634,N_13615);
xor U13990 (N_13990,N_13601,N_13690);
and U13991 (N_13991,N_13685,N_13728);
or U13992 (N_13992,N_13768,N_13621);
or U13993 (N_13993,N_13734,N_13673);
and U13994 (N_13994,N_13693,N_13700);
xnor U13995 (N_13995,N_13648,N_13638);
nand U13996 (N_13996,N_13709,N_13621);
or U13997 (N_13997,N_13666,N_13601);
xnor U13998 (N_13998,N_13653,N_13705);
or U13999 (N_13999,N_13609,N_13701);
or U14000 (N_14000,N_13927,N_13916);
and U14001 (N_14001,N_13900,N_13819);
xor U14002 (N_14002,N_13961,N_13970);
nor U14003 (N_14003,N_13836,N_13918);
or U14004 (N_14004,N_13937,N_13920);
nor U14005 (N_14005,N_13911,N_13817);
nor U14006 (N_14006,N_13865,N_13827);
and U14007 (N_14007,N_13960,N_13886);
and U14008 (N_14008,N_13824,N_13832);
or U14009 (N_14009,N_13830,N_13958);
or U14010 (N_14010,N_13909,N_13852);
nor U14011 (N_14011,N_13975,N_13919);
nor U14012 (N_14012,N_13985,N_13972);
xor U14013 (N_14013,N_13947,N_13866);
or U14014 (N_14014,N_13899,N_13914);
xor U14015 (N_14015,N_13987,N_13984);
and U14016 (N_14016,N_13951,N_13854);
or U14017 (N_14017,N_13870,N_13890);
or U14018 (N_14018,N_13946,N_13889);
and U14019 (N_14019,N_13912,N_13989);
and U14020 (N_14020,N_13897,N_13873);
nor U14021 (N_14021,N_13986,N_13954);
nand U14022 (N_14022,N_13839,N_13996);
xnor U14023 (N_14023,N_13877,N_13885);
and U14024 (N_14024,N_13833,N_13853);
nor U14025 (N_14025,N_13935,N_13879);
nand U14026 (N_14026,N_13803,N_13862);
nor U14027 (N_14027,N_13808,N_13843);
nand U14028 (N_14028,N_13904,N_13962);
nand U14029 (N_14029,N_13829,N_13901);
nand U14030 (N_14030,N_13814,N_13851);
and U14031 (N_14031,N_13822,N_13867);
nor U14032 (N_14032,N_13857,N_13856);
nor U14033 (N_14033,N_13915,N_13846);
or U14034 (N_14034,N_13805,N_13974);
and U14035 (N_14035,N_13864,N_13982);
xnor U14036 (N_14036,N_13894,N_13823);
nor U14037 (N_14037,N_13977,N_13903);
nand U14038 (N_14038,N_13991,N_13884);
nor U14039 (N_14039,N_13800,N_13847);
and U14040 (N_14040,N_13922,N_13952);
or U14041 (N_14041,N_13930,N_13995);
nor U14042 (N_14042,N_13921,N_13956);
xor U14043 (N_14043,N_13964,N_13950);
nand U14044 (N_14044,N_13940,N_13845);
nand U14045 (N_14045,N_13831,N_13934);
and U14046 (N_14046,N_13876,N_13992);
nor U14047 (N_14047,N_13926,N_13849);
xor U14048 (N_14048,N_13869,N_13941);
nand U14049 (N_14049,N_13892,N_13932);
nand U14050 (N_14050,N_13931,N_13841);
xor U14051 (N_14051,N_13933,N_13850);
nor U14052 (N_14052,N_13949,N_13907);
xnor U14053 (N_14053,N_13874,N_13888);
nor U14054 (N_14054,N_13871,N_13828);
nor U14055 (N_14055,N_13959,N_13998);
or U14056 (N_14056,N_13968,N_13910);
nor U14057 (N_14057,N_13872,N_13861);
and U14058 (N_14058,N_13801,N_13925);
nand U14059 (N_14059,N_13896,N_13837);
nand U14060 (N_14060,N_13953,N_13955);
or U14061 (N_14061,N_13967,N_13860);
xnor U14062 (N_14062,N_13928,N_13834);
xnor U14063 (N_14063,N_13883,N_13988);
xnor U14064 (N_14064,N_13898,N_13971);
nor U14065 (N_14065,N_13880,N_13936);
xnor U14066 (N_14066,N_13994,N_13878);
and U14067 (N_14067,N_13891,N_13809);
and U14068 (N_14068,N_13939,N_13966);
and U14069 (N_14069,N_13976,N_13844);
nor U14070 (N_14070,N_13806,N_13815);
nand U14071 (N_14071,N_13802,N_13944);
or U14072 (N_14072,N_13980,N_13875);
or U14073 (N_14073,N_13842,N_13997);
or U14074 (N_14074,N_13826,N_13979);
nor U14075 (N_14075,N_13825,N_13923);
and U14076 (N_14076,N_13859,N_13948);
nand U14077 (N_14077,N_13821,N_13812);
nand U14078 (N_14078,N_13990,N_13908);
or U14079 (N_14079,N_13999,N_13973);
and U14080 (N_14080,N_13835,N_13863);
or U14081 (N_14081,N_13945,N_13993);
xnor U14082 (N_14082,N_13848,N_13820);
xor U14083 (N_14083,N_13813,N_13881);
nand U14084 (N_14084,N_13858,N_13868);
or U14085 (N_14085,N_13807,N_13840);
nor U14086 (N_14086,N_13917,N_13804);
xor U14087 (N_14087,N_13981,N_13882);
xor U14088 (N_14088,N_13895,N_13816);
or U14089 (N_14089,N_13963,N_13957);
xor U14090 (N_14090,N_13938,N_13943);
xor U14091 (N_14091,N_13838,N_13929);
nor U14092 (N_14092,N_13942,N_13893);
nand U14093 (N_14093,N_13905,N_13887);
nand U14094 (N_14094,N_13924,N_13855);
nand U14095 (N_14095,N_13983,N_13818);
nor U14096 (N_14096,N_13810,N_13906);
nor U14097 (N_14097,N_13969,N_13965);
xnor U14098 (N_14098,N_13913,N_13978);
nand U14099 (N_14099,N_13902,N_13811);
nor U14100 (N_14100,N_13902,N_13952);
nor U14101 (N_14101,N_13952,N_13869);
and U14102 (N_14102,N_13845,N_13989);
nand U14103 (N_14103,N_13933,N_13877);
xnor U14104 (N_14104,N_13947,N_13850);
or U14105 (N_14105,N_13920,N_13870);
and U14106 (N_14106,N_13811,N_13843);
or U14107 (N_14107,N_13956,N_13996);
nand U14108 (N_14108,N_13919,N_13856);
and U14109 (N_14109,N_13811,N_13906);
or U14110 (N_14110,N_13993,N_13882);
xor U14111 (N_14111,N_13819,N_13850);
nor U14112 (N_14112,N_13917,N_13832);
or U14113 (N_14113,N_13895,N_13946);
or U14114 (N_14114,N_13948,N_13917);
nor U14115 (N_14115,N_13899,N_13996);
xnor U14116 (N_14116,N_13996,N_13801);
and U14117 (N_14117,N_13805,N_13891);
nand U14118 (N_14118,N_13807,N_13812);
and U14119 (N_14119,N_13864,N_13820);
or U14120 (N_14120,N_13885,N_13987);
nor U14121 (N_14121,N_13820,N_13895);
nand U14122 (N_14122,N_13855,N_13860);
and U14123 (N_14123,N_13960,N_13867);
xor U14124 (N_14124,N_13851,N_13897);
or U14125 (N_14125,N_13979,N_13805);
nor U14126 (N_14126,N_13997,N_13865);
and U14127 (N_14127,N_13938,N_13980);
or U14128 (N_14128,N_13899,N_13821);
nand U14129 (N_14129,N_13987,N_13951);
and U14130 (N_14130,N_13969,N_13907);
xor U14131 (N_14131,N_13831,N_13832);
or U14132 (N_14132,N_13842,N_13846);
xnor U14133 (N_14133,N_13933,N_13925);
and U14134 (N_14134,N_13954,N_13942);
and U14135 (N_14135,N_13961,N_13873);
or U14136 (N_14136,N_13834,N_13806);
nand U14137 (N_14137,N_13996,N_13945);
xnor U14138 (N_14138,N_13875,N_13858);
nand U14139 (N_14139,N_13889,N_13845);
nand U14140 (N_14140,N_13916,N_13996);
xor U14141 (N_14141,N_13941,N_13858);
and U14142 (N_14142,N_13928,N_13879);
xor U14143 (N_14143,N_13986,N_13848);
or U14144 (N_14144,N_13960,N_13888);
or U14145 (N_14145,N_13982,N_13866);
or U14146 (N_14146,N_13983,N_13939);
nor U14147 (N_14147,N_13945,N_13965);
or U14148 (N_14148,N_13970,N_13876);
xnor U14149 (N_14149,N_13843,N_13995);
and U14150 (N_14150,N_13845,N_13872);
nand U14151 (N_14151,N_13832,N_13944);
and U14152 (N_14152,N_13995,N_13972);
or U14153 (N_14153,N_13968,N_13980);
nor U14154 (N_14154,N_13954,N_13899);
and U14155 (N_14155,N_13843,N_13989);
and U14156 (N_14156,N_13988,N_13845);
and U14157 (N_14157,N_13929,N_13886);
xor U14158 (N_14158,N_13809,N_13986);
and U14159 (N_14159,N_13878,N_13976);
or U14160 (N_14160,N_13871,N_13838);
xnor U14161 (N_14161,N_13972,N_13978);
nand U14162 (N_14162,N_13810,N_13981);
nand U14163 (N_14163,N_13804,N_13831);
nor U14164 (N_14164,N_13817,N_13864);
and U14165 (N_14165,N_13890,N_13918);
and U14166 (N_14166,N_13889,N_13814);
xor U14167 (N_14167,N_13816,N_13981);
nor U14168 (N_14168,N_13907,N_13901);
and U14169 (N_14169,N_13846,N_13864);
and U14170 (N_14170,N_13804,N_13974);
and U14171 (N_14171,N_13880,N_13997);
and U14172 (N_14172,N_13866,N_13815);
and U14173 (N_14173,N_13910,N_13825);
or U14174 (N_14174,N_13897,N_13824);
xor U14175 (N_14175,N_13918,N_13879);
xor U14176 (N_14176,N_13968,N_13900);
and U14177 (N_14177,N_13840,N_13928);
xnor U14178 (N_14178,N_13903,N_13922);
xor U14179 (N_14179,N_13846,N_13961);
nor U14180 (N_14180,N_13901,N_13849);
xor U14181 (N_14181,N_13828,N_13929);
and U14182 (N_14182,N_13923,N_13955);
xor U14183 (N_14183,N_13934,N_13861);
and U14184 (N_14184,N_13838,N_13963);
xor U14185 (N_14185,N_13860,N_13813);
nand U14186 (N_14186,N_13804,N_13824);
xnor U14187 (N_14187,N_13898,N_13812);
xor U14188 (N_14188,N_13892,N_13943);
and U14189 (N_14189,N_13816,N_13861);
nand U14190 (N_14190,N_13825,N_13891);
nor U14191 (N_14191,N_13923,N_13956);
xor U14192 (N_14192,N_13932,N_13855);
xnor U14193 (N_14193,N_13806,N_13841);
nor U14194 (N_14194,N_13937,N_13832);
and U14195 (N_14195,N_13973,N_13803);
or U14196 (N_14196,N_13908,N_13958);
nor U14197 (N_14197,N_13973,N_13842);
nand U14198 (N_14198,N_13906,N_13860);
xnor U14199 (N_14199,N_13844,N_13927);
xor U14200 (N_14200,N_14183,N_14049);
and U14201 (N_14201,N_14041,N_14014);
nor U14202 (N_14202,N_14081,N_14174);
xor U14203 (N_14203,N_14080,N_14169);
nor U14204 (N_14204,N_14015,N_14153);
xor U14205 (N_14205,N_14085,N_14197);
or U14206 (N_14206,N_14070,N_14179);
or U14207 (N_14207,N_14092,N_14100);
xnor U14208 (N_14208,N_14160,N_14066);
or U14209 (N_14209,N_14019,N_14002);
and U14210 (N_14210,N_14107,N_14123);
or U14211 (N_14211,N_14168,N_14089);
nand U14212 (N_14212,N_14180,N_14039);
nand U14213 (N_14213,N_14155,N_14071);
and U14214 (N_14214,N_14138,N_14053);
or U14215 (N_14215,N_14105,N_14045);
nor U14216 (N_14216,N_14156,N_14158);
or U14217 (N_14217,N_14079,N_14142);
or U14218 (N_14218,N_14109,N_14151);
nand U14219 (N_14219,N_14073,N_14025);
nor U14220 (N_14220,N_14193,N_14150);
nor U14221 (N_14221,N_14046,N_14145);
or U14222 (N_14222,N_14167,N_14044);
or U14223 (N_14223,N_14022,N_14095);
or U14224 (N_14224,N_14139,N_14061);
nor U14225 (N_14225,N_14065,N_14108);
nand U14226 (N_14226,N_14056,N_14106);
nor U14227 (N_14227,N_14072,N_14147);
nor U14228 (N_14228,N_14163,N_14196);
or U14229 (N_14229,N_14128,N_14136);
nand U14230 (N_14230,N_14004,N_14037);
and U14231 (N_14231,N_14067,N_14101);
nor U14232 (N_14232,N_14023,N_14187);
nand U14233 (N_14233,N_14154,N_14047);
or U14234 (N_14234,N_14175,N_14103);
nor U14235 (N_14235,N_14057,N_14199);
nand U14236 (N_14236,N_14190,N_14165);
and U14237 (N_14237,N_14144,N_14000);
or U14238 (N_14238,N_14048,N_14148);
xnor U14239 (N_14239,N_14099,N_14069);
and U14240 (N_14240,N_14192,N_14171);
nor U14241 (N_14241,N_14164,N_14008);
xnor U14242 (N_14242,N_14010,N_14090);
nand U14243 (N_14243,N_14083,N_14119);
and U14244 (N_14244,N_14186,N_14130);
nor U14245 (N_14245,N_14030,N_14093);
and U14246 (N_14246,N_14018,N_14027);
xnor U14247 (N_14247,N_14157,N_14084);
nor U14248 (N_14248,N_14181,N_14137);
and U14249 (N_14249,N_14082,N_14032);
or U14250 (N_14250,N_14110,N_14020);
xnor U14251 (N_14251,N_14117,N_14006);
nand U14252 (N_14252,N_14011,N_14114);
nor U14253 (N_14253,N_14184,N_14098);
or U14254 (N_14254,N_14122,N_14077);
nand U14255 (N_14255,N_14058,N_14176);
nand U14256 (N_14256,N_14104,N_14195);
or U14257 (N_14257,N_14162,N_14013);
nor U14258 (N_14258,N_14116,N_14021);
nor U14259 (N_14259,N_14191,N_14052);
or U14260 (N_14260,N_14097,N_14024);
and U14261 (N_14261,N_14102,N_14173);
or U14262 (N_14262,N_14120,N_14152);
and U14263 (N_14263,N_14003,N_14096);
and U14264 (N_14264,N_14086,N_14185);
and U14265 (N_14265,N_14177,N_14001);
and U14266 (N_14266,N_14055,N_14135);
and U14267 (N_14267,N_14068,N_14031);
or U14268 (N_14268,N_14198,N_14146);
nand U14269 (N_14269,N_14060,N_14087);
nor U14270 (N_14270,N_14188,N_14124);
nor U14271 (N_14271,N_14111,N_14115);
or U14272 (N_14272,N_14009,N_14063);
nor U14273 (N_14273,N_14078,N_14088);
or U14274 (N_14274,N_14182,N_14140);
or U14275 (N_14275,N_14170,N_14189);
xor U14276 (N_14276,N_14118,N_14112);
and U14277 (N_14277,N_14134,N_14178);
xor U14278 (N_14278,N_14133,N_14054);
nand U14279 (N_14279,N_14074,N_14075);
nor U14280 (N_14280,N_14129,N_14035);
nand U14281 (N_14281,N_14029,N_14126);
or U14282 (N_14282,N_14033,N_14149);
xnor U14283 (N_14283,N_14127,N_14043);
and U14284 (N_14284,N_14194,N_14042);
xnor U14285 (N_14285,N_14143,N_14076);
nor U14286 (N_14286,N_14064,N_14017);
or U14287 (N_14287,N_14028,N_14026);
or U14288 (N_14288,N_14036,N_14094);
nand U14289 (N_14289,N_14034,N_14161);
nor U14290 (N_14290,N_14050,N_14005);
or U14291 (N_14291,N_14172,N_14125);
or U14292 (N_14292,N_14091,N_14062);
or U14293 (N_14293,N_14131,N_14113);
nand U14294 (N_14294,N_14051,N_14121);
and U14295 (N_14295,N_14012,N_14038);
or U14296 (N_14296,N_14059,N_14141);
nor U14297 (N_14297,N_14007,N_14132);
and U14298 (N_14298,N_14166,N_14159);
and U14299 (N_14299,N_14040,N_14016);
or U14300 (N_14300,N_14058,N_14165);
xor U14301 (N_14301,N_14038,N_14013);
nand U14302 (N_14302,N_14193,N_14071);
or U14303 (N_14303,N_14110,N_14122);
nor U14304 (N_14304,N_14054,N_14192);
or U14305 (N_14305,N_14172,N_14057);
or U14306 (N_14306,N_14046,N_14083);
nand U14307 (N_14307,N_14105,N_14163);
and U14308 (N_14308,N_14096,N_14184);
nand U14309 (N_14309,N_14024,N_14043);
nand U14310 (N_14310,N_14155,N_14115);
xor U14311 (N_14311,N_14072,N_14162);
xnor U14312 (N_14312,N_14073,N_14108);
nor U14313 (N_14313,N_14171,N_14091);
and U14314 (N_14314,N_14030,N_14151);
and U14315 (N_14315,N_14040,N_14014);
or U14316 (N_14316,N_14186,N_14084);
nor U14317 (N_14317,N_14089,N_14175);
and U14318 (N_14318,N_14194,N_14088);
nand U14319 (N_14319,N_14125,N_14083);
nor U14320 (N_14320,N_14144,N_14107);
nand U14321 (N_14321,N_14105,N_14080);
and U14322 (N_14322,N_14022,N_14194);
nand U14323 (N_14323,N_14130,N_14118);
nor U14324 (N_14324,N_14082,N_14011);
and U14325 (N_14325,N_14009,N_14135);
and U14326 (N_14326,N_14058,N_14152);
and U14327 (N_14327,N_14160,N_14196);
xor U14328 (N_14328,N_14086,N_14085);
and U14329 (N_14329,N_14056,N_14169);
nor U14330 (N_14330,N_14008,N_14099);
nand U14331 (N_14331,N_14156,N_14174);
nor U14332 (N_14332,N_14023,N_14032);
xnor U14333 (N_14333,N_14106,N_14090);
or U14334 (N_14334,N_14026,N_14174);
xor U14335 (N_14335,N_14047,N_14080);
nand U14336 (N_14336,N_14189,N_14103);
nand U14337 (N_14337,N_14031,N_14085);
or U14338 (N_14338,N_14116,N_14043);
and U14339 (N_14339,N_14102,N_14160);
xor U14340 (N_14340,N_14185,N_14161);
nor U14341 (N_14341,N_14096,N_14034);
and U14342 (N_14342,N_14079,N_14014);
xnor U14343 (N_14343,N_14179,N_14195);
nand U14344 (N_14344,N_14105,N_14081);
and U14345 (N_14345,N_14111,N_14154);
or U14346 (N_14346,N_14063,N_14067);
nand U14347 (N_14347,N_14007,N_14143);
nor U14348 (N_14348,N_14017,N_14179);
nand U14349 (N_14349,N_14076,N_14198);
and U14350 (N_14350,N_14066,N_14167);
or U14351 (N_14351,N_14080,N_14160);
or U14352 (N_14352,N_14111,N_14146);
nand U14353 (N_14353,N_14105,N_14187);
nor U14354 (N_14354,N_14080,N_14110);
xnor U14355 (N_14355,N_14028,N_14192);
and U14356 (N_14356,N_14127,N_14187);
nand U14357 (N_14357,N_14114,N_14025);
nor U14358 (N_14358,N_14064,N_14063);
nand U14359 (N_14359,N_14125,N_14003);
nor U14360 (N_14360,N_14130,N_14136);
xnor U14361 (N_14361,N_14105,N_14175);
and U14362 (N_14362,N_14065,N_14040);
or U14363 (N_14363,N_14025,N_14046);
and U14364 (N_14364,N_14051,N_14042);
xor U14365 (N_14365,N_14184,N_14123);
or U14366 (N_14366,N_14004,N_14029);
nor U14367 (N_14367,N_14062,N_14194);
or U14368 (N_14368,N_14066,N_14035);
xor U14369 (N_14369,N_14066,N_14159);
or U14370 (N_14370,N_14067,N_14192);
nand U14371 (N_14371,N_14094,N_14039);
or U14372 (N_14372,N_14007,N_14142);
nand U14373 (N_14373,N_14116,N_14089);
and U14374 (N_14374,N_14073,N_14183);
nor U14375 (N_14375,N_14168,N_14136);
xnor U14376 (N_14376,N_14080,N_14189);
and U14377 (N_14377,N_14078,N_14063);
and U14378 (N_14378,N_14091,N_14086);
and U14379 (N_14379,N_14010,N_14065);
and U14380 (N_14380,N_14110,N_14012);
xnor U14381 (N_14381,N_14048,N_14058);
xnor U14382 (N_14382,N_14162,N_14118);
and U14383 (N_14383,N_14115,N_14173);
and U14384 (N_14384,N_14162,N_14062);
nor U14385 (N_14385,N_14149,N_14010);
nor U14386 (N_14386,N_14047,N_14176);
nand U14387 (N_14387,N_14110,N_14174);
xor U14388 (N_14388,N_14082,N_14175);
nor U14389 (N_14389,N_14191,N_14144);
xor U14390 (N_14390,N_14133,N_14039);
nand U14391 (N_14391,N_14090,N_14005);
xor U14392 (N_14392,N_14198,N_14111);
nor U14393 (N_14393,N_14073,N_14085);
nor U14394 (N_14394,N_14015,N_14107);
xor U14395 (N_14395,N_14046,N_14188);
nor U14396 (N_14396,N_14122,N_14052);
or U14397 (N_14397,N_14089,N_14018);
nor U14398 (N_14398,N_14145,N_14198);
nor U14399 (N_14399,N_14190,N_14043);
and U14400 (N_14400,N_14318,N_14222);
nor U14401 (N_14401,N_14398,N_14319);
or U14402 (N_14402,N_14272,N_14330);
and U14403 (N_14403,N_14366,N_14295);
xnor U14404 (N_14404,N_14375,N_14247);
nand U14405 (N_14405,N_14347,N_14321);
xor U14406 (N_14406,N_14273,N_14244);
and U14407 (N_14407,N_14207,N_14394);
nor U14408 (N_14408,N_14245,N_14221);
or U14409 (N_14409,N_14359,N_14228);
or U14410 (N_14410,N_14266,N_14335);
and U14411 (N_14411,N_14292,N_14201);
nor U14412 (N_14412,N_14215,N_14357);
nand U14413 (N_14413,N_14339,N_14290);
and U14414 (N_14414,N_14233,N_14379);
nor U14415 (N_14415,N_14211,N_14314);
nor U14416 (N_14416,N_14344,N_14315);
and U14417 (N_14417,N_14322,N_14280);
nand U14418 (N_14418,N_14218,N_14332);
nor U14419 (N_14419,N_14348,N_14224);
nand U14420 (N_14420,N_14223,N_14217);
nor U14421 (N_14421,N_14337,N_14310);
nor U14422 (N_14422,N_14238,N_14303);
nand U14423 (N_14423,N_14237,N_14380);
nand U14424 (N_14424,N_14249,N_14267);
nor U14425 (N_14425,N_14283,N_14284);
or U14426 (N_14426,N_14382,N_14216);
and U14427 (N_14427,N_14317,N_14240);
nand U14428 (N_14428,N_14364,N_14376);
nor U14429 (N_14429,N_14235,N_14260);
nor U14430 (N_14430,N_14341,N_14333);
or U14431 (N_14431,N_14316,N_14371);
nand U14432 (N_14432,N_14263,N_14220);
xor U14433 (N_14433,N_14285,N_14386);
or U14434 (N_14434,N_14385,N_14296);
or U14435 (N_14435,N_14309,N_14326);
nand U14436 (N_14436,N_14251,N_14356);
and U14437 (N_14437,N_14200,N_14252);
and U14438 (N_14438,N_14301,N_14354);
nor U14439 (N_14439,N_14368,N_14306);
and U14440 (N_14440,N_14381,N_14350);
or U14441 (N_14441,N_14392,N_14242);
and U14442 (N_14442,N_14325,N_14230);
or U14443 (N_14443,N_14259,N_14313);
nand U14444 (N_14444,N_14231,N_14212);
nand U14445 (N_14445,N_14210,N_14399);
xnor U14446 (N_14446,N_14355,N_14342);
nor U14447 (N_14447,N_14287,N_14391);
nor U14448 (N_14448,N_14320,N_14293);
and U14449 (N_14449,N_14291,N_14214);
or U14450 (N_14450,N_14288,N_14300);
nor U14451 (N_14451,N_14311,N_14329);
or U14452 (N_14452,N_14378,N_14377);
nand U14453 (N_14453,N_14345,N_14387);
or U14454 (N_14454,N_14365,N_14229);
nand U14455 (N_14455,N_14236,N_14390);
nand U14456 (N_14456,N_14261,N_14206);
xor U14457 (N_14457,N_14336,N_14374);
nor U14458 (N_14458,N_14205,N_14395);
nand U14459 (N_14459,N_14270,N_14274);
and U14460 (N_14460,N_14307,N_14393);
nor U14461 (N_14461,N_14369,N_14334);
or U14462 (N_14462,N_14389,N_14268);
and U14463 (N_14463,N_14254,N_14397);
xnor U14464 (N_14464,N_14257,N_14370);
or U14465 (N_14465,N_14256,N_14243);
nor U14466 (N_14466,N_14358,N_14258);
xnor U14467 (N_14467,N_14343,N_14312);
nor U14468 (N_14468,N_14327,N_14227);
nand U14469 (N_14469,N_14362,N_14372);
or U14470 (N_14470,N_14202,N_14250);
or U14471 (N_14471,N_14248,N_14203);
nand U14472 (N_14472,N_14255,N_14352);
or U14473 (N_14473,N_14308,N_14298);
nand U14474 (N_14474,N_14331,N_14384);
xnor U14475 (N_14475,N_14328,N_14351);
nand U14476 (N_14476,N_14367,N_14373);
xnor U14477 (N_14477,N_14294,N_14338);
xnor U14478 (N_14478,N_14253,N_14213);
or U14479 (N_14479,N_14264,N_14246);
and U14480 (N_14480,N_14286,N_14262);
and U14481 (N_14481,N_14208,N_14361);
nor U14482 (N_14482,N_14277,N_14281);
nand U14483 (N_14483,N_14204,N_14226);
xnor U14484 (N_14484,N_14234,N_14219);
nand U14485 (N_14485,N_14271,N_14279);
or U14486 (N_14486,N_14324,N_14278);
nor U14487 (N_14487,N_14349,N_14241);
xor U14488 (N_14488,N_14304,N_14383);
or U14489 (N_14489,N_14225,N_14363);
nand U14490 (N_14490,N_14275,N_14360);
nand U14491 (N_14491,N_14265,N_14340);
xor U14492 (N_14492,N_14232,N_14239);
xnor U14493 (N_14493,N_14282,N_14297);
and U14494 (N_14494,N_14209,N_14299);
or U14495 (N_14495,N_14276,N_14323);
nor U14496 (N_14496,N_14305,N_14353);
and U14497 (N_14497,N_14289,N_14269);
nand U14498 (N_14498,N_14302,N_14396);
and U14499 (N_14499,N_14346,N_14388);
nor U14500 (N_14500,N_14339,N_14299);
xor U14501 (N_14501,N_14346,N_14274);
xnor U14502 (N_14502,N_14325,N_14288);
or U14503 (N_14503,N_14388,N_14207);
nand U14504 (N_14504,N_14398,N_14280);
nand U14505 (N_14505,N_14327,N_14302);
xnor U14506 (N_14506,N_14257,N_14327);
xnor U14507 (N_14507,N_14380,N_14242);
nor U14508 (N_14508,N_14367,N_14314);
and U14509 (N_14509,N_14225,N_14205);
xor U14510 (N_14510,N_14359,N_14284);
xor U14511 (N_14511,N_14395,N_14220);
nor U14512 (N_14512,N_14240,N_14221);
nor U14513 (N_14513,N_14331,N_14215);
xor U14514 (N_14514,N_14274,N_14271);
nand U14515 (N_14515,N_14338,N_14201);
and U14516 (N_14516,N_14218,N_14225);
nand U14517 (N_14517,N_14287,N_14394);
nor U14518 (N_14518,N_14364,N_14361);
nand U14519 (N_14519,N_14293,N_14394);
xnor U14520 (N_14520,N_14355,N_14298);
or U14521 (N_14521,N_14221,N_14348);
or U14522 (N_14522,N_14355,N_14227);
xnor U14523 (N_14523,N_14279,N_14383);
and U14524 (N_14524,N_14256,N_14229);
xor U14525 (N_14525,N_14364,N_14315);
xnor U14526 (N_14526,N_14249,N_14381);
nand U14527 (N_14527,N_14362,N_14204);
xnor U14528 (N_14528,N_14290,N_14336);
xnor U14529 (N_14529,N_14215,N_14355);
and U14530 (N_14530,N_14330,N_14346);
or U14531 (N_14531,N_14297,N_14309);
nor U14532 (N_14532,N_14211,N_14320);
nor U14533 (N_14533,N_14391,N_14267);
and U14534 (N_14534,N_14259,N_14236);
xnor U14535 (N_14535,N_14278,N_14259);
nand U14536 (N_14536,N_14326,N_14211);
nor U14537 (N_14537,N_14237,N_14212);
nor U14538 (N_14538,N_14311,N_14264);
nor U14539 (N_14539,N_14268,N_14393);
and U14540 (N_14540,N_14354,N_14314);
xnor U14541 (N_14541,N_14296,N_14395);
nor U14542 (N_14542,N_14224,N_14271);
nand U14543 (N_14543,N_14200,N_14396);
and U14544 (N_14544,N_14305,N_14294);
xnor U14545 (N_14545,N_14328,N_14392);
and U14546 (N_14546,N_14338,N_14372);
nor U14547 (N_14547,N_14302,N_14212);
or U14548 (N_14548,N_14347,N_14396);
and U14549 (N_14549,N_14355,N_14205);
nor U14550 (N_14550,N_14390,N_14211);
nand U14551 (N_14551,N_14356,N_14202);
and U14552 (N_14552,N_14310,N_14350);
and U14553 (N_14553,N_14206,N_14234);
or U14554 (N_14554,N_14334,N_14320);
nand U14555 (N_14555,N_14219,N_14350);
or U14556 (N_14556,N_14200,N_14381);
xnor U14557 (N_14557,N_14379,N_14352);
nor U14558 (N_14558,N_14305,N_14282);
xor U14559 (N_14559,N_14295,N_14348);
nor U14560 (N_14560,N_14304,N_14288);
nand U14561 (N_14561,N_14354,N_14396);
xnor U14562 (N_14562,N_14312,N_14362);
or U14563 (N_14563,N_14219,N_14344);
and U14564 (N_14564,N_14361,N_14203);
or U14565 (N_14565,N_14274,N_14273);
nand U14566 (N_14566,N_14378,N_14363);
nand U14567 (N_14567,N_14252,N_14367);
or U14568 (N_14568,N_14389,N_14226);
xor U14569 (N_14569,N_14296,N_14266);
or U14570 (N_14570,N_14222,N_14304);
and U14571 (N_14571,N_14218,N_14366);
or U14572 (N_14572,N_14261,N_14256);
nor U14573 (N_14573,N_14284,N_14291);
xor U14574 (N_14574,N_14346,N_14371);
nand U14575 (N_14575,N_14226,N_14258);
nor U14576 (N_14576,N_14254,N_14212);
nor U14577 (N_14577,N_14230,N_14383);
xor U14578 (N_14578,N_14250,N_14274);
and U14579 (N_14579,N_14207,N_14367);
nand U14580 (N_14580,N_14354,N_14224);
xor U14581 (N_14581,N_14318,N_14349);
or U14582 (N_14582,N_14249,N_14379);
nor U14583 (N_14583,N_14377,N_14270);
nor U14584 (N_14584,N_14272,N_14389);
xor U14585 (N_14585,N_14207,N_14222);
and U14586 (N_14586,N_14201,N_14339);
xor U14587 (N_14587,N_14334,N_14268);
nand U14588 (N_14588,N_14270,N_14289);
and U14589 (N_14589,N_14269,N_14283);
xnor U14590 (N_14590,N_14281,N_14207);
nor U14591 (N_14591,N_14371,N_14342);
or U14592 (N_14592,N_14294,N_14251);
nor U14593 (N_14593,N_14336,N_14221);
and U14594 (N_14594,N_14239,N_14364);
xnor U14595 (N_14595,N_14375,N_14264);
and U14596 (N_14596,N_14267,N_14215);
nor U14597 (N_14597,N_14315,N_14258);
or U14598 (N_14598,N_14350,N_14341);
and U14599 (N_14599,N_14286,N_14206);
and U14600 (N_14600,N_14456,N_14459);
nand U14601 (N_14601,N_14559,N_14444);
and U14602 (N_14602,N_14416,N_14438);
nand U14603 (N_14603,N_14534,N_14599);
nand U14604 (N_14604,N_14562,N_14433);
nand U14605 (N_14605,N_14585,N_14569);
nor U14606 (N_14606,N_14463,N_14471);
and U14607 (N_14607,N_14517,N_14451);
nand U14608 (N_14608,N_14485,N_14556);
or U14609 (N_14609,N_14429,N_14504);
nand U14610 (N_14610,N_14401,N_14500);
nor U14611 (N_14611,N_14489,N_14588);
nand U14612 (N_14612,N_14526,N_14494);
and U14613 (N_14613,N_14548,N_14449);
nand U14614 (N_14614,N_14476,N_14593);
nand U14615 (N_14615,N_14483,N_14447);
xor U14616 (N_14616,N_14570,N_14580);
nand U14617 (N_14617,N_14455,N_14521);
or U14618 (N_14618,N_14442,N_14407);
nor U14619 (N_14619,N_14422,N_14430);
xor U14620 (N_14620,N_14568,N_14555);
or U14621 (N_14621,N_14445,N_14481);
nand U14622 (N_14622,N_14540,N_14546);
nand U14623 (N_14623,N_14474,N_14406);
nand U14624 (N_14624,N_14409,N_14598);
and U14625 (N_14625,N_14529,N_14558);
xnor U14626 (N_14626,N_14510,N_14577);
nand U14627 (N_14627,N_14522,N_14520);
and U14628 (N_14628,N_14417,N_14565);
xnor U14629 (N_14629,N_14578,N_14589);
nand U14630 (N_14630,N_14505,N_14590);
nor U14631 (N_14631,N_14424,N_14514);
nor U14632 (N_14632,N_14516,N_14427);
xnor U14633 (N_14633,N_14508,N_14557);
xnor U14634 (N_14634,N_14573,N_14560);
or U14635 (N_14635,N_14426,N_14462);
or U14636 (N_14636,N_14452,N_14423);
nand U14637 (N_14637,N_14566,N_14525);
or U14638 (N_14638,N_14414,N_14428);
nand U14639 (N_14639,N_14403,N_14511);
nand U14640 (N_14640,N_14421,N_14495);
nand U14641 (N_14641,N_14453,N_14480);
nor U14642 (N_14642,N_14402,N_14412);
nand U14643 (N_14643,N_14475,N_14544);
or U14644 (N_14644,N_14575,N_14535);
nand U14645 (N_14645,N_14542,N_14531);
xnor U14646 (N_14646,N_14418,N_14488);
nor U14647 (N_14647,N_14492,N_14572);
nand U14648 (N_14648,N_14594,N_14567);
and U14649 (N_14649,N_14477,N_14581);
nand U14650 (N_14650,N_14579,N_14457);
and U14651 (N_14651,N_14468,N_14530);
xor U14652 (N_14652,N_14491,N_14518);
or U14653 (N_14653,N_14469,N_14503);
xnor U14654 (N_14654,N_14533,N_14490);
xnor U14655 (N_14655,N_14571,N_14400);
nor U14656 (N_14656,N_14596,N_14552);
nand U14657 (N_14657,N_14537,N_14597);
nor U14658 (N_14658,N_14470,N_14524);
nand U14659 (N_14659,N_14528,N_14527);
nand U14660 (N_14660,N_14509,N_14465);
and U14661 (N_14661,N_14461,N_14458);
xor U14662 (N_14662,N_14501,N_14454);
nor U14663 (N_14663,N_14574,N_14419);
xor U14664 (N_14664,N_14415,N_14486);
and U14665 (N_14665,N_14440,N_14595);
nand U14666 (N_14666,N_14432,N_14583);
and U14667 (N_14667,N_14443,N_14413);
nand U14668 (N_14668,N_14434,N_14539);
nand U14669 (N_14669,N_14512,N_14479);
nor U14670 (N_14670,N_14439,N_14435);
or U14671 (N_14671,N_14498,N_14473);
and U14672 (N_14672,N_14446,N_14538);
nand U14673 (N_14673,N_14408,N_14484);
and U14674 (N_14674,N_14515,N_14507);
xnor U14675 (N_14675,N_14591,N_14410);
or U14676 (N_14676,N_14478,N_14543);
nand U14677 (N_14677,N_14441,N_14404);
nor U14678 (N_14678,N_14547,N_14460);
or U14679 (N_14679,N_14493,N_14519);
xnor U14680 (N_14680,N_14466,N_14587);
or U14681 (N_14681,N_14467,N_14405);
and U14682 (N_14682,N_14431,N_14532);
nor U14683 (N_14683,N_14584,N_14545);
nand U14684 (N_14684,N_14561,N_14506);
xnor U14685 (N_14685,N_14563,N_14564);
xnor U14686 (N_14686,N_14448,N_14482);
nand U14687 (N_14687,N_14502,N_14553);
nand U14688 (N_14688,N_14549,N_14464);
and U14689 (N_14689,N_14551,N_14436);
xnor U14690 (N_14690,N_14496,N_14576);
xnor U14691 (N_14691,N_14499,N_14513);
and U14692 (N_14692,N_14592,N_14541);
nand U14693 (N_14693,N_14487,N_14586);
nand U14694 (N_14694,N_14523,N_14497);
or U14695 (N_14695,N_14425,N_14536);
nor U14696 (N_14696,N_14582,N_14550);
or U14697 (N_14697,N_14450,N_14472);
xor U14698 (N_14698,N_14420,N_14411);
or U14699 (N_14699,N_14437,N_14554);
xnor U14700 (N_14700,N_14414,N_14461);
or U14701 (N_14701,N_14425,N_14541);
nor U14702 (N_14702,N_14557,N_14531);
and U14703 (N_14703,N_14415,N_14541);
and U14704 (N_14704,N_14413,N_14594);
xnor U14705 (N_14705,N_14503,N_14523);
or U14706 (N_14706,N_14534,N_14582);
and U14707 (N_14707,N_14523,N_14596);
or U14708 (N_14708,N_14535,N_14529);
or U14709 (N_14709,N_14535,N_14447);
nor U14710 (N_14710,N_14589,N_14525);
or U14711 (N_14711,N_14418,N_14410);
xnor U14712 (N_14712,N_14458,N_14486);
xor U14713 (N_14713,N_14401,N_14490);
nand U14714 (N_14714,N_14461,N_14445);
xor U14715 (N_14715,N_14480,N_14434);
xnor U14716 (N_14716,N_14518,N_14495);
nor U14717 (N_14717,N_14422,N_14558);
nand U14718 (N_14718,N_14508,N_14560);
nand U14719 (N_14719,N_14419,N_14519);
nor U14720 (N_14720,N_14517,N_14420);
and U14721 (N_14721,N_14485,N_14456);
xnor U14722 (N_14722,N_14548,N_14513);
and U14723 (N_14723,N_14443,N_14580);
nor U14724 (N_14724,N_14496,N_14519);
xor U14725 (N_14725,N_14457,N_14435);
nand U14726 (N_14726,N_14497,N_14499);
or U14727 (N_14727,N_14578,N_14403);
nand U14728 (N_14728,N_14407,N_14405);
or U14729 (N_14729,N_14514,N_14418);
or U14730 (N_14730,N_14526,N_14414);
nor U14731 (N_14731,N_14471,N_14527);
or U14732 (N_14732,N_14513,N_14512);
nand U14733 (N_14733,N_14576,N_14483);
xor U14734 (N_14734,N_14464,N_14404);
nand U14735 (N_14735,N_14494,N_14491);
nor U14736 (N_14736,N_14586,N_14441);
nand U14737 (N_14737,N_14419,N_14421);
nand U14738 (N_14738,N_14404,N_14403);
nand U14739 (N_14739,N_14515,N_14418);
or U14740 (N_14740,N_14591,N_14484);
nor U14741 (N_14741,N_14438,N_14519);
and U14742 (N_14742,N_14404,N_14418);
xnor U14743 (N_14743,N_14572,N_14584);
nand U14744 (N_14744,N_14548,N_14516);
xnor U14745 (N_14745,N_14585,N_14446);
or U14746 (N_14746,N_14411,N_14471);
and U14747 (N_14747,N_14566,N_14496);
and U14748 (N_14748,N_14565,N_14570);
or U14749 (N_14749,N_14574,N_14454);
nand U14750 (N_14750,N_14590,N_14426);
nand U14751 (N_14751,N_14511,N_14564);
nor U14752 (N_14752,N_14582,N_14460);
xnor U14753 (N_14753,N_14485,N_14516);
or U14754 (N_14754,N_14561,N_14420);
xor U14755 (N_14755,N_14400,N_14543);
nor U14756 (N_14756,N_14577,N_14589);
and U14757 (N_14757,N_14419,N_14525);
or U14758 (N_14758,N_14425,N_14458);
xor U14759 (N_14759,N_14517,N_14472);
nor U14760 (N_14760,N_14409,N_14522);
nand U14761 (N_14761,N_14454,N_14513);
and U14762 (N_14762,N_14549,N_14436);
nor U14763 (N_14763,N_14439,N_14596);
nand U14764 (N_14764,N_14586,N_14405);
and U14765 (N_14765,N_14598,N_14413);
or U14766 (N_14766,N_14495,N_14537);
xnor U14767 (N_14767,N_14542,N_14465);
and U14768 (N_14768,N_14432,N_14506);
xor U14769 (N_14769,N_14449,N_14408);
nand U14770 (N_14770,N_14577,N_14501);
nor U14771 (N_14771,N_14473,N_14551);
and U14772 (N_14772,N_14585,N_14410);
nor U14773 (N_14773,N_14495,N_14474);
and U14774 (N_14774,N_14489,N_14408);
and U14775 (N_14775,N_14426,N_14455);
xnor U14776 (N_14776,N_14436,N_14524);
or U14777 (N_14777,N_14583,N_14498);
or U14778 (N_14778,N_14517,N_14499);
xor U14779 (N_14779,N_14559,N_14518);
and U14780 (N_14780,N_14495,N_14435);
and U14781 (N_14781,N_14487,N_14436);
and U14782 (N_14782,N_14403,N_14522);
nor U14783 (N_14783,N_14456,N_14409);
and U14784 (N_14784,N_14449,N_14458);
xor U14785 (N_14785,N_14437,N_14563);
nor U14786 (N_14786,N_14417,N_14436);
nor U14787 (N_14787,N_14530,N_14432);
nor U14788 (N_14788,N_14553,N_14495);
xor U14789 (N_14789,N_14563,N_14567);
nand U14790 (N_14790,N_14423,N_14593);
and U14791 (N_14791,N_14493,N_14588);
nand U14792 (N_14792,N_14572,N_14507);
and U14793 (N_14793,N_14487,N_14476);
xnor U14794 (N_14794,N_14577,N_14437);
xnor U14795 (N_14795,N_14512,N_14560);
and U14796 (N_14796,N_14482,N_14528);
xnor U14797 (N_14797,N_14572,N_14451);
xor U14798 (N_14798,N_14458,N_14535);
or U14799 (N_14799,N_14476,N_14546);
nor U14800 (N_14800,N_14689,N_14690);
and U14801 (N_14801,N_14748,N_14738);
xor U14802 (N_14802,N_14661,N_14728);
and U14803 (N_14803,N_14706,N_14607);
nand U14804 (N_14804,N_14609,N_14633);
nor U14805 (N_14805,N_14737,N_14688);
or U14806 (N_14806,N_14751,N_14641);
or U14807 (N_14807,N_14637,N_14698);
or U14808 (N_14808,N_14611,N_14701);
nor U14809 (N_14809,N_14600,N_14775);
nor U14810 (N_14810,N_14782,N_14789);
or U14811 (N_14811,N_14790,N_14615);
nor U14812 (N_14812,N_14765,N_14735);
and U14813 (N_14813,N_14753,N_14696);
nor U14814 (N_14814,N_14713,N_14608);
nand U14815 (N_14815,N_14645,N_14705);
or U14816 (N_14816,N_14653,N_14792);
nor U14817 (N_14817,N_14648,N_14684);
xor U14818 (N_14818,N_14752,N_14694);
or U14819 (N_14819,N_14783,N_14642);
nor U14820 (N_14820,N_14716,N_14750);
xor U14821 (N_14821,N_14766,N_14614);
and U14822 (N_14822,N_14736,N_14606);
nand U14823 (N_14823,N_14733,N_14715);
and U14824 (N_14824,N_14691,N_14649);
xor U14825 (N_14825,N_14763,N_14612);
and U14826 (N_14826,N_14676,N_14699);
xnor U14827 (N_14827,N_14764,N_14620);
nand U14828 (N_14828,N_14788,N_14680);
nand U14829 (N_14829,N_14669,N_14628);
nor U14830 (N_14830,N_14650,N_14762);
nor U14831 (N_14831,N_14602,N_14670);
xor U14832 (N_14832,N_14796,N_14663);
nand U14833 (N_14833,N_14719,N_14786);
nor U14834 (N_14834,N_14603,N_14732);
nor U14835 (N_14835,N_14709,N_14671);
nor U14836 (N_14836,N_14665,N_14793);
and U14837 (N_14837,N_14655,N_14779);
nor U14838 (N_14838,N_14714,N_14743);
or U14839 (N_14839,N_14652,N_14756);
nor U14840 (N_14840,N_14659,N_14619);
nor U14841 (N_14841,N_14629,N_14718);
nor U14842 (N_14842,N_14668,N_14780);
nand U14843 (N_14843,N_14700,N_14730);
nand U14844 (N_14844,N_14623,N_14695);
nand U14845 (N_14845,N_14729,N_14749);
nor U14846 (N_14846,N_14794,N_14744);
or U14847 (N_14847,N_14767,N_14672);
nor U14848 (N_14848,N_14654,N_14673);
or U14849 (N_14849,N_14674,N_14631);
nand U14850 (N_14850,N_14682,N_14687);
xor U14851 (N_14851,N_14664,N_14708);
xor U14852 (N_14852,N_14679,N_14703);
xor U14853 (N_14853,N_14784,N_14635);
nor U14854 (N_14854,N_14772,N_14683);
xor U14855 (N_14855,N_14771,N_14660);
nor U14856 (N_14856,N_14723,N_14798);
or U14857 (N_14857,N_14605,N_14754);
or U14858 (N_14858,N_14702,N_14617);
nor U14859 (N_14859,N_14740,N_14795);
nand U14860 (N_14860,N_14725,N_14681);
nor U14861 (N_14861,N_14746,N_14638);
nand U14862 (N_14862,N_14624,N_14797);
xor U14863 (N_14863,N_14651,N_14710);
and U14864 (N_14864,N_14722,N_14761);
nor U14865 (N_14865,N_14678,N_14768);
and U14866 (N_14866,N_14776,N_14757);
nor U14867 (N_14867,N_14711,N_14777);
and U14868 (N_14868,N_14785,N_14781);
nor U14869 (N_14869,N_14717,N_14656);
nor U14870 (N_14870,N_14747,N_14646);
nand U14871 (N_14871,N_14739,N_14760);
xor U14872 (N_14872,N_14704,N_14741);
nand U14873 (N_14873,N_14657,N_14644);
nor U14874 (N_14874,N_14787,N_14675);
nor U14875 (N_14875,N_14758,N_14692);
or U14876 (N_14876,N_14634,N_14625);
and U14877 (N_14877,N_14724,N_14697);
and U14878 (N_14878,N_14616,N_14791);
nor U14879 (N_14879,N_14770,N_14677);
nand U14880 (N_14880,N_14636,N_14742);
nand U14881 (N_14881,N_14769,N_14621);
or U14882 (N_14882,N_14774,N_14618);
nand U14883 (N_14883,N_14727,N_14632);
and U14884 (N_14884,N_14627,N_14693);
and U14885 (N_14885,N_14726,N_14712);
xnor U14886 (N_14886,N_14755,N_14799);
and U14887 (N_14887,N_14630,N_14666);
nor U14888 (N_14888,N_14731,N_14610);
nor U14889 (N_14889,N_14613,N_14662);
nor U14890 (N_14890,N_14745,N_14601);
and U14891 (N_14891,N_14667,N_14707);
nand U14892 (N_14892,N_14604,N_14647);
or U14893 (N_14893,N_14759,N_14720);
or U14894 (N_14894,N_14626,N_14658);
or U14895 (N_14895,N_14773,N_14640);
nand U14896 (N_14896,N_14639,N_14685);
and U14897 (N_14897,N_14643,N_14778);
or U14898 (N_14898,N_14721,N_14734);
nor U14899 (N_14899,N_14622,N_14686);
or U14900 (N_14900,N_14785,N_14644);
xnor U14901 (N_14901,N_14703,N_14610);
or U14902 (N_14902,N_14702,N_14788);
or U14903 (N_14903,N_14686,N_14714);
nand U14904 (N_14904,N_14602,N_14732);
nor U14905 (N_14905,N_14709,N_14613);
nand U14906 (N_14906,N_14776,N_14606);
xor U14907 (N_14907,N_14687,N_14797);
nand U14908 (N_14908,N_14697,N_14631);
nand U14909 (N_14909,N_14767,N_14738);
xnor U14910 (N_14910,N_14780,N_14792);
nor U14911 (N_14911,N_14737,N_14650);
xor U14912 (N_14912,N_14755,N_14650);
or U14913 (N_14913,N_14635,N_14656);
or U14914 (N_14914,N_14617,N_14649);
nand U14915 (N_14915,N_14703,N_14657);
and U14916 (N_14916,N_14734,N_14751);
nand U14917 (N_14917,N_14784,N_14723);
xor U14918 (N_14918,N_14671,N_14678);
or U14919 (N_14919,N_14618,N_14711);
nand U14920 (N_14920,N_14604,N_14607);
or U14921 (N_14921,N_14611,N_14773);
or U14922 (N_14922,N_14651,N_14727);
and U14923 (N_14923,N_14616,N_14619);
or U14924 (N_14924,N_14792,N_14683);
xnor U14925 (N_14925,N_14638,N_14656);
xor U14926 (N_14926,N_14621,N_14624);
xor U14927 (N_14927,N_14719,N_14669);
and U14928 (N_14928,N_14692,N_14634);
or U14929 (N_14929,N_14799,N_14785);
xor U14930 (N_14930,N_14691,N_14607);
nor U14931 (N_14931,N_14669,N_14699);
nand U14932 (N_14932,N_14677,N_14702);
xnor U14933 (N_14933,N_14687,N_14741);
nor U14934 (N_14934,N_14665,N_14718);
xnor U14935 (N_14935,N_14678,N_14659);
xor U14936 (N_14936,N_14704,N_14728);
nor U14937 (N_14937,N_14650,N_14793);
nor U14938 (N_14938,N_14740,N_14726);
and U14939 (N_14939,N_14658,N_14600);
xor U14940 (N_14940,N_14777,N_14675);
nand U14941 (N_14941,N_14717,N_14678);
or U14942 (N_14942,N_14662,N_14706);
xnor U14943 (N_14943,N_14675,N_14721);
nor U14944 (N_14944,N_14720,N_14631);
xnor U14945 (N_14945,N_14694,N_14683);
xor U14946 (N_14946,N_14732,N_14649);
xor U14947 (N_14947,N_14638,N_14681);
nand U14948 (N_14948,N_14608,N_14609);
nor U14949 (N_14949,N_14787,N_14781);
xor U14950 (N_14950,N_14611,N_14757);
or U14951 (N_14951,N_14642,N_14676);
or U14952 (N_14952,N_14600,N_14630);
and U14953 (N_14953,N_14676,N_14691);
or U14954 (N_14954,N_14784,N_14672);
and U14955 (N_14955,N_14651,N_14617);
xor U14956 (N_14956,N_14689,N_14620);
xor U14957 (N_14957,N_14721,N_14749);
and U14958 (N_14958,N_14766,N_14749);
and U14959 (N_14959,N_14741,N_14787);
xnor U14960 (N_14960,N_14621,N_14651);
nor U14961 (N_14961,N_14644,N_14635);
nor U14962 (N_14962,N_14614,N_14667);
or U14963 (N_14963,N_14764,N_14627);
xor U14964 (N_14964,N_14623,N_14631);
nand U14965 (N_14965,N_14735,N_14712);
nand U14966 (N_14966,N_14769,N_14614);
nor U14967 (N_14967,N_14732,N_14693);
nand U14968 (N_14968,N_14761,N_14667);
nor U14969 (N_14969,N_14716,N_14688);
and U14970 (N_14970,N_14605,N_14718);
nand U14971 (N_14971,N_14683,N_14749);
nor U14972 (N_14972,N_14786,N_14745);
or U14973 (N_14973,N_14614,N_14753);
nor U14974 (N_14974,N_14691,N_14761);
nand U14975 (N_14975,N_14738,N_14673);
and U14976 (N_14976,N_14670,N_14633);
or U14977 (N_14977,N_14729,N_14747);
xor U14978 (N_14978,N_14608,N_14747);
nand U14979 (N_14979,N_14797,N_14772);
nand U14980 (N_14980,N_14796,N_14702);
xor U14981 (N_14981,N_14782,N_14753);
or U14982 (N_14982,N_14691,N_14609);
xor U14983 (N_14983,N_14628,N_14733);
xor U14984 (N_14984,N_14681,N_14639);
nor U14985 (N_14985,N_14721,N_14708);
xnor U14986 (N_14986,N_14750,N_14652);
nor U14987 (N_14987,N_14770,N_14640);
nor U14988 (N_14988,N_14743,N_14657);
nor U14989 (N_14989,N_14671,N_14665);
and U14990 (N_14990,N_14753,N_14642);
nor U14991 (N_14991,N_14604,N_14635);
xor U14992 (N_14992,N_14680,N_14692);
or U14993 (N_14993,N_14782,N_14665);
or U14994 (N_14994,N_14738,N_14601);
xnor U14995 (N_14995,N_14600,N_14744);
nand U14996 (N_14996,N_14763,N_14647);
nor U14997 (N_14997,N_14706,N_14612);
nor U14998 (N_14998,N_14619,N_14724);
nor U14999 (N_14999,N_14683,N_14606);
xnor U15000 (N_15000,N_14990,N_14930);
and U15001 (N_15001,N_14850,N_14981);
and U15002 (N_15002,N_14826,N_14817);
and U15003 (N_15003,N_14909,N_14805);
or U15004 (N_15004,N_14941,N_14828);
nor U15005 (N_15005,N_14814,N_14873);
and U15006 (N_15006,N_14834,N_14924);
and U15007 (N_15007,N_14988,N_14951);
xnor U15008 (N_15008,N_14827,N_14907);
xor U15009 (N_15009,N_14878,N_14986);
or U15010 (N_15010,N_14855,N_14995);
nor U15011 (N_15011,N_14962,N_14892);
nor U15012 (N_15012,N_14838,N_14932);
nor U15013 (N_15013,N_14968,N_14852);
nor U15014 (N_15014,N_14865,N_14920);
xor U15015 (N_15015,N_14959,N_14969);
xor U15016 (N_15016,N_14897,N_14845);
xor U15017 (N_15017,N_14934,N_14812);
nand U15018 (N_15018,N_14862,N_14867);
nor U15019 (N_15019,N_14877,N_14872);
nor U15020 (N_15020,N_14844,N_14821);
and U15021 (N_15021,N_14957,N_14960);
and U15022 (N_15022,N_14996,N_14964);
xnor U15023 (N_15023,N_14980,N_14836);
xnor U15024 (N_15024,N_14938,N_14992);
nand U15025 (N_15025,N_14857,N_14880);
nand U15026 (N_15026,N_14854,N_14953);
or U15027 (N_15027,N_14984,N_14918);
xnor U15028 (N_15028,N_14835,N_14853);
or U15029 (N_15029,N_14816,N_14856);
nor U15030 (N_15030,N_14923,N_14888);
xor U15031 (N_15031,N_14802,N_14985);
or U15032 (N_15032,N_14917,N_14851);
or U15033 (N_15033,N_14848,N_14913);
and U15034 (N_15034,N_14824,N_14815);
xnor U15035 (N_15035,N_14806,N_14931);
or U15036 (N_15036,N_14879,N_14868);
or U15037 (N_15037,N_14894,N_14881);
nor U15038 (N_15038,N_14900,N_14846);
and U15039 (N_15039,N_14808,N_14874);
or U15040 (N_15040,N_14961,N_14978);
nor U15041 (N_15041,N_14926,N_14803);
or U15042 (N_15042,N_14963,N_14983);
or U15043 (N_15043,N_14970,N_14809);
nor U15044 (N_15044,N_14993,N_14869);
or U15045 (N_15045,N_14893,N_14940);
xnor U15046 (N_15046,N_14936,N_14921);
nand U15047 (N_15047,N_14819,N_14820);
nor U15048 (N_15048,N_14883,N_14863);
or U15049 (N_15049,N_14870,N_14991);
and U15050 (N_15050,N_14947,N_14801);
nor U15051 (N_15051,N_14825,N_14840);
or U15052 (N_15052,N_14967,N_14974);
nand U15053 (N_15053,N_14823,N_14939);
and U15054 (N_15054,N_14989,N_14858);
or U15055 (N_15055,N_14911,N_14837);
or U15056 (N_15056,N_14998,N_14922);
nor U15057 (N_15057,N_14833,N_14979);
nand U15058 (N_15058,N_14908,N_14891);
or U15059 (N_15059,N_14914,N_14800);
nor U15060 (N_15060,N_14899,N_14842);
nand U15061 (N_15061,N_14956,N_14860);
nor U15062 (N_15062,N_14935,N_14876);
xor U15063 (N_15063,N_14927,N_14937);
and U15064 (N_15064,N_14866,N_14919);
xnor U15065 (N_15065,N_14952,N_14902);
or U15066 (N_15066,N_14889,N_14822);
nand U15067 (N_15067,N_14955,N_14942);
and U15068 (N_15068,N_14906,N_14977);
or U15069 (N_15069,N_14903,N_14829);
nor U15070 (N_15070,N_14949,N_14886);
or U15071 (N_15071,N_14975,N_14841);
or U15072 (N_15072,N_14948,N_14915);
nand U15073 (N_15073,N_14813,N_14925);
xor U15074 (N_15074,N_14896,N_14933);
or U15075 (N_15075,N_14861,N_14832);
xor U15076 (N_15076,N_14944,N_14849);
nand U15077 (N_15077,N_14811,N_14972);
nand U15078 (N_15078,N_14839,N_14898);
nand U15079 (N_15079,N_14904,N_14982);
and U15080 (N_15080,N_14966,N_14958);
nor U15081 (N_15081,N_14987,N_14994);
xor U15082 (N_15082,N_14895,N_14831);
and U15083 (N_15083,N_14916,N_14875);
nor U15084 (N_15084,N_14804,N_14830);
or U15085 (N_15085,N_14954,N_14971);
or U15086 (N_15086,N_14928,N_14871);
xnor U15087 (N_15087,N_14818,N_14999);
nor U15088 (N_15088,N_14843,N_14810);
and U15089 (N_15089,N_14887,N_14890);
nor U15090 (N_15090,N_14910,N_14864);
nand U15091 (N_15091,N_14946,N_14929);
or U15092 (N_15092,N_14905,N_14973);
nor U15093 (N_15093,N_14965,N_14976);
xor U15094 (N_15094,N_14943,N_14885);
nand U15095 (N_15095,N_14884,N_14859);
or U15096 (N_15096,N_14847,N_14882);
and U15097 (N_15097,N_14997,N_14950);
and U15098 (N_15098,N_14945,N_14901);
nand U15099 (N_15099,N_14807,N_14912);
nor U15100 (N_15100,N_14970,N_14873);
or U15101 (N_15101,N_14947,N_14919);
nand U15102 (N_15102,N_14993,N_14910);
or U15103 (N_15103,N_14985,N_14941);
nand U15104 (N_15104,N_14815,N_14935);
xor U15105 (N_15105,N_14815,N_14878);
xor U15106 (N_15106,N_14964,N_14959);
nand U15107 (N_15107,N_14977,N_14883);
nor U15108 (N_15108,N_14933,N_14829);
xor U15109 (N_15109,N_14982,N_14886);
or U15110 (N_15110,N_14911,N_14826);
and U15111 (N_15111,N_14800,N_14960);
or U15112 (N_15112,N_14961,N_14936);
nor U15113 (N_15113,N_14860,N_14821);
nand U15114 (N_15114,N_14993,N_14828);
and U15115 (N_15115,N_14869,N_14969);
nand U15116 (N_15116,N_14822,N_14873);
xnor U15117 (N_15117,N_14931,N_14856);
nand U15118 (N_15118,N_14882,N_14839);
nand U15119 (N_15119,N_14894,N_14855);
nand U15120 (N_15120,N_14991,N_14819);
and U15121 (N_15121,N_14807,N_14874);
and U15122 (N_15122,N_14952,N_14809);
and U15123 (N_15123,N_14836,N_14930);
and U15124 (N_15124,N_14880,N_14877);
nand U15125 (N_15125,N_14835,N_14843);
and U15126 (N_15126,N_14952,N_14931);
and U15127 (N_15127,N_14807,N_14820);
xor U15128 (N_15128,N_14909,N_14835);
nor U15129 (N_15129,N_14987,N_14810);
and U15130 (N_15130,N_14839,N_14911);
nor U15131 (N_15131,N_14840,N_14811);
or U15132 (N_15132,N_14872,N_14917);
or U15133 (N_15133,N_14814,N_14872);
or U15134 (N_15134,N_14843,N_14820);
or U15135 (N_15135,N_14989,N_14883);
and U15136 (N_15136,N_14900,N_14988);
nand U15137 (N_15137,N_14840,N_14834);
and U15138 (N_15138,N_14841,N_14981);
nand U15139 (N_15139,N_14818,N_14834);
or U15140 (N_15140,N_14926,N_14869);
nor U15141 (N_15141,N_14854,N_14906);
nand U15142 (N_15142,N_14890,N_14990);
or U15143 (N_15143,N_14938,N_14804);
nand U15144 (N_15144,N_14821,N_14902);
and U15145 (N_15145,N_14924,N_14829);
and U15146 (N_15146,N_14918,N_14897);
nand U15147 (N_15147,N_14859,N_14865);
nand U15148 (N_15148,N_14805,N_14955);
nand U15149 (N_15149,N_14941,N_14819);
nor U15150 (N_15150,N_14950,N_14831);
nand U15151 (N_15151,N_14824,N_14958);
and U15152 (N_15152,N_14922,N_14902);
and U15153 (N_15153,N_14975,N_14980);
nand U15154 (N_15154,N_14921,N_14812);
xor U15155 (N_15155,N_14811,N_14964);
nand U15156 (N_15156,N_14928,N_14872);
or U15157 (N_15157,N_14975,N_14877);
nand U15158 (N_15158,N_14901,N_14827);
xor U15159 (N_15159,N_14822,N_14870);
nand U15160 (N_15160,N_14877,N_14937);
xor U15161 (N_15161,N_14947,N_14913);
and U15162 (N_15162,N_14926,N_14905);
or U15163 (N_15163,N_14974,N_14851);
or U15164 (N_15164,N_14882,N_14812);
and U15165 (N_15165,N_14816,N_14984);
xnor U15166 (N_15166,N_14830,N_14825);
nor U15167 (N_15167,N_14832,N_14880);
nand U15168 (N_15168,N_14885,N_14959);
nand U15169 (N_15169,N_14943,N_14820);
nor U15170 (N_15170,N_14897,N_14844);
or U15171 (N_15171,N_14828,N_14827);
or U15172 (N_15172,N_14927,N_14824);
xnor U15173 (N_15173,N_14970,N_14949);
or U15174 (N_15174,N_14982,N_14898);
and U15175 (N_15175,N_14859,N_14923);
nor U15176 (N_15176,N_14946,N_14965);
nand U15177 (N_15177,N_14830,N_14813);
nor U15178 (N_15178,N_14944,N_14934);
and U15179 (N_15179,N_14876,N_14809);
or U15180 (N_15180,N_14808,N_14922);
or U15181 (N_15181,N_14942,N_14883);
xor U15182 (N_15182,N_14818,N_14821);
xor U15183 (N_15183,N_14827,N_14871);
nand U15184 (N_15184,N_14933,N_14934);
and U15185 (N_15185,N_14956,N_14835);
and U15186 (N_15186,N_14930,N_14813);
nor U15187 (N_15187,N_14895,N_14890);
or U15188 (N_15188,N_14889,N_14960);
xnor U15189 (N_15189,N_14971,N_14943);
xnor U15190 (N_15190,N_14896,N_14811);
and U15191 (N_15191,N_14855,N_14821);
nand U15192 (N_15192,N_14959,N_14838);
nand U15193 (N_15193,N_14978,N_14901);
nand U15194 (N_15194,N_14919,N_14954);
and U15195 (N_15195,N_14948,N_14849);
nand U15196 (N_15196,N_14974,N_14861);
nor U15197 (N_15197,N_14979,N_14828);
or U15198 (N_15198,N_14877,N_14961);
or U15199 (N_15199,N_14892,N_14956);
nand U15200 (N_15200,N_15108,N_15153);
nand U15201 (N_15201,N_15087,N_15188);
xnor U15202 (N_15202,N_15023,N_15024);
nor U15203 (N_15203,N_15102,N_15010);
or U15204 (N_15204,N_15114,N_15140);
xnor U15205 (N_15205,N_15058,N_15062);
xor U15206 (N_15206,N_15176,N_15131);
nand U15207 (N_15207,N_15029,N_15044);
xnor U15208 (N_15208,N_15132,N_15015);
xnor U15209 (N_15209,N_15152,N_15118);
nand U15210 (N_15210,N_15097,N_15175);
nand U15211 (N_15211,N_15103,N_15060);
or U15212 (N_15212,N_15159,N_15178);
nor U15213 (N_15213,N_15122,N_15196);
nand U15214 (N_15214,N_15038,N_15170);
nor U15215 (N_15215,N_15162,N_15180);
nor U15216 (N_15216,N_15068,N_15027);
and U15217 (N_15217,N_15005,N_15107);
nor U15218 (N_15218,N_15165,N_15158);
nor U15219 (N_15219,N_15066,N_15173);
nor U15220 (N_15220,N_15112,N_15128);
and U15221 (N_15221,N_15033,N_15148);
or U15222 (N_15222,N_15046,N_15021);
or U15223 (N_15223,N_15047,N_15067);
and U15224 (N_15224,N_15077,N_15166);
and U15225 (N_15225,N_15056,N_15028);
nor U15226 (N_15226,N_15111,N_15126);
xnor U15227 (N_15227,N_15019,N_15093);
xor U15228 (N_15228,N_15041,N_15163);
nand U15229 (N_15229,N_15187,N_15115);
xnor U15230 (N_15230,N_15133,N_15013);
nor U15231 (N_15231,N_15138,N_15117);
and U15232 (N_15232,N_15141,N_15052);
and U15233 (N_15233,N_15098,N_15048);
and U15234 (N_15234,N_15084,N_15139);
and U15235 (N_15235,N_15150,N_15085);
nand U15236 (N_15236,N_15185,N_15151);
or U15237 (N_15237,N_15104,N_15020);
nor U15238 (N_15238,N_15080,N_15168);
xor U15239 (N_15239,N_15040,N_15161);
or U15240 (N_15240,N_15078,N_15130);
nand U15241 (N_15241,N_15169,N_15149);
nand U15242 (N_15242,N_15094,N_15183);
and U15243 (N_15243,N_15042,N_15039);
and U15244 (N_15244,N_15069,N_15123);
or U15245 (N_15245,N_15120,N_15092);
nor U15246 (N_15246,N_15177,N_15003);
nand U15247 (N_15247,N_15086,N_15194);
or U15248 (N_15248,N_15171,N_15125);
xor U15249 (N_15249,N_15006,N_15025);
nand U15250 (N_15250,N_15018,N_15109);
or U15251 (N_15251,N_15053,N_15106);
or U15252 (N_15252,N_15026,N_15037);
xnor U15253 (N_15253,N_15129,N_15195);
xor U15254 (N_15254,N_15030,N_15070);
or U15255 (N_15255,N_15082,N_15181);
xor U15256 (N_15256,N_15049,N_15124);
and U15257 (N_15257,N_15009,N_15096);
nand U15258 (N_15258,N_15014,N_15136);
and U15259 (N_15259,N_15075,N_15121);
xor U15260 (N_15260,N_15184,N_15045);
and U15261 (N_15261,N_15190,N_15011);
nor U15262 (N_15262,N_15189,N_15105);
and U15263 (N_15263,N_15000,N_15007);
nand U15264 (N_15264,N_15182,N_15101);
or U15265 (N_15265,N_15032,N_15100);
nand U15266 (N_15266,N_15160,N_15031);
xor U15267 (N_15267,N_15065,N_15193);
and U15268 (N_15268,N_15147,N_15074);
nand U15269 (N_15269,N_15008,N_15076);
or U15270 (N_15270,N_15017,N_15157);
or U15271 (N_15271,N_15199,N_15002);
nor U15272 (N_15272,N_15034,N_15051);
and U15273 (N_15273,N_15089,N_15146);
or U15274 (N_15274,N_15036,N_15119);
or U15275 (N_15275,N_15197,N_15135);
or U15276 (N_15276,N_15144,N_15063);
nand U15277 (N_15277,N_15154,N_15088);
or U15278 (N_15278,N_15155,N_15116);
and U15279 (N_15279,N_15061,N_15016);
and U15280 (N_15280,N_15050,N_15143);
nor U15281 (N_15281,N_15137,N_15057);
and U15282 (N_15282,N_15172,N_15073);
and U15283 (N_15283,N_15095,N_15145);
nor U15284 (N_15284,N_15055,N_15127);
xnor U15285 (N_15285,N_15079,N_15186);
and U15286 (N_15286,N_15179,N_15164);
or U15287 (N_15287,N_15156,N_15099);
xnor U15288 (N_15288,N_15090,N_15001);
xnor U15289 (N_15289,N_15174,N_15192);
xnor U15290 (N_15290,N_15198,N_15167);
and U15291 (N_15291,N_15191,N_15043);
or U15292 (N_15292,N_15091,N_15134);
and U15293 (N_15293,N_15110,N_15113);
xor U15294 (N_15294,N_15064,N_15081);
and U15295 (N_15295,N_15083,N_15054);
nor U15296 (N_15296,N_15004,N_15071);
or U15297 (N_15297,N_15012,N_15059);
nand U15298 (N_15298,N_15142,N_15072);
xnor U15299 (N_15299,N_15035,N_15022);
xnor U15300 (N_15300,N_15050,N_15170);
and U15301 (N_15301,N_15176,N_15034);
or U15302 (N_15302,N_15022,N_15183);
xor U15303 (N_15303,N_15148,N_15166);
or U15304 (N_15304,N_15196,N_15040);
and U15305 (N_15305,N_15021,N_15078);
and U15306 (N_15306,N_15133,N_15179);
nor U15307 (N_15307,N_15079,N_15116);
xor U15308 (N_15308,N_15083,N_15185);
xor U15309 (N_15309,N_15148,N_15124);
and U15310 (N_15310,N_15178,N_15143);
nor U15311 (N_15311,N_15188,N_15004);
or U15312 (N_15312,N_15106,N_15176);
nand U15313 (N_15313,N_15083,N_15146);
nor U15314 (N_15314,N_15163,N_15051);
or U15315 (N_15315,N_15053,N_15092);
nor U15316 (N_15316,N_15105,N_15035);
nand U15317 (N_15317,N_15119,N_15066);
xnor U15318 (N_15318,N_15007,N_15081);
or U15319 (N_15319,N_15121,N_15067);
or U15320 (N_15320,N_15012,N_15099);
or U15321 (N_15321,N_15019,N_15098);
nand U15322 (N_15322,N_15011,N_15070);
xor U15323 (N_15323,N_15068,N_15183);
or U15324 (N_15324,N_15182,N_15040);
and U15325 (N_15325,N_15180,N_15002);
nand U15326 (N_15326,N_15084,N_15186);
and U15327 (N_15327,N_15121,N_15197);
or U15328 (N_15328,N_15067,N_15055);
nand U15329 (N_15329,N_15183,N_15121);
xnor U15330 (N_15330,N_15083,N_15148);
or U15331 (N_15331,N_15155,N_15052);
nand U15332 (N_15332,N_15123,N_15114);
or U15333 (N_15333,N_15185,N_15166);
and U15334 (N_15334,N_15038,N_15052);
or U15335 (N_15335,N_15004,N_15018);
xnor U15336 (N_15336,N_15038,N_15004);
nor U15337 (N_15337,N_15173,N_15108);
xnor U15338 (N_15338,N_15138,N_15091);
nor U15339 (N_15339,N_15042,N_15087);
and U15340 (N_15340,N_15017,N_15019);
xnor U15341 (N_15341,N_15131,N_15136);
nand U15342 (N_15342,N_15069,N_15028);
nor U15343 (N_15343,N_15195,N_15092);
or U15344 (N_15344,N_15093,N_15064);
xor U15345 (N_15345,N_15134,N_15132);
or U15346 (N_15346,N_15107,N_15184);
and U15347 (N_15347,N_15155,N_15042);
and U15348 (N_15348,N_15116,N_15173);
or U15349 (N_15349,N_15067,N_15079);
nor U15350 (N_15350,N_15127,N_15014);
xnor U15351 (N_15351,N_15070,N_15056);
or U15352 (N_15352,N_15119,N_15055);
xnor U15353 (N_15353,N_15187,N_15077);
or U15354 (N_15354,N_15122,N_15045);
or U15355 (N_15355,N_15022,N_15047);
or U15356 (N_15356,N_15065,N_15113);
xor U15357 (N_15357,N_15193,N_15138);
nand U15358 (N_15358,N_15031,N_15010);
and U15359 (N_15359,N_15014,N_15149);
xor U15360 (N_15360,N_15037,N_15094);
xor U15361 (N_15361,N_15134,N_15195);
and U15362 (N_15362,N_15087,N_15155);
xor U15363 (N_15363,N_15115,N_15156);
nor U15364 (N_15364,N_15187,N_15138);
nor U15365 (N_15365,N_15069,N_15174);
nor U15366 (N_15366,N_15082,N_15097);
xor U15367 (N_15367,N_15155,N_15102);
nor U15368 (N_15368,N_15181,N_15132);
nor U15369 (N_15369,N_15080,N_15111);
xnor U15370 (N_15370,N_15005,N_15154);
or U15371 (N_15371,N_15163,N_15155);
xnor U15372 (N_15372,N_15131,N_15078);
or U15373 (N_15373,N_15127,N_15098);
xnor U15374 (N_15374,N_15134,N_15085);
nor U15375 (N_15375,N_15185,N_15029);
nor U15376 (N_15376,N_15036,N_15086);
xor U15377 (N_15377,N_15162,N_15111);
nand U15378 (N_15378,N_15119,N_15155);
and U15379 (N_15379,N_15068,N_15010);
nand U15380 (N_15380,N_15133,N_15106);
or U15381 (N_15381,N_15191,N_15095);
or U15382 (N_15382,N_15109,N_15136);
nand U15383 (N_15383,N_15124,N_15131);
nand U15384 (N_15384,N_15065,N_15061);
xor U15385 (N_15385,N_15028,N_15038);
nand U15386 (N_15386,N_15177,N_15142);
nor U15387 (N_15387,N_15010,N_15082);
nand U15388 (N_15388,N_15176,N_15141);
nor U15389 (N_15389,N_15195,N_15012);
or U15390 (N_15390,N_15033,N_15093);
and U15391 (N_15391,N_15172,N_15111);
and U15392 (N_15392,N_15106,N_15179);
nor U15393 (N_15393,N_15172,N_15126);
nor U15394 (N_15394,N_15094,N_15079);
and U15395 (N_15395,N_15084,N_15013);
nand U15396 (N_15396,N_15182,N_15187);
nor U15397 (N_15397,N_15116,N_15081);
nand U15398 (N_15398,N_15072,N_15108);
xor U15399 (N_15399,N_15078,N_15014);
nor U15400 (N_15400,N_15282,N_15314);
xor U15401 (N_15401,N_15368,N_15238);
or U15402 (N_15402,N_15395,N_15394);
and U15403 (N_15403,N_15366,N_15256);
or U15404 (N_15404,N_15278,N_15398);
or U15405 (N_15405,N_15287,N_15353);
nand U15406 (N_15406,N_15369,N_15304);
or U15407 (N_15407,N_15355,N_15244);
and U15408 (N_15408,N_15214,N_15333);
xor U15409 (N_15409,N_15228,N_15266);
xor U15410 (N_15410,N_15286,N_15220);
and U15411 (N_15411,N_15272,N_15247);
or U15412 (N_15412,N_15391,N_15240);
nand U15413 (N_15413,N_15271,N_15281);
nand U15414 (N_15414,N_15312,N_15218);
and U15415 (N_15415,N_15237,N_15385);
or U15416 (N_15416,N_15322,N_15372);
and U15417 (N_15417,N_15248,N_15300);
nand U15418 (N_15418,N_15309,N_15345);
or U15419 (N_15419,N_15306,N_15340);
nand U15420 (N_15420,N_15359,N_15207);
xor U15421 (N_15421,N_15364,N_15202);
and U15422 (N_15422,N_15234,N_15362);
nor U15423 (N_15423,N_15283,N_15373);
or U15424 (N_15424,N_15386,N_15363);
and U15425 (N_15425,N_15379,N_15332);
nor U15426 (N_15426,N_15310,N_15260);
and U15427 (N_15427,N_15375,N_15224);
or U15428 (N_15428,N_15290,N_15239);
nand U15429 (N_15429,N_15251,N_15381);
nor U15430 (N_15430,N_15325,N_15273);
nor U15431 (N_15431,N_15201,N_15250);
nor U15432 (N_15432,N_15370,N_15219);
and U15433 (N_15433,N_15227,N_15280);
nor U15434 (N_15434,N_15261,N_15299);
and U15435 (N_15435,N_15213,N_15380);
xnor U15436 (N_15436,N_15377,N_15296);
and U15437 (N_15437,N_15285,N_15317);
and U15438 (N_15438,N_15324,N_15265);
xnor U15439 (N_15439,N_15230,N_15326);
and U15440 (N_15440,N_15242,N_15327);
or U15441 (N_15441,N_15390,N_15259);
and U15442 (N_15442,N_15216,N_15357);
and U15443 (N_15443,N_15222,N_15378);
xor U15444 (N_15444,N_15335,N_15307);
xor U15445 (N_15445,N_15245,N_15262);
nand U15446 (N_15446,N_15315,N_15305);
nand U15447 (N_15447,N_15293,N_15376);
nor U15448 (N_15448,N_15269,N_15204);
xor U15449 (N_15449,N_15252,N_15212);
nor U15450 (N_15450,N_15383,N_15288);
xor U15451 (N_15451,N_15387,N_15267);
and U15452 (N_15452,N_15263,N_15343);
nor U15453 (N_15453,N_15298,N_15399);
nand U15454 (N_15454,N_15336,N_15384);
or U15455 (N_15455,N_15257,N_15330);
nand U15456 (N_15456,N_15302,N_15389);
nand U15457 (N_15457,N_15253,N_15291);
nand U15458 (N_15458,N_15348,N_15374);
and U15459 (N_15459,N_15349,N_15270);
xnor U15460 (N_15460,N_15277,N_15241);
nor U15461 (N_15461,N_15208,N_15221);
nand U15462 (N_15462,N_15382,N_15276);
nor U15463 (N_15463,N_15354,N_15249);
nand U15464 (N_15464,N_15225,N_15279);
nand U15465 (N_15465,N_15297,N_15226);
xnor U15466 (N_15466,N_15331,N_15284);
nor U15467 (N_15467,N_15210,N_15223);
xnor U15468 (N_15468,N_15308,N_15255);
and U15469 (N_15469,N_15342,N_15209);
and U15470 (N_15470,N_15393,N_15352);
xnor U15471 (N_15471,N_15318,N_15231);
xnor U15472 (N_15472,N_15360,N_15320);
nand U15473 (N_15473,N_15346,N_15264);
or U15474 (N_15474,N_15396,N_15323);
or U15475 (N_15475,N_15350,N_15339);
xor U15476 (N_15476,N_15301,N_15367);
nand U15477 (N_15477,N_15258,N_15321);
or U15478 (N_15478,N_15217,N_15206);
and U15479 (N_15479,N_15356,N_15211);
xnor U15480 (N_15480,N_15254,N_15337);
or U15481 (N_15481,N_15294,N_15313);
nor U15482 (N_15482,N_15200,N_15338);
xnor U15483 (N_15483,N_15246,N_15347);
nand U15484 (N_15484,N_15397,N_15229);
or U15485 (N_15485,N_15236,N_15361);
and U15486 (N_15486,N_15295,N_15316);
nor U15487 (N_15487,N_15392,N_15235);
nand U15488 (N_15488,N_15388,N_15205);
nor U15489 (N_15489,N_15232,N_15289);
and U15490 (N_15490,N_15371,N_15334);
nor U15491 (N_15491,N_15329,N_15344);
or U15492 (N_15492,N_15351,N_15328);
nor U15493 (N_15493,N_15303,N_15311);
nor U15494 (N_15494,N_15233,N_15268);
xor U15495 (N_15495,N_15275,N_15243);
and U15496 (N_15496,N_15358,N_15319);
nor U15497 (N_15497,N_15365,N_15341);
nor U15498 (N_15498,N_15203,N_15292);
or U15499 (N_15499,N_15215,N_15274);
and U15500 (N_15500,N_15236,N_15216);
and U15501 (N_15501,N_15222,N_15225);
and U15502 (N_15502,N_15276,N_15324);
xnor U15503 (N_15503,N_15202,N_15200);
nand U15504 (N_15504,N_15385,N_15290);
nor U15505 (N_15505,N_15279,N_15258);
xnor U15506 (N_15506,N_15318,N_15222);
or U15507 (N_15507,N_15378,N_15204);
and U15508 (N_15508,N_15397,N_15244);
nand U15509 (N_15509,N_15251,N_15332);
or U15510 (N_15510,N_15261,N_15399);
or U15511 (N_15511,N_15327,N_15366);
and U15512 (N_15512,N_15344,N_15373);
nand U15513 (N_15513,N_15291,N_15293);
nor U15514 (N_15514,N_15247,N_15325);
or U15515 (N_15515,N_15339,N_15280);
nor U15516 (N_15516,N_15325,N_15292);
and U15517 (N_15517,N_15375,N_15321);
nor U15518 (N_15518,N_15303,N_15355);
nor U15519 (N_15519,N_15347,N_15391);
and U15520 (N_15520,N_15268,N_15274);
nand U15521 (N_15521,N_15337,N_15282);
nor U15522 (N_15522,N_15204,N_15386);
xor U15523 (N_15523,N_15245,N_15258);
and U15524 (N_15524,N_15205,N_15237);
nand U15525 (N_15525,N_15236,N_15224);
and U15526 (N_15526,N_15278,N_15319);
nor U15527 (N_15527,N_15397,N_15277);
and U15528 (N_15528,N_15335,N_15370);
and U15529 (N_15529,N_15259,N_15212);
or U15530 (N_15530,N_15354,N_15340);
or U15531 (N_15531,N_15217,N_15267);
and U15532 (N_15532,N_15236,N_15369);
and U15533 (N_15533,N_15265,N_15373);
xnor U15534 (N_15534,N_15393,N_15223);
nor U15535 (N_15535,N_15242,N_15378);
or U15536 (N_15536,N_15292,N_15372);
xor U15537 (N_15537,N_15333,N_15275);
xor U15538 (N_15538,N_15246,N_15224);
or U15539 (N_15539,N_15201,N_15242);
and U15540 (N_15540,N_15399,N_15306);
nand U15541 (N_15541,N_15227,N_15333);
nor U15542 (N_15542,N_15390,N_15362);
xnor U15543 (N_15543,N_15340,N_15310);
nor U15544 (N_15544,N_15275,N_15283);
nand U15545 (N_15545,N_15250,N_15298);
and U15546 (N_15546,N_15202,N_15373);
and U15547 (N_15547,N_15344,N_15260);
nor U15548 (N_15548,N_15381,N_15202);
nor U15549 (N_15549,N_15205,N_15395);
or U15550 (N_15550,N_15377,N_15300);
nand U15551 (N_15551,N_15343,N_15306);
or U15552 (N_15552,N_15202,N_15358);
nand U15553 (N_15553,N_15345,N_15249);
xor U15554 (N_15554,N_15323,N_15384);
and U15555 (N_15555,N_15363,N_15316);
nand U15556 (N_15556,N_15220,N_15294);
xor U15557 (N_15557,N_15337,N_15341);
or U15558 (N_15558,N_15240,N_15215);
nand U15559 (N_15559,N_15213,N_15334);
and U15560 (N_15560,N_15203,N_15216);
or U15561 (N_15561,N_15285,N_15257);
nand U15562 (N_15562,N_15380,N_15282);
nor U15563 (N_15563,N_15252,N_15329);
and U15564 (N_15564,N_15219,N_15302);
or U15565 (N_15565,N_15226,N_15322);
and U15566 (N_15566,N_15360,N_15230);
or U15567 (N_15567,N_15202,N_15372);
xor U15568 (N_15568,N_15369,N_15339);
nand U15569 (N_15569,N_15330,N_15214);
or U15570 (N_15570,N_15251,N_15327);
and U15571 (N_15571,N_15244,N_15388);
nor U15572 (N_15572,N_15370,N_15347);
xor U15573 (N_15573,N_15303,N_15307);
xor U15574 (N_15574,N_15327,N_15248);
and U15575 (N_15575,N_15311,N_15334);
nand U15576 (N_15576,N_15213,N_15336);
nand U15577 (N_15577,N_15253,N_15343);
or U15578 (N_15578,N_15308,N_15296);
nor U15579 (N_15579,N_15224,N_15311);
nor U15580 (N_15580,N_15247,N_15237);
and U15581 (N_15581,N_15375,N_15263);
and U15582 (N_15582,N_15219,N_15337);
and U15583 (N_15583,N_15305,N_15203);
nand U15584 (N_15584,N_15243,N_15294);
or U15585 (N_15585,N_15250,N_15324);
and U15586 (N_15586,N_15373,N_15316);
and U15587 (N_15587,N_15223,N_15341);
or U15588 (N_15588,N_15347,N_15249);
xor U15589 (N_15589,N_15342,N_15297);
or U15590 (N_15590,N_15249,N_15337);
nor U15591 (N_15591,N_15328,N_15297);
nand U15592 (N_15592,N_15219,N_15397);
nor U15593 (N_15593,N_15364,N_15376);
xor U15594 (N_15594,N_15217,N_15254);
nand U15595 (N_15595,N_15359,N_15334);
or U15596 (N_15596,N_15368,N_15272);
nand U15597 (N_15597,N_15322,N_15309);
xor U15598 (N_15598,N_15337,N_15247);
nand U15599 (N_15599,N_15292,N_15326);
and U15600 (N_15600,N_15460,N_15565);
and U15601 (N_15601,N_15439,N_15455);
nor U15602 (N_15602,N_15464,N_15427);
or U15603 (N_15603,N_15531,N_15471);
and U15604 (N_15604,N_15507,N_15503);
nand U15605 (N_15605,N_15418,N_15404);
nor U15606 (N_15606,N_15473,N_15413);
and U15607 (N_15607,N_15433,N_15533);
nor U15608 (N_15608,N_15461,N_15514);
nor U15609 (N_15609,N_15526,N_15478);
nor U15610 (N_15610,N_15434,N_15489);
nand U15611 (N_15611,N_15571,N_15578);
or U15612 (N_15612,N_15568,N_15538);
or U15613 (N_15613,N_15591,N_15562);
xnor U15614 (N_15614,N_15549,N_15415);
nand U15615 (N_15615,N_15414,N_15468);
or U15616 (N_15616,N_15465,N_15534);
or U15617 (N_15617,N_15444,N_15518);
nand U15618 (N_15618,N_15492,N_15546);
nor U15619 (N_15619,N_15522,N_15419);
or U15620 (N_15620,N_15457,N_15594);
and U15621 (N_15621,N_15564,N_15520);
and U15622 (N_15622,N_15490,N_15502);
and U15623 (N_15623,N_15596,N_15530);
and U15624 (N_15624,N_15482,N_15409);
nor U15625 (N_15625,N_15459,N_15437);
xnor U15626 (N_15626,N_15428,N_15481);
nand U15627 (N_15627,N_15550,N_15510);
xnor U15628 (N_15628,N_15528,N_15402);
and U15629 (N_15629,N_15424,N_15500);
or U15630 (N_15630,N_15488,N_15451);
or U15631 (N_15631,N_15569,N_15576);
nand U15632 (N_15632,N_15494,N_15421);
xnor U15633 (N_15633,N_15512,N_15506);
and U15634 (N_15634,N_15570,N_15430);
or U15635 (N_15635,N_15472,N_15560);
xnor U15636 (N_15636,N_15516,N_15475);
nor U15637 (N_15637,N_15498,N_15479);
or U15638 (N_15638,N_15499,N_15483);
nand U15639 (N_15639,N_15417,N_15599);
and U15640 (N_15640,N_15521,N_15448);
nand U15641 (N_15641,N_15412,N_15420);
nor U15642 (N_15642,N_15575,N_15524);
and U15643 (N_15643,N_15429,N_15504);
or U15644 (N_15644,N_15443,N_15519);
xor U15645 (N_15645,N_15441,N_15501);
or U15646 (N_15646,N_15541,N_15553);
xnor U15647 (N_15647,N_15497,N_15535);
xnor U15648 (N_15648,N_15410,N_15551);
and U15649 (N_15649,N_15480,N_15401);
nor U15650 (N_15650,N_15435,N_15505);
nand U15651 (N_15651,N_15496,N_15595);
nor U15652 (N_15652,N_15580,N_15563);
and U15653 (N_15653,N_15432,N_15508);
or U15654 (N_15654,N_15452,N_15540);
nand U15655 (N_15655,N_15423,N_15573);
or U15656 (N_15656,N_15405,N_15527);
or U15657 (N_15657,N_15467,N_15539);
or U15658 (N_15658,N_15511,N_15403);
or U15659 (N_15659,N_15436,N_15545);
xor U15660 (N_15660,N_15566,N_15487);
nor U15661 (N_15661,N_15583,N_15582);
xnor U15662 (N_15662,N_15552,N_15416);
or U15663 (N_15663,N_15556,N_15548);
nor U15664 (N_15664,N_15593,N_15588);
xor U15665 (N_15665,N_15598,N_15589);
or U15666 (N_15666,N_15581,N_15485);
and U15667 (N_15667,N_15529,N_15561);
and U15668 (N_15668,N_15400,N_15543);
nor U15669 (N_15669,N_15567,N_15585);
nor U15670 (N_15670,N_15513,N_15532);
and U15671 (N_15671,N_15584,N_15442);
nor U15672 (N_15672,N_15574,N_15446);
nand U15673 (N_15673,N_15542,N_15440);
nor U15674 (N_15674,N_15476,N_15597);
or U15675 (N_15675,N_15537,N_15557);
xnor U15676 (N_15676,N_15491,N_15450);
or U15677 (N_15677,N_15408,N_15453);
nor U15678 (N_15678,N_15462,N_15454);
nand U15679 (N_15679,N_15447,N_15525);
xnor U15680 (N_15680,N_15523,N_15592);
and U15681 (N_15681,N_15579,N_15463);
nand U15682 (N_15682,N_15559,N_15486);
and U15683 (N_15683,N_15572,N_15558);
nand U15684 (N_15684,N_15431,N_15466);
or U15685 (N_15685,N_15515,N_15426);
xor U15686 (N_15686,N_15445,N_15438);
or U15687 (N_15687,N_15411,N_15536);
xor U15688 (N_15688,N_15587,N_15458);
or U15689 (N_15689,N_15470,N_15544);
nand U15690 (N_15690,N_15469,N_15547);
and U15691 (N_15691,N_15449,N_15407);
xor U15692 (N_15692,N_15456,N_15484);
nand U15693 (N_15693,N_15493,N_15474);
nor U15694 (N_15694,N_15577,N_15425);
and U15695 (N_15695,N_15555,N_15590);
or U15696 (N_15696,N_15517,N_15495);
or U15697 (N_15697,N_15509,N_15422);
or U15698 (N_15698,N_15586,N_15477);
or U15699 (N_15699,N_15554,N_15406);
or U15700 (N_15700,N_15513,N_15515);
nor U15701 (N_15701,N_15461,N_15404);
nor U15702 (N_15702,N_15563,N_15541);
nor U15703 (N_15703,N_15447,N_15502);
and U15704 (N_15704,N_15590,N_15566);
or U15705 (N_15705,N_15475,N_15584);
and U15706 (N_15706,N_15415,N_15459);
nand U15707 (N_15707,N_15426,N_15597);
or U15708 (N_15708,N_15445,N_15572);
xor U15709 (N_15709,N_15589,N_15479);
xor U15710 (N_15710,N_15411,N_15596);
nand U15711 (N_15711,N_15413,N_15552);
nand U15712 (N_15712,N_15536,N_15551);
nor U15713 (N_15713,N_15523,N_15415);
nand U15714 (N_15714,N_15495,N_15405);
nor U15715 (N_15715,N_15510,N_15519);
xnor U15716 (N_15716,N_15591,N_15486);
nor U15717 (N_15717,N_15456,N_15523);
nor U15718 (N_15718,N_15571,N_15436);
nor U15719 (N_15719,N_15438,N_15466);
nor U15720 (N_15720,N_15569,N_15469);
nand U15721 (N_15721,N_15411,N_15482);
nand U15722 (N_15722,N_15406,N_15430);
or U15723 (N_15723,N_15481,N_15507);
or U15724 (N_15724,N_15565,N_15499);
xor U15725 (N_15725,N_15459,N_15593);
and U15726 (N_15726,N_15434,N_15541);
nor U15727 (N_15727,N_15437,N_15573);
or U15728 (N_15728,N_15554,N_15474);
and U15729 (N_15729,N_15423,N_15593);
and U15730 (N_15730,N_15551,N_15470);
and U15731 (N_15731,N_15428,N_15442);
nor U15732 (N_15732,N_15409,N_15517);
and U15733 (N_15733,N_15401,N_15516);
and U15734 (N_15734,N_15567,N_15590);
xnor U15735 (N_15735,N_15581,N_15575);
nand U15736 (N_15736,N_15513,N_15536);
and U15737 (N_15737,N_15519,N_15540);
nand U15738 (N_15738,N_15452,N_15551);
and U15739 (N_15739,N_15507,N_15529);
xor U15740 (N_15740,N_15580,N_15577);
or U15741 (N_15741,N_15518,N_15481);
nand U15742 (N_15742,N_15420,N_15527);
nand U15743 (N_15743,N_15503,N_15592);
or U15744 (N_15744,N_15455,N_15547);
xor U15745 (N_15745,N_15448,N_15519);
xnor U15746 (N_15746,N_15462,N_15405);
xnor U15747 (N_15747,N_15411,N_15571);
xor U15748 (N_15748,N_15468,N_15535);
xor U15749 (N_15749,N_15477,N_15543);
nand U15750 (N_15750,N_15471,N_15422);
nand U15751 (N_15751,N_15566,N_15589);
nor U15752 (N_15752,N_15516,N_15451);
nor U15753 (N_15753,N_15563,N_15443);
and U15754 (N_15754,N_15420,N_15405);
or U15755 (N_15755,N_15568,N_15416);
or U15756 (N_15756,N_15451,N_15526);
nor U15757 (N_15757,N_15453,N_15465);
and U15758 (N_15758,N_15437,N_15598);
nand U15759 (N_15759,N_15563,N_15428);
nand U15760 (N_15760,N_15410,N_15541);
xor U15761 (N_15761,N_15437,N_15540);
or U15762 (N_15762,N_15537,N_15471);
nor U15763 (N_15763,N_15599,N_15446);
nand U15764 (N_15764,N_15517,N_15417);
nand U15765 (N_15765,N_15541,N_15466);
or U15766 (N_15766,N_15427,N_15567);
xnor U15767 (N_15767,N_15460,N_15453);
or U15768 (N_15768,N_15482,N_15500);
and U15769 (N_15769,N_15537,N_15447);
nor U15770 (N_15770,N_15413,N_15439);
or U15771 (N_15771,N_15424,N_15597);
nor U15772 (N_15772,N_15521,N_15579);
xor U15773 (N_15773,N_15564,N_15424);
nor U15774 (N_15774,N_15597,N_15432);
nor U15775 (N_15775,N_15568,N_15419);
or U15776 (N_15776,N_15425,N_15418);
xor U15777 (N_15777,N_15445,N_15545);
nand U15778 (N_15778,N_15522,N_15404);
and U15779 (N_15779,N_15409,N_15416);
nor U15780 (N_15780,N_15525,N_15470);
or U15781 (N_15781,N_15505,N_15416);
xor U15782 (N_15782,N_15589,N_15480);
and U15783 (N_15783,N_15437,N_15476);
or U15784 (N_15784,N_15491,N_15472);
nor U15785 (N_15785,N_15578,N_15524);
or U15786 (N_15786,N_15433,N_15423);
or U15787 (N_15787,N_15488,N_15527);
nand U15788 (N_15788,N_15412,N_15483);
nor U15789 (N_15789,N_15405,N_15594);
xor U15790 (N_15790,N_15448,N_15504);
xnor U15791 (N_15791,N_15552,N_15567);
xor U15792 (N_15792,N_15447,N_15408);
xor U15793 (N_15793,N_15410,N_15405);
nor U15794 (N_15794,N_15513,N_15553);
nand U15795 (N_15795,N_15441,N_15489);
nand U15796 (N_15796,N_15450,N_15548);
and U15797 (N_15797,N_15576,N_15596);
nor U15798 (N_15798,N_15462,N_15559);
xnor U15799 (N_15799,N_15497,N_15476);
and U15800 (N_15800,N_15739,N_15650);
nor U15801 (N_15801,N_15679,N_15705);
and U15802 (N_15802,N_15724,N_15667);
nand U15803 (N_15803,N_15777,N_15764);
and U15804 (N_15804,N_15653,N_15771);
and U15805 (N_15805,N_15775,N_15701);
or U15806 (N_15806,N_15695,N_15628);
nor U15807 (N_15807,N_15692,N_15772);
xnor U15808 (N_15808,N_15728,N_15799);
nor U15809 (N_15809,N_15652,N_15608);
nor U15810 (N_15810,N_15688,N_15614);
nor U15811 (N_15811,N_15713,N_15673);
and U15812 (N_15812,N_15716,N_15649);
nand U15813 (N_15813,N_15745,N_15657);
nor U15814 (N_15814,N_15788,N_15662);
and U15815 (N_15815,N_15618,N_15605);
xnor U15816 (N_15816,N_15754,N_15674);
and U15817 (N_15817,N_15795,N_15699);
nor U15818 (N_15818,N_15635,N_15714);
or U15819 (N_15819,N_15619,N_15759);
nor U15820 (N_15820,N_15742,N_15791);
xor U15821 (N_15821,N_15607,N_15768);
xnor U15822 (N_15822,N_15735,N_15664);
nand U15823 (N_15823,N_15779,N_15686);
nor U15824 (N_15824,N_15661,N_15634);
nor U15825 (N_15825,N_15610,N_15697);
nor U15826 (N_15826,N_15659,N_15606);
and U15827 (N_15827,N_15602,N_15633);
nor U15828 (N_15828,N_15785,N_15647);
nor U15829 (N_15829,N_15601,N_15797);
nor U15830 (N_15830,N_15763,N_15696);
and U15831 (N_15831,N_15672,N_15694);
xnor U15832 (N_15832,N_15636,N_15725);
and U15833 (N_15833,N_15668,N_15729);
nor U15834 (N_15834,N_15769,N_15639);
nor U15835 (N_15835,N_15641,N_15637);
or U15836 (N_15836,N_15625,N_15762);
nand U15837 (N_15837,N_15717,N_15616);
and U15838 (N_15838,N_15770,N_15669);
and U15839 (N_15839,N_15689,N_15784);
and U15840 (N_15840,N_15645,N_15684);
nor U15841 (N_15841,N_15741,N_15747);
or U15842 (N_15842,N_15629,N_15700);
or U15843 (N_15843,N_15773,N_15737);
and U15844 (N_15844,N_15767,N_15613);
nand U15845 (N_15845,N_15743,N_15726);
xnor U15846 (N_15846,N_15603,N_15627);
xnor U15847 (N_15847,N_15656,N_15703);
nor U15848 (N_15848,N_15660,N_15732);
nor U15849 (N_15849,N_15707,N_15709);
or U15850 (N_15850,N_15632,N_15758);
and U15851 (N_15851,N_15630,N_15793);
nor U15852 (N_15852,N_15794,N_15731);
or U15853 (N_15853,N_15727,N_15680);
or U15854 (N_15854,N_15796,N_15658);
or U15855 (N_15855,N_15644,N_15786);
nor U15856 (N_15856,N_15774,N_15761);
nand U15857 (N_15857,N_15612,N_15609);
nor U15858 (N_15858,N_15787,N_15704);
nor U15859 (N_15859,N_15710,N_15666);
or U15860 (N_15860,N_15783,N_15623);
nand U15861 (N_15861,N_15631,N_15626);
or U15862 (N_15862,N_15755,N_15746);
and U15863 (N_15863,N_15722,N_15624);
nor U15864 (N_15864,N_15654,N_15676);
and U15865 (N_15865,N_15675,N_15789);
nor U15866 (N_15866,N_15778,N_15611);
and U15867 (N_15867,N_15749,N_15685);
nor U15868 (N_15868,N_15604,N_15643);
or U15869 (N_15869,N_15708,N_15723);
nand U15870 (N_15870,N_15691,N_15780);
and U15871 (N_15871,N_15646,N_15698);
nor U15872 (N_15872,N_15766,N_15663);
nand U15873 (N_15873,N_15782,N_15690);
xor U15874 (N_15874,N_15733,N_15744);
nor U15875 (N_15875,N_15621,N_15740);
xnor U15876 (N_15876,N_15715,N_15752);
nor U15877 (N_15877,N_15702,N_15677);
nand U15878 (N_15878,N_15681,N_15756);
or U15879 (N_15879,N_15718,N_15781);
xor U15880 (N_15880,N_15670,N_15753);
or U15881 (N_15881,N_15719,N_15665);
nand U15882 (N_15882,N_15671,N_15687);
xnor U15883 (N_15883,N_15738,N_15734);
or U15884 (N_15884,N_15757,N_15638);
or U15885 (N_15885,N_15678,N_15711);
or U15886 (N_15886,N_15760,N_15776);
xor U15887 (N_15887,N_15736,N_15790);
and U15888 (N_15888,N_15642,N_15620);
or U15889 (N_15889,N_15765,N_15683);
xnor U15890 (N_15890,N_15748,N_15648);
xor U15891 (N_15891,N_15798,N_15615);
nor U15892 (N_15892,N_15750,N_15721);
and U15893 (N_15893,N_15693,N_15720);
or U15894 (N_15894,N_15617,N_15730);
or U15895 (N_15895,N_15622,N_15751);
nor U15896 (N_15896,N_15712,N_15655);
or U15897 (N_15897,N_15600,N_15792);
nor U15898 (N_15898,N_15640,N_15706);
xor U15899 (N_15899,N_15682,N_15651);
and U15900 (N_15900,N_15731,N_15688);
nand U15901 (N_15901,N_15712,N_15747);
or U15902 (N_15902,N_15764,N_15687);
and U15903 (N_15903,N_15644,N_15642);
or U15904 (N_15904,N_15732,N_15688);
and U15905 (N_15905,N_15714,N_15621);
nor U15906 (N_15906,N_15634,N_15737);
or U15907 (N_15907,N_15729,N_15771);
or U15908 (N_15908,N_15699,N_15752);
and U15909 (N_15909,N_15761,N_15637);
nor U15910 (N_15910,N_15766,N_15755);
xor U15911 (N_15911,N_15605,N_15704);
and U15912 (N_15912,N_15742,N_15697);
nand U15913 (N_15913,N_15653,N_15791);
or U15914 (N_15914,N_15795,N_15709);
or U15915 (N_15915,N_15689,N_15629);
and U15916 (N_15916,N_15697,N_15601);
and U15917 (N_15917,N_15738,N_15603);
and U15918 (N_15918,N_15721,N_15684);
nand U15919 (N_15919,N_15683,N_15727);
and U15920 (N_15920,N_15604,N_15639);
or U15921 (N_15921,N_15619,N_15651);
nor U15922 (N_15922,N_15686,N_15663);
and U15923 (N_15923,N_15799,N_15790);
xor U15924 (N_15924,N_15749,N_15766);
nand U15925 (N_15925,N_15672,N_15767);
xnor U15926 (N_15926,N_15695,N_15743);
nand U15927 (N_15927,N_15793,N_15774);
nand U15928 (N_15928,N_15642,N_15704);
and U15929 (N_15929,N_15605,N_15784);
and U15930 (N_15930,N_15607,N_15783);
nor U15931 (N_15931,N_15785,N_15652);
and U15932 (N_15932,N_15748,N_15610);
and U15933 (N_15933,N_15652,N_15791);
xor U15934 (N_15934,N_15709,N_15668);
nand U15935 (N_15935,N_15663,N_15649);
and U15936 (N_15936,N_15651,N_15686);
and U15937 (N_15937,N_15675,N_15776);
or U15938 (N_15938,N_15714,N_15651);
nor U15939 (N_15939,N_15734,N_15634);
xor U15940 (N_15940,N_15772,N_15781);
nand U15941 (N_15941,N_15708,N_15669);
nor U15942 (N_15942,N_15707,N_15633);
xor U15943 (N_15943,N_15737,N_15699);
xor U15944 (N_15944,N_15600,N_15666);
or U15945 (N_15945,N_15769,N_15730);
nand U15946 (N_15946,N_15648,N_15785);
or U15947 (N_15947,N_15671,N_15646);
nor U15948 (N_15948,N_15676,N_15666);
xnor U15949 (N_15949,N_15770,N_15753);
and U15950 (N_15950,N_15721,N_15797);
nand U15951 (N_15951,N_15685,N_15620);
nor U15952 (N_15952,N_15786,N_15791);
and U15953 (N_15953,N_15720,N_15788);
or U15954 (N_15954,N_15729,N_15791);
xnor U15955 (N_15955,N_15785,N_15672);
or U15956 (N_15956,N_15762,N_15685);
xnor U15957 (N_15957,N_15601,N_15791);
xor U15958 (N_15958,N_15742,N_15702);
nand U15959 (N_15959,N_15707,N_15720);
and U15960 (N_15960,N_15694,N_15750);
or U15961 (N_15961,N_15752,N_15799);
xor U15962 (N_15962,N_15646,N_15651);
or U15963 (N_15963,N_15664,N_15600);
xnor U15964 (N_15964,N_15694,N_15671);
or U15965 (N_15965,N_15653,N_15745);
or U15966 (N_15966,N_15743,N_15719);
and U15967 (N_15967,N_15658,N_15729);
nand U15968 (N_15968,N_15732,N_15731);
or U15969 (N_15969,N_15701,N_15629);
nor U15970 (N_15970,N_15738,N_15675);
nor U15971 (N_15971,N_15727,N_15761);
and U15972 (N_15972,N_15685,N_15768);
or U15973 (N_15973,N_15719,N_15684);
xnor U15974 (N_15974,N_15673,N_15676);
and U15975 (N_15975,N_15620,N_15737);
nor U15976 (N_15976,N_15661,N_15751);
nand U15977 (N_15977,N_15624,N_15726);
and U15978 (N_15978,N_15690,N_15700);
or U15979 (N_15979,N_15787,N_15707);
xor U15980 (N_15980,N_15622,N_15678);
nand U15981 (N_15981,N_15614,N_15713);
nand U15982 (N_15982,N_15751,N_15746);
nand U15983 (N_15983,N_15746,N_15662);
nor U15984 (N_15984,N_15696,N_15675);
nor U15985 (N_15985,N_15691,N_15718);
nor U15986 (N_15986,N_15730,N_15778);
nand U15987 (N_15987,N_15652,N_15766);
nor U15988 (N_15988,N_15642,N_15645);
nor U15989 (N_15989,N_15644,N_15799);
nor U15990 (N_15990,N_15609,N_15714);
xnor U15991 (N_15991,N_15744,N_15755);
nand U15992 (N_15992,N_15750,N_15744);
and U15993 (N_15993,N_15615,N_15767);
nand U15994 (N_15994,N_15605,N_15703);
or U15995 (N_15995,N_15766,N_15678);
nand U15996 (N_15996,N_15648,N_15640);
and U15997 (N_15997,N_15603,N_15776);
and U15998 (N_15998,N_15619,N_15673);
and U15999 (N_15999,N_15655,N_15799);
nor U16000 (N_16000,N_15840,N_15911);
xor U16001 (N_16001,N_15916,N_15877);
and U16002 (N_16002,N_15930,N_15892);
or U16003 (N_16003,N_15874,N_15879);
nor U16004 (N_16004,N_15897,N_15983);
nor U16005 (N_16005,N_15806,N_15862);
nor U16006 (N_16006,N_15981,N_15949);
or U16007 (N_16007,N_15999,N_15923);
nor U16008 (N_16008,N_15912,N_15827);
nor U16009 (N_16009,N_15984,N_15814);
and U16010 (N_16010,N_15952,N_15944);
or U16011 (N_16011,N_15993,N_15948);
nand U16012 (N_16012,N_15951,N_15808);
and U16013 (N_16013,N_15873,N_15919);
nor U16014 (N_16014,N_15924,N_15917);
and U16015 (N_16015,N_15933,N_15907);
and U16016 (N_16016,N_15964,N_15990);
and U16017 (N_16017,N_15885,N_15967);
and U16018 (N_16018,N_15958,N_15953);
or U16019 (N_16019,N_15970,N_15868);
xor U16020 (N_16020,N_15973,N_15909);
xnor U16021 (N_16021,N_15800,N_15826);
nand U16022 (N_16022,N_15894,N_15977);
nor U16023 (N_16023,N_15942,N_15856);
nand U16024 (N_16024,N_15957,N_15927);
nor U16025 (N_16025,N_15838,N_15902);
nor U16026 (N_16026,N_15881,N_15857);
xor U16027 (N_16027,N_15809,N_15830);
nor U16028 (N_16028,N_15979,N_15985);
nor U16029 (N_16029,N_15893,N_15899);
xnor U16030 (N_16030,N_15928,N_15929);
nor U16031 (N_16031,N_15986,N_15849);
and U16032 (N_16032,N_15935,N_15974);
or U16033 (N_16033,N_15834,N_15965);
or U16034 (N_16034,N_15988,N_15898);
and U16035 (N_16035,N_15835,N_15864);
nor U16036 (N_16036,N_15804,N_15900);
nand U16037 (N_16037,N_15847,N_15869);
nor U16038 (N_16038,N_15908,N_15971);
xnor U16039 (N_16039,N_15829,N_15836);
and U16040 (N_16040,N_15817,N_15956);
nor U16041 (N_16041,N_15853,N_15807);
nor U16042 (N_16042,N_15878,N_15882);
and U16043 (N_16043,N_15833,N_15914);
xor U16044 (N_16044,N_15889,N_15926);
nand U16045 (N_16045,N_15931,N_15921);
nand U16046 (N_16046,N_15896,N_15866);
xor U16047 (N_16047,N_15996,N_15821);
nor U16048 (N_16048,N_15904,N_15987);
nor U16049 (N_16049,N_15858,N_15962);
nor U16050 (N_16050,N_15811,N_15850);
and U16051 (N_16051,N_15888,N_15870);
nor U16052 (N_16052,N_15844,N_15815);
or U16053 (N_16053,N_15876,N_15887);
and U16054 (N_16054,N_15854,N_15901);
nor U16055 (N_16055,N_15867,N_15803);
nor U16056 (N_16056,N_15960,N_15820);
nor U16057 (N_16057,N_15913,N_15954);
nand U16058 (N_16058,N_15805,N_15972);
and U16059 (N_16059,N_15824,N_15802);
and U16060 (N_16060,N_15975,N_15968);
or U16061 (N_16061,N_15890,N_15946);
xor U16062 (N_16062,N_15825,N_15910);
nand U16063 (N_16063,N_15991,N_15891);
nand U16064 (N_16064,N_15925,N_15855);
and U16065 (N_16065,N_15920,N_15872);
xor U16066 (N_16066,N_15841,N_15831);
nor U16067 (N_16067,N_15819,N_15934);
nor U16068 (N_16068,N_15932,N_15915);
nand U16069 (N_16069,N_15801,N_15851);
xor U16070 (N_16070,N_15846,N_15976);
nand U16071 (N_16071,N_15837,N_15884);
xnor U16072 (N_16072,N_15939,N_15950);
or U16073 (N_16073,N_15816,N_15980);
nor U16074 (N_16074,N_15848,N_15998);
xnor U16075 (N_16075,N_15959,N_15832);
nor U16076 (N_16076,N_15865,N_15883);
nor U16077 (N_16077,N_15886,N_15940);
nand U16078 (N_16078,N_15843,N_15969);
and U16079 (N_16079,N_15812,N_15992);
and U16080 (N_16080,N_15905,N_15938);
nand U16081 (N_16081,N_15828,N_15936);
nor U16082 (N_16082,N_15839,N_15852);
nor U16083 (N_16083,N_15861,N_15966);
xor U16084 (N_16084,N_15994,N_15810);
and U16085 (N_16085,N_15863,N_15842);
and U16086 (N_16086,N_15859,N_15903);
xor U16087 (N_16087,N_15982,N_15823);
xnor U16088 (N_16088,N_15922,N_15963);
nand U16089 (N_16089,N_15906,N_15871);
and U16090 (N_16090,N_15978,N_15989);
nand U16091 (N_16091,N_15845,N_15955);
nor U16092 (N_16092,N_15813,N_15947);
and U16093 (N_16093,N_15818,N_15918);
xor U16094 (N_16094,N_15822,N_15875);
xor U16095 (N_16095,N_15945,N_15860);
or U16096 (N_16096,N_15937,N_15895);
or U16097 (N_16097,N_15880,N_15997);
nor U16098 (N_16098,N_15943,N_15995);
xor U16099 (N_16099,N_15941,N_15961);
nor U16100 (N_16100,N_15970,N_15922);
nand U16101 (N_16101,N_15991,N_15867);
or U16102 (N_16102,N_15867,N_15895);
xor U16103 (N_16103,N_15810,N_15843);
or U16104 (N_16104,N_15836,N_15906);
nand U16105 (N_16105,N_15960,N_15991);
or U16106 (N_16106,N_15859,N_15863);
or U16107 (N_16107,N_15906,N_15843);
nor U16108 (N_16108,N_15951,N_15836);
xor U16109 (N_16109,N_15950,N_15858);
and U16110 (N_16110,N_15883,N_15964);
nor U16111 (N_16111,N_15802,N_15998);
or U16112 (N_16112,N_15802,N_15873);
and U16113 (N_16113,N_15882,N_15872);
nand U16114 (N_16114,N_15821,N_15964);
and U16115 (N_16115,N_15837,N_15811);
nand U16116 (N_16116,N_15860,N_15953);
nor U16117 (N_16117,N_15879,N_15860);
nand U16118 (N_16118,N_15925,N_15919);
xor U16119 (N_16119,N_15979,N_15870);
nand U16120 (N_16120,N_15827,N_15900);
nand U16121 (N_16121,N_15826,N_15854);
xor U16122 (N_16122,N_15854,N_15913);
xnor U16123 (N_16123,N_15902,N_15904);
xnor U16124 (N_16124,N_15874,N_15872);
and U16125 (N_16125,N_15963,N_15917);
or U16126 (N_16126,N_15991,N_15842);
xor U16127 (N_16127,N_15977,N_15989);
nand U16128 (N_16128,N_15935,N_15905);
nand U16129 (N_16129,N_15933,N_15978);
or U16130 (N_16130,N_15880,N_15961);
nor U16131 (N_16131,N_15977,N_15952);
or U16132 (N_16132,N_15844,N_15956);
nor U16133 (N_16133,N_15998,N_15912);
or U16134 (N_16134,N_15899,N_15909);
or U16135 (N_16135,N_15897,N_15846);
or U16136 (N_16136,N_15881,N_15844);
nand U16137 (N_16137,N_15962,N_15888);
xnor U16138 (N_16138,N_15996,N_15867);
nor U16139 (N_16139,N_15821,N_15907);
nand U16140 (N_16140,N_15928,N_15967);
and U16141 (N_16141,N_15865,N_15994);
xnor U16142 (N_16142,N_15891,N_15987);
nor U16143 (N_16143,N_15837,N_15916);
and U16144 (N_16144,N_15916,N_15909);
xor U16145 (N_16145,N_15867,N_15995);
and U16146 (N_16146,N_15888,N_15839);
and U16147 (N_16147,N_15896,N_15945);
and U16148 (N_16148,N_15840,N_15993);
nor U16149 (N_16149,N_15946,N_15863);
or U16150 (N_16150,N_15855,N_15928);
nand U16151 (N_16151,N_15823,N_15886);
nor U16152 (N_16152,N_15803,N_15802);
nor U16153 (N_16153,N_15837,N_15865);
and U16154 (N_16154,N_15934,N_15942);
or U16155 (N_16155,N_15951,N_15974);
nand U16156 (N_16156,N_15934,N_15923);
xnor U16157 (N_16157,N_15866,N_15874);
or U16158 (N_16158,N_15979,N_15824);
xnor U16159 (N_16159,N_15902,N_15944);
and U16160 (N_16160,N_15829,N_15889);
or U16161 (N_16161,N_15848,N_15821);
xor U16162 (N_16162,N_15929,N_15879);
and U16163 (N_16163,N_15836,N_15884);
nand U16164 (N_16164,N_15926,N_15947);
or U16165 (N_16165,N_15932,N_15978);
and U16166 (N_16166,N_15943,N_15841);
xnor U16167 (N_16167,N_15820,N_15806);
nor U16168 (N_16168,N_15897,N_15962);
and U16169 (N_16169,N_15812,N_15841);
or U16170 (N_16170,N_15868,N_15958);
or U16171 (N_16171,N_15953,N_15934);
or U16172 (N_16172,N_15949,N_15852);
nand U16173 (N_16173,N_15918,N_15967);
xor U16174 (N_16174,N_15819,N_15904);
nor U16175 (N_16175,N_15838,N_15990);
or U16176 (N_16176,N_15966,N_15997);
nor U16177 (N_16177,N_15876,N_15824);
nor U16178 (N_16178,N_15923,N_15930);
and U16179 (N_16179,N_15811,N_15869);
xor U16180 (N_16180,N_15961,N_15848);
xor U16181 (N_16181,N_15994,N_15878);
nand U16182 (N_16182,N_15896,N_15893);
or U16183 (N_16183,N_15871,N_15900);
nand U16184 (N_16184,N_15839,N_15939);
nand U16185 (N_16185,N_15859,N_15933);
xnor U16186 (N_16186,N_15847,N_15857);
or U16187 (N_16187,N_15870,N_15952);
and U16188 (N_16188,N_15918,N_15844);
nand U16189 (N_16189,N_15947,N_15830);
nor U16190 (N_16190,N_15945,N_15913);
xor U16191 (N_16191,N_15827,N_15956);
nand U16192 (N_16192,N_15986,N_15829);
nand U16193 (N_16193,N_15891,N_15813);
and U16194 (N_16194,N_15906,N_15911);
nand U16195 (N_16195,N_15822,N_15829);
or U16196 (N_16196,N_15860,N_15920);
and U16197 (N_16197,N_15948,N_15842);
nor U16198 (N_16198,N_15997,N_15976);
nor U16199 (N_16199,N_15846,N_15923);
nand U16200 (N_16200,N_16183,N_16148);
nand U16201 (N_16201,N_16061,N_16080);
nor U16202 (N_16202,N_16024,N_16012);
nand U16203 (N_16203,N_16090,N_16190);
nor U16204 (N_16204,N_16164,N_16182);
nand U16205 (N_16205,N_16097,N_16195);
xnor U16206 (N_16206,N_16197,N_16055);
or U16207 (N_16207,N_16101,N_16115);
xnor U16208 (N_16208,N_16196,N_16033);
nor U16209 (N_16209,N_16153,N_16152);
or U16210 (N_16210,N_16037,N_16116);
nor U16211 (N_16211,N_16056,N_16089);
xnor U16212 (N_16212,N_16135,N_16021);
and U16213 (N_16213,N_16181,N_16006);
nand U16214 (N_16214,N_16188,N_16150);
or U16215 (N_16215,N_16078,N_16099);
or U16216 (N_16216,N_16005,N_16067);
and U16217 (N_16217,N_16002,N_16134);
xnor U16218 (N_16218,N_16034,N_16088);
nor U16219 (N_16219,N_16167,N_16041);
xor U16220 (N_16220,N_16048,N_16103);
or U16221 (N_16221,N_16118,N_16193);
and U16222 (N_16222,N_16136,N_16100);
and U16223 (N_16223,N_16051,N_16120);
nor U16224 (N_16224,N_16156,N_16066);
nand U16225 (N_16225,N_16072,N_16062);
nand U16226 (N_16226,N_16003,N_16171);
nor U16227 (N_16227,N_16032,N_16146);
nand U16228 (N_16228,N_16054,N_16151);
and U16229 (N_16229,N_16198,N_16069);
nor U16230 (N_16230,N_16023,N_16045);
or U16231 (N_16231,N_16036,N_16165);
or U16232 (N_16232,N_16064,N_16191);
or U16233 (N_16233,N_16141,N_16137);
nand U16234 (N_16234,N_16176,N_16119);
nand U16235 (N_16235,N_16076,N_16029);
or U16236 (N_16236,N_16145,N_16144);
and U16237 (N_16237,N_16170,N_16113);
or U16238 (N_16238,N_16149,N_16169);
xnor U16239 (N_16239,N_16194,N_16060);
or U16240 (N_16240,N_16059,N_16063);
nor U16241 (N_16241,N_16026,N_16044);
nor U16242 (N_16242,N_16070,N_16157);
and U16243 (N_16243,N_16073,N_16123);
nand U16244 (N_16244,N_16093,N_16128);
and U16245 (N_16245,N_16187,N_16178);
nand U16246 (N_16246,N_16175,N_16142);
and U16247 (N_16247,N_16022,N_16143);
or U16248 (N_16248,N_16081,N_16160);
or U16249 (N_16249,N_16018,N_16052);
xor U16250 (N_16250,N_16130,N_16140);
nor U16251 (N_16251,N_16106,N_16016);
and U16252 (N_16252,N_16091,N_16105);
xor U16253 (N_16253,N_16071,N_16192);
or U16254 (N_16254,N_16065,N_16031);
or U16255 (N_16255,N_16108,N_16043);
nor U16256 (N_16256,N_16083,N_16138);
nor U16257 (N_16257,N_16008,N_16098);
nand U16258 (N_16258,N_16102,N_16132);
or U16259 (N_16259,N_16011,N_16030);
nor U16260 (N_16260,N_16049,N_16110);
nand U16261 (N_16261,N_16094,N_16161);
and U16262 (N_16262,N_16035,N_16058);
and U16263 (N_16263,N_16082,N_16040);
and U16264 (N_16264,N_16117,N_16177);
nand U16265 (N_16265,N_16075,N_16010);
nand U16266 (N_16266,N_16154,N_16086);
and U16267 (N_16267,N_16028,N_16050);
nor U16268 (N_16268,N_16185,N_16020);
nor U16269 (N_16269,N_16009,N_16111);
or U16270 (N_16270,N_16074,N_16166);
or U16271 (N_16271,N_16159,N_16168);
nand U16272 (N_16272,N_16077,N_16184);
and U16273 (N_16273,N_16158,N_16155);
and U16274 (N_16274,N_16122,N_16085);
xor U16275 (N_16275,N_16133,N_16096);
nand U16276 (N_16276,N_16027,N_16124);
and U16277 (N_16277,N_16047,N_16025);
nor U16278 (N_16278,N_16104,N_16125);
or U16279 (N_16279,N_16019,N_16095);
nand U16280 (N_16280,N_16147,N_16053);
xor U16281 (N_16281,N_16180,N_16189);
and U16282 (N_16282,N_16179,N_16084);
or U16283 (N_16283,N_16042,N_16107);
nand U16284 (N_16284,N_16017,N_16014);
or U16285 (N_16285,N_16127,N_16109);
nand U16286 (N_16286,N_16092,N_16199);
or U16287 (N_16287,N_16163,N_16173);
nor U16288 (N_16288,N_16007,N_16114);
nor U16289 (N_16289,N_16057,N_16013);
nand U16290 (N_16290,N_16129,N_16015);
nor U16291 (N_16291,N_16039,N_16038);
and U16292 (N_16292,N_16004,N_16131);
nand U16293 (N_16293,N_16139,N_16046);
nor U16294 (N_16294,N_16162,N_16186);
nor U16295 (N_16295,N_16001,N_16079);
nand U16296 (N_16296,N_16174,N_16000);
and U16297 (N_16297,N_16121,N_16172);
and U16298 (N_16298,N_16087,N_16068);
or U16299 (N_16299,N_16126,N_16112);
nand U16300 (N_16300,N_16047,N_16137);
and U16301 (N_16301,N_16021,N_16083);
or U16302 (N_16302,N_16060,N_16155);
nor U16303 (N_16303,N_16066,N_16003);
nand U16304 (N_16304,N_16037,N_16199);
and U16305 (N_16305,N_16076,N_16032);
and U16306 (N_16306,N_16087,N_16031);
nand U16307 (N_16307,N_16092,N_16033);
or U16308 (N_16308,N_16196,N_16104);
nand U16309 (N_16309,N_16176,N_16017);
or U16310 (N_16310,N_16005,N_16053);
or U16311 (N_16311,N_16156,N_16024);
xnor U16312 (N_16312,N_16028,N_16199);
or U16313 (N_16313,N_16178,N_16163);
or U16314 (N_16314,N_16116,N_16010);
and U16315 (N_16315,N_16059,N_16078);
nor U16316 (N_16316,N_16045,N_16153);
nor U16317 (N_16317,N_16134,N_16032);
or U16318 (N_16318,N_16190,N_16170);
xnor U16319 (N_16319,N_16061,N_16144);
nor U16320 (N_16320,N_16116,N_16036);
nor U16321 (N_16321,N_16046,N_16189);
nand U16322 (N_16322,N_16052,N_16186);
nand U16323 (N_16323,N_16005,N_16190);
xnor U16324 (N_16324,N_16044,N_16076);
nor U16325 (N_16325,N_16124,N_16160);
xnor U16326 (N_16326,N_16056,N_16145);
or U16327 (N_16327,N_16020,N_16036);
or U16328 (N_16328,N_16128,N_16163);
nand U16329 (N_16329,N_16185,N_16129);
or U16330 (N_16330,N_16149,N_16054);
and U16331 (N_16331,N_16097,N_16096);
nand U16332 (N_16332,N_16031,N_16111);
or U16333 (N_16333,N_16008,N_16129);
xor U16334 (N_16334,N_16037,N_16048);
or U16335 (N_16335,N_16098,N_16068);
xor U16336 (N_16336,N_16017,N_16152);
nand U16337 (N_16337,N_16111,N_16059);
or U16338 (N_16338,N_16124,N_16146);
xor U16339 (N_16339,N_16097,N_16141);
nor U16340 (N_16340,N_16081,N_16151);
xor U16341 (N_16341,N_16024,N_16120);
and U16342 (N_16342,N_16082,N_16049);
nand U16343 (N_16343,N_16048,N_16124);
nor U16344 (N_16344,N_16134,N_16067);
nor U16345 (N_16345,N_16025,N_16064);
xnor U16346 (N_16346,N_16069,N_16066);
or U16347 (N_16347,N_16024,N_16197);
and U16348 (N_16348,N_16139,N_16012);
nor U16349 (N_16349,N_16085,N_16017);
nor U16350 (N_16350,N_16110,N_16029);
nor U16351 (N_16351,N_16104,N_16053);
nor U16352 (N_16352,N_16110,N_16131);
nor U16353 (N_16353,N_16091,N_16006);
nand U16354 (N_16354,N_16060,N_16189);
nand U16355 (N_16355,N_16196,N_16101);
and U16356 (N_16356,N_16129,N_16186);
nand U16357 (N_16357,N_16015,N_16111);
or U16358 (N_16358,N_16109,N_16090);
and U16359 (N_16359,N_16008,N_16156);
or U16360 (N_16360,N_16139,N_16075);
xor U16361 (N_16361,N_16135,N_16170);
and U16362 (N_16362,N_16123,N_16085);
nand U16363 (N_16363,N_16159,N_16020);
and U16364 (N_16364,N_16169,N_16112);
xor U16365 (N_16365,N_16119,N_16180);
xor U16366 (N_16366,N_16019,N_16168);
and U16367 (N_16367,N_16155,N_16030);
and U16368 (N_16368,N_16176,N_16171);
nor U16369 (N_16369,N_16106,N_16028);
or U16370 (N_16370,N_16041,N_16115);
and U16371 (N_16371,N_16045,N_16046);
nand U16372 (N_16372,N_16066,N_16036);
and U16373 (N_16373,N_16112,N_16003);
or U16374 (N_16374,N_16072,N_16043);
nand U16375 (N_16375,N_16173,N_16175);
nand U16376 (N_16376,N_16080,N_16069);
nand U16377 (N_16377,N_16072,N_16138);
xor U16378 (N_16378,N_16093,N_16118);
nand U16379 (N_16379,N_16030,N_16109);
nand U16380 (N_16380,N_16113,N_16097);
nand U16381 (N_16381,N_16023,N_16168);
nand U16382 (N_16382,N_16062,N_16156);
or U16383 (N_16383,N_16112,N_16120);
or U16384 (N_16384,N_16115,N_16177);
xor U16385 (N_16385,N_16019,N_16050);
nor U16386 (N_16386,N_16163,N_16157);
xnor U16387 (N_16387,N_16049,N_16140);
or U16388 (N_16388,N_16193,N_16161);
or U16389 (N_16389,N_16015,N_16090);
nand U16390 (N_16390,N_16153,N_16007);
and U16391 (N_16391,N_16186,N_16016);
nand U16392 (N_16392,N_16100,N_16101);
xnor U16393 (N_16393,N_16015,N_16087);
and U16394 (N_16394,N_16199,N_16023);
or U16395 (N_16395,N_16152,N_16180);
nor U16396 (N_16396,N_16082,N_16015);
nand U16397 (N_16397,N_16063,N_16069);
and U16398 (N_16398,N_16165,N_16133);
xnor U16399 (N_16399,N_16077,N_16005);
xor U16400 (N_16400,N_16310,N_16250);
nor U16401 (N_16401,N_16242,N_16215);
xnor U16402 (N_16402,N_16344,N_16369);
or U16403 (N_16403,N_16354,N_16239);
or U16404 (N_16404,N_16333,N_16346);
xnor U16405 (N_16405,N_16229,N_16325);
or U16406 (N_16406,N_16359,N_16349);
xor U16407 (N_16407,N_16307,N_16218);
nor U16408 (N_16408,N_16247,N_16353);
nand U16409 (N_16409,N_16249,N_16201);
nand U16410 (N_16410,N_16306,N_16213);
nand U16411 (N_16411,N_16328,N_16235);
or U16412 (N_16412,N_16308,N_16278);
xor U16413 (N_16413,N_16205,N_16206);
nand U16414 (N_16414,N_16331,N_16287);
nor U16415 (N_16415,N_16329,N_16236);
nand U16416 (N_16416,N_16208,N_16350);
nand U16417 (N_16417,N_16383,N_16355);
and U16418 (N_16418,N_16232,N_16364);
nand U16419 (N_16419,N_16298,N_16253);
or U16420 (N_16420,N_16280,N_16202);
and U16421 (N_16421,N_16334,N_16291);
or U16422 (N_16422,N_16382,N_16342);
nor U16423 (N_16423,N_16246,N_16300);
or U16424 (N_16424,N_16252,N_16376);
xor U16425 (N_16425,N_16389,N_16332);
and U16426 (N_16426,N_16375,N_16319);
or U16427 (N_16427,N_16204,N_16343);
and U16428 (N_16428,N_16267,N_16245);
and U16429 (N_16429,N_16323,N_16279);
and U16430 (N_16430,N_16394,N_16297);
or U16431 (N_16431,N_16301,N_16288);
xor U16432 (N_16432,N_16220,N_16203);
nand U16433 (N_16433,N_16295,N_16385);
xor U16434 (N_16434,N_16263,N_16387);
nand U16435 (N_16435,N_16289,N_16209);
xor U16436 (N_16436,N_16338,N_16207);
and U16437 (N_16437,N_16221,N_16374);
xnor U16438 (N_16438,N_16224,N_16282);
and U16439 (N_16439,N_16260,N_16339);
nor U16440 (N_16440,N_16284,N_16251);
xor U16441 (N_16441,N_16276,N_16372);
nor U16442 (N_16442,N_16360,N_16371);
nand U16443 (N_16443,N_16366,N_16399);
and U16444 (N_16444,N_16351,N_16368);
and U16445 (N_16445,N_16322,N_16258);
nor U16446 (N_16446,N_16214,N_16378);
nor U16447 (N_16447,N_16271,N_16233);
or U16448 (N_16448,N_16261,N_16290);
or U16449 (N_16449,N_16379,N_16316);
nor U16450 (N_16450,N_16226,N_16317);
nand U16451 (N_16451,N_16238,N_16315);
nand U16452 (N_16452,N_16200,N_16391);
and U16453 (N_16453,N_16286,N_16318);
xnor U16454 (N_16454,N_16259,N_16227);
and U16455 (N_16455,N_16277,N_16324);
or U16456 (N_16456,N_16393,N_16386);
or U16457 (N_16457,N_16269,N_16312);
or U16458 (N_16458,N_16381,N_16212);
and U16459 (N_16459,N_16268,N_16241);
xor U16460 (N_16460,N_16257,N_16348);
xnor U16461 (N_16461,N_16356,N_16330);
xnor U16462 (N_16462,N_16272,N_16255);
or U16463 (N_16463,N_16262,N_16222);
nand U16464 (N_16464,N_16390,N_16217);
xnor U16465 (N_16465,N_16345,N_16370);
nor U16466 (N_16466,N_16377,N_16304);
and U16467 (N_16467,N_16347,N_16311);
xnor U16468 (N_16468,N_16231,N_16243);
xnor U16469 (N_16469,N_16216,N_16327);
xnor U16470 (N_16470,N_16223,N_16293);
and U16471 (N_16471,N_16309,N_16321);
or U16472 (N_16472,N_16285,N_16367);
and U16473 (N_16473,N_16303,N_16361);
nor U16474 (N_16474,N_16275,N_16283);
or U16475 (N_16475,N_16294,N_16395);
xor U16476 (N_16476,N_16388,N_16398);
xor U16477 (N_16477,N_16392,N_16266);
xor U16478 (N_16478,N_16320,N_16337);
xnor U16479 (N_16479,N_16335,N_16274);
nand U16480 (N_16480,N_16256,N_16254);
and U16481 (N_16481,N_16365,N_16305);
nand U16482 (N_16482,N_16336,N_16230);
and U16483 (N_16483,N_16237,N_16373);
and U16484 (N_16484,N_16397,N_16219);
or U16485 (N_16485,N_16384,N_16281);
and U16486 (N_16486,N_16228,N_16362);
nand U16487 (N_16487,N_16244,N_16314);
xor U16488 (N_16488,N_16225,N_16248);
and U16489 (N_16489,N_16380,N_16299);
nand U16490 (N_16490,N_16313,N_16264);
nor U16491 (N_16491,N_16352,N_16326);
and U16492 (N_16492,N_16340,N_16357);
nor U16493 (N_16493,N_16296,N_16210);
nor U16494 (N_16494,N_16270,N_16273);
or U16495 (N_16495,N_16240,N_16211);
nor U16496 (N_16496,N_16234,N_16396);
nor U16497 (N_16497,N_16292,N_16363);
and U16498 (N_16498,N_16358,N_16265);
xnor U16499 (N_16499,N_16341,N_16302);
nand U16500 (N_16500,N_16291,N_16239);
nor U16501 (N_16501,N_16260,N_16396);
nand U16502 (N_16502,N_16371,N_16290);
xnor U16503 (N_16503,N_16387,N_16369);
or U16504 (N_16504,N_16268,N_16336);
nor U16505 (N_16505,N_16392,N_16347);
or U16506 (N_16506,N_16223,N_16326);
nor U16507 (N_16507,N_16331,N_16280);
xnor U16508 (N_16508,N_16275,N_16245);
nor U16509 (N_16509,N_16368,N_16203);
xor U16510 (N_16510,N_16221,N_16280);
and U16511 (N_16511,N_16320,N_16216);
xor U16512 (N_16512,N_16281,N_16301);
nand U16513 (N_16513,N_16268,N_16331);
or U16514 (N_16514,N_16315,N_16328);
nand U16515 (N_16515,N_16262,N_16322);
nor U16516 (N_16516,N_16388,N_16202);
xor U16517 (N_16517,N_16242,N_16254);
and U16518 (N_16518,N_16306,N_16347);
nor U16519 (N_16519,N_16360,N_16283);
and U16520 (N_16520,N_16382,N_16397);
and U16521 (N_16521,N_16299,N_16200);
nor U16522 (N_16522,N_16279,N_16251);
or U16523 (N_16523,N_16287,N_16321);
nor U16524 (N_16524,N_16377,N_16397);
nand U16525 (N_16525,N_16244,N_16379);
nand U16526 (N_16526,N_16303,N_16360);
nor U16527 (N_16527,N_16223,N_16242);
nand U16528 (N_16528,N_16232,N_16257);
xnor U16529 (N_16529,N_16206,N_16215);
xor U16530 (N_16530,N_16342,N_16388);
xor U16531 (N_16531,N_16294,N_16298);
or U16532 (N_16532,N_16229,N_16279);
nor U16533 (N_16533,N_16270,N_16242);
and U16534 (N_16534,N_16226,N_16249);
nor U16535 (N_16535,N_16322,N_16398);
xnor U16536 (N_16536,N_16308,N_16306);
or U16537 (N_16537,N_16396,N_16304);
or U16538 (N_16538,N_16285,N_16221);
and U16539 (N_16539,N_16292,N_16341);
nand U16540 (N_16540,N_16323,N_16321);
nand U16541 (N_16541,N_16220,N_16260);
or U16542 (N_16542,N_16285,N_16222);
nand U16543 (N_16543,N_16270,N_16393);
nor U16544 (N_16544,N_16217,N_16285);
nand U16545 (N_16545,N_16353,N_16275);
nor U16546 (N_16546,N_16294,N_16223);
and U16547 (N_16547,N_16242,N_16284);
and U16548 (N_16548,N_16253,N_16220);
nand U16549 (N_16549,N_16287,N_16300);
xor U16550 (N_16550,N_16245,N_16237);
xnor U16551 (N_16551,N_16346,N_16309);
nor U16552 (N_16552,N_16341,N_16254);
and U16553 (N_16553,N_16255,N_16329);
and U16554 (N_16554,N_16271,N_16343);
xnor U16555 (N_16555,N_16216,N_16386);
nand U16556 (N_16556,N_16232,N_16205);
xor U16557 (N_16557,N_16316,N_16210);
or U16558 (N_16558,N_16275,N_16205);
xnor U16559 (N_16559,N_16269,N_16342);
or U16560 (N_16560,N_16349,N_16371);
xnor U16561 (N_16561,N_16328,N_16301);
xnor U16562 (N_16562,N_16253,N_16254);
xor U16563 (N_16563,N_16331,N_16211);
or U16564 (N_16564,N_16336,N_16202);
xnor U16565 (N_16565,N_16305,N_16288);
or U16566 (N_16566,N_16325,N_16344);
nor U16567 (N_16567,N_16286,N_16320);
nor U16568 (N_16568,N_16215,N_16391);
or U16569 (N_16569,N_16397,N_16228);
nand U16570 (N_16570,N_16306,N_16357);
xor U16571 (N_16571,N_16330,N_16277);
and U16572 (N_16572,N_16324,N_16222);
and U16573 (N_16573,N_16365,N_16334);
xnor U16574 (N_16574,N_16225,N_16328);
nand U16575 (N_16575,N_16320,N_16393);
and U16576 (N_16576,N_16212,N_16343);
xor U16577 (N_16577,N_16292,N_16399);
nor U16578 (N_16578,N_16307,N_16260);
and U16579 (N_16579,N_16307,N_16257);
nand U16580 (N_16580,N_16218,N_16292);
nand U16581 (N_16581,N_16250,N_16387);
and U16582 (N_16582,N_16384,N_16250);
nand U16583 (N_16583,N_16392,N_16220);
and U16584 (N_16584,N_16325,N_16360);
xor U16585 (N_16585,N_16345,N_16331);
and U16586 (N_16586,N_16210,N_16294);
nand U16587 (N_16587,N_16296,N_16213);
and U16588 (N_16588,N_16274,N_16324);
and U16589 (N_16589,N_16204,N_16235);
and U16590 (N_16590,N_16250,N_16353);
nand U16591 (N_16591,N_16372,N_16290);
nor U16592 (N_16592,N_16237,N_16308);
nor U16593 (N_16593,N_16395,N_16397);
or U16594 (N_16594,N_16306,N_16364);
and U16595 (N_16595,N_16238,N_16379);
nor U16596 (N_16596,N_16282,N_16290);
nor U16597 (N_16597,N_16376,N_16286);
nand U16598 (N_16598,N_16204,N_16355);
or U16599 (N_16599,N_16250,N_16317);
nand U16600 (N_16600,N_16571,N_16511);
nand U16601 (N_16601,N_16443,N_16583);
nand U16602 (N_16602,N_16427,N_16457);
and U16603 (N_16603,N_16445,N_16595);
xnor U16604 (N_16604,N_16548,N_16472);
nand U16605 (N_16605,N_16426,N_16522);
xnor U16606 (N_16606,N_16565,N_16534);
and U16607 (N_16607,N_16581,N_16491);
nor U16608 (N_16608,N_16418,N_16417);
or U16609 (N_16609,N_16579,N_16588);
xnor U16610 (N_16610,N_16529,N_16598);
and U16611 (N_16611,N_16509,N_16596);
nand U16612 (N_16612,N_16449,N_16451);
nand U16613 (N_16613,N_16513,N_16495);
and U16614 (N_16614,N_16585,N_16433);
or U16615 (N_16615,N_16458,N_16554);
or U16616 (N_16616,N_16514,N_16436);
nand U16617 (N_16617,N_16525,N_16544);
xnor U16618 (N_16618,N_16424,N_16599);
nand U16619 (N_16619,N_16448,N_16488);
nand U16620 (N_16620,N_16504,N_16453);
or U16621 (N_16621,N_16532,N_16425);
and U16622 (N_16622,N_16429,N_16582);
or U16623 (N_16623,N_16414,N_16493);
and U16624 (N_16624,N_16465,N_16401);
or U16625 (N_16625,N_16528,N_16478);
or U16626 (N_16626,N_16573,N_16503);
or U16627 (N_16627,N_16570,N_16586);
nand U16628 (N_16628,N_16408,N_16479);
nor U16629 (N_16629,N_16428,N_16410);
and U16630 (N_16630,N_16496,N_16468);
nand U16631 (N_16631,N_16407,N_16560);
xor U16632 (N_16632,N_16537,N_16421);
xor U16633 (N_16633,N_16405,N_16473);
nor U16634 (N_16634,N_16489,N_16439);
xor U16635 (N_16635,N_16430,N_16461);
nor U16636 (N_16636,N_16557,N_16447);
nor U16637 (N_16637,N_16476,N_16477);
xor U16638 (N_16638,N_16467,N_16523);
or U16639 (N_16639,N_16597,N_16454);
and U16640 (N_16640,N_16535,N_16515);
nor U16641 (N_16641,N_16484,N_16575);
or U16642 (N_16642,N_16568,N_16475);
or U16643 (N_16643,N_16577,N_16552);
nand U16644 (N_16644,N_16482,N_16555);
and U16645 (N_16645,N_16463,N_16438);
or U16646 (N_16646,N_16563,N_16416);
nand U16647 (N_16647,N_16527,N_16497);
nand U16648 (N_16648,N_16512,N_16492);
or U16649 (N_16649,N_16580,N_16593);
nor U16650 (N_16650,N_16481,N_16494);
nor U16651 (N_16651,N_16508,N_16402);
and U16652 (N_16652,N_16499,N_16569);
xnor U16653 (N_16653,N_16466,N_16412);
or U16654 (N_16654,N_16591,N_16530);
nand U16655 (N_16655,N_16538,N_16558);
xnor U16656 (N_16656,N_16441,N_16413);
nor U16657 (N_16657,N_16450,N_16422);
nor U16658 (N_16658,N_16432,N_16498);
nand U16659 (N_16659,N_16406,N_16531);
nor U16660 (N_16660,N_16400,N_16455);
nand U16661 (N_16661,N_16415,N_16431);
xor U16662 (N_16662,N_16546,N_16584);
xor U16663 (N_16663,N_16470,N_16442);
nand U16664 (N_16664,N_16519,N_16517);
and U16665 (N_16665,N_16462,N_16556);
or U16666 (N_16666,N_16549,N_16423);
nor U16667 (N_16667,N_16490,N_16516);
nor U16668 (N_16668,N_16592,N_16404);
xor U16669 (N_16669,N_16435,N_16550);
xnor U16670 (N_16670,N_16566,N_16589);
nand U16671 (N_16671,N_16460,N_16561);
xnor U16672 (N_16672,N_16510,N_16419);
nand U16673 (N_16673,N_16437,N_16456);
or U16674 (N_16674,N_16409,N_16403);
or U16675 (N_16675,N_16553,N_16444);
or U16676 (N_16676,N_16551,N_16594);
nor U16677 (N_16677,N_16420,N_16480);
or U16678 (N_16678,N_16543,N_16520);
xnor U16679 (N_16679,N_16567,N_16471);
nand U16680 (N_16680,N_16464,N_16452);
or U16681 (N_16681,N_16590,N_16434);
xnor U16682 (N_16682,N_16486,N_16540);
and U16683 (N_16683,N_16483,N_16505);
xor U16684 (N_16684,N_16564,N_16501);
or U16685 (N_16685,N_16459,N_16578);
xnor U16686 (N_16686,N_16411,N_16545);
nor U16687 (N_16687,N_16507,N_16572);
nor U16688 (N_16688,N_16539,N_16542);
or U16689 (N_16689,N_16487,N_16521);
and U16690 (N_16690,N_16485,N_16562);
nor U16691 (N_16691,N_16559,N_16500);
or U16692 (N_16692,N_16518,N_16502);
nand U16693 (N_16693,N_16536,N_16533);
or U16694 (N_16694,N_16547,N_16526);
nor U16695 (N_16695,N_16474,N_16524);
nor U16696 (N_16696,N_16440,N_16587);
and U16697 (N_16697,N_16506,N_16576);
nand U16698 (N_16698,N_16446,N_16469);
xor U16699 (N_16699,N_16541,N_16574);
or U16700 (N_16700,N_16422,N_16491);
nor U16701 (N_16701,N_16561,N_16463);
and U16702 (N_16702,N_16470,N_16559);
nor U16703 (N_16703,N_16412,N_16459);
nor U16704 (N_16704,N_16570,N_16493);
nand U16705 (N_16705,N_16569,N_16547);
nor U16706 (N_16706,N_16470,N_16505);
or U16707 (N_16707,N_16458,N_16576);
nand U16708 (N_16708,N_16564,N_16484);
xnor U16709 (N_16709,N_16525,N_16547);
and U16710 (N_16710,N_16426,N_16507);
xor U16711 (N_16711,N_16470,N_16463);
xnor U16712 (N_16712,N_16554,N_16478);
and U16713 (N_16713,N_16549,N_16517);
nor U16714 (N_16714,N_16429,N_16481);
xor U16715 (N_16715,N_16429,N_16439);
and U16716 (N_16716,N_16496,N_16545);
and U16717 (N_16717,N_16507,N_16493);
xor U16718 (N_16718,N_16490,N_16429);
nand U16719 (N_16719,N_16533,N_16553);
or U16720 (N_16720,N_16508,N_16501);
nand U16721 (N_16721,N_16543,N_16521);
nand U16722 (N_16722,N_16597,N_16508);
and U16723 (N_16723,N_16504,N_16497);
xnor U16724 (N_16724,N_16555,N_16551);
xor U16725 (N_16725,N_16516,N_16446);
or U16726 (N_16726,N_16532,N_16444);
and U16727 (N_16727,N_16533,N_16476);
or U16728 (N_16728,N_16578,N_16535);
xor U16729 (N_16729,N_16595,N_16524);
xnor U16730 (N_16730,N_16424,N_16519);
and U16731 (N_16731,N_16572,N_16503);
or U16732 (N_16732,N_16444,N_16410);
or U16733 (N_16733,N_16572,N_16430);
nor U16734 (N_16734,N_16587,N_16547);
or U16735 (N_16735,N_16400,N_16582);
nand U16736 (N_16736,N_16476,N_16548);
nor U16737 (N_16737,N_16544,N_16446);
or U16738 (N_16738,N_16421,N_16483);
nand U16739 (N_16739,N_16412,N_16469);
and U16740 (N_16740,N_16403,N_16502);
xor U16741 (N_16741,N_16541,N_16598);
nor U16742 (N_16742,N_16554,N_16519);
and U16743 (N_16743,N_16555,N_16576);
xnor U16744 (N_16744,N_16406,N_16465);
xnor U16745 (N_16745,N_16554,N_16491);
and U16746 (N_16746,N_16512,N_16534);
or U16747 (N_16747,N_16507,N_16527);
or U16748 (N_16748,N_16481,N_16495);
nor U16749 (N_16749,N_16524,N_16594);
nand U16750 (N_16750,N_16584,N_16586);
xnor U16751 (N_16751,N_16485,N_16470);
nor U16752 (N_16752,N_16466,N_16470);
or U16753 (N_16753,N_16412,N_16454);
and U16754 (N_16754,N_16503,N_16438);
or U16755 (N_16755,N_16412,N_16529);
and U16756 (N_16756,N_16405,N_16569);
and U16757 (N_16757,N_16556,N_16499);
xnor U16758 (N_16758,N_16428,N_16487);
and U16759 (N_16759,N_16461,N_16522);
or U16760 (N_16760,N_16567,N_16534);
xor U16761 (N_16761,N_16467,N_16404);
xor U16762 (N_16762,N_16515,N_16408);
xor U16763 (N_16763,N_16485,N_16456);
nor U16764 (N_16764,N_16496,N_16447);
nor U16765 (N_16765,N_16487,N_16583);
nand U16766 (N_16766,N_16422,N_16559);
nor U16767 (N_16767,N_16503,N_16486);
nor U16768 (N_16768,N_16535,N_16503);
or U16769 (N_16769,N_16537,N_16517);
xnor U16770 (N_16770,N_16493,N_16429);
xor U16771 (N_16771,N_16561,N_16407);
nand U16772 (N_16772,N_16450,N_16514);
nand U16773 (N_16773,N_16471,N_16444);
or U16774 (N_16774,N_16416,N_16570);
xor U16775 (N_16775,N_16583,N_16509);
and U16776 (N_16776,N_16582,N_16503);
xnor U16777 (N_16777,N_16429,N_16499);
xor U16778 (N_16778,N_16444,N_16454);
nand U16779 (N_16779,N_16554,N_16512);
nor U16780 (N_16780,N_16591,N_16595);
xor U16781 (N_16781,N_16539,N_16409);
or U16782 (N_16782,N_16430,N_16423);
xor U16783 (N_16783,N_16573,N_16570);
xor U16784 (N_16784,N_16565,N_16517);
xor U16785 (N_16785,N_16519,N_16500);
xor U16786 (N_16786,N_16427,N_16581);
and U16787 (N_16787,N_16507,N_16504);
nor U16788 (N_16788,N_16483,N_16564);
nand U16789 (N_16789,N_16546,N_16556);
xnor U16790 (N_16790,N_16402,N_16449);
xor U16791 (N_16791,N_16566,N_16590);
nand U16792 (N_16792,N_16528,N_16544);
or U16793 (N_16793,N_16487,N_16572);
nor U16794 (N_16794,N_16523,N_16556);
nand U16795 (N_16795,N_16504,N_16443);
nand U16796 (N_16796,N_16409,N_16447);
nand U16797 (N_16797,N_16411,N_16435);
and U16798 (N_16798,N_16572,N_16520);
and U16799 (N_16799,N_16454,N_16456);
nor U16800 (N_16800,N_16629,N_16678);
or U16801 (N_16801,N_16774,N_16752);
and U16802 (N_16802,N_16672,N_16631);
nand U16803 (N_16803,N_16753,N_16600);
xor U16804 (N_16804,N_16708,N_16755);
or U16805 (N_16805,N_16662,N_16691);
nor U16806 (N_16806,N_16716,N_16741);
or U16807 (N_16807,N_16659,N_16642);
nand U16808 (N_16808,N_16761,N_16685);
nand U16809 (N_16809,N_16735,N_16737);
or U16810 (N_16810,N_16732,N_16689);
nor U16811 (N_16811,N_16791,N_16698);
xnor U16812 (N_16812,N_16632,N_16617);
xor U16813 (N_16813,N_16707,N_16713);
xor U16814 (N_16814,N_16663,N_16609);
and U16815 (N_16815,N_16696,N_16683);
nor U16816 (N_16816,N_16602,N_16718);
or U16817 (N_16817,N_16789,N_16643);
and U16818 (N_16818,N_16766,N_16613);
nand U16819 (N_16819,N_16796,N_16606);
xor U16820 (N_16820,N_16799,N_16701);
or U16821 (N_16821,N_16675,N_16736);
and U16822 (N_16822,N_16773,N_16775);
and U16823 (N_16823,N_16769,N_16618);
nor U16824 (N_16824,N_16762,N_16624);
nor U16825 (N_16825,N_16634,N_16792);
xnor U16826 (N_16826,N_16740,N_16654);
and U16827 (N_16827,N_16640,N_16649);
nand U16828 (N_16828,N_16754,N_16627);
or U16829 (N_16829,N_16699,N_16616);
and U16830 (N_16830,N_16730,N_16610);
nor U16831 (N_16831,N_16676,N_16767);
or U16832 (N_16832,N_16619,N_16648);
or U16833 (N_16833,N_16666,N_16763);
or U16834 (N_16834,N_16725,N_16668);
xnor U16835 (N_16835,N_16615,N_16650);
or U16836 (N_16836,N_16694,N_16623);
nor U16837 (N_16837,N_16681,N_16744);
xnor U16838 (N_16838,N_16720,N_16651);
nor U16839 (N_16839,N_16787,N_16630);
nand U16840 (N_16840,N_16764,N_16690);
and U16841 (N_16841,N_16751,N_16715);
nor U16842 (N_16842,N_16680,N_16779);
xnor U16843 (N_16843,N_16729,N_16622);
nor U16844 (N_16844,N_16717,N_16728);
nor U16845 (N_16845,N_16709,N_16727);
nor U16846 (N_16846,N_16750,N_16652);
and U16847 (N_16847,N_16626,N_16684);
or U16848 (N_16848,N_16679,N_16778);
and U16849 (N_16849,N_16719,N_16757);
or U16850 (N_16850,N_16661,N_16781);
xor U16851 (N_16851,N_16790,N_16658);
nor U16852 (N_16852,N_16771,N_16747);
or U16853 (N_16853,N_16768,N_16703);
and U16854 (N_16854,N_16697,N_16759);
nand U16855 (N_16855,N_16743,N_16693);
nor U16856 (N_16856,N_16611,N_16797);
nand U16857 (N_16857,N_16625,N_16635);
or U16858 (N_16858,N_16667,N_16734);
or U16859 (N_16859,N_16655,N_16682);
nand U16860 (N_16860,N_16704,N_16620);
xnor U16861 (N_16861,N_16653,N_16772);
nor U16862 (N_16862,N_16669,N_16601);
nor U16863 (N_16863,N_16656,N_16665);
or U16864 (N_16864,N_16687,N_16639);
or U16865 (N_16865,N_16657,N_16636);
and U16866 (N_16866,N_16786,N_16795);
and U16867 (N_16867,N_16603,N_16738);
xnor U16868 (N_16868,N_16641,N_16758);
and U16869 (N_16869,N_16793,N_16628);
and U16870 (N_16870,N_16777,N_16645);
nor U16871 (N_16871,N_16695,N_16608);
and U16872 (N_16872,N_16660,N_16670);
nand U16873 (N_16873,N_16726,N_16712);
xnor U16874 (N_16874,N_16702,N_16794);
nor U16875 (N_16875,N_16692,N_16760);
xor U16876 (N_16876,N_16674,N_16722);
xnor U16877 (N_16877,N_16783,N_16788);
nand U16878 (N_16878,N_16677,N_16780);
nor U16879 (N_16879,N_16765,N_16646);
nand U16880 (N_16880,N_16721,N_16671);
and U16881 (N_16881,N_16798,N_16733);
or U16882 (N_16882,N_16664,N_16705);
nand U16883 (N_16883,N_16605,N_16724);
nor U16884 (N_16884,N_16700,N_16749);
nor U16885 (N_16885,N_16745,N_16607);
and U16886 (N_16886,N_16673,N_16644);
and U16887 (N_16887,N_16647,N_16637);
and U16888 (N_16888,N_16621,N_16710);
nand U16889 (N_16889,N_16784,N_16612);
or U16890 (N_16890,N_16688,N_16785);
or U16891 (N_16891,N_16686,N_16614);
nor U16892 (N_16892,N_16723,N_16748);
nand U16893 (N_16893,N_16782,N_16746);
nor U16894 (N_16894,N_16714,N_16633);
or U16895 (N_16895,N_16776,N_16638);
nand U16896 (N_16896,N_16756,N_16742);
or U16897 (N_16897,N_16711,N_16770);
nand U16898 (N_16898,N_16731,N_16739);
nand U16899 (N_16899,N_16604,N_16706);
xnor U16900 (N_16900,N_16755,N_16789);
and U16901 (N_16901,N_16631,N_16653);
or U16902 (N_16902,N_16779,N_16750);
nor U16903 (N_16903,N_16728,N_16605);
nor U16904 (N_16904,N_16782,N_16671);
xor U16905 (N_16905,N_16750,N_16655);
xor U16906 (N_16906,N_16620,N_16773);
and U16907 (N_16907,N_16761,N_16633);
nor U16908 (N_16908,N_16676,N_16723);
nand U16909 (N_16909,N_16682,N_16672);
xnor U16910 (N_16910,N_16617,N_16641);
or U16911 (N_16911,N_16642,N_16612);
nand U16912 (N_16912,N_16606,N_16627);
xnor U16913 (N_16913,N_16649,N_16799);
nor U16914 (N_16914,N_16666,N_16796);
nor U16915 (N_16915,N_16677,N_16683);
nor U16916 (N_16916,N_16608,N_16779);
or U16917 (N_16917,N_16657,N_16647);
or U16918 (N_16918,N_16787,N_16773);
nand U16919 (N_16919,N_16604,N_16786);
and U16920 (N_16920,N_16752,N_16649);
xor U16921 (N_16921,N_16749,N_16746);
xor U16922 (N_16922,N_16735,N_16648);
xnor U16923 (N_16923,N_16626,N_16787);
and U16924 (N_16924,N_16682,N_16711);
or U16925 (N_16925,N_16777,N_16691);
nand U16926 (N_16926,N_16683,N_16734);
xor U16927 (N_16927,N_16615,N_16722);
or U16928 (N_16928,N_16686,N_16621);
nand U16929 (N_16929,N_16654,N_16752);
nor U16930 (N_16930,N_16743,N_16771);
or U16931 (N_16931,N_16654,N_16785);
or U16932 (N_16932,N_16602,N_16666);
nand U16933 (N_16933,N_16722,N_16793);
or U16934 (N_16934,N_16604,N_16713);
xnor U16935 (N_16935,N_16756,N_16690);
nand U16936 (N_16936,N_16678,N_16673);
and U16937 (N_16937,N_16708,N_16746);
nand U16938 (N_16938,N_16737,N_16685);
nor U16939 (N_16939,N_16686,N_16714);
or U16940 (N_16940,N_16698,N_16719);
and U16941 (N_16941,N_16714,N_16738);
and U16942 (N_16942,N_16669,N_16646);
xnor U16943 (N_16943,N_16700,N_16678);
or U16944 (N_16944,N_16610,N_16680);
and U16945 (N_16945,N_16784,N_16693);
and U16946 (N_16946,N_16748,N_16653);
and U16947 (N_16947,N_16654,N_16718);
nand U16948 (N_16948,N_16692,N_16747);
xnor U16949 (N_16949,N_16607,N_16661);
or U16950 (N_16950,N_16640,N_16670);
xor U16951 (N_16951,N_16731,N_16782);
xnor U16952 (N_16952,N_16697,N_16639);
nor U16953 (N_16953,N_16661,N_16629);
nor U16954 (N_16954,N_16790,N_16623);
and U16955 (N_16955,N_16702,N_16738);
nand U16956 (N_16956,N_16626,N_16695);
and U16957 (N_16957,N_16713,N_16709);
and U16958 (N_16958,N_16691,N_16627);
nor U16959 (N_16959,N_16656,N_16724);
or U16960 (N_16960,N_16708,N_16799);
nand U16961 (N_16961,N_16796,N_16733);
or U16962 (N_16962,N_16661,N_16619);
or U16963 (N_16963,N_16652,N_16651);
and U16964 (N_16964,N_16708,N_16663);
nor U16965 (N_16965,N_16719,N_16752);
or U16966 (N_16966,N_16644,N_16694);
xor U16967 (N_16967,N_16784,N_16787);
xnor U16968 (N_16968,N_16661,N_16655);
or U16969 (N_16969,N_16686,N_16699);
or U16970 (N_16970,N_16641,N_16674);
or U16971 (N_16971,N_16687,N_16648);
xnor U16972 (N_16972,N_16741,N_16728);
nor U16973 (N_16973,N_16607,N_16725);
nor U16974 (N_16974,N_16625,N_16741);
nor U16975 (N_16975,N_16779,N_16762);
xor U16976 (N_16976,N_16794,N_16723);
xor U16977 (N_16977,N_16736,N_16782);
xnor U16978 (N_16978,N_16632,N_16780);
and U16979 (N_16979,N_16791,N_16714);
nor U16980 (N_16980,N_16650,N_16794);
nor U16981 (N_16981,N_16663,N_16686);
or U16982 (N_16982,N_16728,N_16782);
nand U16983 (N_16983,N_16704,N_16789);
xor U16984 (N_16984,N_16693,N_16728);
nand U16985 (N_16985,N_16776,N_16685);
nand U16986 (N_16986,N_16665,N_16705);
nor U16987 (N_16987,N_16633,N_16728);
nor U16988 (N_16988,N_16703,N_16641);
nor U16989 (N_16989,N_16618,N_16722);
and U16990 (N_16990,N_16633,N_16767);
xor U16991 (N_16991,N_16636,N_16654);
and U16992 (N_16992,N_16784,N_16708);
nand U16993 (N_16993,N_16661,N_16670);
and U16994 (N_16994,N_16622,N_16797);
nand U16995 (N_16995,N_16617,N_16679);
nor U16996 (N_16996,N_16764,N_16777);
xor U16997 (N_16997,N_16780,N_16703);
or U16998 (N_16998,N_16616,N_16744);
and U16999 (N_16999,N_16637,N_16741);
or U17000 (N_17000,N_16924,N_16861);
and U17001 (N_17001,N_16853,N_16919);
nand U17002 (N_17002,N_16979,N_16994);
xnor U17003 (N_17003,N_16995,N_16887);
xnor U17004 (N_17004,N_16841,N_16940);
xnor U17005 (N_17005,N_16873,N_16825);
nor U17006 (N_17006,N_16933,N_16833);
xnor U17007 (N_17007,N_16848,N_16943);
and U17008 (N_17008,N_16954,N_16870);
and U17009 (N_17009,N_16883,N_16959);
nand U17010 (N_17010,N_16880,N_16991);
nand U17011 (N_17011,N_16829,N_16903);
and U17012 (N_17012,N_16847,N_16857);
or U17013 (N_17013,N_16818,N_16850);
xor U17014 (N_17014,N_16974,N_16914);
and U17015 (N_17015,N_16926,N_16865);
nor U17016 (N_17016,N_16863,N_16931);
nand U17017 (N_17017,N_16891,N_16920);
and U17018 (N_17018,N_16886,N_16872);
nor U17019 (N_17019,N_16814,N_16937);
nor U17020 (N_17020,N_16821,N_16837);
or U17021 (N_17021,N_16985,N_16882);
xor U17022 (N_17022,N_16980,N_16934);
nor U17023 (N_17023,N_16961,N_16955);
xor U17024 (N_17024,N_16810,N_16942);
nor U17025 (N_17025,N_16984,N_16976);
and U17026 (N_17026,N_16944,N_16905);
nor U17027 (N_17027,N_16913,N_16827);
or U17028 (N_17028,N_16808,N_16895);
and U17029 (N_17029,N_16904,N_16890);
or U17030 (N_17030,N_16912,N_16845);
nor U17031 (N_17031,N_16909,N_16977);
xor U17032 (N_17032,N_16947,N_16932);
nor U17033 (N_17033,N_16978,N_16908);
nand U17034 (N_17034,N_16851,N_16876);
nor U17035 (N_17035,N_16982,N_16892);
xor U17036 (N_17036,N_16869,N_16800);
and U17037 (N_17037,N_16815,N_16889);
or U17038 (N_17038,N_16971,N_16834);
and U17039 (N_17039,N_16875,N_16826);
nor U17040 (N_17040,N_16948,N_16981);
xnor U17041 (N_17041,N_16806,N_16881);
or U17042 (N_17042,N_16956,N_16992);
xnor U17043 (N_17043,N_16858,N_16811);
nor U17044 (N_17044,N_16925,N_16813);
and U17045 (N_17045,N_16840,N_16949);
xor U17046 (N_17046,N_16824,N_16807);
nand U17047 (N_17047,N_16804,N_16987);
nand U17048 (N_17048,N_16859,N_16900);
or U17049 (N_17049,N_16822,N_16838);
or U17050 (N_17050,N_16816,N_16911);
nor U17051 (N_17051,N_16849,N_16820);
xor U17052 (N_17052,N_16953,N_16988);
nand U17053 (N_17053,N_16910,N_16965);
xnor U17054 (N_17054,N_16819,N_16832);
and U17055 (N_17055,N_16894,N_16946);
nand U17056 (N_17056,N_16999,N_16866);
nand U17057 (N_17057,N_16983,N_16964);
nor U17058 (N_17058,N_16868,N_16962);
nor U17059 (N_17059,N_16996,N_16916);
xor U17060 (N_17060,N_16823,N_16902);
xnor U17061 (N_17061,N_16839,N_16835);
xnor U17062 (N_17062,N_16852,N_16828);
xnor U17063 (N_17063,N_16855,N_16950);
nor U17064 (N_17064,N_16939,N_16836);
nor U17065 (N_17065,N_16871,N_16960);
nand U17066 (N_17066,N_16896,N_16930);
or U17067 (N_17067,N_16862,N_16923);
or U17068 (N_17068,N_16997,N_16990);
and U17069 (N_17069,N_16938,N_16812);
and U17070 (N_17070,N_16958,N_16975);
nand U17071 (N_17071,N_16805,N_16936);
nor U17072 (N_17072,N_16972,N_16879);
and U17073 (N_17073,N_16941,N_16856);
nor U17074 (N_17074,N_16921,N_16884);
xnor U17075 (N_17075,N_16901,N_16830);
nor U17076 (N_17076,N_16998,N_16952);
nand U17077 (N_17077,N_16842,N_16893);
or U17078 (N_17078,N_16802,N_16969);
or U17079 (N_17079,N_16877,N_16951);
and U17080 (N_17080,N_16973,N_16967);
nor U17081 (N_17081,N_16929,N_16957);
xor U17082 (N_17082,N_16915,N_16898);
nand U17083 (N_17083,N_16846,N_16945);
nand U17084 (N_17084,N_16809,N_16899);
xor U17085 (N_17085,N_16843,N_16888);
or U17086 (N_17086,N_16854,N_16803);
and U17087 (N_17087,N_16917,N_16860);
nand U17088 (N_17088,N_16966,N_16993);
nand U17089 (N_17089,N_16927,N_16844);
or U17090 (N_17090,N_16831,N_16864);
nand U17091 (N_17091,N_16986,N_16878);
xnor U17092 (N_17092,N_16970,N_16867);
and U17093 (N_17093,N_16906,N_16928);
nor U17094 (N_17094,N_16989,N_16874);
nor U17095 (N_17095,N_16968,N_16963);
nor U17096 (N_17096,N_16801,N_16922);
xnor U17097 (N_17097,N_16907,N_16935);
nor U17098 (N_17098,N_16885,N_16897);
and U17099 (N_17099,N_16817,N_16918);
nand U17100 (N_17100,N_16840,N_16973);
nor U17101 (N_17101,N_16945,N_16801);
nor U17102 (N_17102,N_16895,N_16993);
xor U17103 (N_17103,N_16964,N_16974);
or U17104 (N_17104,N_16914,N_16894);
and U17105 (N_17105,N_16888,N_16821);
xor U17106 (N_17106,N_16939,N_16829);
nor U17107 (N_17107,N_16997,N_16949);
or U17108 (N_17108,N_16939,N_16886);
or U17109 (N_17109,N_16929,N_16976);
or U17110 (N_17110,N_16860,N_16913);
or U17111 (N_17111,N_16832,N_16803);
nor U17112 (N_17112,N_16936,N_16806);
nor U17113 (N_17113,N_16937,N_16874);
xor U17114 (N_17114,N_16828,N_16880);
nor U17115 (N_17115,N_16820,N_16869);
nand U17116 (N_17116,N_16892,N_16852);
or U17117 (N_17117,N_16830,N_16874);
nor U17118 (N_17118,N_16930,N_16916);
and U17119 (N_17119,N_16999,N_16831);
or U17120 (N_17120,N_16860,N_16870);
nor U17121 (N_17121,N_16847,N_16885);
nand U17122 (N_17122,N_16977,N_16949);
or U17123 (N_17123,N_16960,N_16832);
xor U17124 (N_17124,N_16891,N_16968);
nor U17125 (N_17125,N_16850,N_16860);
nand U17126 (N_17126,N_16833,N_16845);
xor U17127 (N_17127,N_16927,N_16926);
nand U17128 (N_17128,N_16942,N_16927);
and U17129 (N_17129,N_16973,N_16890);
nand U17130 (N_17130,N_16947,N_16906);
xor U17131 (N_17131,N_16961,N_16943);
and U17132 (N_17132,N_16979,N_16876);
or U17133 (N_17133,N_16804,N_16999);
or U17134 (N_17134,N_16984,N_16850);
nor U17135 (N_17135,N_16977,N_16843);
nor U17136 (N_17136,N_16800,N_16851);
nor U17137 (N_17137,N_16862,N_16853);
or U17138 (N_17138,N_16939,N_16974);
and U17139 (N_17139,N_16953,N_16963);
nand U17140 (N_17140,N_16863,N_16895);
nand U17141 (N_17141,N_16865,N_16869);
or U17142 (N_17142,N_16945,N_16875);
and U17143 (N_17143,N_16948,N_16989);
and U17144 (N_17144,N_16987,N_16872);
nor U17145 (N_17145,N_16924,N_16841);
xor U17146 (N_17146,N_16996,N_16838);
and U17147 (N_17147,N_16948,N_16902);
or U17148 (N_17148,N_16825,N_16920);
nand U17149 (N_17149,N_16880,N_16893);
nand U17150 (N_17150,N_16896,N_16921);
and U17151 (N_17151,N_16867,N_16918);
nand U17152 (N_17152,N_16965,N_16985);
xor U17153 (N_17153,N_16857,N_16819);
nor U17154 (N_17154,N_16833,N_16964);
and U17155 (N_17155,N_16860,N_16886);
and U17156 (N_17156,N_16826,N_16857);
nand U17157 (N_17157,N_16984,N_16816);
or U17158 (N_17158,N_16822,N_16841);
and U17159 (N_17159,N_16829,N_16882);
nor U17160 (N_17160,N_16973,N_16969);
xnor U17161 (N_17161,N_16883,N_16906);
nand U17162 (N_17162,N_16871,N_16969);
xor U17163 (N_17163,N_16949,N_16815);
xor U17164 (N_17164,N_16818,N_16851);
xor U17165 (N_17165,N_16893,N_16920);
or U17166 (N_17166,N_16912,N_16873);
and U17167 (N_17167,N_16840,N_16948);
and U17168 (N_17168,N_16876,N_16939);
nand U17169 (N_17169,N_16865,N_16975);
or U17170 (N_17170,N_16812,N_16952);
and U17171 (N_17171,N_16960,N_16849);
nor U17172 (N_17172,N_16854,N_16945);
nor U17173 (N_17173,N_16981,N_16808);
and U17174 (N_17174,N_16959,N_16966);
nor U17175 (N_17175,N_16850,N_16979);
nor U17176 (N_17176,N_16878,N_16815);
xnor U17177 (N_17177,N_16952,N_16835);
xnor U17178 (N_17178,N_16903,N_16825);
and U17179 (N_17179,N_16966,N_16834);
and U17180 (N_17180,N_16935,N_16820);
or U17181 (N_17181,N_16817,N_16995);
xor U17182 (N_17182,N_16901,N_16940);
xnor U17183 (N_17183,N_16894,N_16834);
and U17184 (N_17184,N_16896,N_16940);
nand U17185 (N_17185,N_16919,N_16802);
or U17186 (N_17186,N_16896,N_16916);
nand U17187 (N_17187,N_16949,N_16982);
or U17188 (N_17188,N_16936,N_16809);
or U17189 (N_17189,N_16951,N_16815);
or U17190 (N_17190,N_16952,N_16831);
and U17191 (N_17191,N_16846,N_16821);
xnor U17192 (N_17192,N_16978,N_16882);
nand U17193 (N_17193,N_16868,N_16978);
nor U17194 (N_17194,N_16943,N_16860);
nor U17195 (N_17195,N_16982,N_16935);
nor U17196 (N_17196,N_16930,N_16966);
nand U17197 (N_17197,N_16917,N_16838);
xnor U17198 (N_17198,N_16993,N_16936);
nand U17199 (N_17199,N_16932,N_16898);
xnor U17200 (N_17200,N_17094,N_17035);
nand U17201 (N_17201,N_17073,N_17087);
nor U17202 (N_17202,N_17173,N_17186);
and U17203 (N_17203,N_17164,N_17066);
nor U17204 (N_17204,N_17093,N_17109);
or U17205 (N_17205,N_17132,N_17058);
nand U17206 (N_17206,N_17020,N_17004);
and U17207 (N_17207,N_17133,N_17027);
xor U17208 (N_17208,N_17131,N_17114);
nor U17209 (N_17209,N_17144,N_17100);
or U17210 (N_17210,N_17012,N_17129);
or U17211 (N_17211,N_17101,N_17130);
xor U17212 (N_17212,N_17134,N_17189);
nor U17213 (N_17213,N_17149,N_17019);
nand U17214 (N_17214,N_17167,N_17174);
xor U17215 (N_17215,N_17053,N_17067);
nor U17216 (N_17216,N_17071,N_17034);
nand U17217 (N_17217,N_17108,N_17003);
nor U17218 (N_17218,N_17143,N_17104);
nor U17219 (N_17219,N_17128,N_17113);
nand U17220 (N_17220,N_17013,N_17043);
and U17221 (N_17221,N_17054,N_17184);
nor U17222 (N_17222,N_17048,N_17115);
nand U17223 (N_17223,N_17009,N_17146);
or U17224 (N_17224,N_17086,N_17153);
or U17225 (N_17225,N_17060,N_17162);
nand U17226 (N_17226,N_17088,N_17148);
nand U17227 (N_17227,N_17125,N_17171);
nor U17228 (N_17228,N_17039,N_17092);
or U17229 (N_17229,N_17187,N_17000);
or U17230 (N_17230,N_17118,N_17036);
nor U17231 (N_17231,N_17079,N_17180);
nand U17232 (N_17232,N_17098,N_17029);
and U17233 (N_17233,N_17028,N_17191);
and U17234 (N_17234,N_17031,N_17078);
or U17235 (N_17235,N_17002,N_17007);
nand U17236 (N_17236,N_17099,N_17181);
xnor U17237 (N_17237,N_17001,N_17006);
and U17238 (N_17238,N_17188,N_17110);
and U17239 (N_17239,N_17056,N_17119);
xor U17240 (N_17240,N_17177,N_17135);
and U17241 (N_17241,N_17150,N_17089);
nand U17242 (N_17242,N_17175,N_17050);
nor U17243 (N_17243,N_17102,N_17084);
or U17244 (N_17244,N_17082,N_17085);
or U17245 (N_17245,N_17139,N_17185);
and U17246 (N_17246,N_17055,N_17192);
nor U17247 (N_17247,N_17011,N_17168);
and U17248 (N_17248,N_17198,N_17199);
nor U17249 (N_17249,N_17136,N_17033);
nand U17250 (N_17250,N_17176,N_17190);
nor U17251 (N_17251,N_17062,N_17025);
or U17252 (N_17252,N_17170,N_17010);
nor U17253 (N_17253,N_17091,N_17140);
or U17254 (N_17254,N_17122,N_17103);
or U17255 (N_17255,N_17074,N_17160);
nand U17256 (N_17256,N_17116,N_17032);
xnor U17257 (N_17257,N_17141,N_17106);
nand U17258 (N_17258,N_17080,N_17005);
and U17259 (N_17259,N_17037,N_17157);
xnor U17260 (N_17260,N_17096,N_17169);
nand U17261 (N_17261,N_17017,N_17016);
or U17262 (N_17262,N_17194,N_17156);
or U17263 (N_17263,N_17163,N_17166);
or U17264 (N_17264,N_17059,N_17142);
or U17265 (N_17265,N_17069,N_17138);
xor U17266 (N_17266,N_17161,N_17197);
or U17267 (N_17267,N_17049,N_17112);
or U17268 (N_17268,N_17018,N_17117);
nand U17269 (N_17269,N_17022,N_17083);
nor U17270 (N_17270,N_17057,N_17038);
or U17271 (N_17271,N_17145,N_17026);
or U17272 (N_17272,N_17076,N_17095);
xnor U17273 (N_17273,N_17172,N_17123);
xor U17274 (N_17274,N_17014,N_17042);
or U17275 (N_17275,N_17051,N_17024);
xnor U17276 (N_17276,N_17178,N_17147);
nor U17277 (N_17277,N_17030,N_17137);
nor U17278 (N_17278,N_17158,N_17040);
and U17279 (N_17279,N_17183,N_17068);
nor U17280 (N_17280,N_17107,N_17075);
or U17281 (N_17281,N_17070,N_17193);
nor U17282 (N_17282,N_17120,N_17121);
and U17283 (N_17283,N_17023,N_17111);
xnor U17284 (N_17284,N_17063,N_17195);
xnor U17285 (N_17285,N_17151,N_17090);
and U17286 (N_17286,N_17044,N_17061);
nor U17287 (N_17287,N_17196,N_17124);
and U17288 (N_17288,N_17152,N_17165);
or U17289 (N_17289,N_17081,N_17041);
nor U17290 (N_17290,N_17155,N_17072);
or U17291 (N_17291,N_17015,N_17179);
nand U17292 (N_17292,N_17046,N_17008);
or U17293 (N_17293,N_17047,N_17045);
or U17294 (N_17294,N_17182,N_17105);
xor U17295 (N_17295,N_17052,N_17077);
and U17296 (N_17296,N_17126,N_17065);
nand U17297 (N_17297,N_17154,N_17021);
nand U17298 (N_17298,N_17159,N_17097);
xnor U17299 (N_17299,N_17064,N_17127);
or U17300 (N_17300,N_17151,N_17191);
nor U17301 (N_17301,N_17176,N_17089);
or U17302 (N_17302,N_17090,N_17189);
xnor U17303 (N_17303,N_17111,N_17113);
xnor U17304 (N_17304,N_17046,N_17001);
xnor U17305 (N_17305,N_17048,N_17165);
xnor U17306 (N_17306,N_17113,N_17066);
or U17307 (N_17307,N_17005,N_17061);
nor U17308 (N_17308,N_17177,N_17100);
or U17309 (N_17309,N_17076,N_17049);
or U17310 (N_17310,N_17187,N_17121);
nor U17311 (N_17311,N_17063,N_17106);
xnor U17312 (N_17312,N_17091,N_17086);
nand U17313 (N_17313,N_17106,N_17171);
nand U17314 (N_17314,N_17085,N_17197);
nand U17315 (N_17315,N_17094,N_17195);
and U17316 (N_17316,N_17106,N_17008);
nor U17317 (N_17317,N_17112,N_17091);
or U17318 (N_17318,N_17001,N_17079);
nor U17319 (N_17319,N_17007,N_17056);
or U17320 (N_17320,N_17096,N_17057);
xnor U17321 (N_17321,N_17002,N_17074);
and U17322 (N_17322,N_17129,N_17075);
xor U17323 (N_17323,N_17102,N_17034);
nand U17324 (N_17324,N_17008,N_17069);
nand U17325 (N_17325,N_17008,N_17007);
and U17326 (N_17326,N_17088,N_17147);
nand U17327 (N_17327,N_17099,N_17138);
nand U17328 (N_17328,N_17058,N_17019);
or U17329 (N_17329,N_17039,N_17163);
or U17330 (N_17330,N_17175,N_17092);
or U17331 (N_17331,N_17087,N_17148);
or U17332 (N_17332,N_17115,N_17095);
nand U17333 (N_17333,N_17036,N_17153);
and U17334 (N_17334,N_17142,N_17164);
nor U17335 (N_17335,N_17133,N_17185);
and U17336 (N_17336,N_17079,N_17022);
nand U17337 (N_17337,N_17191,N_17195);
and U17338 (N_17338,N_17113,N_17092);
or U17339 (N_17339,N_17025,N_17054);
and U17340 (N_17340,N_17056,N_17141);
and U17341 (N_17341,N_17154,N_17070);
nor U17342 (N_17342,N_17153,N_17171);
or U17343 (N_17343,N_17121,N_17053);
nor U17344 (N_17344,N_17084,N_17077);
and U17345 (N_17345,N_17024,N_17169);
xnor U17346 (N_17346,N_17054,N_17046);
xnor U17347 (N_17347,N_17060,N_17075);
or U17348 (N_17348,N_17188,N_17073);
xnor U17349 (N_17349,N_17104,N_17019);
and U17350 (N_17350,N_17139,N_17103);
nor U17351 (N_17351,N_17180,N_17099);
nand U17352 (N_17352,N_17072,N_17149);
and U17353 (N_17353,N_17127,N_17070);
and U17354 (N_17354,N_17071,N_17110);
or U17355 (N_17355,N_17130,N_17168);
or U17356 (N_17356,N_17185,N_17106);
nor U17357 (N_17357,N_17072,N_17015);
or U17358 (N_17358,N_17069,N_17091);
and U17359 (N_17359,N_17132,N_17174);
nand U17360 (N_17360,N_17098,N_17004);
or U17361 (N_17361,N_17037,N_17170);
nor U17362 (N_17362,N_17042,N_17146);
or U17363 (N_17363,N_17102,N_17041);
xor U17364 (N_17364,N_17141,N_17132);
nor U17365 (N_17365,N_17073,N_17008);
xor U17366 (N_17366,N_17034,N_17020);
or U17367 (N_17367,N_17025,N_17005);
or U17368 (N_17368,N_17042,N_17114);
and U17369 (N_17369,N_17171,N_17090);
or U17370 (N_17370,N_17066,N_17156);
nor U17371 (N_17371,N_17146,N_17114);
nor U17372 (N_17372,N_17080,N_17191);
xnor U17373 (N_17373,N_17018,N_17152);
and U17374 (N_17374,N_17180,N_17167);
or U17375 (N_17375,N_17073,N_17047);
xor U17376 (N_17376,N_17018,N_17070);
and U17377 (N_17377,N_17000,N_17135);
nand U17378 (N_17378,N_17035,N_17198);
nand U17379 (N_17379,N_17140,N_17045);
xnor U17380 (N_17380,N_17001,N_17196);
nor U17381 (N_17381,N_17057,N_17172);
nand U17382 (N_17382,N_17161,N_17004);
xnor U17383 (N_17383,N_17015,N_17174);
nor U17384 (N_17384,N_17166,N_17030);
nor U17385 (N_17385,N_17174,N_17001);
and U17386 (N_17386,N_17078,N_17002);
nor U17387 (N_17387,N_17158,N_17077);
nor U17388 (N_17388,N_17071,N_17067);
nand U17389 (N_17389,N_17097,N_17092);
xor U17390 (N_17390,N_17129,N_17196);
nor U17391 (N_17391,N_17045,N_17026);
xnor U17392 (N_17392,N_17144,N_17119);
and U17393 (N_17393,N_17094,N_17051);
or U17394 (N_17394,N_17067,N_17063);
xor U17395 (N_17395,N_17140,N_17117);
or U17396 (N_17396,N_17070,N_17087);
nand U17397 (N_17397,N_17088,N_17142);
and U17398 (N_17398,N_17115,N_17098);
nor U17399 (N_17399,N_17086,N_17143);
xor U17400 (N_17400,N_17297,N_17236);
and U17401 (N_17401,N_17293,N_17295);
nand U17402 (N_17402,N_17288,N_17228);
and U17403 (N_17403,N_17243,N_17253);
nor U17404 (N_17404,N_17357,N_17309);
nand U17405 (N_17405,N_17338,N_17366);
nor U17406 (N_17406,N_17242,N_17279);
nor U17407 (N_17407,N_17300,N_17394);
nor U17408 (N_17408,N_17377,N_17212);
or U17409 (N_17409,N_17238,N_17332);
and U17410 (N_17410,N_17375,N_17321);
xor U17411 (N_17411,N_17319,N_17251);
nor U17412 (N_17412,N_17213,N_17223);
xor U17413 (N_17413,N_17203,N_17362);
nor U17414 (N_17414,N_17388,N_17313);
xnor U17415 (N_17415,N_17361,N_17214);
xor U17416 (N_17416,N_17344,N_17372);
and U17417 (N_17417,N_17327,N_17235);
xor U17418 (N_17418,N_17356,N_17333);
nand U17419 (N_17419,N_17353,N_17283);
nor U17420 (N_17420,N_17368,N_17285);
or U17421 (N_17421,N_17200,N_17231);
and U17422 (N_17422,N_17320,N_17264);
or U17423 (N_17423,N_17281,N_17289);
xnor U17424 (N_17424,N_17227,N_17343);
nand U17425 (N_17425,N_17269,N_17380);
nor U17426 (N_17426,N_17350,N_17364);
xnor U17427 (N_17427,N_17382,N_17329);
or U17428 (N_17428,N_17303,N_17294);
or U17429 (N_17429,N_17337,N_17274);
nor U17430 (N_17430,N_17229,N_17325);
or U17431 (N_17431,N_17314,N_17389);
nor U17432 (N_17432,N_17206,N_17399);
xnor U17433 (N_17433,N_17221,N_17345);
or U17434 (N_17434,N_17205,N_17398);
nor U17435 (N_17435,N_17275,N_17230);
nand U17436 (N_17436,N_17324,N_17347);
nor U17437 (N_17437,N_17348,N_17312);
nor U17438 (N_17438,N_17370,N_17385);
xor U17439 (N_17439,N_17260,N_17201);
xor U17440 (N_17440,N_17359,N_17298);
nor U17441 (N_17441,N_17393,N_17244);
nand U17442 (N_17442,N_17257,N_17373);
and U17443 (N_17443,N_17308,N_17358);
and U17444 (N_17444,N_17266,N_17277);
nor U17445 (N_17445,N_17261,N_17280);
or U17446 (N_17446,N_17323,N_17371);
or U17447 (N_17447,N_17392,N_17250);
or U17448 (N_17448,N_17255,N_17249);
xor U17449 (N_17449,N_17225,N_17335);
nand U17450 (N_17450,N_17349,N_17395);
xnor U17451 (N_17451,N_17219,N_17374);
nand U17452 (N_17452,N_17387,N_17311);
or U17453 (N_17453,N_17306,N_17384);
and U17454 (N_17454,N_17381,N_17296);
xnor U17455 (N_17455,N_17216,N_17322);
nand U17456 (N_17456,N_17271,N_17259);
nand U17457 (N_17457,N_17316,N_17270);
nand U17458 (N_17458,N_17217,N_17273);
or U17459 (N_17459,N_17352,N_17254);
nand U17460 (N_17460,N_17237,N_17367);
or U17461 (N_17461,N_17208,N_17334);
or U17462 (N_17462,N_17202,N_17272);
nor U17463 (N_17463,N_17252,N_17258);
or U17464 (N_17464,N_17204,N_17286);
and U17465 (N_17465,N_17376,N_17268);
and U17466 (N_17466,N_17310,N_17292);
nand U17467 (N_17467,N_17299,N_17224);
and U17468 (N_17468,N_17351,N_17354);
or U17469 (N_17469,N_17317,N_17207);
nand U17470 (N_17470,N_17397,N_17331);
nor U17471 (N_17471,N_17304,N_17276);
nand U17472 (N_17472,N_17226,N_17301);
nand U17473 (N_17473,N_17256,N_17302);
and U17474 (N_17474,N_17233,N_17247);
or U17475 (N_17475,N_17391,N_17278);
or U17476 (N_17476,N_17355,N_17220);
xor U17477 (N_17477,N_17383,N_17234);
and U17478 (N_17478,N_17318,N_17267);
and U17479 (N_17479,N_17240,N_17290);
xnor U17480 (N_17480,N_17379,N_17218);
and U17481 (N_17481,N_17239,N_17284);
xor U17482 (N_17482,N_17241,N_17291);
xnor U17483 (N_17483,N_17378,N_17246);
nand U17484 (N_17484,N_17328,N_17210);
xnor U17485 (N_17485,N_17330,N_17336);
nor U17486 (N_17486,N_17360,N_17307);
or U17487 (N_17487,N_17262,N_17396);
nor U17488 (N_17488,N_17211,N_17248);
nor U17489 (N_17489,N_17342,N_17369);
and U17490 (N_17490,N_17287,N_17365);
nand U17491 (N_17491,N_17245,N_17315);
nor U17492 (N_17492,N_17390,N_17340);
nor U17493 (N_17493,N_17232,N_17222);
or U17494 (N_17494,N_17282,N_17209);
or U17495 (N_17495,N_17363,N_17346);
or U17496 (N_17496,N_17215,N_17305);
or U17497 (N_17497,N_17265,N_17263);
nor U17498 (N_17498,N_17341,N_17339);
xnor U17499 (N_17499,N_17326,N_17386);
xor U17500 (N_17500,N_17258,N_17268);
nor U17501 (N_17501,N_17326,N_17286);
and U17502 (N_17502,N_17320,N_17378);
or U17503 (N_17503,N_17260,N_17262);
or U17504 (N_17504,N_17315,N_17287);
nand U17505 (N_17505,N_17263,N_17302);
and U17506 (N_17506,N_17347,N_17358);
and U17507 (N_17507,N_17227,N_17213);
and U17508 (N_17508,N_17200,N_17311);
or U17509 (N_17509,N_17267,N_17214);
or U17510 (N_17510,N_17229,N_17338);
or U17511 (N_17511,N_17227,N_17228);
nand U17512 (N_17512,N_17310,N_17232);
or U17513 (N_17513,N_17202,N_17283);
xor U17514 (N_17514,N_17300,N_17335);
xnor U17515 (N_17515,N_17233,N_17367);
xor U17516 (N_17516,N_17346,N_17244);
nand U17517 (N_17517,N_17373,N_17335);
nor U17518 (N_17518,N_17327,N_17350);
or U17519 (N_17519,N_17378,N_17211);
or U17520 (N_17520,N_17383,N_17302);
or U17521 (N_17521,N_17385,N_17294);
nand U17522 (N_17522,N_17304,N_17335);
or U17523 (N_17523,N_17382,N_17297);
or U17524 (N_17524,N_17205,N_17346);
nor U17525 (N_17525,N_17292,N_17398);
and U17526 (N_17526,N_17223,N_17241);
nor U17527 (N_17527,N_17237,N_17264);
nand U17528 (N_17528,N_17291,N_17367);
or U17529 (N_17529,N_17325,N_17235);
or U17530 (N_17530,N_17291,N_17285);
nor U17531 (N_17531,N_17350,N_17378);
nor U17532 (N_17532,N_17383,N_17318);
nor U17533 (N_17533,N_17267,N_17262);
xnor U17534 (N_17534,N_17362,N_17201);
and U17535 (N_17535,N_17224,N_17273);
and U17536 (N_17536,N_17302,N_17390);
nor U17537 (N_17537,N_17347,N_17221);
and U17538 (N_17538,N_17209,N_17338);
nand U17539 (N_17539,N_17221,N_17259);
nand U17540 (N_17540,N_17293,N_17247);
and U17541 (N_17541,N_17261,N_17339);
xor U17542 (N_17542,N_17244,N_17335);
xnor U17543 (N_17543,N_17351,N_17284);
nand U17544 (N_17544,N_17344,N_17258);
nand U17545 (N_17545,N_17351,N_17335);
nor U17546 (N_17546,N_17327,N_17385);
nor U17547 (N_17547,N_17356,N_17361);
xor U17548 (N_17548,N_17248,N_17363);
and U17549 (N_17549,N_17312,N_17217);
or U17550 (N_17550,N_17376,N_17246);
or U17551 (N_17551,N_17330,N_17239);
or U17552 (N_17552,N_17237,N_17390);
xor U17553 (N_17553,N_17378,N_17306);
and U17554 (N_17554,N_17292,N_17213);
or U17555 (N_17555,N_17298,N_17213);
nor U17556 (N_17556,N_17317,N_17235);
or U17557 (N_17557,N_17353,N_17218);
nand U17558 (N_17558,N_17311,N_17358);
nand U17559 (N_17559,N_17307,N_17378);
xnor U17560 (N_17560,N_17282,N_17229);
or U17561 (N_17561,N_17242,N_17272);
xor U17562 (N_17562,N_17280,N_17278);
nor U17563 (N_17563,N_17337,N_17369);
xor U17564 (N_17564,N_17376,N_17297);
nor U17565 (N_17565,N_17379,N_17281);
nand U17566 (N_17566,N_17325,N_17357);
and U17567 (N_17567,N_17322,N_17298);
nor U17568 (N_17568,N_17374,N_17202);
nand U17569 (N_17569,N_17274,N_17373);
nor U17570 (N_17570,N_17389,N_17228);
or U17571 (N_17571,N_17244,N_17275);
and U17572 (N_17572,N_17311,N_17208);
xnor U17573 (N_17573,N_17379,N_17239);
xor U17574 (N_17574,N_17326,N_17319);
and U17575 (N_17575,N_17262,N_17241);
and U17576 (N_17576,N_17214,N_17230);
nor U17577 (N_17577,N_17366,N_17396);
nand U17578 (N_17578,N_17289,N_17328);
or U17579 (N_17579,N_17389,N_17264);
nand U17580 (N_17580,N_17302,N_17227);
nand U17581 (N_17581,N_17205,N_17336);
or U17582 (N_17582,N_17340,N_17299);
nand U17583 (N_17583,N_17301,N_17375);
nor U17584 (N_17584,N_17377,N_17394);
nand U17585 (N_17585,N_17237,N_17284);
and U17586 (N_17586,N_17242,N_17232);
nor U17587 (N_17587,N_17335,N_17307);
and U17588 (N_17588,N_17298,N_17358);
xnor U17589 (N_17589,N_17376,N_17226);
or U17590 (N_17590,N_17296,N_17292);
or U17591 (N_17591,N_17332,N_17210);
and U17592 (N_17592,N_17307,N_17274);
and U17593 (N_17593,N_17236,N_17368);
and U17594 (N_17594,N_17268,N_17275);
nor U17595 (N_17595,N_17351,N_17313);
nand U17596 (N_17596,N_17245,N_17343);
and U17597 (N_17597,N_17207,N_17371);
nand U17598 (N_17598,N_17386,N_17399);
or U17599 (N_17599,N_17342,N_17282);
or U17600 (N_17600,N_17529,N_17460);
xor U17601 (N_17601,N_17519,N_17517);
or U17602 (N_17602,N_17575,N_17548);
nor U17603 (N_17603,N_17549,N_17560);
nand U17604 (N_17604,N_17562,N_17432);
or U17605 (N_17605,N_17435,N_17457);
xor U17606 (N_17606,N_17415,N_17459);
nand U17607 (N_17607,N_17533,N_17550);
nor U17608 (N_17608,N_17480,N_17443);
xnor U17609 (N_17609,N_17586,N_17483);
nor U17610 (N_17610,N_17447,N_17574);
nor U17611 (N_17611,N_17495,N_17493);
xor U17612 (N_17612,N_17425,N_17518);
or U17613 (N_17613,N_17451,N_17478);
nor U17614 (N_17614,N_17589,N_17405);
or U17615 (N_17615,N_17564,N_17458);
and U17616 (N_17616,N_17546,N_17410);
or U17617 (N_17617,N_17462,N_17540);
or U17618 (N_17618,N_17472,N_17416);
and U17619 (N_17619,N_17568,N_17599);
nand U17620 (N_17620,N_17565,N_17521);
or U17621 (N_17621,N_17542,N_17563);
and U17622 (N_17622,N_17488,N_17404);
or U17623 (N_17623,N_17492,N_17487);
nand U17624 (N_17624,N_17592,N_17406);
xor U17625 (N_17625,N_17420,N_17491);
nor U17626 (N_17626,N_17547,N_17580);
and U17627 (N_17627,N_17513,N_17531);
nor U17628 (N_17628,N_17584,N_17428);
nand U17629 (N_17629,N_17448,N_17507);
nand U17630 (N_17630,N_17494,N_17468);
nor U17631 (N_17631,N_17477,N_17515);
and U17632 (N_17632,N_17528,N_17411);
xnor U17633 (N_17633,N_17496,N_17409);
nor U17634 (N_17634,N_17585,N_17572);
xor U17635 (N_17635,N_17538,N_17421);
and U17636 (N_17636,N_17543,N_17536);
nand U17637 (N_17637,N_17429,N_17467);
nor U17638 (N_17638,N_17427,N_17583);
nand U17639 (N_17639,N_17527,N_17441);
xor U17640 (N_17640,N_17469,N_17481);
nor U17641 (N_17641,N_17530,N_17449);
or U17642 (N_17642,N_17401,N_17407);
nand U17643 (N_17643,N_17524,N_17578);
nor U17644 (N_17644,N_17450,N_17553);
or U17645 (N_17645,N_17556,N_17473);
and U17646 (N_17646,N_17593,N_17471);
nand U17647 (N_17647,N_17474,N_17512);
xor U17648 (N_17648,N_17508,N_17456);
and U17649 (N_17649,N_17567,N_17440);
nand U17650 (N_17650,N_17541,N_17596);
xor U17651 (N_17651,N_17412,N_17579);
xnor U17652 (N_17652,N_17511,N_17453);
nand U17653 (N_17653,N_17434,N_17597);
and U17654 (N_17654,N_17557,N_17402);
nor U17655 (N_17655,N_17506,N_17479);
xor U17656 (N_17656,N_17485,N_17570);
nor U17657 (N_17657,N_17582,N_17501);
xor U17658 (N_17658,N_17532,N_17475);
or U17659 (N_17659,N_17446,N_17523);
nor U17660 (N_17660,N_17516,N_17445);
xor U17661 (N_17661,N_17484,N_17490);
xnor U17662 (N_17662,N_17413,N_17520);
nand U17663 (N_17663,N_17418,N_17439);
xnor U17664 (N_17664,N_17559,N_17417);
or U17665 (N_17665,N_17577,N_17590);
xor U17666 (N_17666,N_17414,N_17576);
nand U17667 (N_17667,N_17482,N_17423);
xnor U17668 (N_17668,N_17581,N_17525);
xnor U17669 (N_17669,N_17499,N_17545);
or U17670 (N_17670,N_17424,N_17470);
nor U17671 (N_17671,N_17452,N_17500);
nand U17672 (N_17672,N_17408,N_17598);
xor U17673 (N_17673,N_17573,N_17505);
xnor U17674 (N_17674,N_17537,N_17431);
or U17675 (N_17675,N_17587,N_17438);
xor U17676 (N_17676,N_17403,N_17437);
and U17677 (N_17677,N_17498,N_17461);
nand U17678 (N_17678,N_17514,N_17558);
xor U17679 (N_17679,N_17509,N_17588);
nor U17680 (N_17680,N_17522,N_17463);
xnor U17681 (N_17681,N_17419,N_17486);
or U17682 (N_17682,N_17430,N_17426);
nand U17683 (N_17683,N_17534,N_17569);
xnor U17684 (N_17684,N_17489,N_17510);
nor U17685 (N_17685,N_17554,N_17442);
nor U17686 (N_17686,N_17552,N_17465);
nand U17687 (N_17687,N_17476,N_17535);
and U17688 (N_17688,N_17466,N_17455);
or U17689 (N_17689,N_17444,N_17591);
or U17690 (N_17690,N_17571,N_17561);
nor U17691 (N_17691,N_17551,N_17539);
nand U17692 (N_17692,N_17526,N_17503);
and U17693 (N_17693,N_17497,N_17436);
nand U17694 (N_17694,N_17502,N_17422);
nand U17695 (N_17695,N_17555,N_17400);
nand U17696 (N_17696,N_17544,N_17504);
xnor U17697 (N_17697,N_17566,N_17433);
nand U17698 (N_17698,N_17464,N_17454);
nor U17699 (N_17699,N_17594,N_17595);
xor U17700 (N_17700,N_17415,N_17544);
nor U17701 (N_17701,N_17486,N_17431);
nand U17702 (N_17702,N_17594,N_17546);
nand U17703 (N_17703,N_17438,N_17514);
or U17704 (N_17704,N_17481,N_17586);
nor U17705 (N_17705,N_17466,N_17458);
or U17706 (N_17706,N_17407,N_17400);
nand U17707 (N_17707,N_17422,N_17546);
xnor U17708 (N_17708,N_17501,N_17551);
and U17709 (N_17709,N_17584,N_17434);
nand U17710 (N_17710,N_17452,N_17481);
xnor U17711 (N_17711,N_17467,N_17413);
or U17712 (N_17712,N_17472,N_17442);
xnor U17713 (N_17713,N_17523,N_17531);
nand U17714 (N_17714,N_17526,N_17480);
and U17715 (N_17715,N_17491,N_17498);
and U17716 (N_17716,N_17456,N_17518);
and U17717 (N_17717,N_17503,N_17561);
or U17718 (N_17718,N_17425,N_17401);
nand U17719 (N_17719,N_17447,N_17529);
nor U17720 (N_17720,N_17581,N_17411);
xor U17721 (N_17721,N_17520,N_17442);
nor U17722 (N_17722,N_17442,N_17413);
or U17723 (N_17723,N_17547,N_17540);
and U17724 (N_17724,N_17458,N_17409);
xor U17725 (N_17725,N_17487,N_17534);
nor U17726 (N_17726,N_17592,N_17403);
xnor U17727 (N_17727,N_17411,N_17534);
nand U17728 (N_17728,N_17564,N_17445);
or U17729 (N_17729,N_17452,N_17430);
nand U17730 (N_17730,N_17490,N_17572);
nand U17731 (N_17731,N_17443,N_17477);
and U17732 (N_17732,N_17517,N_17501);
nor U17733 (N_17733,N_17598,N_17402);
and U17734 (N_17734,N_17453,N_17578);
and U17735 (N_17735,N_17541,N_17551);
nor U17736 (N_17736,N_17569,N_17540);
nor U17737 (N_17737,N_17429,N_17478);
or U17738 (N_17738,N_17421,N_17599);
nor U17739 (N_17739,N_17473,N_17464);
xnor U17740 (N_17740,N_17533,N_17421);
nand U17741 (N_17741,N_17596,N_17501);
or U17742 (N_17742,N_17429,N_17423);
xnor U17743 (N_17743,N_17568,N_17535);
and U17744 (N_17744,N_17424,N_17429);
nor U17745 (N_17745,N_17444,N_17539);
xor U17746 (N_17746,N_17585,N_17420);
nor U17747 (N_17747,N_17567,N_17546);
nand U17748 (N_17748,N_17400,N_17424);
nor U17749 (N_17749,N_17527,N_17489);
or U17750 (N_17750,N_17530,N_17596);
and U17751 (N_17751,N_17525,N_17462);
and U17752 (N_17752,N_17460,N_17568);
nand U17753 (N_17753,N_17421,N_17505);
and U17754 (N_17754,N_17541,N_17467);
xor U17755 (N_17755,N_17486,N_17577);
nand U17756 (N_17756,N_17582,N_17584);
xnor U17757 (N_17757,N_17445,N_17599);
nor U17758 (N_17758,N_17497,N_17443);
nand U17759 (N_17759,N_17583,N_17512);
xnor U17760 (N_17760,N_17586,N_17414);
or U17761 (N_17761,N_17550,N_17562);
or U17762 (N_17762,N_17562,N_17401);
and U17763 (N_17763,N_17498,N_17455);
and U17764 (N_17764,N_17423,N_17418);
or U17765 (N_17765,N_17544,N_17521);
xor U17766 (N_17766,N_17422,N_17541);
xnor U17767 (N_17767,N_17516,N_17528);
nor U17768 (N_17768,N_17406,N_17568);
nand U17769 (N_17769,N_17462,N_17581);
nand U17770 (N_17770,N_17449,N_17485);
or U17771 (N_17771,N_17402,N_17560);
nor U17772 (N_17772,N_17549,N_17484);
nand U17773 (N_17773,N_17570,N_17500);
xnor U17774 (N_17774,N_17494,N_17511);
or U17775 (N_17775,N_17505,N_17501);
xor U17776 (N_17776,N_17442,N_17458);
xnor U17777 (N_17777,N_17599,N_17475);
nor U17778 (N_17778,N_17444,N_17577);
nand U17779 (N_17779,N_17459,N_17554);
nor U17780 (N_17780,N_17533,N_17417);
and U17781 (N_17781,N_17412,N_17472);
nor U17782 (N_17782,N_17509,N_17440);
nand U17783 (N_17783,N_17532,N_17524);
and U17784 (N_17784,N_17553,N_17525);
or U17785 (N_17785,N_17476,N_17528);
nor U17786 (N_17786,N_17420,N_17507);
and U17787 (N_17787,N_17514,N_17489);
nor U17788 (N_17788,N_17406,N_17566);
or U17789 (N_17789,N_17477,N_17500);
or U17790 (N_17790,N_17485,N_17520);
or U17791 (N_17791,N_17536,N_17556);
nand U17792 (N_17792,N_17440,N_17540);
nand U17793 (N_17793,N_17590,N_17531);
or U17794 (N_17794,N_17481,N_17554);
and U17795 (N_17795,N_17420,N_17479);
nand U17796 (N_17796,N_17422,N_17412);
nand U17797 (N_17797,N_17458,N_17400);
and U17798 (N_17798,N_17575,N_17449);
and U17799 (N_17799,N_17405,N_17436);
nor U17800 (N_17800,N_17712,N_17747);
nor U17801 (N_17801,N_17622,N_17628);
or U17802 (N_17802,N_17771,N_17750);
and U17803 (N_17803,N_17710,N_17656);
nor U17804 (N_17804,N_17647,N_17705);
or U17805 (N_17805,N_17767,N_17641);
or U17806 (N_17806,N_17753,N_17607);
or U17807 (N_17807,N_17620,N_17789);
nor U17808 (N_17808,N_17758,N_17794);
and U17809 (N_17809,N_17681,N_17650);
xor U17810 (N_17810,N_17701,N_17602);
and U17811 (N_17811,N_17693,N_17636);
and U17812 (N_17812,N_17691,N_17670);
nand U17813 (N_17813,N_17726,N_17736);
nor U17814 (N_17814,N_17665,N_17731);
and U17815 (N_17815,N_17743,N_17612);
nor U17816 (N_17816,N_17708,N_17796);
nor U17817 (N_17817,N_17611,N_17734);
nand U17818 (N_17818,N_17741,N_17654);
nand U17819 (N_17819,N_17615,N_17746);
or U17820 (N_17820,N_17661,N_17754);
nand U17821 (N_17821,N_17777,N_17763);
and U17822 (N_17822,N_17732,N_17711);
nand U17823 (N_17823,N_17713,N_17660);
nand U17824 (N_17824,N_17694,N_17793);
xnor U17825 (N_17825,N_17677,N_17755);
nor U17826 (N_17826,N_17621,N_17657);
nor U17827 (N_17827,N_17652,N_17798);
or U17828 (N_17828,N_17604,N_17601);
xor U17829 (N_17829,N_17672,N_17630);
nor U17830 (N_17830,N_17714,N_17737);
nor U17831 (N_17831,N_17759,N_17724);
nor U17832 (N_17832,N_17618,N_17649);
or U17833 (N_17833,N_17664,N_17745);
nor U17834 (N_17834,N_17653,N_17682);
xor U17835 (N_17835,N_17686,N_17679);
or U17836 (N_17836,N_17678,N_17651);
and U17837 (N_17837,N_17695,N_17752);
and U17838 (N_17838,N_17613,N_17748);
and U17839 (N_17839,N_17709,N_17627);
nor U17840 (N_17840,N_17799,N_17716);
nand U17841 (N_17841,N_17635,N_17697);
or U17842 (N_17842,N_17676,N_17662);
nand U17843 (N_17843,N_17783,N_17603);
nand U17844 (N_17844,N_17766,N_17634);
nand U17845 (N_17845,N_17663,N_17778);
nor U17846 (N_17846,N_17702,N_17655);
nand U17847 (N_17847,N_17617,N_17614);
xnor U17848 (N_17848,N_17659,N_17648);
nor U17849 (N_17849,N_17623,N_17785);
nor U17850 (N_17850,N_17756,N_17715);
nand U17851 (N_17851,N_17761,N_17626);
nor U17852 (N_17852,N_17795,N_17770);
nor U17853 (N_17853,N_17768,N_17773);
or U17854 (N_17854,N_17674,N_17646);
nand U17855 (N_17855,N_17645,N_17772);
and U17856 (N_17856,N_17619,N_17669);
xnor U17857 (N_17857,N_17762,N_17632);
and U17858 (N_17858,N_17742,N_17703);
nand U17859 (N_17859,N_17722,N_17683);
nand U17860 (N_17860,N_17719,N_17718);
nor U17861 (N_17861,N_17675,N_17658);
nor U17862 (N_17862,N_17727,N_17765);
xnor U17863 (N_17863,N_17788,N_17775);
xor U17864 (N_17864,N_17606,N_17725);
nand U17865 (N_17865,N_17744,N_17738);
nand U17866 (N_17866,N_17637,N_17616);
nor U17867 (N_17867,N_17704,N_17690);
and U17868 (N_17868,N_17721,N_17642);
nor U17869 (N_17869,N_17685,N_17684);
nor U17870 (N_17870,N_17638,N_17720);
or U17871 (N_17871,N_17760,N_17643);
nor U17872 (N_17872,N_17780,N_17733);
and U17873 (N_17873,N_17740,N_17764);
nand U17874 (N_17874,N_17644,N_17781);
or U17875 (N_17875,N_17791,N_17605);
nand U17876 (N_17876,N_17739,N_17776);
xnor U17877 (N_17877,N_17728,N_17757);
and U17878 (N_17878,N_17609,N_17699);
or U17879 (N_17879,N_17717,N_17666);
nor U17880 (N_17880,N_17730,N_17784);
xor U17881 (N_17881,N_17625,N_17698);
nand U17882 (N_17882,N_17687,N_17729);
nand U17883 (N_17883,N_17797,N_17787);
xor U17884 (N_17884,N_17749,N_17610);
and U17885 (N_17885,N_17774,N_17782);
or U17886 (N_17886,N_17600,N_17786);
xor U17887 (N_17887,N_17671,N_17696);
nor U17888 (N_17888,N_17769,N_17629);
nand U17889 (N_17889,N_17790,N_17688);
and U17890 (N_17890,N_17633,N_17792);
nand U17891 (N_17891,N_17779,N_17706);
nand U17892 (N_17892,N_17667,N_17673);
nor U17893 (N_17893,N_17735,N_17668);
xor U17894 (N_17894,N_17608,N_17640);
nand U17895 (N_17895,N_17751,N_17723);
or U17896 (N_17896,N_17624,N_17631);
nand U17897 (N_17897,N_17700,N_17707);
or U17898 (N_17898,N_17692,N_17680);
or U17899 (N_17899,N_17639,N_17689);
nand U17900 (N_17900,N_17609,N_17679);
xnor U17901 (N_17901,N_17733,N_17661);
nand U17902 (N_17902,N_17616,N_17629);
and U17903 (N_17903,N_17712,N_17672);
nand U17904 (N_17904,N_17774,N_17606);
or U17905 (N_17905,N_17600,N_17693);
nand U17906 (N_17906,N_17628,N_17704);
and U17907 (N_17907,N_17653,N_17600);
and U17908 (N_17908,N_17601,N_17626);
and U17909 (N_17909,N_17696,N_17730);
xor U17910 (N_17910,N_17675,N_17770);
nor U17911 (N_17911,N_17683,N_17690);
nand U17912 (N_17912,N_17733,N_17727);
or U17913 (N_17913,N_17718,N_17706);
or U17914 (N_17914,N_17680,N_17793);
or U17915 (N_17915,N_17607,N_17773);
and U17916 (N_17916,N_17672,N_17601);
and U17917 (N_17917,N_17693,N_17627);
nand U17918 (N_17918,N_17628,N_17678);
nand U17919 (N_17919,N_17620,N_17626);
nand U17920 (N_17920,N_17644,N_17737);
xor U17921 (N_17921,N_17646,N_17706);
or U17922 (N_17922,N_17770,N_17643);
and U17923 (N_17923,N_17728,N_17775);
nand U17924 (N_17924,N_17792,N_17636);
nand U17925 (N_17925,N_17733,N_17747);
and U17926 (N_17926,N_17689,N_17634);
nand U17927 (N_17927,N_17602,N_17785);
xor U17928 (N_17928,N_17778,N_17752);
xor U17929 (N_17929,N_17719,N_17678);
and U17930 (N_17930,N_17719,N_17617);
or U17931 (N_17931,N_17721,N_17768);
nor U17932 (N_17932,N_17622,N_17755);
or U17933 (N_17933,N_17698,N_17700);
xor U17934 (N_17934,N_17674,N_17799);
or U17935 (N_17935,N_17631,N_17636);
or U17936 (N_17936,N_17658,N_17707);
nand U17937 (N_17937,N_17734,N_17717);
or U17938 (N_17938,N_17796,N_17606);
or U17939 (N_17939,N_17765,N_17651);
xnor U17940 (N_17940,N_17633,N_17728);
nor U17941 (N_17941,N_17609,N_17669);
nand U17942 (N_17942,N_17730,N_17642);
nand U17943 (N_17943,N_17770,N_17701);
nand U17944 (N_17944,N_17641,N_17739);
and U17945 (N_17945,N_17678,N_17741);
xor U17946 (N_17946,N_17733,N_17608);
and U17947 (N_17947,N_17732,N_17748);
and U17948 (N_17948,N_17724,N_17638);
xor U17949 (N_17949,N_17784,N_17725);
nand U17950 (N_17950,N_17688,N_17760);
xnor U17951 (N_17951,N_17781,N_17745);
nor U17952 (N_17952,N_17600,N_17763);
or U17953 (N_17953,N_17607,N_17755);
and U17954 (N_17954,N_17780,N_17628);
or U17955 (N_17955,N_17656,N_17723);
or U17956 (N_17956,N_17750,N_17773);
and U17957 (N_17957,N_17648,N_17738);
nor U17958 (N_17958,N_17631,N_17608);
xor U17959 (N_17959,N_17783,N_17693);
nor U17960 (N_17960,N_17713,N_17726);
and U17961 (N_17961,N_17678,N_17656);
xnor U17962 (N_17962,N_17677,N_17628);
nand U17963 (N_17963,N_17799,N_17631);
xnor U17964 (N_17964,N_17631,N_17763);
xnor U17965 (N_17965,N_17642,N_17612);
nand U17966 (N_17966,N_17768,N_17654);
nor U17967 (N_17967,N_17677,N_17750);
xnor U17968 (N_17968,N_17674,N_17749);
xor U17969 (N_17969,N_17742,N_17668);
or U17970 (N_17970,N_17692,N_17635);
nor U17971 (N_17971,N_17626,N_17709);
nor U17972 (N_17972,N_17638,N_17791);
xor U17973 (N_17973,N_17618,N_17614);
xnor U17974 (N_17974,N_17604,N_17745);
or U17975 (N_17975,N_17776,N_17635);
nand U17976 (N_17976,N_17608,N_17714);
nor U17977 (N_17977,N_17650,N_17603);
xor U17978 (N_17978,N_17734,N_17744);
nor U17979 (N_17979,N_17736,N_17635);
and U17980 (N_17980,N_17621,N_17663);
nor U17981 (N_17981,N_17657,N_17742);
xnor U17982 (N_17982,N_17745,N_17608);
xor U17983 (N_17983,N_17743,N_17751);
nand U17984 (N_17984,N_17790,N_17725);
nand U17985 (N_17985,N_17777,N_17620);
and U17986 (N_17986,N_17695,N_17763);
or U17987 (N_17987,N_17751,N_17670);
nor U17988 (N_17988,N_17616,N_17727);
xnor U17989 (N_17989,N_17665,N_17785);
and U17990 (N_17990,N_17777,N_17749);
or U17991 (N_17991,N_17671,N_17737);
and U17992 (N_17992,N_17669,N_17633);
and U17993 (N_17993,N_17607,N_17766);
and U17994 (N_17994,N_17623,N_17730);
xnor U17995 (N_17995,N_17716,N_17782);
nand U17996 (N_17996,N_17642,N_17724);
xnor U17997 (N_17997,N_17755,N_17789);
and U17998 (N_17998,N_17676,N_17670);
nand U17999 (N_17999,N_17703,N_17679);
and U18000 (N_18000,N_17872,N_17934);
and U18001 (N_18001,N_17926,N_17947);
nand U18002 (N_18002,N_17827,N_17861);
xor U18003 (N_18003,N_17885,N_17951);
nor U18004 (N_18004,N_17978,N_17937);
nor U18005 (N_18005,N_17830,N_17814);
nand U18006 (N_18006,N_17884,N_17913);
nand U18007 (N_18007,N_17834,N_17836);
or U18008 (N_18008,N_17971,N_17980);
xnor U18009 (N_18009,N_17974,N_17918);
nor U18010 (N_18010,N_17924,N_17805);
or U18011 (N_18011,N_17999,N_17994);
or U18012 (N_18012,N_17869,N_17952);
nand U18013 (N_18013,N_17990,N_17898);
and U18014 (N_18014,N_17929,N_17832);
or U18015 (N_18015,N_17841,N_17863);
xnor U18016 (N_18016,N_17903,N_17874);
or U18017 (N_18017,N_17866,N_17968);
xnor U18018 (N_18018,N_17995,N_17953);
xor U18019 (N_18019,N_17915,N_17916);
xnor U18020 (N_18020,N_17996,N_17993);
nor U18021 (N_18021,N_17960,N_17847);
and U18022 (N_18022,N_17806,N_17852);
nor U18023 (N_18023,N_17857,N_17826);
nor U18024 (N_18024,N_17939,N_17816);
nor U18025 (N_18025,N_17803,N_17901);
or U18026 (N_18026,N_17928,N_17844);
xor U18027 (N_18027,N_17867,N_17983);
xnor U18028 (N_18028,N_17908,N_17845);
and U18029 (N_18029,N_17919,N_17940);
nand U18030 (N_18030,N_17855,N_17840);
and U18031 (N_18031,N_17849,N_17865);
and U18032 (N_18032,N_17879,N_17900);
nand U18033 (N_18033,N_17889,N_17975);
nor U18034 (N_18034,N_17967,N_17820);
or U18035 (N_18035,N_17887,N_17818);
or U18036 (N_18036,N_17813,N_17949);
nand U18037 (N_18037,N_17970,N_17933);
and U18038 (N_18038,N_17808,N_17800);
nand U18039 (N_18039,N_17899,N_17930);
xor U18040 (N_18040,N_17810,N_17981);
nand U18041 (N_18041,N_17821,N_17833);
and U18042 (N_18042,N_17936,N_17911);
nor U18043 (N_18043,N_17825,N_17829);
xnor U18044 (N_18044,N_17846,N_17877);
nand U18045 (N_18045,N_17906,N_17895);
xnor U18046 (N_18046,N_17894,N_17956);
nand U18047 (N_18047,N_17853,N_17902);
or U18048 (N_18048,N_17905,N_17907);
and U18049 (N_18049,N_17950,N_17969);
and U18050 (N_18050,N_17858,N_17987);
or U18051 (N_18051,N_17946,N_17997);
or U18052 (N_18052,N_17988,N_17882);
and U18053 (N_18053,N_17839,N_17938);
or U18054 (N_18054,N_17973,N_17965);
and U18055 (N_18055,N_17864,N_17870);
or U18056 (N_18056,N_17896,N_17986);
xnor U18057 (N_18057,N_17977,N_17878);
nor U18058 (N_18058,N_17935,N_17961);
nand U18059 (N_18059,N_17881,N_17955);
nor U18060 (N_18060,N_17823,N_17860);
or U18061 (N_18061,N_17944,N_17850);
or U18062 (N_18062,N_17856,N_17972);
nand U18063 (N_18063,N_17912,N_17876);
or U18064 (N_18064,N_17809,N_17959);
xnor U18065 (N_18065,N_17835,N_17851);
nor U18066 (N_18066,N_17824,N_17875);
and U18067 (N_18067,N_17942,N_17848);
nor U18068 (N_18068,N_17931,N_17893);
nand U18069 (N_18069,N_17957,N_17910);
nand U18070 (N_18070,N_17843,N_17892);
nor U18071 (N_18071,N_17891,N_17802);
xor U18072 (N_18072,N_17964,N_17862);
nand U18073 (N_18073,N_17941,N_17932);
nand U18074 (N_18074,N_17925,N_17917);
xnor U18075 (N_18075,N_17914,N_17909);
or U18076 (N_18076,N_17812,N_17945);
xor U18077 (N_18077,N_17831,N_17963);
or U18078 (N_18078,N_17958,N_17948);
xor U18079 (N_18079,N_17991,N_17871);
or U18080 (N_18080,N_17854,N_17927);
and U18081 (N_18081,N_17920,N_17888);
nor U18082 (N_18082,N_17897,N_17837);
or U18083 (N_18083,N_17859,N_17998);
and U18084 (N_18084,N_17966,N_17890);
nor U18085 (N_18085,N_17904,N_17842);
nand U18086 (N_18086,N_17868,N_17984);
and U18087 (N_18087,N_17828,N_17807);
nor U18088 (N_18088,N_17979,N_17943);
and U18089 (N_18089,N_17886,N_17822);
nand U18090 (N_18090,N_17954,N_17982);
xor U18091 (N_18091,N_17922,N_17819);
and U18092 (N_18092,N_17985,N_17815);
and U18093 (N_18093,N_17811,N_17804);
nor U18094 (N_18094,N_17817,N_17989);
nand U18095 (N_18095,N_17801,N_17873);
xnor U18096 (N_18096,N_17976,N_17992);
and U18097 (N_18097,N_17838,N_17880);
nor U18098 (N_18098,N_17923,N_17962);
nor U18099 (N_18099,N_17921,N_17883);
nor U18100 (N_18100,N_17832,N_17942);
and U18101 (N_18101,N_17998,N_17847);
or U18102 (N_18102,N_17889,N_17910);
xnor U18103 (N_18103,N_17920,N_17813);
or U18104 (N_18104,N_17930,N_17889);
xor U18105 (N_18105,N_17971,N_17999);
and U18106 (N_18106,N_17990,N_17979);
nand U18107 (N_18107,N_17814,N_17844);
nand U18108 (N_18108,N_17813,N_17892);
and U18109 (N_18109,N_17877,N_17890);
nor U18110 (N_18110,N_17969,N_17889);
and U18111 (N_18111,N_17878,N_17852);
nor U18112 (N_18112,N_17956,N_17939);
or U18113 (N_18113,N_17952,N_17923);
nor U18114 (N_18114,N_17916,N_17803);
xnor U18115 (N_18115,N_17865,N_17809);
nand U18116 (N_18116,N_17844,N_17936);
or U18117 (N_18117,N_17851,N_17907);
xnor U18118 (N_18118,N_17818,N_17994);
nor U18119 (N_18119,N_17984,N_17982);
or U18120 (N_18120,N_17809,N_17958);
nor U18121 (N_18121,N_17936,N_17950);
and U18122 (N_18122,N_17856,N_17936);
xnor U18123 (N_18123,N_17896,N_17918);
or U18124 (N_18124,N_17895,N_17891);
nor U18125 (N_18125,N_17975,N_17846);
nand U18126 (N_18126,N_17825,N_17809);
xnor U18127 (N_18127,N_17825,N_17943);
and U18128 (N_18128,N_17926,N_17802);
and U18129 (N_18129,N_17997,N_17847);
nor U18130 (N_18130,N_17912,N_17916);
or U18131 (N_18131,N_17966,N_17807);
and U18132 (N_18132,N_17992,N_17948);
xnor U18133 (N_18133,N_17947,N_17950);
or U18134 (N_18134,N_17833,N_17880);
nand U18135 (N_18135,N_17832,N_17806);
nor U18136 (N_18136,N_17985,N_17964);
xnor U18137 (N_18137,N_17907,N_17818);
or U18138 (N_18138,N_17841,N_17814);
and U18139 (N_18139,N_17924,N_17921);
or U18140 (N_18140,N_17844,N_17884);
nor U18141 (N_18141,N_17836,N_17920);
xor U18142 (N_18142,N_17926,N_17994);
xor U18143 (N_18143,N_17916,N_17987);
xor U18144 (N_18144,N_17902,N_17990);
nor U18145 (N_18145,N_17893,N_17899);
xor U18146 (N_18146,N_17980,N_17817);
and U18147 (N_18147,N_17991,N_17950);
nor U18148 (N_18148,N_17929,N_17800);
and U18149 (N_18149,N_17912,N_17894);
and U18150 (N_18150,N_17993,N_17979);
nor U18151 (N_18151,N_17908,N_17998);
xnor U18152 (N_18152,N_17886,N_17923);
xnor U18153 (N_18153,N_17983,N_17935);
xnor U18154 (N_18154,N_17865,N_17831);
and U18155 (N_18155,N_17964,N_17969);
nor U18156 (N_18156,N_17815,N_17978);
nand U18157 (N_18157,N_17980,N_17946);
nor U18158 (N_18158,N_17909,N_17930);
nand U18159 (N_18159,N_17929,N_17932);
or U18160 (N_18160,N_17913,N_17839);
or U18161 (N_18161,N_17879,N_17928);
nor U18162 (N_18162,N_17900,N_17803);
and U18163 (N_18163,N_17952,N_17992);
xor U18164 (N_18164,N_17968,N_17999);
nand U18165 (N_18165,N_17926,N_17848);
or U18166 (N_18166,N_17842,N_17955);
and U18167 (N_18167,N_17987,N_17922);
or U18168 (N_18168,N_17978,N_17976);
or U18169 (N_18169,N_17924,N_17945);
nand U18170 (N_18170,N_17838,N_17870);
xnor U18171 (N_18171,N_17964,N_17863);
xor U18172 (N_18172,N_17959,N_17827);
nor U18173 (N_18173,N_17985,N_17855);
xnor U18174 (N_18174,N_17865,N_17961);
nor U18175 (N_18175,N_17844,N_17985);
or U18176 (N_18176,N_17896,N_17833);
and U18177 (N_18177,N_17921,N_17822);
or U18178 (N_18178,N_17830,N_17835);
nand U18179 (N_18179,N_17860,N_17895);
and U18180 (N_18180,N_17948,N_17953);
nor U18181 (N_18181,N_17883,N_17860);
xnor U18182 (N_18182,N_17850,N_17863);
xnor U18183 (N_18183,N_17962,N_17856);
or U18184 (N_18184,N_17968,N_17835);
nor U18185 (N_18185,N_17980,N_17995);
xnor U18186 (N_18186,N_17946,N_17824);
or U18187 (N_18187,N_17981,N_17892);
or U18188 (N_18188,N_17875,N_17852);
or U18189 (N_18189,N_17921,N_17997);
or U18190 (N_18190,N_17886,N_17855);
and U18191 (N_18191,N_17837,N_17951);
and U18192 (N_18192,N_17948,N_17969);
xnor U18193 (N_18193,N_17893,N_17883);
or U18194 (N_18194,N_17855,N_17860);
nor U18195 (N_18195,N_17857,N_17873);
or U18196 (N_18196,N_17941,N_17929);
xor U18197 (N_18197,N_17823,N_17953);
nand U18198 (N_18198,N_17907,N_17801);
or U18199 (N_18199,N_17853,N_17919);
nor U18200 (N_18200,N_18125,N_18192);
or U18201 (N_18201,N_18128,N_18168);
nand U18202 (N_18202,N_18076,N_18098);
or U18203 (N_18203,N_18084,N_18153);
and U18204 (N_18204,N_18010,N_18115);
nor U18205 (N_18205,N_18004,N_18081);
nor U18206 (N_18206,N_18119,N_18180);
nor U18207 (N_18207,N_18034,N_18197);
or U18208 (N_18208,N_18104,N_18056);
or U18209 (N_18209,N_18186,N_18018);
nand U18210 (N_18210,N_18089,N_18090);
nand U18211 (N_18211,N_18059,N_18072);
and U18212 (N_18212,N_18163,N_18091);
or U18213 (N_18213,N_18196,N_18199);
xnor U18214 (N_18214,N_18039,N_18105);
or U18215 (N_18215,N_18130,N_18007);
and U18216 (N_18216,N_18166,N_18177);
or U18217 (N_18217,N_18053,N_18086);
or U18218 (N_18218,N_18013,N_18092);
nand U18219 (N_18219,N_18117,N_18073);
and U18220 (N_18220,N_18055,N_18083);
nand U18221 (N_18221,N_18079,N_18151);
nor U18222 (N_18222,N_18155,N_18139);
or U18223 (N_18223,N_18003,N_18126);
or U18224 (N_18224,N_18001,N_18103);
or U18225 (N_18225,N_18127,N_18148);
or U18226 (N_18226,N_18136,N_18071);
xnor U18227 (N_18227,N_18100,N_18142);
nor U18228 (N_18228,N_18077,N_18191);
nand U18229 (N_18229,N_18044,N_18048);
nor U18230 (N_18230,N_18158,N_18114);
nand U18231 (N_18231,N_18030,N_18016);
xor U18232 (N_18232,N_18164,N_18137);
xnor U18233 (N_18233,N_18135,N_18049);
or U18234 (N_18234,N_18122,N_18012);
and U18235 (N_18235,N_18160,N_18140);
xor U18236 (N_18236,N_18124,N_18096);
xor U18237 (N_18237,N_18069,N_18181);
nand U18238 (N_18238,N_18041,N_18133);
xnor U18239 (N_18239,N_18040,N_18037);
or U18240 (N_18240,N_18015,N_18146);
xor U18241 (N_18241,N_18147,N_18009);
xor U18242 (N_18242,N_18107,N_18198);
nand U18243 (N_18243,N_18029,N_18118);
and U18244 (N_18244,N_18087,N_18052);
xnor U18245 (N_18245,N_18162,N_18167);
and U18246 (N_18246,N_18057,N_18182);
xnor U18247 (N_18247,N_18129,N_18108);
nand U18248 (N_18248,N_18165,N_18102);
nand U18249 (N_18249,N_18141,N_18111);
or U18250 (N_18250,N_18112,N_18033);
or U18251 (N_18251,N_18179,N_18188);
xnor U18252 (N_18252,N_18131,N_18183);
nand U18253 (N_18253,N_18176,N_18157);
or U18254 (N_18254,N_18022,N_18078);
nor U18255 (N_18255,N_18132,N_18085);
nor U18256 (N_18256,N_18043,N_18035);
nor U18257 (N_18257,N_18050,N_18047);
xor U18258 (N_18258,N_18144,N_18066);
and U18259 (N_18259,N_18194,N_18024);
and U18260 (N_18260,N_18099,N_18193);
and U18261 (N_18261,N_18172,N_18025);
or U18262 (N_18262,N_18045,N_18002);
xnor U18263 (N_18263,N_18110,N_18169);
nor U18264 (N_18264,N_18070,N_18005);
nand U18265 (N_18265,N_18143,N_18171);
nor U18266 (N_18266,N_18145,N_18011);
xnor U18267 (N_18267,N_18093,N_18095);
nand U18268 (N_18268,N_18082,N_18021);
and U18269 (N_18269,N_18152,N_18051);
or U18270 (N_18270,N_18074,N_18195);
and U18271 (N_18271,N_18032,N_18097);
or U18272 (N_18272,N_18116,N_18189);
nand U18273 (N_18273,N_18062,N_18170);
and U18274 (N_18274,N_18088,N_18138);
nand U18275 (N_18275,N_18161,N_18064);
xor U18276 (N_18276,N_18023,N_18065);
nor U18277 (N_18277,N_18101,N_18113);
nand U18278 (N_18278,N_18067,N_18061);
xor U18279 (N_18279,N_18121,N_18173);
nand U18280 (N_18280,N_18075,N_18109);
and U18281 (N_18281,N_18185,N_18080);
nand U18282 (N_18282,N_18017,N_18054);
nor U18283 (N_18283,N_18038,N_18019);
nor U18284 (N_18284,N_18031,N_18175);
nand U18285 (N_18285,N_18008,N_18150);
nand U18286 (N_18286,N_18026,N_18159);
nand U18287 (N_18287,N_18058,N_18094);
nand U18288 (N_18288,N_18027,N_18106);
nand U18289 (N_18289,N_18174,N_18000);
xnor U18290 (N_18290,N_18156,N_18120);
or U18291 (N_18291,N_18006,N_18068);
xor U18292 (N_18292,N_18187,N_18014);
or U18293 (N_18293,N_18020,N_18184);
nor U18294 (N_18294,N_18134,N_18046);
and U18295 (N_18295,N_18060,N_18154);
nand U18296 (N_18296,N_18190,N_18028);
or U18297 (N_18297,N_18042,N_18123);
or U18298 (N_18298,N_18149,N_18178);
nor U18299 (N_18299,N_18036,N_18063);
xnor U18300 (N_18300,N_18143,N_18007);
nand U18301 (N_18301,N_18000,N_18139);
nor U18302 (N_18302,N_18004,N_18022);
nand U18303 (N_18303,N_18142,N_18038);
nand U18304 (N_18304,N_18176,N_18113);
nand U18305 (N_18305,N_18155,N_18041);
and U18306 (N_18306,N_18065,N_18056);
nand U18307 (N_18307,N_18050,N_18152);
nand U18308 (N_18308,N_18003,N_18048);
and U18309 (N_18309,N_18154,N_18096);
or U18310 (N_18310,N_18139,N_18168);
nand U18311 (N_18311,N_18183,N_18198);
xor U18312 (N_18312,N_18015,N_18071);
nor U18313 (N_18313,N_18040,N_18005);
and U18314 (N_18314,N_18175,N_18081);
and U18315 (N_18315,N_18178,N_18107);
nand U18316 (N_18316,N_18020,N_18149);
nand U18317 (N_18317,N_18084,N_18051);
and U18318 (N_18318,N_18066,N_18077);
or U18319 (N_18319,N_18132,N_18035);
nor U18320 (N_18320,N_18113,N_18053);
nor U18321 (N_18321,N_18126,N_18093);
xor U18322 (N_18322,N_18121,N_18096);
and U18323 (N_18323,N_18142,N_18163);
and U18324 (N_18324,N_18127,N_18074);
or U18325 (N_18325,N_18124,N_18108);
xnor U18326 (N_18326,N_18046,N_18056);
or U18327 (N_18327,N_18135,N_18095);
or U18328 (N_18328,N_18193,N_18179);
and U18329 (N_18329,N_18085,N_18086);
nand U18330 (N_18330,N_18097,N_18096);
or U18331 (N_18331,N_18039,N_18056);
xor U18332 (N_18332,N_18056,N_18165);
nand U18333 (N_18333,N_18130,N_18096);
nor U18334 (N_18334,N_18177,N_18064);
xor U18335 (N_18335,N_18045,N_18001);
nand U18336 (N_18336,N_18176,N_18017);
nand U18337 (N_18337,N_18136,N_18146);
and U18338 (N_18338,N_18157,N_18181);
or U18339 (N_18339,N_18167,N_18004);
nand U18340 (N_18340,N_18042,N_18002);
nand U18341 (N_18341,N_18109,N_18140);
or U18342 (N_18342,N_18071,N_18120);
or U18343 (N_18343,N_18090,N_18087);
nand U18344 (N_18344,N_18073,N_18155);
nor U18345 (N_18345,N_18153,N_18194);
nor U18346 (N_18346,N_18010,N_18094);
nor U18347 (N_18347,N_18184,N_18025);
or U18348 (N_18348,N_18096,N_18161);
and U18349 (N_18349,N_18127,N_18184);
and U18350 (N_18350,N_18091,N_18071);
nand U18351 (N_18351,N_18199,N_18075);
or U18352 (N_18352,N_18073,N_18088);
or U18353 (N_18353,N_18066,N_18175);
xnor U18354 (N_18354,N_18018,N_18019);
or U18355 (N_18355,N_18024,N_18170);
xnor U18356 (N_18356,N_18006,N_18198);
or U18357 (N_18357,N_18107,N_18042);
xor U18358 (N_18358,N_18060,N_18043);
nor U18359 (N_18359,N_18012,N_18175);
or U18360 (N_18360,N_18179,N_18091);
nor U18361 (N_18361,N_18165,N_18180);
xnor U18362 (N_18362,N_18118,N_18192);
and U18363 (N_18363,N_18038,N_18108);
nor U18364 (N_18364,N_18071,N_18059);
nor U18365 (N_18365,N_18006,N_18060);
nand U18366 (N_18366,N_18197,N_18093);
or U18367 (N_18367,N_18008,N_18067);
xnor U18368 (N_18368,N_18184,N_18166);
and U18369 (N_18369,N_18048,N_18006);
or U18370 (N_18370,N_18034,N_18141);
xnor U18371 (N_18371,N_18067,N_18108);
or U18372 (N_18372,N_18097,N_18040);
nand U18373 (N_18373,N_18103,N_18071);
nor U18374 (N_18374,N_18085,N_18154);
xor U18375 (N_18375,N_18029,N_18153);
xnor U18376 (N_18376,N_18082,N_18061);
nand U18377 (N_18377,N_18118,N_18088);
xnor U18378 (N_18378,N_18139,N_18055);
nor U18379 (N_18379,N_18143,N_18081);
or U18380 (N_18380,N_18152,N_18073);
nand U18381 (N_18381,N_18085,N_18184);
and U18382 (N_18382,N_18092,N_18018);
nand U18383 (N_18383,N_18104,N_18021);
and U18384 (N_18384,N_18128,N_18163);
or U18385 (N_18385,N_18123,N_18076);
xnor U18386 (N_18386,N_18112,N_18020);
xor U18387 (N_18387,N_18036,N_18009);
nor U18388 (N_18388,N_18064,N_18123);
and U18389 (N_18389,N_18196,N_18065);
xor U18390 (N_18390,N_18037,N_18151);
xor U18391 (N_18391,N_18043,N_18183);
or U18392 (N_18392,N_18176,N_18065);
nor U18393 (N_18393,N_18131,N_18181);
xor U18394 (N_18394,N_18044,N_18011);
xnor U18395 (N_18395,N_18039,N_18098);
nor U18396 (N_18396,N_18086,N_18126);
xnor U18397 (N_18397,N_18140,N_18039);
or U18398 (N_18398,N_18166,N_18125);
nor U18399 (N_18399,N_18031,N_18083);
or U18400 (N_18400,N_18201,N_18323);
and U18401 (N_18401,N_18292,N_18215);
and U18402 (N_18402,N_18342,N_18280);
nand U18403 (N_18403,N_18209,N_18336);
nand U18404 (N_18404,N_18243,N_18312);
and U18405 (N_18405,N_18377,N_18208);
nor U18406 (N_18406,N_18315,N_18265);
or U18407 (N_18407,N_18356,N_18269);
and U18408 (N_18408,N_18255,N_18233);
nand U18409 (N_18409,N_18277,N_18373);
xnor U18410 (N_18410,N_18202,N_18392);
nor U18411 (N_18411,N_18319,N_18311);
and U18412 (N_18412,N_18276,N_18262);
and U18413 (N_18413,N_18317,N_18388);
xnor U18414 (N_18414,N_18258,N_18338);
or U18415 (N_18415,N_18207,N_18318);
xor U18416 (N_18416,N_18221,N_18264);
nor U18417 (N_18417,N_18223,N_18375);
xor U18418 (N_18418,N_18306,N_18217);
nand U18419 (N_18419,N_18297,N_18316);
and U18420 (N_18420,N_18353,N_18372);
or U18421 (N_18421,N_18250,N_18396);
nor U18422 (N_18422,N_18352,N_18256);
or U18423 (N_18423,N_18299,N_18349);
nor U18424 (N_18424,N_18360,N_18385);
and U18425 (N_18425,N_18290,N_18273);
nor U18426 (N_18426,N_18357,N_18270);
xnor U18427 (N_18427,N_18218,N_18259);
nand U18428 (N_18428,N_18206,N_18278);
or U18429 (N_18429,N_18271,N_18231);
xnor U18430 (N_18430,N_18399,N_18298);
nor U18431 (N_18431,N_18252,N_18241);
nor U18432 (N_18432,N_18322,N_18348);
nand U18433 (N_18433,N_18397,N_18267);
or U18434 (N_18434,N_18227,N_18328);
nor U18435 (N_18435,N_18331,N_18314);
nand U18436 (N_18436,N_18393,N_18275);
nor U18437 (N_18437,N_18214,N_18367);
nand U18438 (N_18438,N_18391,N_18358);
xnor U18439 (N_18439,N_18390,N_18324);
and U18440 (N_18440,N_18363,N_18370);
xor U18441 (N_18441,N_18347,N_18237);
xor U18442 (N_18442,N_18309,N_18302);
xor U18443 (N_18443,N_18266,N_18220);
and U18444 (N_18444,N_18283,N_18383);
nand U18445 (N_18445,N_18253,N_18350);
and U18446 (N_18446,N_18320,N_18313);
nand U18447 (N_18447,N_18294,N_18282);
xor U18448 (N_18448,N_18235,N_18288);
xnor U18449 (N_18449,N_18395,N_18242);
xor U18450 (N_18450,N_18291,N_18389);
xnor U18451 (N_18451,N_18329,N_18210);
xnor U18452 (N_18452,N_18268,N_18371);
or U18453 (N_18453,N_18248,N_18272);
nand U18454 (N_18454,N_18339,N_18226);
and U18455 (N_18455,N_18335,N_18213);
xnor U18456 (N_18456,N_18257,N_18244);
nor U18457 (N_18457,N_18364,N_18378);
or U18458 (N_18458,N_18310,N_18216);
nand U18459 (N_18459,N_18366,N_18200);
nor U18460 (N_18460,N_18379,N_18344);
and U18461 (N_18461,N_18254,N_18212);
nand U18462 (N_18462,N_18387,N_18345);
or U18463 (N_18463,N_18332,N_18203);
xor U18464 (N_18464,N_18238,N_18304);
nor U18465 (N_18465,N_18308,N_18260);
nand U18466 (N_18466,N_18285,N_18386);
and U18467 (N_18467,N_18205,N_18251);
xor U18468 (N_18468,N_18307,N_18239);
nor U18469 (N_18469,N_18296,N_18263);
xnor U18470 (N_18470,N_18368,N_18230);
and U18471 (N_18471,N_18279,N_18204);
nand U18472 (N_18472,N_18382,N_18362);
nor U18473 (N_18473,N_18384,N_18234);
or U18474 (N_18474,N_18289,N_18359);
nand U18475 (N_18475,N_18274,N_18327);
and U18476 (N_18476,N_18346,N_18249);
and U18477 (N_18477,N_18246,N_18343);
and U18478 (N_18478,N_18240,N_18295);
nand U18479 (N_18479,N_18337,N_18380);
xor U18480 (N_18480,N_18224,N_18355);
or U18481 (N_18481,N_18376,N_18361);
and U18482 (N_18482,N_18287,N_18281);
or U18483 (N_18483,N_18333,N_18398);
and U18484 (N_18484,N_18219,N_18301);
xor U18485 (N_18485,N_18341,N_18284);
or U18486 (N_18486,N_18225,N_18365);
nand U18487 (N_18487,N_18245,N_18330);
nor U18488 (N_18488,N_18293,N_18228);
and U18489 (N_18489,N_18286,N_18229);
nor U18490 (N_18490,N_18222,N_18305);
nand U18491 (N_18491,N_18232,N_18381);
nand U18492 (N_18492,N_18340,N_18334);
xor U18493 (N_18493,N_18351,N_18321);
xnor U18494 (N_18494,N_18374,N_18303);
nor U18495 (N_18495,N_18325,N_18236);
and U18496 (N_18496,N_18354,N_18394);
nand U18497 (N_18497,N_18300,N_18326);
xnor U18498 (N_18498,N_18369,N_18211);
nand U18499 (N_18499,N_18247,N_18261);
nor U18500 (N_18500,N_18244,N_18383);
nor U18501 (N_18501,N_18325,N_18371);
xnor U18502 (N_18502,N_18372,N_18367);
nand U18503 (N_18503,N_18214,N_18372);
xnor U18504 (N_18504,N_18270,N_18221);
xor U18505 (N_18505,N_18395,N_18256);
nand U18506 (N_18506,N_18378,N_18357);
and U18507 (N_18507,N_18281,N_18283);
and U18508 (N_18508,N_18218,N_18221);
nor U18509 (N_18509,N_18255,N_18239);
and U18510 (N_18510,N_18236,N_18385);
or U18511 (N_18511,N_18399,N_18379);
xnor U18512 (N_18512,N_18306,N_18300);
and U18513 (N_18513,N_18337,N_18395);
nand U18514 (N_18514,N_18247,N_18206);
xor U18515 (N_18515,N_18287,N_18376);
xnor U18516 (N_18516,N_18386,N_18206);
nand U18517 (N_18517,N_18271,N_18370);
nand U18518 (N_18518,N_18215,N_18369);
nand U18519 (N_18519,N_18340,N_18289);
xor U18520 (N_18520,N_18261,N_18348);
or U18521 (N_18521,N_18365,N_18255);
xnor U18522 (N_18522,N_18386,N_18299);
xor U18523 (N_18523,N_18319,N_18231);
nand U18524 (N_18524,N_18347,N_18329);
nand U18525 (N_18525,N_18200,N_18258);
and U18526 (N_18526,N_18343,N_18298);
nand U18527 (N_18527,N_18285,N_18224);
or U18528 (N_18528,N_18285,N_18207);
and U18529 (N_18529,N_18283,N_18227);
xnor U18530 (N_18530,N_18264,N_18265);
xor U18531 (N_18531,N_18311,N_18369);
nand U18532 (N_18532,N_18335,N_18324);
or U18533 (N_18533,N_18223,N_18243);
xor U18534 (N_18534,N_18392,N_18215);
and U18535 (N_18535,N_18230,N_18277);
and U18536 (N_18536,N_18248,N_18256);
xnor U18537 (N_18537,N_18256,N_18226);
nor U18538 (N_18538,N_18222,N_18256);
nand U18539 (N_18539,N_18248,N_18334);
or U18540 (N_18540,N_18247,N_18283);
xnor U18541 (N_18541,N_18296,N_18343);
nor U18542 (N_18542,N_18208,N_18232);
and U18543 (N_18543,N_18304,N_18351);
and U18544 (N_18544,N_18298,N_18360);
nand U18545 (N_18545,N_18258,N_18321);
xor U18546 (N_18546,N_18317,N_18328);
nand U18547 (N_18547,N_18308,N_18227);
xnor U18548 (N_18548,N_18211,N_18206);
nor U18549 (N_18549,N_18202,N_18273);
and U18550 (N_18550,N_18228,N_18277);
nor U18551 (N_18551,N_18394,N_18385);
xor U18552 (N_18552,N_18264,N_18201);
nand U18553 (N_18553,N_18315,N_18280);
nor U18554 (N_18554,N_18206,N_18257);
nor U18555 (N_18555,N_18297,N_18386);
or U18556 (N_18556,N_18316,N_18293);
xor U18557 (N_18557,N_18358,N_18285);
and U18558 (N_18558,N_18266,N_18340);
and U18559 (N_18559,N_18332,N_18323);
xor U18560 (N_18560,N_18227,N_18302);
nand U18561 (N_18561,N_18218,N_18217);
or U18562 (N_18562,N_18349,N_18341);
nor U18563 (N_18563,N_18247,N_18274);
nor U18564 (N_18564,N_18331,N_18317);
xnor U18565 (N_18565,N_18320,N_18264);
nor U18566 (N_18566,N_18354,N_18326);
nor U18567 (N_18567,N_18263,N_18214);
or U18568 (N_18568,N_18393,N_18380);
nand U18569 (N_18569,N_18239,N_18327);
nor U18570 (N_18570,N_18391,N_18339);
nor U18571 (N_18571,N_18319,N_18304);
xor U18572 (N_18572,N_18333,N_18276);
and U18573 (N_18573,N_18275,N_18247);
or U18574 (N_18574,N_18352,N_18381);
xnor U18575 (N_18575,N_18331,N_18348);
nand U18576 (N_18576,N_18292,N_18367);
nor U18577 (N_18577,N_18393,N_18316);
xor U18578 (N_18578,N_18276,N_18368);
xnor U18579 (N_18579,N_18370,N_18231);
nor U18580 (N_18580,N_18356,N_18279);
or U18581 (N_18581,N_18209,N_18237);
xnor U18582 (N_18582,N_18302,N_18351);
or U18583 (N_18583,N_18202,N_18220);
nor U18584 (N_18584,N_18351,N_18336);
nand U18585 (N_18585,N_18238,N_18303);
nand U18586 (N_18586,N_18395,N_18398);
or U18587 (N_18587,N_18290,N_18261);
xor U18588 (N_18588,N_18362,N_18270);
nor U18589 (N_18589,N_18307,N_18304);
nand U18590 (N_18590,N_18374,N_18309);
and U18591 (N_18591,N_18333,N_18273);
and U18592 (N_18592,N_18332,N_18276);
or U18593 (N_18593,N_18316,N_18244);
or U18594 (N_18594,N_18263,N_18211);
and U18595 (N_18595,N_18398,N_18241);
nand U18596 (N_18596,N_18399,N_18340);
nor U18597 (N_18597,N_18344,N_18295);
nor U18598 (N_18598,N_18243,N_18266);
or U18599 (N_18599,N_18345,N_18227);
and U18600 (N_18600,N_18455,N_18436);
nand U18601 (N_18601,N_18437,N_18491);
nor U18602 (N_18602,N_18500,N_18459);
xor U18603 (N_18603,N_18441,N_18496);
and U18604 (N_18604,N_18516,N_18514);
nand U18605 (N_18605,N_18428,N_18470);
xor U18606 (N_18606,N_18530,N_18536);
nor U18607 (N_18607,N_18414,N_18505);
nor U18608 (N_18608,N_18576,N_18597);
xnor U18609 (N_18609,N_18484,N_18445);
nor U18610 (N_18610,N_18583,N_18545);
xnor U18611 (N_18611,N_18430,N_18547);
or U18612 (N_18612,N_18562,N_18497);
and U18613 (N_18613,N_18580,N_18490);
nand U18614 (N_18614,N_18570,N_18543);
nand U18615 (N_18615,N_18418,N_18524);
nor U18616 (N_18616,N_18555,N_18568);
nand U18617 (N_18617,N_18458,N_18498);
or U18618 (N_18618,N_18477,N_18599);
and U18619 (N_18619,N_18573,N_18566);
and U18620 (N_18620,N_18564,N_18529);
nor U18621 (N_18621,N_18577,N_18457);
xnor U18622 (N_18622,N_18433,N_18575);
or U18623 (N_18623,N_18557,N_18535);
or U18624 (N_18624,N_18410,N_18434);
or U18625 (N_18625,N_18501,N_18537);
nand U18626 (N_18626,N_18587,N_18439);
nand U18627 (N_18627,N_18559,N_18469);
xor U18628 (N_18628,N_18413,N_18453);
nand U18629 (N_18629,N_18549,N_18526);
nor U18630 (N_18630,N_18493,N_18572);
xnor U18631 (N_18631,N_18412,N_18542);
xnor U18632 (N_18632,N_18594,N_18423);
or U18633 (N_18633,N_18591,N_18520);
nand U18634 (N_18634,N_18539,N_18478);
nor U18635 (N_18635,N_18528,N_18534);
xnor U18636 (N_18636,N_18421,N_18533);
or U18637 (N_18637,N_18510,N_18476);
xnor U18638 (N_18638,N_18460,N_18485);
nand U18639 (N_18639,N_18585,N_18574);
or U18640 (N_18640,N_18468,N_18554);
and U18641 (N_18641,N_18584,N_18517);
or U18642 (N_18642,N_18451,N_18563);
xor U18643 (N_18643,N_18512,N_18513);
nand U18644 (N_18644,N_18571,N_18425);
nor U18645 (N_18645,N_18400,N_18544);
nand U18646 (N_18646,N_18409,N_18552);
nor U18647 (N_18647,N_18443,N_18569);
xor U18648 (N_18648,N_18595,N_18408);
or U18649 (N_18649,N_18466,N_18593);
nand U18650 (N_18650,N_18567,N_18427);
and U18651 (N_18651,N_18407,N_18411);
nor U18652 (N_18652,N_18452,N_18503);
nor U18653 (N_18653,N_18463,N_18483);
and U18654 (N_18654,N_18507,N_18442);
or U18655 (N_18655,N_18474,N_18426);
or U18656 (N_18656,N_18481,N_18487);
nor U18657 (N_18657,N_18472,N_18588);
xor U18658 (N_18658,N_18590,N_18489);
nand U18659 (N_18659,N_18448,N_18471);
xor U18660 (N_18660,N_18419,N_18581);
or U18661 (N_18661,N_18431,N_18565);
nand U18662 (N_18662,N_18465,N_18582);
or U18663 (N_18663,N_18515,N_18446);
or U18664 (N_18664,N_18589,N_18444);
xor U18665 (N_18665,N_18415,N_18420);
and U18666 (N_18666,N_18461,N_18447);
nor U18667 (N_18667,N_18531,N_18422);
nand U18668 (N_18668,N_18553,N_18416);
nand U18669 (N_18669,N_18479,N_18550);
and U18670 (N_18670,N_18435,N_18521);
and U18671 (N_18671,N_18432,N_18586);
nand U18672 (N_18672,N_18502,N_18538);
nand U18673 (N_18673,N_18551,N_18509);
or U18674 (N_18674,N_18417,N_18405);
xor U18675 (N_18675,N_18525,N_18473);
nor U18676 (N_18676,N_18532,N_18523);
xnor U18677 (N_18677,N_18527,N_18519);
nor U18678 (N_18678,N_18561,N_18401);
nor U18679 (N_18679,N_18438,N_18506);
and U18680 (N_18680,N_18540,N_18504);
nand U18681 (N_18681,N_18546,N_18456);
or U18682 (N_18682,N_18486,N_18450);
nand U18683 (N_18683,N_18548,N_18592);
xnor U18684 (N_18684,N_18522,N_18402);
xor U18685 (N_18685,N_18482,N_18429);
nor U18686 (N_18686,N_18454,N_18560);
nor U18687 (N_18687,N_18541,N_18403);
or U18688 (N_18688,N_18556,N_18492);
nand U18689 (N_18689,N_18467,N_18596);
nand U18690 (N_18690,N_18578,N_18579);
nor U18691 (N_18691,N_18440,N_18424);
or U18692 (N_18692,N_18598,N_18464);
nor U18693 (N_18693,N_18518,N_18495);
or U18694 (N_18694,N_18558,N_18511);
and U18695 (N_18695,N_18480,N_18508);
nand U18696 (N_18696,N_18499,N_18449);
nor U18697 (N_18697,N_18488,N_18462);
nor U18698 (N_18698,N_18406,N_18475);
xor U18699 (N_18699,N_18404,N_18494);
or U18700 (N_18700,N_18456,N_18485);
nand U18701 (N_18701,N_18508,N_18457);
nor U18702 (N_18702,N_18541,N_18498);
and U18703 (N_18703,N_18550,N_18561);
or U18704 (N_18704,N_18558,N_18556);
or U18705 (N_18705,N_18482,N_18462);
or U18706 (N_18706,N_18497,N_18540);
and U18707 (N_18707,N_18427,N_18431);
xnor U18708 (N_18708,N_18496,N_18450);
nor U18709 (N_18709,N_18520,N_18590);
nand U18710 (N_18710,N_18511,N_18424);
and U18711 (N_18711,N_18541,N_18575);
nor U18712 (N_18712,N_18414,N_18532);
or U18713 (N_18713,N_18592,N_18447);
or U18714 (N_18714,N_18469,N_18532);
xor U18715 (N_18715,N_18437,N_18571);
and U18716 (N_18716,N_18590,N_18409);
or U18717 (N_18717,N_18588,N_18547);
and U18718 (N_18718,N_18448,N_18461);
or U18719 (N_18719,N_18548,N_18511);
nand U18720 (N_18720,N_18598,N_18542);
nor U18721 (N_18721,N_18579,N_18561);
or U18722 (N_18722,N_18512,N_18476);
nand U18723 (N_18723,N_18408,N_18431);
and U18724 (N_18724,N_18574,N_18478);
nor U18725 (N_18725,N_18450,N_18519);
or U18726 (N_18726,N_18409,N_18570);
nand U18727 (N_18727,N_18413,N_18449);
or U18728 (N_18728,N_18529,N_18463);
xor U18729 (N_18729,N_18499,N_18550);
or U18730 (N_18730,N_18492,N_18418);
nand U18731 (N_18731,N_18426,N_18506);
xnor U18732 (N_18732,N_18557,N_18538);
nand U18733 (N_18733,N_18418,N_18585);
xor U18734 (N_18734,N_18598,N_18487);
or U18735 (N_18735,N_18479,N_18409);
and U18736 (N_18736,N_18557,N_18476);
xor U18737 (N_18737,N_18404,N_18455);
nor U18738 (N_18738,N_18489,N_18453);
nand U18739 (N_18739,N_18510,N_18567);
nor U18740 (N_18740,N_18483,N_18482);
xnor U18741 (N_18741,N_18417,N_18411);
and U18742 (N_18742,N_18470,N_18498);
xor U18743 (N_18743,N_18531,N_18448);
nand U18744 (N_18744,N_18414,N_18488);
or U18745 (N_18745,N_18421,N_18598);
nand U18746 (N_18746,N_18438,N_18496);
or U18747 (N_18747,N_18579,N_18401);
nand U18748 (N_18748,N_18598,N_18419);
nand U18749 (N_18749,N_18556,N_18482);
xnor U18750 (N_18750,N_18574,N_18533);
or U18751 (N_18751,N_18598,N_18555);
or U18752 (N_18752,N_18500,N_18592);
and U18753 (N_18753,N_18578,N_18550);
and U18754 (N_18754,N_18546,N_18583);
and U18755 (N_18755,N_18423,N_18595);
and U18756 (N_18756,N_18560,N_18407);
xnor U18757 (N_18757,N_18523,N_18472);
xor U18758 (N_18758,N_18506,N_18419);
and U18759 (N_18759,N_18576,N_18535);
and U18760 (N_18760,N_18553,N_18576);
xnor U18761 (N_18761,N_18577,N_18559);
or U18762 (N_18762,N_18465,N_18559);
xnor U18763 (N_18763,N_18423,N_18520);
nor U18764 (N_18764,N_18447,N_18469);
nand U18765 (N_18765,N_18503,N_18569);
nor U18766 (N_18766,N_18435,N_18551);
or U18767 (N_18767,N_18581,N_18428);
xnor U18768 (N_18768,N_18569,N_18555);
nor U18769 (N_18769,N_18552,N_18592);
or U18770 (N_18770,N_18553,N_18572);
and U18771 (N_18771,N_18464,N_18438);
nor U18772 (N_18772,N_18544,N_18579);
nor U18773 (N_18773,N_18407,N_18450);
and U18774 (N_18774,N_18409,N_18507);
nor U18775 (N_18775,N_18401,N_18540);
nand U18776 (N_18776,N_18434,N_18477);
nor U18777 (N_18777,N_18507,N_18462);
nor U18778 (N_18778,N_18515,N_18433);
and U18779 (N_18779,N_18534,N_18425);
or U18780 (N_18780,N_18416,N_18479);
xnor U18781 (N_18781,N_18569,N_18498);
xor U18782 (N_18782,N_18536,N_18529);
nand U18783 (N_18783,N_18466,N_18574);
nand U18784 (N_18784,N_18567,N_18468);
nand U18785 (N_18785,N_18418,N_18446);
xnor U18786 (N_18786,N_18532,N_18425);
nor U18787 (N_18787,N_18527,N_18526);
nand U18788 (N_18788,N_18465,N_18412);
or U18789 (N_18789,N_18415,N_18424);
nand U18790 (N_18790,N_18511,N_18405);
nor U18791 (N_18791,N_18423,N_18458);
and U18792 (N_18792,N_18519,N_18400);
xor U18793 (N_18793,N_18553,N_18491);
xor U18794 (N_18794,N_18471,N_18540);
nand U18795 (N_18795,N_18431,N_18537);
or U18796 (N_18796,N_18546,N_18558);
nand U18797 (N_18797,N_18586,N_18572);
nand U18798 (N_18798,N_18514,N_18508);
and U18799 (N_18799,N_18428,N_18504);
nor U18800 (N_18800,N_18706,N_18755);
nor U18801 (N_18801,N_18635,N_18723);
nand U18802 (N_18802,N_18752,N_18680);
nor U18803 (N_18803,N_18776,N_18783);
xor U18804 (N_18804,N_18756,N_18773);
xor U18805 (N_18805,N_18616,N_18622);
nor U18806 (N_18806,N_18711,N_18623);
or U18807 (N_18807,N_18660,N_18639);
nor U18808 (N_18808,N_18770,N_18748);
nand U18809 (N_18809,N_18712,N_18787);
and U18810 (N_18810,N_18628,N_18619);
nor U18811 (N_18811,N_18797,N_18676);
and U18812 (N_18812,N_18688,N_18689);
nor U18813 (N_18813,N_18761,N_18775);
nor U18814 (N_18814,N_18701,N_18603);
xor U18815 (N_18815,N_18644,N_18699);
xor U18816 (N_18816,N_18789,N_18741);
nand U18817 (N_18817,N_18719,N_18790);
xor U18818 (N_18818,N_18700,N_18665);
and U18819 (N_18819,N_18772,N_18663);
or U18820 (N_18820,N_18664,N_18602);
nand U18821 (N_18821,N_18698,N_18679);
nand U18822 (N_18822,N_18725,N_18740);
nor U18823 (N_18823,N_18788,N_18657);
nand U18824 (N_18824,N_18794,N_18684);
and U18825 (N_18825,N_18738,N_18716);
nor U18826 (N_18826,N_18627,N_18702);
or U18827 (N_18827,N_18781,N_18754);
xnor U18828 (N_18828,N_18746,N_18724);
xor U18829 (N_18829,N_18737,N_18708);
and U18830 (N_18830,N_18734,N_18796);
nor U18831 (N_18831,N_18693,N_18733);
or U18832 (N_18832,N_18624,N_18611);
nor U18833 (N_18833,N_18604,N_18681);
and U18834 (N_18834,N_18631,N_18726);
xor U18835 (N_18835,N_18732,N_18717);
xnor U18836 (N_18836,N_18714,N_18601);
or U18837 (N_18837,N_18784,N_18605);
xor U18838 (N_18838,N_18697,N_18682);
and U18839 (N_18839,N_18728,N_18786);
or U18840 (N_18840,N_18769,N_18764);
nor U18841 (N_18841,N_18718,N_18650);
xor U18842 (N_18842,N_18600,N_18767);
xnor U18843 (N_18843,N_18606,N_18648);
nor U18844 (N_18844,N_18656,N_18675);
or U18845 (N_18845,N_18651,N_18638);
or U18846 (N_18846,N_18791,N_18653);
nor U18847 (N_18847,N_18743,N_18713);
and U18848 (N_18848,N_18694,N_18760);
nand U18849 (N_18849,N_18710,N_18780);
xnor U18850 (N_18850,N_18670,N_18795);
xor U18851 (N_18851,N_18690,N_18612);
xor U18852 (N_18852,N_18739,N_18799);
and U18853 (N_18853,N_18695,N_18729);
nor U18854 (N_18854,N_18641,N_18652);
or U18855 (N_18855,N_18659,N_18685);
xnor U18856 (N_18856,N_18637,N_18722);
and U18857 (N_18857,N_18666,N_18704);
and U18858 (N_18858,N_18610,N_18662);
xnor U18859 (N_18859,N_18766,N_18793);
xnor U18860 (N_18860,N_18674,N_18747);
xnor U18861 (N_18861,N_18765,N_18646);
xor U18862 (N_18862,N_18720,N_18687);
nor U18863 (N_18863,N_18757,N_18762);
and U18864 (N_18864,N_18671,N_18613);
nor U18865 (N_18865,N_18705,N_18751);
or U18866 (N_18866,N_18614,N_18771);
or U18867 (N_18867,N_18615,N_18759);
or U18868 (N_18868,N_18750,N_18655);
xnor U18869 (N_18869,N_18745,N_18792);
xor U18870 (N_18870,N_18620,N_18749);
nand U18871 (N_18871,N_18621,N_18763);
or U18872 (N_18872,N_18617,N_18625);
xnor U18873 (N_18873,N_18645,N_18785);
or U18874 (N_18874,N_18735,N_18721);
nor U18875 (N_18875,N_18633,N_18742);
and U18876 (N_18876,N_18715,N_18683);
and U18877 (N_18877,N_18658,N_18632);
xnor U18878 (N_18878,N_18649,N_18608);
nand U18879 (N_18879,N_18629,N_18609);
and U18880 (N_18880,N_18636,N_18677);
nor U18881 (N_18881,N_18777,N_18707);
nor U18882 (N_18882,N_18630,N_18691);
and U18883 (N_18883,N_18768,N_18774);
xnor U18884 (N_18884,N_18753,N_18642);
nand U18885 (N_18885,N_18703,N_18626);
or U18886 (N_18886,N_18647,N_18730);
nor U18887 (N_18887,N_18778,N_18744);
nand U18888 (N_18888,N_18709,N_18686);
xnor U18889 (N_18889,N_18779,N_18798);
nand U18890 (N_18890,N_18618,N_18668);
nor U18891 (N_18891,N_18640,N_18672);
or U18892 (N_18892,N_18782,N_18736);
nand U18893 (N_18893,N_18661,N_18654);
nand U18894 (N_18894,N_18696,N_18607);
and U18895 (N_18895,N_18634,N_18678);
or U18896 (N_18896,N_18669,N_18692);
and U18897 (N_18897,N_18727,N_18731);
xor U18898 (N_18898,N_18643,N_18667);
nor U18899 (N_18899,N_18673,N_18758);
and U18900 (N_18900,N_18731,N_18711);
nor U18901 (N_18901,N_18641,N_18640);
xor U18902 (N_18902,N_18754,N_18742);
and U18903 (N_18903,N_18651,N_18672);
xnor U18904 (N_18904,N_18644,N_18648);
xor U18905 (N_18905,N_18669,N_18749);
or U18906 (N_18906,N_18623,N_18672);
nor U18907 (N_18907,N_18632,N_18681);
nand U18908 (N_18908,N_18687,N_18641);
and U18909 (N_18909,N_18720,N_18734);
nand U18910 (N_18910,N_18746,N_18603);
or U18911 (N_18911,N_18644,N_18709);
xor U18912 (N_18912,N_18715,N_18720);
nand U18913 (N_18913,N_18634,N_18750);
xor U18914 (N_18914,N_18635,N_18627);
nand U18915 (N_18915,N_18695,N_18765);
and U18916 (N_18916,N_18694,N_18785);
and U18917 (N_18917,N_18659,N_18737);
xor U18918 (N_18918,N_18753,N_18696);
or U18919 (N_18919,N_18726,N_18774);
xor U18920 (N_18920,N_18787,N_18767);
xor U18921 (N_18921,N_18794,N_18704);
xnor U18922 (N_18922,N_18647,N_18699);
or U18923 (N_18923,N_18693,N_18746);
nor U18924 (N_18924,N_18785,N_18708);
nor U18925 (N_18925,N_18783,N_18793);
and U18926 (N_18926,N_18639,N_18771);
xnor U18927 (N_18927,N_18764,N_18733);
xnor U18928 (N_18928,N_18745,N_18687);
xor U18929 (N_18929,N_18770,N_18698);
xnor U18930 (N_18930,N_18684,N_18760);
and U18931 (N_18931,N_18792,N_18726);
nor U18932 (N_18932,N_18633,N_18658);
nand U18933 (N_18933,N_18630,N_18766);
and U18934 (N_18934,N_18679,N_18658);
nand U18935 (N_18935,N_18627,N_18660);
nor U18936 (N_18936,N_18629,N_18666);
and U18937 (N_18937,N_18608,N_18700);
xor U18938 (N_18938,N_18666,N_18773);
and U18939 (N_18939,N_18649,N_18688);
nor U18940 (N_18940,N_18755,N_18601);
nand U18941 (N_18941,N_18794,N_18783);
nand U18942 (N_18942,N_18770,N_18746);
and U18943 (N_18943,N_18723,N_18757);
nor U18944 (N_18944,N_18617,N_18668);
xor U18945 (N_18945,N_18798,N_18725);
xor U18946 (N_18946,N_18641,N_18775);
nand U18947 (N_18947,N_18642,N_18647);
and U18948 (N_18948,N_18779,N_18734);
xor U18949 (N_18949,N_18681,N_18682);
nand U18950 (N_18950,N_18776,N_18702);
xnor U18951 (N_18951,N_18722,N_18621);
or U18952 (N_18952,N_18688,N_18684);
and U18953 (N_18953,N_18741,N_18616);
and U18954 (N_18954,N_18617,N_18719);
nor U18955 (N_18955,N_18636,N_18752);
or U18956 (N_18956,N_18721,N_18712);
or U18957 (N_18957,N_18771,N_18738);
xor U18958 (N_18958,N_18734,N_18667);
and U18959 (N_18959,N_18756,N_18749);
nor U18960 (N_18960,N_18678,N_18630);
xnor U18961 (N_18961,N_18761,N_18624);
or U18962 (N_18962,N_18653,N_18766);
and U18963 (N_18963,N_18664,N_18767);
or U18964 (N_18964,N_18615,N_18738);
or U18965 (N_18965,N_18747,N_18699);
and U18966 (N_18966,N_18723,N_18706);
or U18967 (N_18967,N_18709,N_18758);
and U18968 (N_18968,N_18761,N_18760);
nor U18969 (N_18969,N_18746,N_18656);
nor U18970 (N_18970,N_18779,N_18755);
and U18971 (N_18971,N_18706,N_18607);
or U18972 (N_18972,N_18709,N_18761);
or U18973 (N_18973,N_18618,N_18603);
nor U18974 (N_18974,N_18708,N_18605);
and U18975 (N_18975,N_18747,N_18718);
or U18976 (N_18976,N_18695,N_18721);
and U18977 (N_18977,N_18795,N_18713);
and U18978 (N_18978,N_18789,N_18632);
or U18979 (N_18979,N_18609,N_18736);
nand U18980 (N_18980,N_18779,N_18677);
and U18981 (N_18981,N_18629,N_18783);
and U18982 (N_18982,N_18745,N_18631);
xnor U18983 (N_18983,N_18652,N_18709);
and U18984 (N_18984,N_18651,N_18792);
xnor U18985 (N_18985,N_18669,N_18788);
or U18986 (N_18986,N_18625,N_18740);
and U18987 (N_18987,N_18675,N_18750);
nand U18988 (N_18988,N_18655,N_18788);
and U18989 (N_18989,N_18770,N_18707);
xor U18990 (N_18990,N_18626,N_18697);
xnor U18991 (N_18991,N_18788,N_18674);
xor U18992 (N_18992,N_18690,N_18787);
and U18993 (N_18993,N_18701,N_18691);
xor U18994 (N_18994,N_18673,N_18643);
xnor U18995 (N_18995,N_18617,N_18730);
xnor U18996 (N_18996,N_18661,N_18713);
or U18997 (N_18997,N_18796,N_18676);
and U18998 (N_18998,N_18695,N_18606);
and U18999 (N_18999,N_18787,N_18744);
nor U19000 (N_19000,N_18827,N_18893);
or U19001 (N_19001,N_18917,N_18916);
nand U19002 (N_19002,N_18975,N_18962);
xor U19003 (N_19003,N_18853,N_18802);
and U19004 (N_19004,N_18836,N_18904);
nor U19005 (N_19005,N_18929,N_18877);
or U19006 (N_19006,N_18932,N_18841);
nand U19007 (N_19007,N_18983,N_18808);
nor U19008 (N_19008,N_18870,N_18990);
or U19009 (N_19009,N_18812,N_18866);
and U19010 (N_19010,N_18847,N_18928);
xnor U19011 (N_19011,N_18944,N_18986);
and U19012 (N_19012,N_18833,N_18897);
xnor U19013 (N_19013,N_18997,N_18855);
nor U19014 (N_19014,N_18807,N_18989);
or U19015 (N_19015,N_18822,N_18942);
or U19016 (N_19016,N_18820,N_18839);
nand U19017 (N_19017,N_18919,N_18940);
nor U19018 (N_19018,N_18909,N_18834);
nand U19019 (N_19019,N_18949,N_18843);
or U19020 (N_19020,N_18814,N_18939);
nor U19021 (N_19021,N_18838,N_18850);
or U19022 (N_19022,N_18824,N_18806);
and U19023 (N_19023,N_18885,N_18801);
or U19024 (N_19024,N_18943,N_18846);
and U19025 (N_19025,N_18869,N_18800);
xnor U19026 (N_19026,N_18988,N_18972);
nand U19027 (N_19027,N_18921,N_18970);
and U19028 (N_19028,N_18871,N_18809);
or U19029 (N_19029,N_18813,N_18856);
nand U19030 (N_19030,N_18920,N_18964);
xnor U19031 (N_19031,N_18922,N_18933);
nand U19032 (N_19032,N_18828,N_18858);
nand U19033 (N_19033,N_18954,N_18927);
nor U19034 (N_19034,N_18882,N_18886);
or U19035 (N_19035,N_18965,N_18831);
xor U19036 (N_19036,N_18947,N_18938);
or U19037 (N_19037,N_18840,N_18819);
xor U19038 (N_19038,N_18914,N_18832);
nor U19039 (N_19039,N_18875,N_18905);
xor U19040 (N_19040,N_18851,N_18896);
or U19041 (N_19041,N_18995,N_18883);
xor U19042 (N_19042,N_18823,N_18992);
nor U19043 (N_19043,N_18966,N_18811);
xnor U19044 (N_19044,N_18815,N_18874);
or U19045 (N_19045,N_18898,N_18979);
or U19046 (N_19046,N_18977,N_18956);
xnor U19047 (N_19047,N_18830,N_18907);
nand U19048 (N_19048,N_18901,N_18993);
or U19049 (N_19049,N_18931,N_18980);
or U19050 (N_19050,N_18961,N_18888);
nor U19051 (N_19051,N_18941,N_18890);
nor U19052 (N_19052,N_18984,N_18881);
nor U19053 (N_19053,N_18996,N_18889);
nor U19054 (N_19054,N_18926,N_18878);
or U19055 (N_19055,N_18844,N_18887);
nor U19056 (N_19056,N_18987,N_18911);
xor U19057 (N_19057,N_18842,N_18973);
xnor U19058 (N_19058,N_18835,N_18810);
xnor U19059 (N_19059,N_18976,N_18994);
or U19060 (N_19060,N_18860,N_18952);
or U19061 (N_19061,N_18955,N_18934);
xnor U19062 (N_19062,N_18857,N_18978);
xnor U19063 (N_19063,N_18868,N_18859);
and U19064 (N_19064,N_18872,N_18937);
or U19065 (N_19065,N_18957,N_18968);
nor U19066 (N_19066,N_18879,N_18908);
xor U19067 (N_19067,N_18865,N_18826);
or U19068 (N_19068,N_18991,N_18825);
nand U19069 (N_19069,N_18912,N_18910);
or U19070 (N_19070,N_18948,N_18924);
nor U19071 (N_19071,N_18903,N_18891);
or U19072 (N_19072,N_18817,N_18845);
nand U19073 (N_19073,N_18894,N_18915);
nand U19074 (N_19074,N_18863,N_18818);
nand U19075 (N_19075,N_18960,N_18963);
and U19076 (N_19076,N_18899,N_18852);
or U19077 (N_19077,N_18945,N_18959);
and U19078 (N_19078,N_18950,N_18829);
nand U19079 (N_19079,N_18935,N_18876);
and U19080 (N_19080,N_18864,N_18805);
nand U19081 (N_19081,N_18946,N_18862);
xor U19082 (N_19082,N_18998,N_18985);
nand U19083 (N_19083,N_18923,N_18974);
xnor U19084 (N_19084,N_18913,N_18902);
or U19085 (N_19085,N_18873,N_18804);
xnor U19086 (N_19086,N_18999,N_18981);
xnor U19087 (N_19087,N_18895,N_18953);
nor U19088 (N_19088,N_18854,N_18861);
and U19089 (N_19089,N_18867,N_18918);
nand U19090 (N_19090,N_18892,N_18971);
xor U19091 (N_19091,N_18967,N_18803);
nand U19092 (N_19092,N_18880,N_18925);
nor U19093 (N_19093,N_18982,N_18900);
and U19094 (N_19094,N_18906,N_18849);
and U19095 (N_19095,N_18848,N_18821);
xor U19096 (N_19096,N_18951,N_18958);
and U19097 (N_19097,N_18837,N_18930);
xor U19098 (N_19098,N_18969,N_18816);
and U19099 (N_19099,N_18936,N_18884);
nand U19100 (N_19100,N_18944,N_18871);
nand U19101 (N_19101,N_18881,N_18870);
nor U19102 (N_19102,N_18811,N_18924);
or U19103 (N_19103,N_18970,N_18815);
or U19104 (N_19104,N_18849,N_18830);
xor U19105 (N_19105,N_18954,N_18914);
xnor U19106 (N_19106,N_18964,N_18889);
or U19107 (N_19107,N_18972,N_18982);
or U19108 (N_19108,N_18867,N_18842);
or U19109 (N_19109,N_18880,N_18862);
xor U19110 (N_19110,N_18816,N_18851);
nand U19111 (N_19111,N_18854,N_18883);
or U19112 (N_19112,N_18948,N_18821);
and U19113 (N_19113,N_18817,N_18977);
and U19114 (N_19114,N_18806,N_18948);
xnor U19115 (N_19115,N_18953,N_18856);
and U19116 (N_19116,N_18970,N_18886);
or U19117 (N_19117,N_18860,N_18820);
xor U19118 (N_19118,N_18838,N_18826);
or U19119 (N_19119,N_18883,N_18916);
nand U19120 (N_19120,N_18935,N_18864);
nor U19121 (N_19121,N_18876,N_18895);
xnor U19122 (N_19122,N_18985,N_18921);
and U19123 (N_19123,N_18997,N_18926);
nand U19124 (N_19124,N_18937,N_18920);
and U19125 (N_19125,N_18889,N_18868);
and U19126 (N_19126,N_18875,N_18949);
nand U19127 (N_19127,N_18958,N_18967);
or U19128 (N_19128,N_18838,N_18987);
xor U19129 (N_19129,N_18892,N_18840);
and U19130 (N_19130,N_18864,N_18959);
nor U19131 (N_19131,N_18903,N_18829);
nor U19132 (N_19132,N_18892,N_18985);
nor U19133 (N_19133,N_18830,N_18820);
xnor U19134 (N_19134,N_18998,N_18987);
and U19135 (N_19135,N_18807,N_18866);
and U19136 (N_19136,N_18933,N_18858);
xnor U19137 (N_19137,N_18929,N_18907);
xnor U19138 (N_19138,N_18914,N_18957);
nor U19139 (N_19139,N_18833,N_18892);
xnor U19140 (N_19140,N_18938,N_18859);
nand U19141 (N_19141,N_18922,N_18834);
nor U19142 (N_19142,N_18805,N_18823);
and U19143 (N_19143,N_18868,N_18995);
xnor U19144 (N_19144,N_18949,N_18854);
xnor U19145 (N_19145,N_18803,N_18884);
nand U19146 (N_19146,N_18916,N_18821);
nor U19147 (N_19147,N_18879,N_18900);
xor U19148 (N_19148,N_18903,N_18873);
and U19149 (N_19149,N_18938,N_18925);
xor U19150 (N_19150,N_18867,N_18826);
nor U19151 (N_19151,N_18978,N_18959);
xor U19152 (N_19152,N_18830,N_18840);
xnor U19153 (N_19153,N_18803,N_18838);
or U19154 (N_19154,N_18915,N_18911);
and U19155 (N_19155,N_18868,N_18811);
nor U19156 (N_19156,N_18838,N_18879);
xnor U19157 (N_19157,N_18973,N_18829);
and U19158 (N_19158,N_18926,N_18965);
nand U19159 (N_19159,N_18879,N_18938);
nand U19160 (N_19160,N_18967,N_18941);
and U19161 (N_19161,N_18806,N_18961);
and U19162 (N_19162,N_18820,N_18986);
or U19163 (N_19163,N_18861,N_18868);
xnor U19164 (N_19164,N_18966,N_18823);
nand U19165 (N_19165,N_18934,N_18995);
nor U19166 (N_19166,N_18891,N_18990);
or U19167 (N_19167,N_18979,N_18881);
and U19168 (N_19168,N_18860,N_18897);
nor U19169 (N_19169,N_18859,N_18944);
and U19170 (N_19170,N_18995,N_18938);
nand U19171 (N_19171,N_18992,N_18951);
or U19172 (N_19172,N_18999,N_18808);
nand U19173 (N_19173,N_18968,N_18930);
and U19174 (N_19174,N_18831,N_18816);
xnor U19175 (N_19175,N_18890,N_18971);
nor U19176 (N_19176,N_18998,N_18963);
or U19177 (N_19177,N_18812,N_18901);
xor U19178 (N_19178,N_18802,N_18938);
nor U19179 (N_19179,N_18804,N_18846);
or U19180 (N_19180,N_18893,N_18970);
nand U19181 (N_19181,N_18968,N_18808);
xor U19182 (N_19182,N_18893,N_18824);
or U19183 (N_19183,N_18901,N_18836);
or U19184 (N_19184,N_18892,N_18962);
nand U19185 (N_19185,N_18830,N_18873);
or U19186 (N_19186,N_18869,N_18848);
xnor U19187 (N_19187,N_18949,N_18921);
or U19188 (N_19188,N_18856,N_18952);
nor U19189 (N_19189,N_18974,N_18819);
nand U19190 (N_19190,N_18830,N_18918);
xnor U19191 (N_19191,N_18923,N_18943);
nor U19192 (N_19192,N_18905,N_18854);
nand U19193 (N_19193,N_18920,N_18853);
xor U19194 (N_19194,N_18841,N_18826);
nor U19195 (N_19195,N_18851,N_18960);
xnor U19196 (N_19196,N_18880,N_18854);
xnor U19197 (N_19197,N_18978,N_18896);
and U19198 (N_19198,N_18823,N_18861);
or U19199 (N_19199,N_18951,N_18934);
and U19200 (N_19200,N_19090,N_19045);
and U19201 (N_19201,N_19001,N_19165);
and U19202 (N_19202,N_19124,N_19093);
nand U19203 (N_19203,N_19163,N_19027);
nand U19204 (N_19204,N_19009,N_19138);
xor U19205 (N_19205,N_19117,N_19031);
xor U19206 (N_19206,N_19129,N_19144);
or U19207 (N_19207,N_19136,N_19169);
nor U19208 (N_19208,N_19061,N_19025);
nand U19209 (N_19209,N_19185,N_19076);
nand U19210 (N_19210,N_19033,N_19088);
and U19211 (N_19211,N_19021,N_19114);
and U19212 (N_19212,N_19150,N_19170);
nor U19213 (N_19213,N_19049,N_19123);
and U19214 (N_19214,N_19018,N_19168);
nand U19215 (N_19215,N_19055,N_19089);
or U19216 (N_19216,N_19157,N_19000);
nor U19217 (N_19217,N_19137,N_19042);
and U19218 (N_19218,N_19108,N_19142);
or U19219 (N_19219,N_19162,N_19012);
nand U19220 (N_19220,N_19176,N_19057);
and U19221 (N_19221,N_19128,N_19171);
nor U19222 (N_19222,N_19017,N_19040);
xnor U19223 (N_19223,N_19193,N_19192);
or U19224 (N_19224,N_19036,N_19102);
and U19225 (N_19225,N_19107,N_19004);
or U19226 (N_19226,N_19167,N_19091);
nand U19227 (N_19227,N_19056,N_19007);
nor U19228 (N_19228,N_19189,N_19106);
and U19229 (N_19229,N_19188,N_19131);
nand U19230 (N_19230,N_19191,N_19084);
or U19231 (N_19231,N_19141,N_19153);
and U19232 (N_19232,N_19104,N_19121);
and U19233 (N_19233,N_19183,N_19134);
xnor U19234 (N_19234,N_19066,N_19068);
nor U19235 (N_19235,N_19197,N_19070);
and U19236 (N_19236,N_19135,N_19120);
and U19237 (N_19237,N_19078,N_19133);
nor U19238 (N_19238,N_19010,N_19022);
nand U19239 (N_19239,N_19080,N_19140);
nand U19240 (N_19240,N_19092,N_19047);
nor U19241 (N_19241,N_19072,N_19014);
nand U19242 (N_19242,N_19172,N_19083);
and U19243 (N_19243,N_19166,N_19094);
or U19244 (N_19244,N_19041,N_19154);
and U19245 (N_19245,N_19156,N_19116);
and U19246 (N_19246,N_19071,N_19062);
and U19247 (N_19247,N_19064,N_19160);
xnor U19248 (N_19248,N_19179,N_19074);
xor U19249 (N_19249,N_19186,N_19178);
nor U19250 (N_19250,N_19173,N_19177);
nand U19251 (N_19251,N_19051,N_19037);
or U19252 (N_19252,N_19130,N_19020);
nor U19253 (N_19253,N_19038,N_19075);
and U19254 (N_19254,N_19198,N_19109);
nor U19255 (N_19255,N_19005,N_19028);
and U19256 (N_19256,N_19187,N_19035);
nand U19257 (N_19257,N_19048,N_19063);
nor U19258 (N_19258,N_19043,N_19081);
nor U19259 (N_19259,N_19147,N_19182);
nor U19260 (N_19260,N_19019,N_19161);
xor U19261 (N_19261,N_19155,N_19006);
and U19262 (N_19262,N_19113,N_19032);
xnor U19263 (N_19263,N_19024,N_19199);
nor U19264 (N_19264,N_19099,N_19065);
nand U19265 (N_19265,N_19053,N_19026);
nor U19266 (N_19266,N_19127,N_19149);
nand U19267 (N_19267,N_19175,N_19077);
nor U19268 (N_19268,N_19023,N_19180);
and U19269 (N_19269,N_19122,N_19111);
and U19270 (N_19270,N_19054,N_19101);
nor U19271 (N_19271,N_19146,N_19164);
and U19272 (N_19272,N_19112,N_19139);
and U19273 (N_19273,N_19100,N_19098);
xor U19274 (N_19274,N_19097,N_19152);
nand U19275 (N_19275,N_19159,N_19044);
and U19276 (N_19276,N_19195,N_19050);
nand U19277 (N_19277,N_19151,N_19119);
nor U19278 (N_19278,N_19190,N_19016);
and U19279 (N_19279,N_19034,N_19067);
or U19280 (N_19280,N_19011,N_19030);
xnor U19281 (N_19281,N_19059,N_19015);
nor U19282 (N_19282,N_19052,N_19110);
nor U19283 (N_19283,N_19096,N_19039);
nand U19284 (N_19284,N_19181,N_19115);
and U19285 (N_19285,N_19125,N_19082);
nor U19286 (N_19286,N_19148,N_19085);
or U19287 (N_19287,N_19105,N_19087);
nor U19288 (N_19288,N_19143,N_19196);
and U19289 (N_19289,N_19060,N_19145);
or U19290 (N_19290,N_19003,N_19079);
nor U19291 (N_19291,N_19095,N_19132);
nand U19292 (N_19292,N_19069,N_19029);
nor U19293 (N_19293,N_19103,N_19073);
xnor U19294 (N_19294,N_19184,N_19158);
and U19295 (N_19295,N_19194,N_19086);
nand U19296 (N_19296,N_19118,N_19008);
nand U19297 (N_19297,N_19126,N_19013);
xor U19298 (N_19298,N_19046,N_19174);
nor U19299 (N_19299,N_19058,N_19002);
nand U19300 (N_19300,N_19153,N_19005);
nand U19301 (N_19301,N_19130,N_19059);
or U19302 (N_19302,N_19054,N_19123);
xor U19303 (N_19303,N_19113,N_19110);
nand U19304 (N_19304,N_19151,N_19074);
nor U19305 (N_19305,N_19130,N_19004);
and U19306 (N_19306,N_19161,N_19188);
nor U19307 (N_19307,N_19053,N_19054);
xor U19308 (N_19308,N_19182,N_19114);
or U19309 (N_19309,N_19084,N_19067);
nand U19310 (N_19310,N_19135,N_19055);
nand U19311 (N_19311,N_19063,N_19150);
and U19312 (N_19312,N_19081,N_19083);
nor U19313 (N_19313,N_19162,N_19132);
and U19314 (N_19314,N_19025,N_19072);
or U19315 (N_19315,N_19010,N_19177);
or U19316 (N_19316,N_19196,N_19188);
nand U19317 (N_19317,N_19005,N_19073);
xnor U19318 (N_19318,N_19001,N_19011);
nor U19319 (N_19319,N_19037,N_19098);
and U19320 (N_19320,N_19145,N_19077);
or U19321 (N_19321,N_19170,N_19039);
nor U19322 (N_19322,N_19184,N_19075);
nor U19323 (N_19323,N_19189,N_19007);
or U19324 (N_19324,N_19026,N_19067);
or U19325 (N_19325,N_19069,N_19166);
nand U19326 (N_19326,N_19111,N_19002);
and U19327 (N_19327,N_19132,N_19182);
xnor U19328 (N_19328,N_19057,N_19104);
or U19329 (N_19329,N_19122,N_19104);
or U19330 (N_19330,N_19037,N_19039);
and U19331 (N_19331,N_19086,N_19014);
nor U19332 (N_19332,N_19095,N_19092);
nand U19333 (N_19333,N_19072,N_19185);
nand U19334 (N_19334,N_19067,N_19188);
xnor U19335 (N_19335,N_19040,N_19030);
or U19336 (N_19336,N_19126,N_19019);
and U19337 (N_19337,N_19077,N_19162);
nand U19338 (N_19338,N_19037,N_19192);
nand U19339 (N_19339,N_19185,N_19054);
nor U19340 (N_19340,N_19077,N_19144);
nand U19341 (N_19341,N_19192,N_19149);
or U19342 (N_19342,N_19196,N_19061);
nand U19343 (N_19343,N_19105,N_19092);
nand U19344 (N_19344,N_19057,N_19005);
nor U19345 (N_19345,N_19174,N_19005);
nor U19346 (N_19346,N_19018,N_19097);
nand U19347 (N_19347,N_19110,N_19039);
nor U19348 (N_19348,N_19077,N_19178);
or U19349 (N_19349,N_19180,N_19007);
xor U19350 (N_19350,N_19195,N_19051);
nor U19351 (N_19351,N_19184,N_19027);
or U19352 (N_19352,N_19122,N_19139);
nand U19353 (N_19353,N_19008,N_19075);
or U19354 (N_19354,N_19160,N_19104);
nor U19355 (N_19355,N_19044,N_19015);
xnor U19356 (N_19356,N_19014,N_19132);
and U19357 (N_19357,N_19087,N_19030);
xnor U19358 (N_19358,N_19189,N_19178);
xnor U19359 (N_19359,N_19051,N_19149);
and U19360 (N_19360,N_19013,N_19018);
xor U19361 (N_19361,N_19140,N_19018);
xor U19362 (N_19362,N_19168,N_19083);
nand U19363 (N_19363,N_19000,N_19054);
nand U19364 (N_19364,N_19173,N_19064);
or U19365 (N_19365,N_19090,N_19110);
xor U19366 (N_19366,N_19111,N_19141);
nand U19367 (N_19367,N_19089,N_19149);
nor U19368 (N_19368,N_19198,N_19192);
nor U19369 (N_19369,N_19059,N_19166);
or U19370 (N_19370,N_19184,N_19090);
nand U19371 (N_19371,N_19060,N_19024);
nand U19372 (N_19372,N_19136,N_19182);
nand U19373 (N_19373,N_19076,N_19115);
and U19374 (N_19374,N_19174,N_19045);
xor U19375 (N_19375,N_19057,N_19105);
xor U19376 (N_19376,N_19122,N_19006);
nor U19377 (N_19377,N_19163,N_19089);
or U19378 (N_19378,N_19170,N_19080);
nand U19379 (N_19379,N_19181,N_19119);
and U19380 (N_19380,N_19096,N_19189);
nor U19381 (N_19381,N_19166,N_19068);
or U19382 (N_19382,N_19029,N_19048);
nand U19383 (N_19383,N_19099,N_19044);
xor U19384 (N_19384,N_19086,N_19090);
and U19385 (N_19385,N_19008,N_19029);
xor U19386 (N_19386,N_19193,N_19181);
and U19387 (N_19387,N_19076,N_19083);
nand U19388 (N_19388,N_19160,N_19114);
xor U19389 (N_19389,N_19078,N_19173);
nor U19390 (N_19390,N_19016,N_19025);
and U19391 (N_19391,N_19139,N_19117);
nor U19392 (N_19392,N_19178,N_19174);
or U19393 (N_19393,N_19158,N_19090);
nor U19394 (N_19394,N_19153,N_19199);
and U19395 (N_19395,N_19153,N_19064);
nor U19396 (N_19396,N_19104,N_19124);
and U19397 (N_19397,N_19063,N_19034);
or U19398 (N_19398,N_19125,N_19049);
nor U19399 (N_19399,N_19008,N_19049);
or U19400 (N_19400,N_19200,N_19393);
nand U19401 (N_19401,N_19339,N_19267);
xnor U19402 (N_19402,N_19234,N_19381);
or U19403 (N_19403,N_19336,N_19372);
and U19404 (N_19404,N_19209,N_19320);
nand U19405 (N_19405,N_19213,N_19259);
nor U19406 (N_19406,N_19374,N_19379);
nand U19407 (N_19407,N_19331,N_19313);
and U19408 (N_19408,N_19324,N_19323);
nand U19409 (N_19409,N_19342,N_19235);
nor U19410 (N_19410,N_19295,N_19380);
nor U19411 (N_19411,N_19354,N_19304);
xor U19412 (N_19412,N_19226,N_19206);
nand U19413 (N_19413,N_19303,N_19375);
nand U19414 (N_19414,N_19264,N_19256);
and U19415 (N_19415,N_19254,N_19387);
xnor U19416 (N_19416,N_19329,N_19395);
or U19417 (N_19417,N_19203,N_19325);
nor U19418 (N_19418,N_19279,N_19385);
xnor U19419 (N_19419,N_19348,N_19371);
xor U19420 (N_19420,N_19352,N_19221);
and U19421 (N_19421,N_19308,N_19302);
or U19422 (N_19422,N_19390,N_19220);
nand U19423 (N_19423,N_19370,N_19208);
nand U19424 (N_19424,N_19300,N_19346);
and U19425 (N_19425,N_19391,N_19283);
or U19426 (N_19426,N_19305,N_19261);
or U19427 (N_19427,N_19253,N_19289);
xnor U19428 (N_19428,N_19369,N_19260);
nor U19429 (N_19429,N_19232,N_19246);
or U19430 (N_19430,N_19337,N_19312);
nor U19431 (N_19431,N_19201,N_19398);
xor U19432 (N_19432,N_19298,N_19263);
nand U19433 (N_19433,N_19317,N_19316);
or U19434 (N_19434,N_19204,N_19228);
xnor U19435 (N_19435,N_19286,N_19241);
nor U19436 (N_19436,N_19248,N_19242);
xor U19437 (N_19437,N_19255,N_19243);
nor U19438 (N_19438,N_19297,N_19335);
nand U19439 (N_19439,N_19276,N_19377);
nor U19440 (N_19440,N_19363,N_19344);
and U19441 (N_19441,N_19230,N_19207);
or U19442 (N_19442,N_19211,N_19338);
xnor U19443 (N_19443,N_19284,N_19394);
nand U19444 (N_19444,N_19347,N_19291);
nand U19445 (N_19445,N_19265,N_19247);
nor U19446 (N_19446,N_19361,N_19233);
xnor U19447 (N_19447,N_19245,N_19386);
nor U19448 (N_19448,N_19288,N_19210);
nand U19449 (N_19449,N_19307,N_19268);
or U19450 (N_19450,N_19294,N_19357);
or U19451 (N_19451,N_19343,N_19321);
nand U19452 (N_19452,N_19349,N_19319);
xor U19453 (N_19453,N_19306,N_19314);
and U19454 (N_19454,N_19383,N_19388);
and U19455 (N_19455,N_19292,N_19310);
xnor U19456 (N_19456,N_19236,N_19212);
or U19457 (N_19457,N_19205,N_19353);
and U19458 (N_19458,N_19285,N_19287);
and U19459 (N_19459,N_19382,N_19275);
or U19460 (N_19460,N_19277,N_19373);
or U19461 (N_19461,N_19219,N_19367);
nor U19462 (N_19462,N_19223,N_19332);
and U19463 (N_19463,N_19214,N_19315);
xor U19464 (N_19464,N_19397,N_19216);
nor U19465 (N_19465,N_19280,N_19266);
xnor U19466 (N_19466,N_19322,N_19333);
nand U19467 (N_19467,N_19282,N_19202);
nor U19468 (N_19468,N_19258,N_19318);
xnor U19469 (N_19469,N_19237,N_19365);
nand U19470 (N_19470,N_19376,N_19334);
xnor U19471 (N_19471,N_19309,N_19328);
nor U19472 (N_19472,N_19271,N_19351);
nand U19473 (N_19473,N_19366,N_19355);
or U19474 (N_19474,N_19360,N_19399);
and U19475 (N_19475,N_19274,N_19356);
nand U19476 (N_19476,N_19217,N_19227);
nor U19477 (N_19477,N_19341,N_19240);
nor U19478 (N_19478,N_19362,N_19340);
and U19479 (N_19479,N_19225,N_19272);
xor U19480 (N_19480,N_19224,N_19311);
nor U19481 (N_19481,N_19299,N_19270);
and U19482 (N_19482,N_19273,N_19364);
or U19483 (N_19483,N_19350,N_19238);
and U19484 (N_19484,N_19296,N_19293);
or U19485 (N_19485,N_19231,N_19229);
xor U19486 (N_19486,N_19359,N_19345);
nor U19487 (N_19487,N_19326,N_19251);
and U19488 (N_19488,N_19396,N_19215);
nor U19489 (N_19489,N_19368,N_19384);
xor U19490 (N_19490,N_19269,N_19330);
and U19491 (N_19491,N_19257,N_19249);
or U19492 (N_19492,N_19278,N_19301);
or U19493 (N_19493,N_19358,N_19392);
nand U19494 (N_19494,N_19239,N_19222);
nand U19495 (N_19495,N_19327,N_19262);
nor U19496 (N_19496,N_19389,N_19252);
xnor U19497 (N_19497,N_19290,N_19218);
or U19498 (N_19498,N_19250,N_19378);
and U19499 (N_19499,N_19281,N_19244);
nand U19500 (N_19500,N_19293,N_19345);
xor U19501 (N_19501,N_19298,N_19273);
xnor U19502 (N_19502,N_19273,N_19368);
or U19503 (N_19503,N_19376,N_19368);
xnor U19504 (N_19504,N_19231,N_19304);
xnor U19505 (N_19505,N_19322,N_19334);
and U19506 (N_19506,N_19294,N_19281);
or U19507 (N_19507,N_19285,N_19280);
or U19508 (N_19508,N_19303,N_19365);
and U19509 (N_19509,N_19319,N_19317);
and U19510 (N_19510,N_19370,N_19250);
nand U19511 (N_19511,N_19362,N_19269);
nand U19512 (N_19512,N_19302,N_19212);
and U19513 (N_19513,N_19378,N_19286);
xnor U19514 (N_19514,N_19389,N_19233);
or U19515 (N_19515,N_19227,N_19390);
xor U19516 (N_19516,N_19379,N_19325);
nand U19517 (N_19517,N_19251,N_19387);
nor U19518 (N_19518,N_19298,N_19236);
nand U19519 (N_19519,N_19388,N_19291);
nand U19520 (N_19520,N_19366,N_19207);
xnor U19521 (N_19521,N_19264,N_19239);
or U19522 (N_19522,N_19291,N_19267);
and U19523 (N_19523,N_19260,N_19222);
and U19524 (N_19524,N_19313,N_19297);
nor U19525 (N_19525,N_19310,N_19356);
nor U19526 (N_19526,N_19385,N_19345);
nand U19527 (N_19527,N_19300,N_19292);
xnor U19528 (N_19528,N_19351,N_19342);
nor U19529 (N_19529,N_19388,N_19299);
nand U19530 (N_19530,N_19263,N_19243);
and U19531 (N_19531,N_19280,N_19225);
and U19532 (N_19532,N_19249,N_19228);
and U19533 (N_19533,N_19379,N_19252);
or U19534 (N_19534,N_19280,N_19307);
xor U19535 (N_19535,N_19395,N_19251);
nand U19536 (N_19536,N_19246,N_19361);
nand U19537 (N_19537,N_19399,N_19283);
xor U19538 (N_19538,N_19313,N_19252);
and U19539 (N_19539,N_19315,N_19376);
nor U19540 (N_19540,N_19381,N_19311);
nand U19541 (N_19541,N_19330,N_19321);
nand U19542 (N_19542,N_19279,N_19346);
xor U19543 (N_19543,N_19327,N_19235);
xor U19544 (N_19544,N_19313,N_19236);
nor U19545 (N_19545,N_19267,N_19302);
nor U19546 (N_19546,N_19291,N_19264);
and U19547 (N_19547,N_19364,N_19217);
and U19548 (N_19548,N_19247,N_19373);
xnor U19549 (N_19549,N_19315,N_19330);
and U19550 (N_19550,N_19251,N_19206);
or U19551 (N_19551,N_19225,N_19204);
xor U19552 (N_19552,N_19367,N_19321);
nand U19553 (N_19553,N_19296,N_19257);
xor U19554 (N_19554,N_19224,N_19291);
xnor U19555 (N_19555,N_19304,N_19242);
nor U19556 (N_19556,N_19272,N_19333);
or U19557 (N_19557,N_19284,N_19325);
xnor U19558 (N_19558,N_19265,N_19206);
xor U19559 (N_19559,N_19235,N_19344);
xor U19560 (N_19560,N_19279,N_19256);
xor U19561 (N_19561,N_19286,N_19302);
nor U19562 (N_19562,N_19373,N_19275);
nand U19563 (N_19563,N_19364,N_19234);
xor U19564 (N_19564,N_19200,N_19299);
and U19565 (N_19565,N_19288,N_19375);
nor U19566 (N_19566,N_19325,N_19257);
and U19567 (N_19567,N_19237,N_19260);
xnor U19568 (N_19568,N_19246,N_19340);
xor U19569 (N_19569,N_19264,N_19377);
and U19570 (N_19570,N_19342,N_19316);
nand U19571 (N_19571,N_19203,N_19396);
and U19572 (N_19572,N_19315,N_19237);
or U19573 (N_19573,N_19311,N_19376);
or U19574 (N_19574,N_19392,N_19246);
xor U19575 (N_19575,N_19285,N_19330);
nand U19576 (N_19576,N_19312,N_19345);
nor U19577 (N_19577,N_19227,N_19275);
and U19578 (N_19578,N_19208,N_19387);
or U19579 (N_19579,N_19394,N_19324);
and U19580 (N_19580,N_19291,N_19274);
or U19581 (N_19581,N_19363,N_19397);
nand U19582 (N_19582,N_19245,N_19226);
xnor U19583 (N_19583,N_19253,N_19206);
or U19584 (N_19584,N_19365,N_19203);
nor U19585 (N_19585,N_19279,N_19392);
xor U19586 (N_19586,N_19287,N_19276);
and U19587 (N_19587,N_19356,N_19397);
nor U19588 (N_19588,N_19212,N_19260);
nand U19589 (N_19589,N_19342,N_19345);
and U19590 (N_19590,N_19316,N_19399);
nand U19591 (N_19591,N_19348,N_19384);
and U19592 (N_19592,N_19347,N_19219);
nor U19593 (N_19593,N_19227,N_19239);
xor U19594 (N_19594,N_19277,N_19266);
nor U19595 (N_19595,N_19219,N_19205);
nand U19596 (N_19596,N_19293,N_19332);
nand U19597 (N_19597,N_19280,N_19305);
nor U19598 (N_19598,N_19314,N_19254);
and U19599 (N_19599,N_19359,N_19364);
and U19600 (N_19600,N_19558,N_19508);
xor U19601 (N_19601,N_19505,N_19471);
nor U19602 (N_19602,N_19551,N_19559);
or U19603 (N_19603,N_19585,N_19448);
and U19604 (N_19604,N_19475,N_19495);
nand U19605 (N_19605,N_19434,N_19501);
and U19606 (N_19606,N_19599,N_19492);
nor U19607 (N_19607,N_19439,N_19576);
nand U19608 (N_19608,N_19509,N_19442);
xor U19609 (N_19609,N_19420,N_19416);
nand U19610 (N_19610,N_19528,N_19529);
nor U19611 (N_19611,N_19406,N_19484);
xor U19612 (N_19612,N_19487,N_19482);
nand U19613 (N_19613,N_19541,N_19536);
nor U19614 (N_19614,N_19497,N_19400);
nand U19615 (N_19615,N_19423,N_19565);
or U19616 (N_19616,N_19527,N_19514);
xor U19617 (N_19617,N_19555,N_19411);
nand U19618 (N_19618,N_19440,N_19449);
nor U19619 (N_19619,N_19445,N_19459);
and U19620 (N_19620,N_19464,N_19597);
and U19621 (N_19621,N_19590,N_19403);
nor U19622 (N_19622,N_19598,N_19472);
and U19623 (N_19623,N_19593,N_19488);
xnor U19624 (N_19624,N_19455,N_19537);
or U19625 (N_19625,N_19572,N_19580);
nor U19626 (N_19626,N_19534,N_19494);
nor U19627 (N_19627,N_19467,N_19575);
xnor U19628 (N_19628,N_19550,N_19520);
and U19629 (N_19629,N_19502,N_19507);
or U19630 (N_19630,N_19409,N_19594);
and U19631 (N_19631,N_19561,N_19511);
xnor U19632 (N_19632,N_19436,N_19513);
xnor U19633 (N_19633,N_19539,N_19584);
nor U19634 (N_19634,N_19531,N_19457);
nor U19635 (N_19635,N_19540,N_19415);
xnor U19636 (N_19636,N_19557,N_19503);
nor U19637 (N_19637,N_19438,N_19563);
nor U19638 (N_19638,N_19535,N_19553);
or U19639 (N_19639,N_19533,N_19504);
nor U19640 (N_19640,N_19428,N_19463);
or U19641 (N_19641,N_19564,N_19583);
or U19642 (N_19642,N_19491,N_19510);
xnor U19643 (N_19643,N_19515,N_19465);
xor U19644 (N_19644,N_19573,N_19521);
nor U19645 (N_19645,N_19567,N_19595);
xnor U19646 (N_19646,N_19589,N_19413);
and U19647 (N_19647,N_19452,N_19523);
nand U19648 (N_19648,N_19519,N_19405);
nand U19649 (N_19649,N_19419,N_19468);
and U19650 (N_19650,N_19592,N_19454);
nand U19651 (N_19651,N_19493,N_19404);
or U19652 (N_19652,N_19429,N_19532);
nor U19653 (N_19653,N_19435,N_19432);
or U19654 (N_19654,N_19518,N_19500);
or U19655 (N_19655,N_19461,N_19478);
xnor U19656 (N_19656,N_19560,N_19483);
and U19657 (N_19657,N_19542,N_19570);
xor U19658 (N_19658,N_19548,N_19525);
and U19659 (N_19659,N_19506,N_19596);
or U19660 (N_19660,N_19407,N_19422);
nand U19661 (N_19661,N_19552,N_19496);
and U19662 (N_19662,N_19578,N_19517);
or U19663 (N_19663,N_19410,N_19480);
or U19664 (N_19664,N_19425,N_19401);
nand U19665 (N_19665,N_19421,N_19545);
nand U19666 (N_19666,N_19562,N_19577);
nor U19667 (N_19667,N_19469,N_19499);
xor U19668 (N_19668,N_19568,N_19418);
or U19669 (N_19669,N_19498,N_19476);
nand U19670 (N_19670,N_19473,N_19489);
nor U19671 (N_19671,N_19433,N_19543);
or U19672 (N_19672,N_19554,N_19443);
nor U19673 (N_19673,N_19426,N_19530);
xor U19674 (N_19674,N_19450,N_19587);
xnor U19675 (N_19675,N_19477,N_19571);
nand U19676 (N_19676,N_19586,N_19446);
or U19677 (N_19677,N_19430,N_19566);
nor U19678 (N_19678,N_19481,N_19444);
or U19679 (N_19679,N_19547,N_19417);
xnor U19680 (N_19680,N_19574,N_19462);
and U19681 (N_19681,N_19524,N_19538);
xnor U19682 (N_19682,N_19470,N_19437);
or U19683 (N_19683,N_19427,N_19588);
nand U19684 (N_19684,N_19544,N_19581);
nor U19685 (N_19685,N_19451,N_19441);
nand U19686 (N_19686,N_19486,N_19431);
nor U19687 (N_19687,N_19474,N_19582);
xnor U19688 (N_19688,N_19569,N_19424);
xnor U19689 (N_19689,N_19556,N_19412);
and U19690 (N_19690,N_19458,N_19549);
nor U19691 (N_19691,N_19460,N_19479);
or U19692 (N_19692,N_19490,N_19453);
and U19693 (N_19693,N_19516,N_19414);
or U19694 (N_19694,N_19579,N_19526);
and U19695 (N_19695,N_19456,N_19402);
nand U19696 (N_19696,N_19485,N_19512);
nor U19697 (N_19697,N_19466,N_19522);
or U19698 (N_19698,N_19447,N_19408);
nor U19699 (N_19699,N_19591,N_19546);
nor U19700 (N_19700,N_19535,N_19454);
or U19701 (N_19701,N_19596,N_19488);
or U19702 (N_19702,N_19477,N_19476);
xnor U19703 (N_19703,N_19547,N_19563);
and U19704 (N_19704,N_19512,N_19453);
or U19705 (N_19705,N_19485,N_19523);
nor U19706 (N_19706,N_19528,N_19421);
xor U19707 (N_19707,N_19556,N_19453);
and U19708 (N_19708,N_19412,N_19427);
nand U19709 (N_19709,N_19597,N_19567);
xor U19710 (N_19710,N_19461,N_19423);
nand U19711 (N_19711,N_19423,N_19513);
nor U19712 (N_19712,N_19402,N_19455);
or U19713 (N_19713,N_19400,N_19590);
xnor U19714 (N_19714,N_19573,N_19563);
xnor U19715 (N_19715,N_19478,N_19445);
nor U19716 (N_19716,N_19538,N_19493);
nor U19717 (N_19717,N_19483,N_19501);
and U19718 (N_19718,N_19594,N_19566);
and U19719 (N_19719,N_19415,N_19499);
or U19720 (N_19720,N_19581,N_19417);
and U19721 (N_19721,N_19585,N_19465);
and U19722 (N_19722,N_19558,N_19571);
xor U19723 (N_19723,N_19536,N_19533);
nand U19724 (N_19724,N_19583,N_19412);
nor U19725 (N_19725,N_19475,N_19576);
xor U19726 (N_19726,N_19437,N_19408);
and U19727 (N_19727,N_19524,N_19497);
xnor U19728 (N_19728,N_19422,N_19513);
xnor U19729 (N_19729,N_19558,N_19433);
and U19730 (N_19730,N_19484,N_19555);
nand U19731 (N_19731,N_19425,N_19486);
xor U19732 (N_19732,N_19454,N_19489);
nor U19733 (N_19733,N_19521,N_19584);
and U19734 (N_19734,N_19551,N_19525);
and U19735 (N_19735,N_19466,N_19569);
nand U19736 (N_19736,N_19453,N_19440);
or U19737 (N_19737,N_19495,N_19589);
nor U19738 (N_19738,N_19455,N_19480);
or U19739 (N_19739,N_19590,N_19485);
nand U19740 (N_19740,N_19450,N_19584);
nor U19741 (N_19741,N_19443,N_19470);
and U19742 (N_19742,N_19505,N_19426);
nor U19743 (N_19743,N_19449,N_19419);
xor U19744 (N_19744,N_19434,N_19552);
nand U19745 (N_19745,N_19524,N_19443);
and U19746 (N_19746,N_19411,N_19595);
nand U19747 (N_19747,N_19473,N_19478);
nor U19748 (N_19748,N_19413,N_19542);
and U19749 (N_19749,N_19444,N_19437);
nor U19750 (N_19750,N_19572,N_19561);
and U19751 (N_19751,N_19408,N_19464);
nor U19752 (N_19752,N_19536,N_19401);
xnor U19753 (N_19753,N_19434,N_19448);
nand U19754 (N_19754,N_19413,N_19547);
or U19755 (N_19755,N_19474,N_19571);
or U19756 (N_19756,N_19586,N_19444);
xnor U19757 (N_19757,N_19484,N_19541);
nand U19758 (N_19758,N_19591,N_19561);
xor U19759 (N_19759,N_19405,N_19442);
nor U19760 (N_19760,N_19414,N_19568);
nor U19761 (N_19761,N_19522,N_19505);
or U19762 (N_19762,N_19545,N_19588);
or U19763 (N_19763,N_19471,N_19426);
nand U19764 (N_19764,N_19538,N_19502);
and U19765 (N_19765,N_19549,N_19559);
nand U19766 (N_19766,N_19578,N_19407);
xnor U19767 (N_19767,N_19426,N_19554);
or U19768 (N_19768,N_19482,N_19451);
or U19769 (N_19769,N_19406,N_19555);
or U19770 (N_19770,N_19576,N_19543);
or U19771 (N_19771,N_19458,N_19431);
nor U19772 (N_19772,N_19474,N_19518);
and U19773 (N_19773,N_19484,N_19566);
nand U19774 (N_19774,N_19463,N_19545);
xnor U19775 (N_19775,N_19401,N_19414);
nand U19776 (N_19776,N_19544,N_19597);
or U19777 (N_19777,N_19439,N_19456);
and U19778 (N_19778,N_19435,N_19525);
nand U19779 (N_19779,N_19530,N_19457);
xor U19780 (N_19780,N_19523,N_19512);
xor U19781 (N_19781,N_19496,N_19486);
nor U19782 (N_19782,N_19590,N_19464);
nor U19783 (N_19783,N_19594,N_19553);
nor U19784 (N_19784,N_19514,N_19582);
or U19785 (N_19785,N_19478,N_19582);
xor U19786 (N_19786,N_19437,N_19472);
or U19787 (N_19787,N_19406,N_19454);
xnor U19788 (N_19788,N_19467,N_19447);
nor U19789 (N_19789,N_19560,N_19430);
xor U19790 (N_19790,N_19574,N_19561);
or U19791 (N_19791,N_19402,N_19488);
or U19792 (N_19792,N_19520,N_19523);
and U19793 (N_19793,N_19560,N_19407);
xor U19794 (N_19794,N_19413,N_19405);
nor U19795 (N_19795,N_19410,N_19586);
nand U19796 (N_19796,N_19541,N_19456);
nor U19797 (N_19797,N_19465,N_19448);
and U19798 (N_19798,N_19568,N_19500);
and U19799 (N_19799,N_19453,N_19533);
or U19800 (N_19800,N_19682,N_19772);
xnor U19801 (N_19801,N_19604,N_19771);
and U19802 (N_19802,N_19657,N_19736);
xor U19803 (N_19803,N_19670,N_19701);
or U19804 (N_19804,N_19714,N_19763);
nand U19805 (N_19805,N_19602,N_19645);
nand U19806 (N_19806,N_19613,N_19799);
and U19807 (N_19807,N_19655,N_19798);
nor U19808 (N_19808,N_19707,N_19684);
and U19809 (N_19809,N_19713,N_19611);
xnor U19810 (N_19810,N_19717,N_19646);
nand U19811 (N_19811,N_19747,N_19774);
xnor U19812 (N_19812,N_19777,N_19699);
and U19813 (N_19813,N_19695,N_19702);
or U19814 (N_19814,N_19729,N_19737);
or U19815 (N_19815,N_19623,N_19617);
nor U19816 (N_19816,N_19663,N_19756);
nor U19817 (N_19817,N_19744,N_19720);
and U19818 (N_19818,N_19605,N_19638);
nor U19819 (N_19819,N_19625,N_19644);
nor U19820 (N_19820,N_19676,N_19787);
nand U19821 (N_19821,N_19758,N_19706);
nor U19822 (N_19822,N_19710,N_19705);
and U19823 (N_19823,N_19620,N_19641);
xnor U19824 (N_19824,N_19766,N_19603);
nand U19825 (N_19825,N_19656,N_19795);
nor U19826 (N_19826,N_19783,N_19773);
and U19827 (N_19827,N_19750,N_19748);
and U19828 (N_19828,N_19786,N_19688);
and U19829 (N_19829,N_19719,N_19742);
or U19830 (N_19830,N_19722,N_19639);
or U19831 (N_19831,N_19732,N_19768);
or U19832 (N_19832,N_19778,N_19640);
and U19833 (N_19833,N_19793,N_19790);
and U19834 (N_19834,N_19650,N_19739);
xnor U19835 (N_19835,N_19674,N_19660);
nand U19836 (N_19836,N_19609,N_19694);
xnor U19837 (N_19837,N_19712,N_19741);
and U19838 (N_19838,N_19683,N_19653);
nor U19839 (N_19839,N_19607,N_19724);
nor U19840 (N_19840,N_19608,N_19630);
and U19841 (N_19841,N_19631,N_19753);
xnor U19842 (N_19842,N_19696,N_19754);
or U19843 (N_19843,N_19716,N_19691);
nand U19844 (N_19844,N_19654,N_19769);
xnor U19845 (N_19845,N_19785,N_19734);
xor U19846 (N_19846,N_19743,N_19721);
or U19847 (N_19847,N_19619,N_19614);
nor U19848 (N_19848,N_19728,N_19651);
xnor U19849 (N_19849,N_19627,N_19634);
nor U19850 (N_19850,N_19666,N_19697);
or U19851 (N_19851,N_19647,N_19681);
xor U19852 (N_19852,N_19689,N_19711);
nor U19853 (N_19853,N_19709,N_19606);
or U19854 (N_19854,N_19635,N_19735);
nor U19855 (N_19855,N_19708,N_19788);
or U19856 (N_19856,N_19671,N_19703);
nor U19857 (N_19857,N_19621,N_19665);
nor U19858 (N_19858,N_19746,N_19789);
nand U19859 (N_19859,N_19751,N_19610);
and U19860 (N_19860,N_19738,N_19733);
nand U19861 (N_19861,N_19761,N_19755);
nor U19862 (N_19862,N_19797,N_19679);
nand U19863 (N_19863,N_19794,N_19727);
nor U19864 (N_19864,N_19791,N_19661);
nand U19865 (N_19865,N_19775,N_19672);
and U19866 (N_19866,N_19765,N_19675);
nor U19867 (N_19867,N_19680,N_19677);
xor U19868 (N_19868,N_19687,N_19637);
nor U19869 (N_19869,N_19698,N_19669);
or U19870 (N_19870,N_19668,N_19658);
nand U19871 (N_19871,N_19770,N_19678);
or U19872 (N_19872,N_19648,N_19718);
or U19873 (N_19873,N_19726,N_19784);
xor U19874 (N_19874,N_19730,N_19796);
and U19875 (N_19875,N_19624,N_19686);
and U19876 (N_19876,N_19659,N_19779);
or U19877 (N_19877,N_19662,N_19612);
xor U19878 (N_19878,N_19642,N_19749);
nor U19879 (N_19879,N_19780,N_19745);
or U19880 (N_19880,N_19601,N_19685);
nor U19881 (N_19881,N_19664,N_19760);
xor U19882 (N_19882,N_19673,N_19690);
xor U19883 (N_19883,N_19723,N_19782);
xnor U19884 (N_19884,N_19715,N_19626);
and U19885 (N_19885,N_19615,N_19633);
xnor U19886 (N_19886,N_19600,N_19618);
nand U19887 (N_19887,N_19731,N_19652);
xor U19888 (N_19888,N_19752,N_19632);
or U19889 (N_19889,N_19792,N_19643);
nor U19890 (N_19890,N_19776,N_19759);
and U19891 (N_19891,N_19628,N_19692);
or U19892 (N_19892,N_19740,N_19781);
xor U19893 (N_19893,N_19764,N_19649);
nand U19894 (N_19894,N_19767,N_19757);
and U19895 (N_19895,N_19693,N_19616);
nand U19896 (N_19896,N_19700,N_19622);
nand U19897 (N_19897,N_19725,N_19667);
or U19898 (N_19898,N_19629,N_19762);
nand U19899 (N_19899,N_19704,N_19636);
and U19900 (N_19900,N_19789,N_19600);
or U19901 (N_19901,N_19643,N_19702);
or U19902 (N_19902,N_19792,N_19676);
nor U19903 (N_19903,N_19672,N_19675);
and U19904 (N_19904,N_19668,N_19605);
xor U19905 (N_19905,N_19689,N_19780);
nor U19906 (N_19906,N_19600,N_19657);
nor U19907 (N_19907,N_19763,N_19732);
nor U19908 (N_19908,N_19673,N_19765);
xor U19909 (N_19909,N_19654,N_19701);
or U19910 (N_19910,N_19725,N_19611);
or U19911 (N_19911,N_19639,N_19768);
xnor U19912 (N_19912,N_19708,N_19795);
nor U19913 (N_19913,N_19704,N_19612);
nand U19914 (N_19914,N_19722,N_19753);
or U19915 (N_19915,N_19626,N_19784);
nor U19916 (N_19916,N_19785,N_19789);
and U19917 (N_19917,N_19760,N_19734);
nand U19918 (N_19918,N_19670,N_19712);
xor U19919 (N_19919,N_19656,N_19664);
and U19920 (N_19920,N_19642,N_19604);
nor U19921 (N_19921,N_19687,N_19623);
nor U19922 (N_19922,N_19671,N_19734);
and U19923 (N_19923,N_19669,N_19761);
and U19924 (N_19924,N_19693,N_19618);
xnor U19925 (N_19925,N_19770,N_19697);
or U19926 (N_19926,N_19699,N_19601);
nor U19927 (N_19927,N_19673,N_19642);
nor U19928 (N_19928,N_19765,N_19740);
nor U19929 (N_19929,N_19655,N_19747);
nand U19930 (N_19930,N_19682,N_19708);
nor U19931 (N_19931,N_19774,N_19650);
or U19932 (N_19932,N_19668,N_19746);
nand U19933 (N_19933,N_19605,N_19648);
nand U19934 (N_19934,N_19750,N_19610);
nand U19935 (N_19935,N_19607,N_19689);
nand U19936 (N_19936,N_19708,N_19703);
nor U19937 (N_19937,N_19796,N_19600);
or U19938 (N_19938,N_19738,N_19772);
nor U19939 (N_19939,N_19693,N_19781);
nand U19940 (N_19940,N_19614,N_19652);
and U19941 (N_19941,N_19747,N_19711);
or U19942 (N_19942,N_19656,N_19629);
nand U19943 (N_19943,N_19714,N_19631);
or U19944 (N_19944,N_19768,N_19626);
and U19945 (N_19945,N_19773,N_19664);
or U19946 (N_19946,N_19724,N_19714);
and U19947 (N_19947,N_19791,N_19760);
nand U19948 (N_19948,N_19616,N_19624);
or U19949 (N_19949,N_19615,N_19783);
xnor U19950 (N_19950,N_19710,N_19706);
xnor U19951 (N_19951,N_19750,N_19644);
or U19952 (N_19952,N_19797,N_19673);
nor U19953 (N_19953,N_19671,N_19715);
xnor U19954 (N_19954,N_19771,N_19750);
xnor U19955 (N_19955,N_19768,N_19621);
nor U19956 (N_19956,N_19610,N_19790);
or U19957 (N_19957,N_19724,N_19693);
and U19958 (N_19958,N_19692,N_19688);
and U19959 (N_19959,N_19755,N_19757);
or U19960 (N_19960,N_19723,N_19653);
nand U19961 (N_19961,N_19793,N_19768);
and U19962 (N_19962,N_19791,N_19724);
nand U19963 (N_19963,N_19673,N_19712);
xor U19964 (N_19964,N_19660,N_19634);
nand U19965 (N_19965,N_19710,N_19631);
and U19966 (N_19966,N_19782,N_19783);
nand U19967 (N_19967,N_19757,N_19702);
or U19968 (N_19968,N_19665,N_19698);
and U19969 (N_19969,N_19716,N_19778);
xnor U19970 (N_19970,N_19711,N_19686);
and U19971 (N_19971,N_19638,N_19769);
nor U19972 (N_19972,N_19785,N_19761);
and U19973 (N_19973,N_19713,N_19670);
nor U19974 (N_19974,N_19691,N_19674);
or U19975 (N_19975,N_19751,N_19686);
nor U19976 (N_19976,N_19621,N_19640);
xor U19977 (N_19977,N_19621,N_19799);
xnor U19978 (N_19978,N_19654,N_19746);
nor U19979 (N_19979,N_19690,N_19662);
nor U19980 (N_19980,N_19764,N_19650);
or U19981 (N_19981,N_19729,N_19708);
or U19982 (N_19982,N_19665,N_19713);
xor U19983 (N_19983,N_19621,N_19674);
nor U19984 (N_19984,N_19666,N_19607);
or U19985 (N_19985,N_19788,N_19797);
and U19986 (N_19986,N_19618,N_19615);
nand U19987 (N_19987,N_19721,N_19726);
or U19988 (N_19988,N_19629,N_19636);
xor U19989 (N_19989,N_19629,N_19616);
xor U19990 (N_19990,N_19750,N_19672);
nor U19991 (N_19991,N_19657,N_19691);
nor U19992 (N_19992,N_19720,N_19647);
or U19993 (N_19993,N_19656,N_19607);
or U19994 (N_19994,N_19628,N_19664);
or U19995 (N_19995,N_19616,N_19758);
and U19996 (N_19996,N_19774,N_19778);
xor U19997 (N_19997,N_19695,N_19707);
nand U19998 (N_19998,N_19759,N_19794);
nor U19999 (N_19999,N_19689,N_19723);
nand U20000 (N_20000,N_19854,N_19842);
nand U20001 (N_20001,N_19810,N_19834);
xor U20002 (N_20002,N_19926,N_19893);
and U20003 (N_20003,N_19975,N_19802);
nand U20004 (N_20004,N_19901,N_19846);
xnor U20005 (N_20005,N_19980,N_19800);
xor U20006 (N_20006,N_19852,N_19839);
xnor U20007 (N_20007,N_19990,N_19828);
xor U20008 (N_20008,N_19905,N_19821);
xor U20009 (N_20009,N_19909,N_19999);
xnor U20010 (N_20010,N_19914,N_19988);
and U20011 (N_20011,N_19950,N_19819);
or U20012 (N_20012,N_19812,N_19886);
nor U20013 (N_20013,N_19872,N_19835);
and U20014 (N_20014,N_19959,N_19912);
xor U20015 (N_20015,N_19853,N_19836);
xnor U20016 (N_20016,N_19870,N_19978);
xor U20017 (N_20017,N_19813,N_19964);
and U20018 (N_20018,N_19930,N_19936);
nand U20019 (N_20019,N_19941,N_19815);
xnor U20020 (N_20020,N_19894,N_19804);
and U20021 (N_20021,N_19983,N_19885);
xnor U20022 (N_20022,N_19916,N_19991);
nand U20023 (N_20023,N_19951,N_19976);
nand U20024 (N_20024,N_19891,N_19907);
nand U20025 (N_20025,N_19939,N_19972);
or U20026 (N_20026,N_19977,N_19833);
and U20027 (N_20027,N_19995,N_19913);
xnor U20028 (N_20028,N_19859,N_19927);
and U20029 (N_20029,N_19862,N_19957);
nand U20030 (N_20030,N_19860,N_19823);
nand U20031 (N_20031,N_19877,N_19897);
and U20032 (N_20032,N_19963,N_19981);
and U20033 (N_20033,N_19934,N_19933);
nor U20034 (N_20034,N_19806,N_19851);
xnor U20035 (N_20035,N_19944,N_19831);
and U20036 (N_20036,N_19937,N_19974);
nor U20037 (N_20037,N_19884,N_19993);
nor U20038 (N_20038,N_19935,N_19887);
nor U20039 (N_20039,N_19880,N_19899);
xnor U20040 (N_20040,N_19845,N_19841);
xnor U20041 (N_20041,N_19827,N_19917);
xnor U20042 (N_20042,N_19882,N_19896);
xnor U20043 (N_20043,N_19807,N_19921);
and U20044 (N_20044,N_19911,N_19952);
nand U20045 (N_20045,N_19915,N_19902);
nor U20046 (N_20046,N_19816,N_19826);
nor U20047 (N_20047,N_19817,N_19979);
or U20048 (N_20048,N_19879,N_19850);
or U20049 (N_20049,N_19947,N_19892);
nand U20050 (N_20050,N_19918,N_19867);
or U20051 (N_20051,N_19874,N_19970);
nor U20052 (N_20052,N_19861,N_19992);
or U20053 (N_20053,N_19837,N_19994);
or U20054 (N_20054,N_19982,N_19869);
nor U20055 (N_20055,N_19820,N_19903);
xor U20056 (N_20056,N_19946,N_19910);
nand U20057 (N_20057,N_19883,N_19809);
nor U20058 (N_20058,N_19890,N_19920);
nand U20059 (N_20059,N_19945,N_19965);
xor U20060 (N_20060,N_19925,N_19898);
xnor U20061 (N_20061,N_19943,N_19855);
xor U20062 (N_20062,N_19973,N_19829);
or U20063 (N_20063,N_19840,N_19960);
and U20064 (N_20064,N_19923,N_19830);
nand U20065 (N_20065,N_19932,N_19956);
and U20066 (N_20066,N_19811,N_19998);
nor U20067 (N_20067,N_19895,N_19942);
and U20068 (N_20068,N_19888,N_19822);
xor U20069 (N_20069,N_19858,N_19969);
nor U20070 (N_20070,N_19987,N_19863);
nand U20071 (N_20071,N_19843,N_19849);
xnor U20072 (N_20072,N_19856,N_19808);
nor U20073 (N_20073,N_19873,N_19948);
or U20074 (N_20074,N_19967,N_19847);
nor U20075 (N_20075,N_19954,N_19868);
nand U20076 (N_20076,N_19844,N_19838);
nor U20077 (N_20077,N_19984,N_19878);
and U20078 (N_20078,N_19924,N_19958);
nor U20079 (N_20079,N_19966,N_19881);
or U20080 (N_20080,N_19938,N_19929);
xnor U20081 (N_20081,N_19803,N_19928);
xnor U20082 (N_20082,N_19922,N_19961);
xnor U20083 (N_20083,N_19876,N_19997);
or U20084 (N_20084,N_19814,N_19900);
and U20085 (N_20085,N_19871,N_19919);
and U20086 (N_20086,N_19818,N_19989);
nor U20087 (N_20087,N_19824,N_19832);
nand U20088 (N_20088,N_19971,N_19857);
nand U20089 (N_20089,N_19904,N_19825);
nor U20090 (N_20090,N_19865,N_19968);
xnor U20091 (N_20091,N_19875,N_19866);
nor U20092 (N_20092,N_19940,N_19953);
nand U20093 (N_20093,N_19931,N_19986);
nand U20094 (N_20094,N_19996,N_19801);
nand U20095 (N_20095,N_19906,N_19985);
nand U20096 (N_20096,N_19962,N_19955);
nand U20097 (N_20097,N_19908,N_19805);
or U20098 (N_20098,N_19949,N_19864);
and U20099 (N_20099,N_19848,N_19889);
or U20100 (N_20100,N_19815,N_19801);
xnor U20101 (N_20101,N_19894,N_19850);
nor U20102 (N_20102,N_19941,N_19947);
and U20103 (N_20103,N_19894,N_19851);
xor U20104 (N_20104,N_19851,N_19979);
or U20105 (N_20105,N_19977,N_19819);
nand U20106 (N_20106,N_19818,N_19827);
or U20107 (N_20107,N_19940,N_19992);
xor U20108 (N_20108,N_19950,N_19912);
xor U20109 (N_20109,N_19865,N_19819);
and U20110 (N_20110,N_19973,N_19825);
nor U20111 (N_20111,N_19956,N_19964);
or U20112 (N_20112,N_19814,N_19842);
nor U20113 (N_20113,N_19811,N_19877);
xor U20114 (N_20114,N_19994,N_19909);
nand U20115 (N_20115,N_19891,N_19966);
and U20116 (N_20116,N_19890,N_19993);
and U20117 (N_20117,N_19923,N_19970);
or U20118 (N_20118,N_19983,N_19844);
xor U20119 (N_20119,N_19967,N_19851);
and U20120 (N_20120,N_19848,N_19993);
xor U20121 (N_20121,N_19923,N_19889);
and U20122 (N_20122,N_19890,N_19871);
and U20123 (N_20123,N_19952,N_19983);
nand U20124 (N_20124,N_19949,N_19818);
or U20125 (N_20125,N_19852,N_19872);
xnor U20126 (N_20126,N_19922,N_19855);
and U20127 (N_20127,N_19857,N_19907);
nor U20128 (N_20128,N_19829,N_19970);
nor U20129 (N_20129,N_19904,N_19917);
nand U20130 (N_20130,N_19818,N_19978);
and U20131 (N_20131,N_19938,N_19981);
nor U20132 (N_20132,N_19818,N_19953);
nand U20133 (N_20133,N_19994,N_19857);
or U20134 (N_20134,N_19994,N_19916);
xnor U20135 (N_20135,N_19993,N_19802);
nor U20136 (N_20136,N_19880,N_19898);
and U20137 (N_20137,N_19859,N_19901);
nor U20138 (N_20138,N_19996,N_19919);
xor U20139 (N_20139,N_19914,N_19813);
and U20140 (N_20140,N_19992,N_19968);
xor U20141 (N_20141,N_19940,N_19845);
or U20142 (N_20142,N_19804,N_19951);
nand U20143 (N_20143,N_19816,N_19801);
or U20144 (N_20144,N_19828,N_19982);
or U20145 (N_20145,N_19963,N_19906);
nand U20146 (N_20146,N_19918,N_19813);
and U20147 (N_20147,N_19980,N_19930);
and U20148 (N_20148,N_19885,N_19863);
xnor U20149 (N_20149,N_19843,N_19961);
xnor U20150 (N_20150,N_19913,N_19899);
nor U20151 (N_20151,N_19925,N_19880);
nand U20152 (N_20152,N_19962,N_19884);
xnor U20153 (N_20153,N_19843,N_19883);
and U20154 (N_20154,N_19986,N_19912);
and U20155 (N_20155,N_19824,N_19868);
and U20156 (N_20156,N_19929,N_19848);
xor U20157 (N_20157,N_19999,N_19872);
nand U20158 (N_20158,N_19892,N_19932);
or U20159 (N_20159,N_19814,N_19877);
nor U20160 (N_20160,N_19943,N_19848);
and U20161 (N_20161,N_19873,N_19943);
nand U20162 (N_20162,N_19831,N_19981);
nor U20163 (N_20163,N_19809,N_19861);
and U20164 (N_20164,N_19835,N_19930);
xnor U20165 (N_20165,N_19861,N_19985);
nand U20166 (N_20166,N_19812,N_19976);
nand U20167 (N_20167,N_19888,N_19871);
nor U20168 (N_20168,N_19833,N_19992);
nor U20169 (N_20169,N_19832,N_19940);
xor U20170 (N_20170,N_19808,N_19879);
nor U20171 (N_20171,N_19959,N_19910);
and U20172 (N_20172,N_19929,N_19871);
nand U20173 (N_20173,N_19975,N_19941);
and U20174 (N_20174,N_19954,N_19915);
nand U20175 (N_20175,N_19931,N_19969);
nand U20176 (N_20176,N_19866,N_19836);
and U20177 (N_20177,N_19951,N_19947);
nor U20178 (N_20178,N_19883,N_19808);
nand U20179 (N_20179,N_19834,N_19877);
xnor U20180 (N_20180,N_19918,N_19972);
or U20181 (N_20181,N_19905,N_19837);
nand U20182 (N_20182,N_19859,N_19972);
nor U20183 (N_20183,N_19950,N_19810);
or U20184 (N_20184,N_19992,N_19917);
and U20185 (N_20185,N_19960,N_19938);
nor U20186 (N_20186,N_19873,N_19934);
or U20187 (N_20187,N_19983,N_19969);
nand U20188 (N_20188,N_19880,N_19852);
nand U20189 (N_20189,N_19848,N_19926);
nand U20190 (N_20190,N_19833,N_19943);
and U20191 (N_20191,N_19966,N_19947);
xnor U20192 (N_20192,N_19846,N_19928);
nand U20193 (N_20193,N_19881,N_19942);
nor U20194 (N_20194,N_19835,N_19976);
nor U20195 (N_20195,N_19982,N_19852);
xnor U20196 (N_20196,N_19955,N_19850);
and U20197 (N_20197,N_19963,N_19822);
or U20198 (N_20198,N_19883,N_19928);
nand U20199 (N_20199,N_19871,N_19853);
or U20200 (N_20200,N_20154,N_20158);
nand U20201 (N_20201,N_20053,N_20060);
nand U20202 (N_20202,N_20162,N_20124);
xnor U20203 (N_20203,N_20132,N_20136);
nor U20204 (N_20204,N_20073,N_20172);
nand U20205 (N_20205,N_20174,N_20098);
xor U20206 (N_20206,N_20010,N_20156);
and U20207 (N_20207,N_20102,N_20085);
and U20208 (N_20208,N_20051,N_20077);
nand U20209 (N_20209,N_20028,N_20128);
or U20210 (N_20210,N_20161,N_20067);
or U20211 (N_20211,N_20117,N_20061);
or U20212 (N_20212,N_20034,N_20152);
or U20213 (N_20213,N_20182,N_20000);
nand U20214 (N_20214,N_20122,N_20116);
nor U20215 (N_20215,N_20047,N_20026);
or U20216 (N_20216,N_20090,N_20168);
nand U20217 (N_20217,N_20138,N_20181);
or U20218 (N_20218,N_20107,N_20140);
xnor U20219 (N_20219,N_20044,N_20105);
nand U20220 (N_20220,N_20036,N_20069);
nor U20221 (N_20221,N_20032,N_20127);
or U20222 (N_20222,N_20015,N_20103);
and U20223 (N_20223,N_20176,N_20184);
xnor U20224 (N_20224,N_20003,N_20120);
or U20225 (N_20225,N_20088,N_20066);
and U20226 (N_20226,N_20106,N_20057);
nor U20227 (N_20227,N_20079,N_20133);
nand U20228 (N_20228,N_20006,N_20005);
or U20229 (N_20229,N_20074,N_20039);
and U20230 (N_20230,N_20040,N_20011);
nand U20231 (N_20231,N_20087,N_20144);
nor U20232 (N_20232,N_20141,N_20110);
nand U20233 (N_20233,N_20020,N_20056);
nand U20234 (N_20234,N_20025,N_20153);
xnor U20235 (N_20235,N_20062,N_20049);
nand U20236 (N_20236,N_20052,N_20163);
and U20237 (N_20237,N_20129,N_20022);
or U20238 (N_20238,N_20197,N_20188);
or U20239 (N_20239,N_20119,N_20097);
or U20240 (N_20240,N_20021,N_20109);
and U20241 (N_20241,N_20091,N_20075);
and U20242 (N_20242,N_20198,N_20179);
xor U20243 (N_20243,N_20167,N_20121);
xor U20244 (N_20244,N_20150,N_20001);
nor U20245 (N_20245,N_20186,N_20046);
nor U20246 (N_20246,N_20007,N_20092);
nor U20247 (N_20247,N_20094,N_20166);
xnor U20248 (N_20248,N_20089,N_20035);
or U20249 (N_20249,N_20112,N_20135);
xor U20250 (N_20250,N_20169,N_20175);
xor U20251 (N_20251,N_20042,N_20063);
or U20252 (N_20252,N_20160,N_20123);
and U20253 (N_20253,N_20023,N_20159);
and U20254 (N_20254,N_20031,N_20195);
nand U20255 (N_20255,N_20148,N_20126);
and U20256 (N_20256,N_20180,N_20083);
and U20257 (N_20257,N_20134,N_20113);
xor U20258 (N_20258,N_20037,N_20157);
xnor U20259 (N_20259,N_20139,N_20002);
or U20260 (N_20260,N_20095,N_20165);
or U20261 (N_20261,N_20178,N_20050);
xor U20262 (N_20262,N_20187,N_20142);
and U20263 (N_20263,N_20016,N_20014);
and U20264 (N_20264,N_20177,N_20170);
or U20265 (N_20265,N_20009,N_20108);
nand U20266 (N_20266,N_20076,N_20072);
nand U20267 (N_20267,N_20071,N_20093);
and U20268 (N_20268,N_20008,N_20143);
nand U20269 (N_20269,N_20084,N_20147);
nand U20270 (N_20270,N_20192,N_20146);
nand U20271 (N_20271,N_20100,N_20058);
and U20272 (N_20272,N_20194,N_20018);
and U20273 (N_20273,N_20081,N_20019);
or U20274 (N_20274,N_20068,N_20078);
xnor U20275 (N_20275,N_20065,N_20099);
xnor U20276 (N_20276,N_20054,N_20125);
nand U20277 (N_20277,N_20012,N_20030);
or U20278 (N_20278,N_20173,N_20013);
xor U20279 (N_20279,N_20191,N_20171);
nand U20280 (N_20280,N_20164,N_20045);
and U20281 (N_20281,N_20183,N_20027);
and U20282 (N_20282,N_20104,N_20190);
nor U20283 (N_20283,N_20082,N_20149);
nand U20284 (N_20284,N_20038,N_20059);
or U20285 (N_20285,N_20004,N_20029);
or U20286 (N_20286,N_20185,N_20086);
and U20287 (N_20287,N_20118,N_20017);
or U20288 (N_20288,N_20070,N_20131);
nor U20289 (N_20289,N_20196,N_20189);
nand U20290 (N_20290,N_20111,N_20080);
and U20291 (N_20291,N_20137,N_20064);
or U20292 (N_20292,N_20199,N_20041);
nand U20293 (N_20293,N_20155,N_20024);
xor U20294 (N_20294,N_20145,N_20115);
or U20295 (N_20295,N_20043,N_20101);
nor U20296 (N_20296,N_20055,N_20114);
nand U20297 (N_20297,N_20033,N_20096);
and U20298 (N_20298,N_20048,N_20151);
or U20299 (N_20299,N_20193,N_20130);
nor U20300 (N_20300,N_20105,N_20176);
and U20301 (N_20301,N_20177,N_20097);
xor U20302 (N_20302,N_20001,N_20178);
xnor U20303 (N_20303,N_20120,N_20133);
and U20304 (N_20304,N_20162,N_20008);
nor U20305 (N_20305,N_20068,N_20023);
nor U20306 (N_20306,N_20048,N_20154);
or U20307 (N_20307,N_20034,N_20095);
and U20308 (N_20308,N_20007,N_20018);
nor U20309 (N_20309,N_20026,N_20111);
nand U20310 (N_20310,N_20157,N_20126);
or U20311 (N_20311,N_20075,N_20107);
and U20312 (N_20312,N_20196,N_20043);
xor U20313 (N_20313,N_20175,N_20130);
nand U20314 (N_20314,N_20155,N_20124);
xor U20315 (N_20315,N_20059,N_20043);
xnor U20316 (N_20316,N_20040,N_20080);
or U20317 (N_20317,N_20162,N_20048);
and U20318 (N_20318,N_20134,N_20069);
or U20319 (N_20319,N_20089,N_20019);
xor U20320 (N_20320,N_20031,N_20008);
and U20321 (N_20321,N_20034,N_20160);
or U20322 (N_20322,N_20046,N_20096);
and U20323 (N_20323,N_20066,N_20152);
nor U20324 (N_20324,N_20179,N_20082);
nand U20325 (N_20325,N_20156,N_20182);
or U20326 (N_20326,N_20130,N_20068);
nor U20327 (N_20327,N_20166,N_20002);
nand U20328 (N_20328,N_20015,N_20009);
and U20329 (N_20329,N_20125,N_20017);
nand U20330 (N_20330,N_20051,N_20172);
and U20331 (N_20331,N_20190,N_20035);
xor U20332 (N_20332,N_20052,N_20134);
nand U20333 (N_20333,N_20013,N_20102);
nor U20334 (N_20334,N_20112,N_20053);
xor U20335 (N_20335,N_20026,N_20144);
nand U20336 (N_20336,N_20141,N_20101);
xnor U20337 (N_20337,N_20118,N_20078);
and U20338 (N_20338,N_20070,N_20081);
nor U20339 (N_20339,N_20197,N_20027);
xnor U20340 (N_20340,N_20168,N_20094);
or U20341 (N_20341,N_20163,N_20133);
and U20342 (N_20342,N_20159,N_20115);
xnor U20343 (N_20343,N_20041,N_20049);
and U20344 (N_20344,N_20087,N_20017);
nor U20345 (N_20345,N_20037,N_20026);
and U20346 (N_20346,N_20014,N_20067);
nor U20347 (N_20347,N_20134,N_20070);
nand U20348 (N_20348,N_20011,N_20037);
nand U20349 (N_20349,N_20017,N_20098);
xor U20350 (N_20350,N_20044,N_20003);
nor U20351 (N_20351,N_20135,N_20118);
and U20352 (N_20352,N_20112,N_20065);
nand U20353 (N_20353,N_20159,N_20096);
or U20354 (N_20354,N_20170,N_20092);
nand U20355 (N_20355,N_20032,N_20110);
nand U20356 (N_20356,N_20015,N_20173);
nor U20357 (N_20357,N_20127,N_20039);
or U20358 (N_20358,N_20088,N_20030);
or U20359 (N_20359,N_20083,N_20077);
nand U20360 (N_20360,N_20083,N_20082);
nor U20361 (N_20361,N_20111,N_20077);
or U20362 (N_20362,N_20134,N_20032);
nor U20363 (N_20363,N_20176,N_20177);
nand U20364 (N_20364,N_20073,N_20037);
nor U20365 (N_20365,N_20091,N_20138);
nand U20366 (N_20366,N_20109,N_20046);
and U20367 (N_20367,N_20085,N_20149);
and U20368 (N_20368,N_20169,N_20039);
xnor U20369 (N_20369,N_20133,N_20105);
xnor U20370 (N_20370,N_20045,N_20137);
nor U20371 (N_20371,N_20140,N_20040);
xnor U20372 (N_20372,N_20135,N_20104);
nor U20373 (N_20373,N_20111,N_20116);
nand U20374 (N_20374,N_20070,N_20117);
and U20375 (N_20375,N_20184,N_20002);
or U20376 (N_20376,N_20037,N_20133);
nand U20377 (N_20377,N_20110,N_20107);
nand U20378 (N_20378,N_20100,N_20147);
xnor U20379 (N_20379,N_20075,N_20142);
nor U20380 (N_20380,N_20076,N_20059);
nor U20381 (N_20381,N_20112,N_20198);
or U20382 (N_20382,N_20091,N_20013);
nor U20383 (N_20383,N_20118,N_20024);
or U20384 (N_20384,N_20000,N_20122);
nor U20385 (N_20385,N_20126,N_20185);
xor U20386 (N_20386,N_20174,N_20043);
nand U20387 (N_20387,N_20109,N_20181);
nor U20388 (N_20388,N_20083,N_20137);
nor U20389 (N_20389,N_20004,N_20160);
nor U20390 (N_20390,N_20041,N_20154);
nor U20391 (N_20391,N_20002,N_20164);
nor U20392 (N_20392,N_20076,N_20086);
or U20393 (N_20393,N_20193,N_20005);
xor U20394 (N_20394,N_20004,N_20111);
xnor U20395 (N_20395,N_20125,N_20038);
nand U20396 (N_20396,N_20040,N_20093);
nor U20397 (N_20397,N_20051,N_20143);
xnor U20398 (N_20398,N_20095,N_20055);
nand U20399 (N_20399,N_20106,N_20054);
nor U20400 (N_20400,N_20391,N_20298);
or U20401 (N_20401,N_20330,N_20299);
nor U20402 (N_20402,N_20293,N_20275);
nand U20403 (N_20403,N_20237,N_20214);
and U20404 (N_20404,N_20282,N_20390);
nor U20405 (N_20405,N_20397,N_20232);
xor U20406 (N_20406,N_20253,N_20383);
and U20407 (N_20407,N_20315,N_20318);
nor U20408 (N_20408,N_20382,N_20358);
xnor U20409 (N_20409,N_20277,N_20262);
nor U20410 (N_20410,N_20288,N_20221);
and U20411 (N_20411,N_20331,N_20393);
or U20412 (N_20412,N_20226,N_20233);
nor U20413 (N_20413,N_20270,N_20323);
xnor U20414 (N_20414,N_20376,N_20324);
or U20415 (N_20415,N_20377,N_20244);
and U20416 (N_20416,N_20285,N_20261);
or U20417 (N_20417,N_20335,N_20268);
or U20418 (N_20418,N_20272,N_20290);
nand U20419 (N_20419,N_20364,N_20291);
nor U20420 (N_20420,N_20276,N_20368);
and U20421 (N_20421,N_20248,N_20325);
nand U20422 (N_20422,N_20337,N_20314);
nand U20423 (N_20423,N_20217,N_20338);
nor U20424 (N_20424,N_20235,N_20342);
or U20425 (N_20425,N_20267,N_20225);
nand U20426 (N_20426,N_20212,N_20273);
nand U20427 (N_20427,N_20359,N_20300);
xor U20428 (N_20428,N_20230,N_20200);
nand U20429 (N_20429,N_20387,N_20327);
nor U20430 (N_20430,N_20220,N_20210);
nand U20431 (N_20431,N_20381,N_20329);
xor U20432 (N_20432,N_20295,N_20341);
nand U20433 (N_20433,N_20375,N_20252);
nor U20434 (N_20434,N_20351,N_20355);
and U20435 (N_20435,N_20336,N_20208);
and U20436 (N_20436,N_20245,N_20322);
and U20437 (N_20437,N_20392,N_20348);
and U20438 (N_20438,N_20339,N_20398);
nor U20439 (N_20439,N_20216,N_20205);
xor U20440 (N_20440,N_20287,N_20242);
nor U20441 (N_20441,N_20345,N_20274);
nor U20442 (N_20442,N_20384,N_20241);
and U20443 (N_20443,N_20257,N_20250);
nor U20444 (N_20444,N_20296,N_20306);
nand U20445 (N_20445,N_20304,N_20349);
nor U20446 (N_20446,N_20334,N_20215);
or U20447 (N_20447,N_20254,N_20307);
nor U20448 (N_20448,N_20260,N_20258);
and U20449 (N_20449,N_20326,N_20309);
and U20450 (N_20450,N_20256,N_20265);
nand U20451 (N_20451,N_20389,N_20302);
or U20452 (N_20452,N_20380,N_20363);
or U20453 (N_20453,N_20366,N_20222);
or U20454 (N_20454,N_20281,N_20350);
nor U20455 (N_20455,N_20319,N_20347);
and U20456 (N_20456,N_20247,N_20206);
and U20457 (N_20457,N_20357,N_20213);
xor U20458 (N_20458,N_20246,N_20316);
nand U20459 (N_20459,N_20279,N_20228);
or U20460 (N_20460,N_20255,N_20388);
and U20461 (N_20461,N_20238,N_20310);
nor U20462 (N_20462,N_20223,N_20289);
nand U20463 (N_20463,N_20374,N_20385);
and U20464 (N_20464,N_20311,N_20394);
nor U20465 (N_20465,N_20263,N_20367);
and U20466 (N_20466,N_20356,N_20399);
and U20467 (N_20467,N_20224,N_20305);
or U20468 (N_20468,N_20202,N_20264);
nor U20469 (N_20469,N_20353,N_20209);
or U20470 (N_20470,N_20231,N_20239);
nand U20471 (N_20471,N_20271,N_20211);
nor U20472 (N_20472,N_20328,N_20371);
xor U20473 (N_20473,N_20284,N_20301);
xnor U20474 (N_20474,N_20266,N_20249);
nor U20475 (N_20475,N_20379,N_20219);
xnor U20476 (N_20476,N_20251,N_20346);
and U20477 (N_20477,N_20372,N_20343);
nand U20478 (N_20478,N_20373,N_20369);
and U20479 (N_20479,N_20236,N_20286);
xor U20480 (N_20480,N_20204,N_20297);
xor U20481 (N_20481,N_20229,N_20292);
or U20482 (N_20482,N_20283,N_20344);
nor U20483 (N_20483,N_20278,N_20378);
xnor U20484 (N_20484,N_20308,N_20320);
nor U20485 (N_20485,N_20361,N_20321);
nand U20486 (N_20486,N_20243,N_20313);
or U20487 (N_20487,N_20294,N_20259);
xnor U20488 (N_20488,N_20386,N_20365);
nor U20489 (N_20489,N_20240,N_20333);
or U20490 (N_20490,N_20218,N_20360);
and U20491 (N_20491,N_20201,N_20207);
nand U20492 (N_20492,N_20396,N_20362);
nor U20493 (N_20493,N_20340,N_20395);
and U20494 (N_20494,N_20354,N_20317);
xor U20495 (N_20495,N_20227,N_20269);
nand U20496 (N_20496,N_20332,N_20234);
and U20497 (N_20497,N_20312,N_20352);
or U20498 (N_20498,N_20370,N_20203);
nand U20499 (N_20499,N_20303,N_20280);
or U20500 (N_20500,N_20381,N_20207);
and U20501 (N_20501,N_20238,N_20233);
nor U20502 (N_20502,N_20377,N_20259);
nor U20503 (N_20503,N_20354,N_20370);
nor U20504 (N_20504,N_20304,N_20275);
xor U20505 (N_20505,N_20201,N_20317);
and U20506 (N_20506,N_20360,N_20247);
or U20507 (N_20507,N_20250,N_20312);
or U20508 (N_20508,N_20204,N_20267);
nand U20509 (N_20509,N_20377,N_20357);
or U20510 (N_20510,N_20241,N_20247);
nand U20511 (N_20511,N_20350,N_20217);
or U20512 (N_20512,N_20308,N_20224);
nor U20513 (N_20513,N_20366,N_20384);
nand U20514 (N_20514,N_20265,N_20232);
xnor U20515 (N_20515,N_20245,N_20217);
nor U20516 (N_20516,N_20337,N_20266);
and U20517 (N_20517,N_20322,N_20274);
xor U20518 (N_20518,N_20259,N_20372);
xnor U20519 (N_20519,N_20373,N_20275);
nand U20520 (N_20520,N_20343,N_20210);
nor U20521 (N_20521,N_20259,N_20242);
nand U20522 (N_20522,N_20347,N_20242);
or U20523 (N_20523,N_20208,N_20366);
or U20524 (N_20524,N_20306,N_20389);
and U20525 (N_20525,N_20305,N_20351);
nand U20526 (N_20526,N_20369,N_20305);
nor U20527 (N_20527,N_20281,N_20289);
and U20528 (N_20528,N_20271,N_20326);
nand U20529 (N_20529,N_20247,N_20372);
xnor U20530 (N_20530,N_20385,N_20281);
xnor U20531 (N_20531,N_20383,N_20256);
and U20532 (N_20532,N_20352,N_20230);
xnor U20533 (N_20533,N_20329,N_20227);
or U20534 (N_20534,N_20310,N_20218);
nand U20535 (N_20535,N_20348,N_20218);
xor U20536 (N_20536,N_20267,N_20242);
xnor U20537 (N_20537,N_20338,N_20381);
nor U20538 (N_20538,N_20342,N_20288);
nor U20539 (N_20539,N_20210,N_20258);
nor U20540 (N_20540,N_20203,N_20251);
nor U20541 (N_20541,N_20273,N_20225);
and U20542 (N_20542,N_20385,N_20335);
nand U20543 (N_20543,N_20377,N_20266);
nor U20544 (N_20544,N_20297,N_20214);
nor U20545 (N_20545,N_20310,N_20313);
or U20546 (N_20546,N_20308,N_20314);
nand U20547 (N_20547,N_20318,N_20258);
xor U20548 (N_20548,N_20228,N_20359);
nor U20549 (N_20549,N_20269,N_20294);
or U20550 (N_20550,N_20332,N_20395);
nand U20551 (N_20551,N_20326,N_20376);
and U20552 (N_20552,N_20207,N_20253);
nor U20553 (N_20553,N_20294,N_20252);
or U20554 (N_20554,N_20304,N_20395);
xor U20555 (N_20555,N_20377,N_20221);
and U20556 (N_20556,N_20311,N_20397);
and U20557 (N_20557,N_20363,N_20365);
nor U20558 (N_20558,N_20303,N_20317);
nand U20559 (N_20559,N_20286,N_20372);
xor U20560 (N_20560,N_20212,N_20295);
nand U20561 (N_20561,N_20224,N_20314);
nand U20562 (N_20562,N_20273,N_20299);
or U20563 (N_20563,N_20214,N_20350);
nor U20564 (N_20564,N_20237,N_20315);
nor U20565 (N_20565,N_20333,N_20298);
or U20566 (N_20566,N_20331,N_20319);
nand U20567 (N_20567,N_20266,N_20231);
nand U20568 (N_20568,N_20251,N_20293);
and U20569 (N_20569,N_20361,N_20332);
or U20570 (N_20570,N_20286,N_20342);
nor U20571 (N_20571,N_20320,N_20354);
or U20572 (N_20572,N_20389,N_20295);
nor U20573 (N_20573,N_20262,N_20207);
xnor U20574 (N_20574,N_20283,N_20289);
and U20575 (N_20575,N_20341,N_20238);
or U20576 (N_20576,N_20211,N_20270);
nor U20577 (N_20577,N_20233,N_20386);
xnor U20578 (N_20578,N_20392,N_20263);
nor U20579 (N_20579,N_20336,N_20276);
nand U20580 (N_20580,N_20375,N_20340);
or U20581 (N_20581,N_20332,N_20297);
or U20582 (N_20582,N_20322,N_20395);
nand U20583 (N_20583,N_20301,N_20279);
nand U20584 (N_20584,N_20275,N_20259);
xor U20585 (N_20585,N_20315,N_20338);
nand U20586 (N_20586,N_20356,N_20203);
or U20587 (N_20587,N_20294,N_20332);
xor U20588 (N_20588,N_20389,N_20220);
nand U20589 (N_20589,N_20314,N_20268);
nor U20590 (N_20590,N_20305,N_20342);
or U20591 (N_20591,N_20391,N_20378);
or U20592 (N_20592,N_20353,N_20231);
or U20593 (N_20593,N_20391,N_20314);
or U20594 (N_20594,N_20344,N_20398);
nand U20595 (N_20595,N_20377,N_20337);
and U20596 (N_20596,N_20250,N_20231);
nor U20597 (N_20597,N_20267,N_20300);
nand U20598 (N_20598,N_20336,N_20250);
and U20599 (N_20599,N_20254,N_20238);
nand U20600 (N_20600,N_20500,N_20510);
xnor U20601 (N_20601,N_20451,N_20537);
nand U20602 (N_20602,N_20579,N_20525);
xor U20603 (N_20603,N_20488,N_20582);
nand U20604 (N_20604,N_20462,N_20529);
and U20605 (N_20605,N_20505,N_20499);
and U20606 (N_20606,N_20434,N_20531);
and U20607 (N_20607,N_20543,N_20435);
and U20608 (N_20608,N_20503,N_20568);
xor U20609 (N_20609,N_20493,N_20418);
or U20610 (N_20610,N_20518,N_20452);
xor U20611 (N_20611,N_20477,N_20420);
nor U20612 (N_20612,N_20547,N_20482);
nor U20613 (N_20613,N_20437,N_20442);
or U20614 (N_20614,N_20599,N_20522);
or U20615 (N_20615,N_20570,N_20440);
and U20616 (N_20616,N_20551,N_20564);
nor U20617 (N_20617,N_20586,N_20517);
and U20618 (N_20618,N_20436,N_20466);
and U20619 (N_20619,N_20456,N_20526);
and U20620 (N_20620,N_20511,N_20595);
or U20621 (N_20621,N_20560,N_20559);
and U20622 (N_20622,N_20561,N_20578);
xnor U20623 (N_20623,N_20485,N_20457);
nor U20624 (N_20624,N_20405,N_20430);
and U20625 (N_20625,N_20447,N_20494);
xnor U20626 (N_20626,N_20549,N_20577);
and U20627 (N_20627,N_20541,N_20489);
or U20628 (N_20628,N_20557,N_20453);
xor U20629 (N_20629,N_20567,N_20514);
and U20630 (N_20630,N_20438,N_20546);
and U20631 (N_20631,N_20449,N_20473);
nand U20632 (N_20632,N_20539,N_20474);
and U20633 (N_20633,N_20492,N_20501);
and U20634 (N_20634,N_20433,N_20571);
nand U20635 (N_20635,N_20454,N_20523);
and U20636 (N_20636,N_20417,N_20475);
or U20637 (N_20637,N_20544,N_20556);
nor U20638 (N_20638,N_20515,N_20536);
nor U20639 (N_20639,N_20471,N_20520);
nand U20640 (N_20640,N_20480,N_20455);
nand U20641 (N_20641,N_20583,N_20572);
nand U20642 (N_20642,N_20598,N_20575);
nand U20643 (N_20643,N_20444,N_20469);
and U20644 (N_20644,N_20465,N_20507);
and U20645 (N_20645,N_20472,N_20461);
nand U20646 (N_20646,N_20594,N_20502);
xnor U20647 (N_20647,N_20450,N_20519);
xor U20648 (N_20648,N_20470,N_20592);
xor U20649 (N_20649,N_20468,N_20552);
and U20650 (N_20650,N_20506,N_20497);
xnor U20651 (N_20651,N_20459,N_20584);
or U20652 (N_20652,N_20413,N_20597);
and U20653 (N_20653,N_20576,N_20425);
xor U20654 (N_20654,N_20402,N_20481);
nor U20655 (N_20655,N_20408,N_20423);
or U20656 (N_20656,N_20508,N_20491);
or U20657 (N_20657,N_20439,N_20590);
nor U20658 (N_20658,N_20504,N_20591);
and U20659 (N_20659,N_20589,N_20458);
xnor U20660 (N_20660,N_20587,N_20407);
and U20661 (N_20661,N_20479,N_20527);
or U20662 (N_20662,N_20463,N_20464);
or U20663 (N_20663,N_20476,N_20445);
and U20664 (N_20664,N_20562,N_20460);
or U20665 (N_20665,N_20534,N_20569);
nand U20666 (N_20666,N_20431,N_20580);
xor U20667 (N_20667,N_20496,N_20404);
and U20668 (N_20668,N_20409,N_20516);
or U20669 (N_20669,N_20446,N_20528);
nor U20670 (N_20670,N_20530,N_20415);
and U20671 (N_20671,N_20540,N_20513);
and U20672 (N_20672,N_20422,N_20448);
or U20673 (N_20673,N_20410,N_20588);
nor U20674 (N_20674,N_20484,N_20424);
and U20675 (N_20675,N_20574,N_20558);
xnor U20676 (N_20676,N_20532,N_20406);
and U20677 (N_20677,N_20535,N_20512);
or U20678 (N_20678,N_20566,N_20432);
or U20679 (N_20679,N_20443,N_20401);
xor U20680 (N_20680,N_20538,N_20550);
xnor U20681 (N_20681,N_20553,N_20585);
and U20682 (N_20682,N_20596,N_20467);
nor U20683 (N_20683,N_20581,N_20483);
xnor U20684 (N_20684,N_20419,N_20486);
nand U20685 (N_20685,N_20555,N_20542);
nor U20686 (N_20686,N_20545,N_20563);
and U20687 (N_20687,N_20490,N_20428);
xor U20688 (N_20688,N_20509,N_20421);
nor U20689 (N_20689,N_20521,N_20487);
nand U20690 (N_20690,N_20427,N_20414);
xnor U20691 (N_20691,N_20403,N_20412);
or U20692 (N_20692,N_20441,N_20593);
nand U20693 (N_20693,N_20478,N_20573);
nand U20694 (N_20694,N_20495,N_20498);
or U20695 (N_20695,N_20554,N_20565);
or U20696 (N_20696,N_20426,N_20411);
nand U20697 (N_20697,N_20429,N_20416);
and U20698 (N_20698,N_20548,N_20400);
nand U20699 (N_20699,N_20524,N_20533);
and U20700 (N_20700,N_20578,N_20574);
and U20701 (N_20701,N_20554,N_20475);
nor U20702 (N_20702,N_20407,N_20513);
or U20703 (N_20703,N_20581,N_20475);
nand U20704 (N_20704,N_20585,N_20470);
or U20705 (N_20705,N_20463,N_20440);
nand U20706 (N_20706,N_20432,N_20583);
or U20707 (N_20707,N_20584,N_20567);
or U20708 (N_20708,N_20403,N_20538);
nand U20709 (N_20709,N_20532,N_20507);
nand U20710 (N_20710,N_20420,N_20577);
nor U20711 (N_20711,N_20584,N_20571);
nor U20712 (N_20712,N_20523,N_20404);
or U20713 (N_20713,N_20464,N_20571);
or U20714 (N_20714,N_20482,N_20575);
or U20715 (N_20715,N_20461,N_20576);
nand U20716 (N_20716,N_20405,N_20568);
xnor U20717 (N_20717,N_20580,N_20528);
nor U20718 (N_20718,N_20530,N_20594);
xor U20719 (N_20719,N_20569,N_20564);
and U20720 (N_20720,N_20501,N_20570);
nand U20721 (N_20721,N_20423,N_20504);
xnor U20722 (N_20722,N_20438,N_20541);
xor U20723 (N_20723,N_20412,N_20449);
or U20724 (N_20724,N_20434,N_20408);
nand U20725 (N_20725,N_20540,N_20586);
or U20726 (N_20726,N_20434,N_20424);
xnor U20727 (N_20727,N_20437,N_20456);
or U20728 (N_20728,N_20582,N_20481);
xor U20729 (N_20729,N_20481,N_20534);
and U20730 (N_20730,N_20561,N_20457);
or U20731 (N_20731,N_20526,N_20528);
xor U20732 (N_20732,N_20433,N_20465);
and U20733 (N_20733,N_20522,N_20416);
nand U20734 (N_20734,N_20408,N_20489);
xor U20735 (N_20735,N_20598,N_20412);
and U20736 (N_20736,N_20427,N_20584);
nand U20737 (N_20737,N_20432,N_20492);
nand U20738 (N_20738,N_20575,N_20524);
nor U20739 (N_20739,N_20427,N_20411);
nand U20740 (N_20740,N_20414,N_20498);
nand U20741 (N_20741,N_20501,N_20548);
or U20742 (N_20742,N_20465,N_20511);
or U20743 (N_20743,N_20516,N_20547);
and U20744 (N_20744,N_20591,N_20540);
xor U20745 (N_20745,N_20490,N_20506);
nand U20746 (N_20746,N_20575,N_20578);
and U20747 (N_20747,N_20597,N_20460);
xor U20748 (N_20748,N_20461,N_20557);
nor U20749 (N_20749,N_20568,N_20462);
nor U20750 (N_20750,N_20593,N_20402);
and U20751 (N_20751,N_20536,N_20571);
or U20752 (N_20752,N_20566,N_20579);
or U20753 (N_20753,N_20479,N_20548);
nor U20754 (N_20754,N_20538,N_20521);
and U20755 (N_20755,N_20517,N_20430);
xnor U20756 (N_20756,N_20548,N_20409);
or U20757 (N_20757,N_20516,N_20562);
xnor U20758 (N_20758,N_20523,N_20562);
nor U20759 (N_20759,N_20564,N_20538);
nor U20760 (N_20760,N_20428,N_20444);
nor U20761 (N_20761,N_20521,N_20436);
xor U20762 (N_20762,N_20532,N_20582);
or U20763 (N_20763,N_20438,N_20588);
or U20764 (N_20764,N_20446,N_20407);
nor U20765 (N_20765,N_20584,N_20529);
and U20766 (N_20766,N_20400,N_20571);
nor U20767 (N_20767,N_20535,N_20562);
and U20768 (N_20768,N_20553,N_20569);
and U20769 (N_20769,N_20437,N_20541);
and U20770 (N_20770,N_20443,N_20591);
or U20771 (N_20771,N_20405,N_20539);
xnor U20772 (N_20772,N_20449,N_20505);
and U20773 (N_20773,N_20424,N_20594);
xor U20774 (N_20774,N_20437,N_20533);
xor U20775 (N_20775,N_20591,N_20528);
xnor U20776 (N_20776,N_20514,N_20565);
and U20777 (N_20777,N_20481,N_20487);
nand U20778 (N_20778,N_20519,N_20430);
nand U20779 (N_20779,N_20585,N_20420);
or U20780 (N_20780,N_20596,N_20445);
nor U20781 (N_20781,N_20494,N_20496);
nand U20782 (N_20782,N_20436,N_20419);
nand U20783 (N_20783,N_20414,N_20505);
xnor U20784 (N_20784,N_20461,N_20436);
xnor U20785 (N_20785,N_20571,N_20436);
or U20786 (N_20786,N_20522,N_20443);
nor U20787 (N_20787,N_20525,N_20476);
or U20788 (N_20788,N_20453,N_20467);
nor U20789 (N_20789,N_20431,N_20529);
nand U20790 (N_20790,N_20447,N_20575);
nor U20791 (N_20791,N_20506,N_20436);
or U20792 (N_20792,N_20548,N_20449);
nand U20793 (N_20793,N_20473,N_20433);
or U20794 (N_20794,N_20553,N_20482);
nand U20795 (N_20795,N_20529,N_20490);
or U20796 (N_20796,N_20524,N_20580);
nand U20797 (N_20797,N_20583,N_20463);
or U20798 (N_20798,N_20545,N_20407);
nand U20799 (N_20799,N_20473,N_20463);
or U20800 (N_20800,N_20608,N_20710);
nor U20801 (N_20801,N_20735,N_20746);
nor U20802 (N_20802,N_20607,N_20727);
xor U20803 (N_20803,N_20669,N_20634);
or U20804 (N_20804,N_20708,N_20676);
nor U20805 (N_20805,N_20650,N_20754);
and U20806 (N_20806,N_20635,N_20796);
or U20807 (N_20807,N_20700,N_20723);
xor U20808 (N_20808,N_20757,N_20756);
nor U20809 (N_20809,N_20680,N_20719);
xor U20810 (N_20810,N_20609,N_20625);
or U20811 (N_20811,N_20622,N_20616);
xnor U20812 (N_20812,N_20658,N_20656);
xnor U20813 (N_20813,N_20627,N_20771);
nor U20814 (N_20814,N_20679,N_20694);
or U20815 (N_20815,N_20624,N_20672);
xnor U20816 (N_20816,N_20766,N_20661);
nor U20817 (N_20817,N_20762,N_20663);
nand U20818 (N_20818,N_20788,N_20652);
nor U20819 (N_20819,N_20779,N_20678);
xnor U20820 (N_20820,N_20686,N_20732);
and U20821 (N_20821,N_20797,N_20740);
xor U20822 (N_20822,N_20665,N_20759);
and U20823 (N_20823,N_20683,N_20602);
xor U20824 (N_20824,N_20783,N_20610);
xor U20825 (N_20825,N_20701,N_20667);
nor U20826 (N_20826,N_20603,N_20617);
xnor U20827 (N_20827,N_20789,N_20659);
nor U20828 (N_20828,N_20688,N_20739);
and U20829 (N_20829,N_20752,N_20628);
nor U20830 (N_20830,N_20720,N_20767);
xnor U20831 (N_20831,N_20798,N_20631);
and U20832 (N_20832,N_20655,N_20793);
nand U20833 (N_20833,N_20773,N_20716);
nor U20834 (N_20834,N_20641,N_20791);
xor U20835 (N_20835,N_20730,N_20612);
nor U20836 (N_20836,N_20760,N_20785);
xor U20837 (N_20837,N_20722,N_20692);
nand U20838 (N_20838,N_20611,N_20668);
nand U20839 (N_20839,N_20690,N_20753);
and U20840 (N_20840,N_20772,N_20613);
xor U20841 (N_20841,N_20750,N_20705);
nor U20842 (N_20842,N_20733,N_20642);
nor U20843 (N_20843,N_20674,N_20709);
and U20844 (N_20844,N_20726,N_20775);
or U20845 (N_20845,N_20729,N_20712);
or U20846 (N_20846,N_20623,N_20749);
nor U20847 (N_20847,N_20687,N_20604);
xor U20848 (N_20848,N_20620,N_20711);
or U20849 (N_20849,N_20643,N_20691);
xor U20850 (N_20850,N_20713,N_20614);
nor U20851 (N_20851,N_20626,N_20706);
and U20852 (N_20852,N_20799,N_20675);
nor U20853 (N_20853,N_20737,N_20619);
nor U20854 (N_20854,N_20751,N_20654);
nor U20855 (N_20855,N_20644,N_20681);
nor U20856 (N_20856,N_20605,N_20638);
xor U20857 (N_20857,N_20606,N_20744);
nand U20858 (N_20858,N_20671,N_20648);
nor U20859 (N_20859,N_20636,N_20728);
xnor U20860 (N_20860,N_20699,N_20715);
nand U20861 (N_20861,N_20697,N_20782);
nor U20862 (N_20862,N_20755,N_20725);
nand U20863 (N_20863,N_20629,N_20600);
and U20864 (N_20864,N_20704,N_20714);
or U20865 (N_20865,N_20790,N_20693);
and U20866 (N_20866,N_20765,N_20670);
nand U20867 (N_20867,N_20768,N_20738);
nand U20868 (N_20868,N_20657,N_20645);
or U20869 (N_20869,N_20781,N_20776);
or U20870 (N_20870,N_20660,N_20795);
or U20871 (N_20871,N_20721,N_20761);
or U20872 (N_20872,N_20615,N_20794);
nor U20873 (N_20873,N_20786,N_20742);
xor U20874 (N_20874,N_20698,N_20770);
xor U20875 (N_20875,N_20633,N_20780);
and U20876 (N_20876,N_20777,N_20618);
and U20877 (N_20877,N_20649,N_20632);
nand U20878 (N_20878,N_20601,N_20731);
and U20879 (N_20879,N_20741,N_20630);
and U20880 (N_20880,N_20651,N_20664);
nand U20881 (N_20881,N_20666,N_20689);
nor U20882 (N_20882,N_20639,N_20695);
or U20883 (N_20883,N_20763,N_20662);
and U20884 (N_20884,N_20673,N_20646);
and U20885 (N_20885,N_20703,N_20764);
xor U20886 (N_20886,N_20717,N_20736);
nor U20887 (N_20887,N_20734,N_20677);
nand U20888 (N_20888,N_20653,N_20784);
or U20889 (N_20889,N_20640,N_20748);
or U20890 (N_20890,N_20647,N_20707);
xor U20891 (N_20891,N_20774,N_20745);
nor U20892 (N_20892,N_20792,N_20718);
and U20893 (N_20893,N_20724,N_20637);
and U20894 (N_20894,N_20682,N_20743);
or U20895 (N_20895,N_20769,N_20621);
nor U20896 (N_20896,N_20702,N_20778);
xor U20897 (N_20897,N_20758,N_20747);
or U20898 (N_20898,N_20685,N_20684);
or U20899 (N_20899,N_20696,N_20787);
or U20900 (N_20900,N_20791,N_20648);
and U20901 (N_20901,N_20709,N_20740);
nand U20902 (N_20902,N_20719,N_20672);
or U20903 (N_20903,N_20626,N_20611);
or U20904 (N_20904,N_20672,N_20766);
and U20905 (N_20905,N_20612,N_20696);
xor U20906 (N_20906,N_20655,N_20658);
or U20907 (N_20907,N_20728,N_20681);
and U20908 (N_20908,N_20635,N_20708);
and U20909 (N_20909,N_20725,N_20794);
xor U20910 (N_20910,N_20790,N_20797);
nand U20911 (N_20911,N_20634,N_20716);
nor U20912 (N_20912,N_20673,N_20679);
nand U20913 (N_20913,N_20798,N_20789);
nor U20914 (N_20914,N_20635,N_20687);
nand U20915 (N_20915,N_20631,N_20745);
and U20916 (N_20916,N_20763,N_20762);
nand U20917 (N_20917,N_20792,N_20660);
nand U20918 (N_20918,N_20699,N_20689);
or U20919 (N_20919,N_20674,N_20688);
nand U20920 (N_20920,N_20742,N_20618);
nand U20921 (N_20921,N_20682,N_20729);
and U20922 (N_20922,N_20664,N_20716);
nor U20923 (N_20923,N_20642,N_20779);
xor U20924 (N_20924,N_20605,N_20677);
xnor U20925 (N_20925,N_20713,N_20720);
nand U20926 (N_20926,N_20606,N_20708);
nand U20927 (N_20927,N_20667,N_20615);
xnor U20928 (N_20928,N_20764,N_20786);
or U20929 (N_20929,N_20709,N_20774);
nand U20930 (N_20930,N_20685,N_20654);
xor U20931 (N_20931,N_20611,N_20618);
xnor U20932 (N_20932,N_20641,N_20734);
nor U20933 (N_20933,N_20756,N_20696);
and U20934 (N_20934,N_20798,N_20681);
xor U20935 (N_20935,N_20790,N_20642);
or U20936 (N_20936,N_20678,N_20761);
xor U20937 (N_20937,N_20713,N_20745);
and U20938 (N_20938,N_20744,N_20784);
xnor U20939 (N_20939,N_20696,N_20728);
nor U20940 (N_20940,N_20693,N_20681);
xnor U20941 (N_20941,N_20618,N_20769);
nor U20942 (N_20942,N_20716,N_20724);
xor U20943 (N_20943,N_20664,N_20656);
nand U20944 (N_20944,N_20722,N_20654);
xor U20945 (N_20945,N_20738,N_20681);
nor U20946 (N_20946,N_20766,N_20641);
xor U20947 (N_20947,N_20796,N_20797);
or U20948 (N_20948,N_20652,N_20662);
and U20949 (N_20949,N_20670,N_20760);
and U20950 (N_20950,N_20636,N_20666);
xnor U20951 (N_20951,N_20765,N_20668);
and U20952 (N_20952,N_20720,N_20689);
or U20953 (N_20953,N_20792,N_20648);
or U20954 (N_20954,N_20615,N_20641);
nor U20955 (N_20955,N_20685,N_20785);
nor U20956 (N_20956,N_20765,N_20607);
xor U20957 (N_20957,N_20649,N_20700);
and U20958 (N_20958,N_20761,N_20700);
nor U20959 (N_20959,N_20702,N_20674);
nand U20960 (N_20960,N_20603,N_20761);
nor U20961 (N_20961,N_20753,N_20651);
or U20962 (N_20962,N_20658,N_20792);
xnor U20963 (N_20963,N_20774,N_20647);
and U20964 (N_20964,N_20666,N_20650);
nor U20965 (N_20965,N_20637,N_20793);
or U20966 (N_20966,N_20667,N_20732);
nand U20967 (N_20967,N_20776,N_20746);
xor U20968 (N_20968,N_20771,N_20750);
nor U20969 (N_20969,N_20656,N_20610);
nor U20970 (N_20970,N_20735,N_20644);
nand U20971 (N_20971,N_20739,N_20721);
nand U20972 (N_20972,N_20619,N_20719);
or U20973 (N_20973,N_20613,N_20677);
xor U20974 (N_20974,N_20629,N_20753);
or U20975 (N_20975,N_20709,N_20699);
xor U20976 (N_20976,N_20769,N_20719);
or U20977 (N_20977,N_20655,N_20611);
nand U20978 (N_20978,N_20741,N_20617);
or U20979 (N_20979,N_20690,N_20726);
xor U20980 (N_20980,N_20674,N_20794);
xnor U20981 (N_20981,N_20704,N_20685);
and U20982 (N_20982,N_20731,N_20798);
or U20983 (N_20983,N_20643,N_20712);
or U20984 (N_20984,N_20791,N_20741);
xnor U20985 (N_20985,N_20617,N_20682);
nand U20986 (N_20986,N_20674,N_20639);
nand U20987 (N_20987,N_20731,N_20715);
nand U20988 (N_20988,N_20671,N_20767);
xor U20989 (N_20989,N_20708,N_20782);
xnor U20990 (N_20990,N_20793,N_20654);
nor U20991 (N_20991,N_20623,N_20798);
and U20992 (N_20992,N_20791,N_20633);
nand U20993 (N_20993,N_20678,N_20702);
nor U20994 (N_20994,N_20678,N_20732);
and U20995 (N_20995,N_20736,N_20695);
or U20996 (N_20996,N_20700,N_20647);
or U20997 (N_20997,N_20624,N_20788);
or U20998 (N_20998,N_20652,N_20729);
nor U20999 (N_20999,N_20620,N_20605);
nand U21000 (N_21000,N_20918,N_20983);
nand U21001 (N_21001,N_20879,N_20864);
nor U21002 (N_21002,N_20847,N_20826);
or U21003 (N_21003,N_20979,N_20809);
or U21004 (N_21004,N_20891,N_20821);
xor U21005 (N_21005,N_20959,N_20938);
or U21006 (N_21006,N_20876,N_20812);
and U21007 (N_21007,N_20892,N_20869);
xor U21008 (N_21008,N_20805,N_20895);
or U21009 (N_21009,N_20957,N_20946);
and U21010 (N_21010,N_20806,N_20834);
nor U21011 (N_21011,N_20940,N_20923);
and U21012 (N_21012,N_20899,N_20916);
nand U21013 (N_21013,N_20935,N_20913);
nor U21014 (N_21014,N_20872,N_20977);
and U21015 (N_21015,N_20816,N_20883);
and U21016 (N_21016,N_20828,N_20944);
nand U21017 (N_21017,N_20819,N_20971);
nand U21018 (N_21018,N_20817,N_20873);
and U21019 (N_21019,N_20880,N_20852);
nor U21020 (N_21020,N_20956,N_20808);
nand U21021 (N_21021,N_20962,N_20877);
and U21022 (N_21022,N_20931,N_20832);
nor U21023 (N_21023,N_20980,N_20922);
xnor U21024 (N_21024,N_20961,N_20998);
and U21025 (N_21025,N_20903,N_20846);
or U21026 (N_21026,N_20898,N_20861);
xnor U21027 (N_21027,N_20815,N_20978);
or U21028 (N_21028,N_20953,N_20972);
or U21029 (N_21029,N_20937,N_20870);
or U21030 (N_21030,N_20884,N_20822);
and U21031 (N_21031,N_20837,N_20800);
or U21032 (N_21032,N_20988,N_20868);
and U21033 (N_21033,N_20995,N_20894);
nand U21034 (N_21034,N_20936,N_20967);
nand U21035 (N_21035,N_20952,N_20849);
nor U21036 (N_21036,N_20802,N_20838);
nor U21037 (N_21037,N_20811,N_20904);
xor U21038 (N_21038,N_20992,N_20910);
xor U21039 (N_21039,N_20885,N_20964);
nor U21040 (N_21040,N_20911,N_20942);
xor U21041 (N_21041,N_20920,N_20853);
nor U21042 (N_21042,N_20839,N_20878);
nand U21043 (N_21043,N_20865,N_20990);
and U21044 (N_21044,N_20941,N_20824);
and U21045 (N_21045,N_20970,N_20845);
nor U21046 (N_21046,N_20874,N_20930);
nand U21047 (N_21047,N_20890,N_20917);
xor U21048 (N_21048,N_20818,N_20875);
nand U21049 (N_21049,N_20833,N_20893);
and U21050 (N_21050,N_20801,N_20825);
nor U21051 (N_21051,N_20888,N_20897);
and U21052 (N_21052,N_20862,N_20827);
nand U21053 (N_21053,N_20943,N_20919);
or U21054 (N_21054,N_20993,N_20803);
nand U21055 (N_21055,N_20968,N_20973);
and U21056 (N_21056,N_20905,N_20850);
xor U21057 (N_21057,N_20831,N_20969);
nor U21058 (N_21058,N_20863,N_20909);
nand U21059 (N_21059,N_20840,N_20939);
xnor U21060 (N_21060,N_20976,N_20814);
nand U21061 (N_21061,N_20948,N_20912);
nor U21062 (N_21062,N_20928,N_20947);
xnor U21063 (N_21063,N_20966,N_20906);
nor U21064 (N_21064,N_20823,N_20830);
nand U21065 (N_21065,N_20857,N_20926);
or U21066 (N_21066,N_20807,N_20933);
and U21067 (N_21067,N_20951,N_20813);
xnor U21068 (N_21068,N_20982,N_20934);
nand U21069 (N_21069,N_20915,N_20986);
and U21070 (N_21070,N_20908,N_20820);
or U21071 (N_21071,N_20987,N_20924);
nor U21072 (N_21072,N_20871,N_20975);
or U21073 (N_21073,N_20925,N_20954);
and U21074 (N_21074,N_20997,N_20914);
nor U21075 (N_21075,N_20985,N_20949);
xor U21076 (N_21076,N_20851,N_20929);
nor U21077 (N_21077,N_20881,N_20841);
nand U21078 (N_21078,N_20984,N_20927);
or U21079 (N_21079,N_20945,N_20974);
nand U21080 (N_21080,N_20842,N_20994);
or U21081 (N_21081,N_20867,N_20889);
nor U21082 (N_21082,N_20960,N_20859);
nand U21083 (N_21083,N_20950,N_20963);
and U21084 (N_21084,N_20902,N_20989);
or U21085 (N_21085,N_20901,N_20844);
or U21086 (N_21086,N_20804,N_20810);
and U21087 (N_21087,N_20958,N_20932);
nand U21088 (N_21088,N_20981,N_20860);
nor U21089 (N_21089,N_20999,N_20887);
and U21090 (N_21090,N_20996,N_20886);
and U21091 (N_21091,N_20836,N_20896);
and U21092 (N_21092,N_20955,N_20855);
xor U21093 (N_21093,N_20843,N_20991);
nor U21094 (N_21094,N_20856,N_20854);
or U21095 (N_21095,N_20829,N_20882);
and U21096 (N_21096,N_20921,N_20835);
nor U21097 (N_21097,N_20907,N_20965);
nand U21098 (N_21098,N_20858,N_20866);
and U21099 (N_21099,N_20848,N_20900);
or U21100 (N_21100,N_20855,N_20820);
xor U21101 (N_21101,N_20971,N_20966);
nor U21102 (N_21102,N_20947,N_20922);
and U21103 (N_21103,N_20823,N_20816);
nand U21104 (N_21104,N_20947,N_20887);
and U21105 (N_21105,N_20880,N_20825);
xnor U21106 (N_21106,N_20927,N_20875);
xor U21107 (N_21107,N_20880,N_20911);
nor U21108 (N_21108,N_20822,N_20928);
and U21109 (N_21109,N_20947,N_20905);
nor U21110 (N_21110,N_20898,N_20819);
nor U21111 (N_21111,N_20892,N_20879);
or U21112 (N_21112,N_20926,N_20891);
and U21113 (N_21113,N_20931,N_20864);
nor U21114 (N_21114,N_20991,N_20999);
and U21115 (N_21115,N_20814,N_20945);
or U21116 (N_21116,N_20843,N_20926);
xor U21117 (N_21117,N_20811,N_20986);
nand U21118 (N_21118,N_20981,N_20811);
nand U21119 (N_21119,N_20823,N_20988);
xnor U21120 (N_21120,N_20860,N_20934);
nand U21121 (N_21121,N_20883,N_20931);
and U21122 (N_21122,N_20836,N_20983);
nand U21123 (N_21123,N_20901,N_20838);
or U21124 (N_21124,N_20979,N_20823);
or U21125 (N_21125,N_20962,N_20956);
or U21126 (N_21126,N_20980,N_20900);
nand U21127 (N_21127,N_20911,N_20876);
nor U21128 (N_21128,N_20887,N_20917);
or U21129 (N_21129,N_20951,N_20944);
nand U21130 (N_21130,N_20932,N_20829);
xnor U21131 (N_21131,N_20860,N_20918);
nand U21132 (N_21132,N_20942,N_20885);
nor U21133 (N_21133,N_20921,N_20936);
nand U21134 (N_21134,N_20842,N_20857);
xnor U21135 (N_21135,N_20882,N_20879);
nor U21136 (N_21136,N_20882,N_20810);
and U21137 (N_21137,N_20895,N_20980);
nor U21138 (N_21138,N_20951,N_20843);
or U21139 (N_21139,N_20931,N_20888);
nand U21140 (N_21140,N_20860,N_20958);
xor U21141 (N_21141,N_20986,N_20963);
or U21142 (N_21142,N_20849,N_20818);
xnor U21143 (N_21143,N_20832,N_20983);
or U21144 (N_21144,N_20970,N_20815);
or U21145 (N_21145,N_20815,N_20871);
and U21146 (N_21146,N_20882,N_20940);
nand U21147 (N_21147,N_20838,N_20813);
nand U21148 (N_21148,N_20902,N_20880);
xor U21149 (N_21149,N_20861,N_20812);
nor U21150 (N_21150,N_20826,N_20944);
and U21151 (N_21151,N_20851,N_20868);
nor U21152 (N_21152,N_20810,N_20985);
and U21153 (N_21153,N_20940,N_20970);
xnor U21154 (N_21154,N_20819,N_20991);
nand U21155 (N_21155,N_20925,N_20870);
nand U21156 (N_21156,N_20809,N_20968);
nand U21157 (N_21157,N_20863,N_20859);
or U21158 (N_21158,N_20941,N_20946);
or U21159 (N_21159,N_20812,N_20810);
xor U21160 (N_21160,N_20955,N_20876);
xor U21161 (N_21161,N_20960,N_20956);
xnor U21162 (N_21162,N_20898,N_20904);
nor U21163 (N_21163,N_20882,N_20852);
or U21164 (N_21164,N_20851,N_20847);
or U21165 (N_21165,N_20866,N_20842);
or U21166 (N_21166,N_20825,N_20853);
nand U21167 (N_21167,N_20910,N_20933);
nor U21168 (N_21168,N_20841,N_20958);
nand U21169 (N_21169,N_20886,N_20987);
and U21170 (N_21170,N_20911,N_20841);
nand U21171 (N_21171,N_20822,N_20929);
or U21172 (N_21172,N_20807,N_20913);
or U21173 (N_21173,N_20826,N_20974);
xnor U21174 (N_21174,N_20847,N_20802);
and U21175 (N_21175,N_20926,N_20884);
nor U21176 (N_21176,N_20865,N_20826);
xor U21177 (N_21177,N_20931,N_20910);
nand U21178 (N_21178,N_20945,N_20881);
nand U21179 (N_21179,N_20934,N_20845);
xnor U21180 (N_21180,N_20898,N_20838);
or U21181 (N_21181,N_20939,N_20964);
nand U21182 (N_21182,N_20838,N_20923);
or U21183 (N_21183,N_20907,N_20978);
xor U21184 (N_21184,N_20998,N_20814);
and U21185 (N_21185,N_20893,N_20862);
nor U21186 (N_21186,N_20816,N_20930);
xnor U21187 (N_21187,N_20945,N_20967);
nand U21188 (N_21188,N_20898,N_20962);
and U21189 (N_21189,N_20875,N_20861);
or U21190 (N_21190,N_20966,N_20941);
nor U21191 (N_21191,N_20840,N_20921);
or U21192 (N_21192,N_20801,N_20805);
nor U21193 (N_21193,N_20871,N_20918);
xor U21194 (N_21194,N_20860,N_20887);
xor U21195 (N_21195,N_20865,N_20846);
nor U21196 (N_21196,N_20949,N_20962);
nor U21197 (N_21197,N_20823,N_20885);
xor U21198 (N_21198,N_20803,N_20928);
nand U21199 (N_21199,N_20919,N_20910);
and U21200 (N_21200,N_21109,N_21145);
xnor U21201 (N_21201,N_21042,N_21192);
nand U21202 (N_21202,N_21060,N_21130);
nor U21203 (N_21203,N_21059,N_21196);
nor U21204 (N_21204,N_21053,N_21088);
nor U21205 (N_21205,N_21076,N_21129);
nor U21206 (N_21206,N_21022,N_21010);
or U21207 (N_21207,N_21075,N_21057);
nor U21208 (N_21208,N_21032,N_21152);
or U21209 (N_21209,N_21068,N_21143);
xor U21210 (N_21210,N_21101,N_21081);
nand U21211 (N_21211,N_21029,N_21124);
or U21212 (N_21212,N_21020,N_21183);
nor U21213 (N_21213,N_21052,N_21110);
xnor U21214 (N_21214,N_21014,N_21131);
or U21215 (N_21215,N_21197,N_21128);
or U21216 (N_21216,N_21037,N_21190);
nand U21217 (N_21217,N_21054,N_21096);
and U21218 (N_21218,N_21033,N_21000);
and U21219 (N_21219,N_21030,N_21168);
nand U21220 (N_21220,N_21174,N_21084);
or U21221 (N_21221,N_21046,N_21195);
nor U21222 (N_21222,N_21074,N_21178);
nand U21223 (N_21223,N_21017,N_21015);
nand U21224 (N_21224,N_21065,N_21188);
or U21225 (N_21225,N_21148,N_21171);
and U21226 (N_21226,N_21159,N_21136);
or U21227 (N_21227,N_21077,N_21189);
nor U21228 (N_21228,N_21001,N_21113);
xnor U21229 (N_21229,N_21169,N_21062);
xor U21230 (N_21230,N_21125,N_21123);
and U21231 (N_21231,N_21170,N_21064);
and U21232 (N_21232,N_21103,N_21194);
nor U21233 (N_21233,N_21126,N_21121);
xor U21234 (N_21234,N_21066,N_21086);
xor U21235 (N_21235,N_21167,N_21161);
nor U21236 (N_21236,N_21082,N_21024);
and U21237 (N_21237,N_21120,N_21091);
nor U21238 (N_21238,N_21184,N_21118);
or U21239 (N_21239,N_21186,N_21108);
and U21240 (N_21240,N_21044,N_21045);
xor U21241 (N_21241,N_21172,N_21034);
and U21242 (N_21242,N_21149,N_21027);
xor U21243 (N_21243,N_21122,N_21102);
nor U21244 (N_21244,N_21049,N_21061);
and U21245 (N_21245,N_21105,N_21090);
nor U21246 (N_21246,N_21011,N_21089);
nand U21247 (N_21247,N_21016,N_21026);
nor U21248 (N_21248,N_21154,N_21008);
xor U21249 (N_21249,N_21115,N_21173);
and U21250 (N_21250,N_21160,N_21112);
nand U21251 (N_21251,N_21006,N_21127);
nor U21252 (N_21252,N_21163,N_21165);
or U21253 (N_21253,N_21083,N_21185);
xor U21254 (N_21254,N_21147,N_21144);
xor U21255 (N_21255,N_21085,N_21141);
nand U21256 (N_21256,N_21080,N_21119);
nand U21257 (N_21257,N_21158,N_21176);
nor U21258 (N_21258,N_21116,N_21199);
nand U21259 (N_21259,N_21013,N_21098);
and U21260 (N_21260,N_21028,N_21050);
nor U21261 (N_21261,N_21092,N_21069);
and U21262 (N_21262,N_21151,N_21004);
and U21263 (N_21263,N_21100,N_21164);
nor U21264 (N_21264,N_21155,N_21031);
nor U21265 (N_21265,N_21019,N_21140);
and U21266 (N_21266,N_21198,N_21104);
nand U21267 (N_21267,N_21079,N_21135);
xor U21268 (N_21268,N_21157,N_21003);
or U21269 (N_21269,N_21041,N_21039);
xor U21270 (N_21270,N_21095,N_21078);
nand U21271 (N_21271,N_21012,N_21021);
or U21272 (N_21272,N_21132,N_21073);
xnor U21273 (N_21273,N_21099,N_21025);
or U21274 (N_21274,N_21181,N_21179);
or U21275 (N_21275,N_21009,N_21051);
or U21276 (N_21276,N_21002,N_21153);
nand U21277 (N_21277,N_21187,N_21007);
xor U21278 (N_21278,N_21139,N_21166);
xnor U21279 (N_21279,N_21036,N_21106);
nor U21280 (N_21280,N_21114,N_21177);
nor U21281 (N_21281,N_21055,N_21087);
xor U21282 (N_21282,N_21134,N_21005);
xor U21283 (N_21283,N_21047,N_21142);
and U21284 (N_21284,N_21117,N_21094);
and U21285 (N_21285,N_21111,N_21156);
or U21286 (N_21286,N_21058,N_21018);
xnor U21287 (N_21287,N_21067,N_21038);
and U21288 (N_21288,N_21150,N_21191);
and U21289 (N_21289,N_21048,N_21193);
nor U21290 (N_21290,N_21138,N_21072);
and U21291 (N_21291,N_21133,N_21093);
nor U21292 (N_21292,N_21097,N_21063);
xnor U21293 (N_21293,N_21040,N_21137);
xor U21294 (N_21294,N_21023,N_21180);
xnor U21295 (N_21295,N_21056,N_21070);
xnor U21296 (N_21296,N_21162,N_21146);
nor U21297 (N_21297,N_21175,N_21043);
and U21298 (N_21298,N_21182,N_21071);
or U21299 (N_21299,N_21107,N_21035);
nand U21300 (N_21300,N_21050,N_21176);
nor U21301 (N_21301,N_21171,N_21046);
nor U21302 (N_21302,N_21136,N_21009);
and U21303 (N_21303,N_21151,N_21176);
nor U21304 (N_21304,N_21038,N_21044);
and U21305 (N_21305,N_21036,N_21074);
nand U21306 (N_21306,N_21036,N_21188);
and U21307 (N_21307,N_21157,N_21042);
or U21308 (N_21308,N_21180,N_21132);
xor U21309 (N_21309,N_21185,N_21154);
nand U21310 (N_21310,N_21128,N_21150);
or U21311 (N_21311,N_21128,N_21007);
xor U21312 (N_21312,N_21026,N_21130);
or U21313 (N_21313,N_21141,N_21042);
nor U21314 (N_21314,N_21005,N_21118);
nand U21315 (N_21315,N_21102,N_21094);
nor U21316 (N_21316,N_21117,N_21198);
xnor U21317 (N_21317,N_21087,N_21108);
xor U21318 (N_21318,N_21078,N_21000);
nor U21319 (N_21319,N_21137,N_21084);
and U21320 (N_21320,N_21160,N_21170);
and U21321 (N_21321,N_21024,N_21093);
or U21322 (N_21322,N_21083,N_21022);
nand U21323 (N_21323,N_21199,N_21118);
nor U21324 (N_21324,N_21016,N_21021);
nand U21325 (N_21325,N_21075,N_21024);
or U21326 (N_21326,N_21018,N_21099);
or U21327 (N_21327,N_21080,N_21016);
and U21328 (N_21328,N_21096,N_21124);
nor U21329 (N_21329,N_21145,N_21113);
nand U21330 (N_21330,N_21142,N_21090);
and U21331 (N_21331,N_21075,N_21145);
xor U21332 (N_21332,N_21130,N_21095);
nor U21333 (N_21333,N_21139,N_21098);
or U21334 (N_21334,N_21038,N_21085);
or U21335 (N_21335,N_21070,N_21064);
and U21336 (N_21336,N_21124,N_21188);
xor U21337 (N_21337,N_21089,N_21021);
and U21338 (N_21338,N_21001,N_21003);
or U21339 (N_21339,N_21104,N_21052);
nand U21340 (N_21340,N_21001,N_21162);
xnor U21341 (N_21341,N_21158,N_21005);
nor U21342 (N_21342,N_21169,N_21142);
xor U21343 (N_21343,N_21066,N_21148);
xnor U21344 (N_21344,N_21068,N_21161);
xor U21345 (N_21345,N_21078,N_21117);
nand U21346 (N_21346,N_21079,N_21033);
nor U21347 (N_21347,N_21053,N_21080);
and U21348 (N_21348,N_21162,N_21000);
nor U21349 (N_21349,N_21015,N_21188);
nor U21350 (N_21350,N_21151,N_21059);
xor U21351 (N_21351,N_21192,N_21029);
xnor U21352 (N_21352,N_21087,N_21123);
nor U21353 (N_21353,N_21186,N_21120);
xor U21354 (N_21354,N_21055,N_21150);
and U21355 (N_21355,N_21177,N_21047);
xnor U21356 (N_21356,N_21054,N_21052);
and U21357 (N_21357,N_21034,N_21173);
or U21358 (N_21358,N_21191,N_21140);
xnor U21359 (N_21359,N_21192,N_21085);
xnor U21360 (N_21360,N_21115,N_21092);
and U21361 (N_21361,N_21162,N_21188);
or U21362 (N_21362,N_21167,N_21184);
xor U21363 (N_21363,N_21129,N_21188);
and U21364 (N_21364,N_21078,N_21086);
and U21365 (N_21365,N_21109,N_21045);
xnor U21366 (N_21366,N_21031,N_21049);
or U21367 (N_21367,N_21061,N_21092);
and U21368 (N_21368,N_21065,N_21145);
nand U21369 (N_21369,N_21152,N_21023);
or U21370 (N_21370,N_21096,N_21007);
or U21371 (N_21371,N_21176,N_21106);
and U21372 (N_21372,N_21128,N_21158);
xor U21373 (N_21373,N_21090,N_21016);
nor U21374 (N_21374,N_21096,N_21088);
and U21375 (N_21375,N_21145,N_21115);
xnor U21376 (N_21376,N_21196,N_21056);
and U21377 (N_21377,N_21067,N_21177);
nor U21378 (N_21378,N_21017,N_21186);
nand U21379 (N_21379,N_21145,N_21077);
nand U21380 (N_21380,N_21066,N_21033);
and U21381 (N_21381,N_21065,N_21047);
and U21382 (N_21382,N_21024,N_21108);
nor U21383 (N_21383,N_21160,N_21182);
or U21384 (N_21384,N_21189,N_21043);
nand U21385 (N_21385,N_21091,N_21198);
nand U21386 (N_21386,N_21187,N_21148);
xor U21387 (N_21387,N_21168,N_21094);
and U21388 (N_21388,N_21141,N_21108);
nand U21389 (N_21389,N_21070,N_21046);
nand U21390 (N_21390,N_21139,N_21125);
and U21391 (N_21391,N_21187,N_21135);
xor U21392 (N_21392,N_21151,N_21125);
or U21393 (N_21393,N_21158,N_21056);
xor U21394 (N_21394,N_21171,N_21047);
nand U21395 (N_21395,N_21191,N_21018);
and U21396 (N_21396,N_21062,N_21162);
or U21397 (N_21397,N_21005,N_21117);
and U21398 (N_21398,N_21026,N_21127);
or U21399 (N_21399,N_21190,N_21031);
nor U21400 (N_21400,N_21387,N_21327);
nor U21401 (N_21401,N_21250,N_21335);
nand U21402 (N_21402,N_21221,N_21396);
nor U21403 (N_21403,N_21201,N_21290);
or U21404 (N_21404,N_21299,N_21237);
xor U21405 (N_21405,N_21224,N_21369);
nor U21406 (N_21406,N_21256,N_21200);
or U21407 (N_21407,N_21296,N_21278);
and U21408 (N_21408,N_21304,N_21264);
xor U21409 (N_21409,N_21223,N_21323);
or U21410 (N_21410,N_21385,N_21381);
and U21411 (N_21411,N_21388,N_21332);
xor U21412 (N_21412,N_21258,N_21271);
xnor U21413 (N_21413,N_21222,N_21282);
xnor U21414 (N_21414,N_21345,N_21215);
and U21415 (N_21415,N_21365,N_21378);
nand U21416 (N_21416,N_21265,N_21230);
xnor U21417 (N_21417,N_21349,N_21359);
xor U21418 (N_21418,N_21247,N_21231);
and U21419 (N_21419,N_21389,N_21269);
nor U21420 (N_21420,N_21322,N_21251);
xnor U21421 (N_21421,N_21288,N_21339);
or U21422 (N_21422,N_21308,N_21391);
xnor U21423 (N_21423,N_21203,N_21210);
nand U21424 (N_21424,N_21228,N_21226);
nand U21425 (N_21425,N_21319,N_21291);
and U21426 (N_21426,N_21374,N_21285);
nor U21427 (N_21427,N_21246,N_21316);
nor U21428 (N_21428,N_21314,N_21384);
and U21429 (N_21429,N_21367,N_21326);
or U21430 (N_21430,N_21350,N_21392);
or U21431 (N_21431,N_21356,N_21383);
and U21432 (N_21432,N_21390,N_21205);
or U21433 (N_21433,N_21270,N_21206);
or U21434 (N_21434,N_21273,N_21238);
nand U21435 (N_21435,N_21245,N_21208);
xnor U21436 (N_21436,N_21253,N_21357);
nor U21437 (N_21437,N_21329,N_21343);
or U21438 (N_21438,N_21204,N_21397);
nand U21439 (N_21439,N_21300,N_21373);
nand U21440 (N_21440,N_21364,N_21235);
or U21441 (N_21441,N_21393,N_21334);
xor U21442 (N_21442,N_21311,N_21340);
nor U21443 (N_21443,N_21274,N_21375);
or U21444 (N_21444,N_21307,N_21280);
or U21445 (N_21445,N_21252,N_21337);
nor U21446 (N_21446,N_21244,N_21289);
xor U21447 (N_21447,N_21255,N_21302);
nor U21448 (N_21448,N_21347,N_21233);
xnor U21449 (N_21449,N_21298,N_21262);
and U21450 (N_21450,N_21361,N_21348);
xnor U21451 (N_21451,N_21313,N_21360);
nor U21452 (N_21452,N_21261,N_21241);
nand U21453 (N_21453,N_21254,N_21212);
xor U21454 (N_21454,N_21305,N_21225);
and U21455 (N_21455,N_21320,N_21234);
or U21456 (N_21456,N_21263,N_21351);
and U21457 (N_21457,N_21287,N_21376);
nand U21458 (N_21458,N_21277,N_21295);
and U21459 (N_21459,N_21260,N_21395);
xnor U21460 (N_21460,N_21294,N_21292);
or U21461 (N_21461,N_21317,N_21267);
nand U21462 (N_21462,N_21276,N_21324);
xor U21463 (N_21463,N_21342,N_21368);
xnor U21464 (N_21464,N_21398,N_21211);
nand U21465 (N_21465,N_21249,N_21257);
or U21466 (N_21466,N_21362,N_21352);
and U21467 (N_21467,N_21399,N_21240);
nor U21468 (N_21468,N_21213,N_21232);
nand U21469 (N_21469,N_21363,N_21328);
or U21470 (N_21470,N_21318,N_21386);
nor U21471 (N_21471,N_21293,N_21279);
and U21472 (N_21472,N_21220,N_21217);
or U21473 (N_21473,N_21333,N_21312);
or U21474 (N_21474,N_21394,N_21214);
xor U21475 (N_21475,N_21336,N_21382);
nor U21476 (N_21476,N_21239,N_21236);
xnor U21477 (N_21477,N_21297,N_21321);
and U21478 (N_21478,N_21366,N_21202);
xnor U21479 (N_21479,N_21330,N_21243);
xnor U21480 (N_21480,N_21331,N_21283);
nand U21481 (N_21481,N_21353,N_21281);
or U21482 (N_21482,N_21227,N_21218);
nor U21483 (N_21483,N_21370,N_21341);
xnor U21484 (N_21484,N_21266,N_21209);
nand U21485 (N_21485,N_21242,N_21207);
and U21486 (N_21486,N_21301,N_21344);
xor U21487 (N_21487,N_21372,N_21219);
nor U21488 (N_21488,N_21229,N_21358);
and U21489 (N_21489,N_21315,N_21371);
xor U21490 (N_21490,N_21377,N_21325);
nand U21491 (N_21491,N_21380,N_21354);
nand U21492 (N_21492,N_21268,N_21216);
and U21493 (N_21493,N_21309,N_21338);
xor U21494 (N_21494,N_21310,N_21284);
nor U21495 (N_21495,N_21303,N_21259);
nor U21496 (N_21496,N_21346,N_21306);
nor U21497 (N_21497,N_21272,N_21379);
or U21498 (N_21498,N_21355,N_21248);
and U21499 (N_21499,N_21275,N_21286);
nand U21500 (N_21500,N_21231,N_21202);
or U21501 (N_21501,N_21313,N_21207);
nand U21502 (N_21502,N_21213,N_21231);
and U21503 (N_21503,N_21274,N_21357);
nor U21504 (N_21504,N_21204,N_21252);
and U21505 (N_21505,N_21395,N_21236);
and U21506 (N_21506,N_21287,N_21375);
nor U21507 (N_21507,N_21257,N_21359);
and U21508 (N_21508,N_21208,N_21364);
nor U21509 (N_21509,N_21394,N_21212);
xnor U21510 (N_21510,N_21279,N_21218);
nor U21511 (N_21511,N_21382,N_21366);
or U21512 (N_21512,N_21277,N_21286);
nand U21513 (N_21513,N_21384,N_21313);
and U21514 (N_21514,N_21241,N_21214);
xnor U21515 (N_21515,N_21375,N_21300);
xnor U21516 (N_21516,N_21353,N_21330);
xnor U21517 (N_21517,N_21328,N_21305);
xor U21518 (N_21518,N_21306,N_21364);
nor U21519 (N_21519,N_21386,N_21274);
xnor U21520 (N_21520,N_21232,N_21305);
nand U21521 (N_21521,N_21217,N_21377);
xnor U21522 (N_21522,N_21306,N_21319);
xor U21523 (N_21523,N_21315,N_21370);
nor U21524 (N_21524,N_21270,N_21220);
or U21525 (N_21525,N_21347,N_21385);
nor U21526 (N_21526,N_21358,N_21278);
xnor U21527 (N_21527,N_21374,N_21329);
nor U21528 (N_21528,N_21303,N_21252);
nor U21529 (N_21529,N_21239,N_21209);
nand U21530 (N_21530,N_21209,N_21201);
or U21531 (N_21531,N_21302,N_21259);
xor U21532 (N_21532,N_21219,N_21258);
and U21533 (N_21533,N_21235,N_21333);
nand U21534 (N_21534,N_21359,N_21392);
nand U21535 (N_21535,N_21280,N_21359);
nand U21536 (N_21536,N_21263,N_21291);
nor U21537 (N_21537,N_21343,N_21390);
nor U21538 (N_21538,N_21349,N_21303);
xnor U21539 (N_21539,N_21215,N_21362);
or U21540 (N_21540,N_21324,N_21217);
xnor U21541 (N_21541,N_21358,N_21269);
nand U21542 (N_21542,N_21214,N_21396);
and U21543 (N_21543,N_21379,N_21372);
nor U21544 (N_21544,N_21203,N_21243);
or U21545 (N_21545,N_21229,N_21369);
and U21546 (N_21546,N_21358,N_21225);
xor U21547 (N_21547,N_21255,N_21286);
nor U21548 (N_21548,N_21384,N_21316);
or U21549 (N_21549,N_21345,N_21232);
nor U21550 (N_21550,N_21201,N_21234);
and U21551 (N_21551,N_21387,N_21352);
or U21552 (N_21552,N_21249,N_21308);
xnor U21553 (N_21553,N_21355,N_21321);
xor U21554 (N_21554,N_21214,N_21311);
xor U21555 (N_21555,N_21399,N_21315);
and U21556 (N_21556,N_21313,N_21369);
nor U21557 (N_21557,N_21330,N_21203);
xor U21558 (N_21558,N_21353,N_21219);
or U21559 (N_21559,N_21320,N_21291);
xor U21560 (N_21560,N_21252,N_21308);
nor U21561 (N_21561,N_21371,N_21386);
and U21562 (N_21562,N_21295,N_21320);
nand U21563 (N_21563,N_21380,N_21255);
nor U21564 (N_21564,N_21309,N_21325);
and U21565 (N_21565,N_21299,N_21339);
nor U21566 (N_21566,N_21243,N_21300);
nor U21567 (N_21567,N_21319,N_21267);
xor U21568 (N_21568,N_21390,N_21260);
xor U21569 (N_21569,N_21304,N_21203);
nand U21570 (N_21570,N_21233,N_21294);
nor U21571 (N_21571,N_21231,N_21300);
and U21572 (N_21572,N_21205,N_21248);
or U21573 (N_21573,N_21203,N_21363);
or U21574 (N_21574,N_21282,N_21315);
and U21575 (N_21575,N_21343,N_21276);
nand U21576 (N_21576,N_21205,N_21218);
and U21577 (N_21577,N_21396,N_21338);
nor U21578 (N_21578,N_21324,N_21245);
or U21579 (N_21579,N_21282,N_21340);
nor U21580 (N_21580,N_21336,N_21221);
and U21581 (N_21581,N_21387,N_21292);
and U21582 (N_21582,N_21280,N_21254);
or U21583 (N_21583,N_21284,N_21389);
or U21584 (N_21584,N_21325,N_21316);
and U21585 (N_21585,N_21355,N_21220);
and U21586 (N_21586,N_21204,N_21386);
or U21587 (N_21587,N_21340,N_21209);
nand U21588 (N_21588,N_21374,N_21247);
nand U21589 (N_21589,N_21251,N_21362);
xnor U21590 (N_21590,N_21330,N_21261);
and U21591 (N_21591,N_21317,N_21345);
and U21592 (N_21592,N_21248,N_21341);
xor U21593 (N_21593,N_21339,N_21216);
nand U21594 (N_21594,N_21326,N_21228);
and U21595 (N_21595,N_21352,N_21203);
nand U21596 (N_21596,N_21358,N_21393);
and U21597 (N_21597,N_21216,N_21307);
or U21598 (N_21598,N_21350,N_21332);
nand U21599 (N_21599,N_21310,N_21303);
nand U21600 (N_21600,N_21423,N_21536);
and U21601 (N_21601,N_21528,N_21428);
nor U21602 (N_21602,N_21509,N_21417);
nor U21603 (N_21603,N_21500,N_21596);
nor U21604 (N_21604,N_21510,N_21525);
nand U21605 (N_21605,N_21405,N_21544);
xor U21606 (N_21606,N_21461,N_21518);
nand U21607 (N_21607,N_21446,N_21571);
and U21608 (N_21608,N_21460,N_21492);
or U21609 (N_21609,N_21523,N_21439);
or U21610 (N_21610,N_21478,N_21447);
xnor U21611 (N_21611,N_21463,N_21402);
nor U21612 (N_21612,N_21441,N_21508);
or U21613 (N_21613,N_21498,N_21579);
xor U21614 (N_21614,N_21457,N_21467);
nor U21615 (N_21615,N_21416,N_21554);
nand U21616 (N_21616,N_21487,N_21502);
nand U21617 (N_21617,N_21421,N_21479);
and U21618 (N_21618,N_21535,N_21513);
nor U21619 (N_21619,N_21520,N_21584);
nand U21620 (N_21620,N_21491,N_21592);
nand U21621 (N_21621,N_21472,N_21533);
nand U21622 (N_21622,N_21473,N_21433);
nor U21623 (N_21623,N_21561,N_21497);
xnor U21624 (N_21624,N_21567,N_21407);
nor U21625 (N_21625,N_21517,N_21477);
xnor U21626 (N_21626,N_21426,N_21539);
or U21627 (N_21627,N_21432,N_21540);
and U21628 (N_21628,N_21551,N_21411);
or U21629 (N_21629,N_21566,N_21522);
and U21630 (N_21630,N_21506,N_21548);
and U21631 (N_21631,N_21430,N_21591);
nor U21632 (N_21632,N_21466,N_21484);
or U21633 (N_21633,N_21422,N_21414);
and U21634 (N_21634,N_21598,N_21437);
and U21635 (N_21635,N_21589,N_21475);
nor U21636 (N_21636,N_21489,N_21538);
or U21637 (N_21637,N_21436,N_21568);
or U21638 (N_21638,N_21454,N_21524);
nor U21639 (N_21639,N_21582,N_21450);
or U21640 (N_21640,N_21403,N_21578);
or U21641 (N_21641,N_21532,N_21575);
nor U21642 (N_21642,N_21462,N_21546);
xor U21643 (N_21643,N_21458,N_21521);
or U21644 (N_21644,N_21552,N_21438);
xnor U21645 (N_21645,N_21440,N_21583);
or U21646 (N_21646,N_21507,N_21541);
and U21647 (N_21647,N_21553,N_21425);
xnor U21648 (N_21648,N_21549,N_21413);
and U21649 (N_21649,N_21499,N_21581);
nand U21650 (N_21650,N_21471,N_21444);
nor U21651 (N_21651,N_21435,N_21555);
xnor U21652 (N_21652,N_21599,N_21486);
or U21653 (N_21653,N_21573,N_21415);
nand U21654 (N_21654,N_21563,N_21576);
xor U21655 (N_21655,N_21419,N_21404);
and U21656 (N_21656,N_21545,N_21455);
nor U21657 (N_21657,N_21501,N_21514);
and U21658 (N_21658,N_21588,N_21485);
nor U21659 (N_21659,N_21559,N_21556);
nand U21660 (N_21660,N_21429,N_21483);
nand U21661 (N_21661,N_21470,N_21488);
or U21662 (N_21662,N_21468,N_21400);
or U21663 (N_21663,N_21476,N_21512);
xor U21664 (N_21664,N_21469,N_21543);
and U21665 (N_21665,N_21442,N_21481);
xnor U21666 (N_21666,N_21443,N_21504);
and U21667 (N_21667,N_21595,N_21557);
nor U21668 (N_21668,N_21562,N_21503);
or U21669 (N_21669,N_21505,N_21564);
nor U21670 (N_21670,N_21570,N_21482);
nand U21671 (N_21671,N_21409,N_21531);
and U21672 (N_21672,N_21445,N_21586);
xnor U21673 (N_21673,N_21537,N_21495);
and U21674 (N_21674,N_21560,N_21448);
or U21675 (N_21675,N_21527,N_21465);
or U21676 (N_21676,N_21585,N_21452);
or U21677 (N_21677,N_21569,N_21558);
or U21678 (N_21678,N_21511,N_21519);
nand U21679 (N_21679,N_21594,N_21453);
nor U21680 (N_21680,N_21449,N_21529);
nor U21681 (N_21681,N_21565,N_21516);
xor U21682 (N_21682,N_21590,N_21412);
nor U21683 (N_21683,N_21572,N_21401);
nand U21684 (N_21684,N_21526,N_21464);
nor U21685 (N_21685,N_21456,N_21547);
nand U21686 (N_21686,N_21593,N_21577);
and U21687 (N_21687,N_21550,N_21480);
xnor U21688 (N_21688,N_21427,N_21597);
nand U21689 (N_21689,N_21493,N_21451);
nor U21690 (N_21690,N_21418,N_21542);
xor U21691 (N_21691,N_21494,N_21406);
or U21692 (N_21692,N_21434,N_21530);
nor U21693 (N_21693,N_21420,N_21459);
nor U21694 (N_21694,N_21515,N_21534);
nand U21695 (N_21695,N_21490,N_21474);
and U21696 (N_21696,N_21574,N_21408);
or U21697 (N_21697,N_21424,N_21580);
nor U21698 (N_21698,N_21431,N_21410);
nor U21699 (N_21699,N_21587,N_21496);
nor U21700 (N_21700,N_21568,N_21423);
nor U21701 (N_21701,N_21548,N_21521);
or U21702 (N_21702,N_21490,N_21536);
and U21703 (N_21703,N_21573,N_21409);
or U21704 (N_21704,N_21465,N_21509);
nor U21705 (N_21705,N_21529,N_21504);
nand U21706 (N_21706,N_21427,N_21522);
xnor U21707 (N_21707,N_21408,N_21462);
nand U21708 (N_21708,N_21432,N_21501);
xnor U21709 (N_21709,N_21519,N_21487);
or U21710 (N_21710,N_21560,N_21480);
xnor U21711 (N_21711,N_21451,N_21477);
nand U21712 (N_21712,N_21524,N_21519);
or U21713 (N_21713,N_21431,N_21552);
nand U21714 (N_21714,N_21578,N_21526);
or U21715 (N_21715,N_21542,N_21539);
nor U21716 (N_21716,N_21504,N_21413);
and U21717 (N_21717,N_21417,N_21457);
or U21718 (N_21718,N_21557,N_21596);
xor U21719 (N_21719,N_21467,N_21406);
nor U21720 (N_21720,N_21466,N_21535);
xor U21721 (N_21721,N_21559,N_21466);
nor U21722 (N_21722,N_21561,N_21526);
and U21723 (N_21723,N_21547,N_21561);
nor U21724 (N_21724,N_21464,N_21436);
nand U21725 (N_21725,N_21590,N_21595);
nand U21726 (N_21726,N_21524,N_21404);
xor U21727 (N_21727,N_21484,N_21495);
and U21728 (N_21728,N_21462,N_21485);
xor U21729 (N_21729,N_21446,N_21405);
or U21730 (N_21730,N_21407,N_21526);
xnor U21731 (N_21731,N_21555,N_21401);
or U21732 (N_21732,N_21494,N_21576);
or U21733 (N_21733,N_21554,N_21463);
xnor U21734 (N_21734,N_21597,N_21419);
or U21735 (N_21735,N_21516,N_21579);
and U21736 (N_21736,N_21554,N_21587);
and U21737 (N_21737,N_21513,N_21530);
nand U21738 (N_21738,N_21410,N_21415);
nand U21739 (N_21739,N_21597,N_21593);
and U21740 (N_21740,N_21477,N_21455);
nand U21741 (N_21741,N_21534,N_21535);
nand U21742 (N_21742,N_21457,N_21505);
or U21743 (N_21743,N_21544,N_21432);
nor U21744 (N_21744,N_21570,N_21553);
nor U21745 (N_21745,N_21542,N_21576);
nand U21746 (N_21746,N_21529,N_21473);
xor U21747 (N_21747,N_21517,N_21534);
nand U21748 (N_21748,N_21539,N_21428);
and U21749 (N_21749,N_21579,N_21461);
and U21750 (N_21750,N_21514,N_21581);
nand U21751 (N_21751,N_21493,N_21514);
nand U21752 (N_21752,N_21491,N_21463);
and U21753 (N_21753,N_21536,N_21554);
nand U21754 (N_21754,N_21565,N_21432);
and U21755 (N_21755,N_21572,N_21496);
and U21756 (N_21756,N_21450,N_21589);
nor U21757 (N_21757,N_21502,N_21584);
xor U21758 (N_21758,N_21505,N_21577);
and U21759 (N_21759,N_21438,N_21410);
nand U21760 (N_21760,N_21585,N_21561);
or U21761 (N_21761,N_21484,N_21534);
nor U21762 (N_21762,N_21434,N_21425);
xor U21763 (N_21763,N_21425,N_21435);
xnor U21764 (N_21764,N_21595,N_21498);
or U21765 (N_21765,N_21565,N_21474);
nand U21766 (N_21766,N_21593,N_21566);
and U21767 (N_21767,N_21571,N_21557);
nor U21768 (N_21768,N_21470,N_21405);
nor U21769 (N_21769,N_21446,N_21573);
and U21770 (N_21770,N_21430,N_21549);
and U21771 (N_21771,N_21501,N_21545);
nand U21772 (N_21772,N_21475,N_21408);
and U21773 (N_21773,N_21593,N_21536);
or U21774 (N_21774,N_21418,N_21584);
or U21775 (N_21775,N_21558,N_21522);
nor U21776 (N_21776,N_21408,N_21522);
xnor U21777 (N_21777,N_21443,N_21494);
and U21778 (N_21778,N_21521,N_21426);
or U21779 (N_21779,N_21597,N_21413);
xnor U21780 (N_21780,N_21594,N_21483);
nand U21781 (N_21781,N_21527,N_21585);
nand U21782 (N_21782,N_21470,N_21548);
or U21783 (N_21783,N_21406,N_21509);
xnor U21784 (N_21784,N_21591,N_21419);
and U21785 (N_21785,N_21408,N_21499);
and U21786 (N_21786,N_21583,N_21544);
nand U21787 (N_21787,N_21532,N_21560);
xor U21788 (N_21788,N_21562,N_21598);
nor U21789 (N_21789,N_21559,N_21511);
nor U21790 (N_21790,N_21471,N_21496);
xor U21791 (N_21791,N_21440,N_21579);
or U21792 (N_21792,N_21480,N_21460);
and U21793 (N_21793,N_21480,N_21484);
and U21794 (N_21794,N_21414,N_21591);
nor U21795 (N_21795,N_21428,N_21556);
and U21796 (N_21796,N_21544,N_21411);
or U21797 (N_21797,N_21471,N_21563);
nand U21798 (N_21798,N_21522,N_21482);
and U21799 (N_21799,N_21500,N_21466);
nand U21800 (N_21800,N_21601,N_21754);
and U21801 (N_21801,N_21764,N_21707);
or U21802 (N_21802,N_21671,N_21664);
xnor U21803 (N_21803,N_21638,N_21680);
xnor U21804 (N_21804,N_21705,N_21727);
nand U21805 (N_21805,N_21686,N_21643);
or U21806 (N_21806,N_21756,N_21688);
nand U21807 (N_21807,N_21616,N_21645);
or U21808 (N_21808,N_21661,N_21783);
nor U21809 (N_21809,N_21769,N_21604);
nor U21810 (N_21810,N_21692,N_21613);
and U21811 (N_21811,N_21749,N_21796);
nand U21812 (N_21812,N_21776,N_21755);
nor U21813 (N_21813,N_21697,N_21672);
nand U21814 (N_21814,N_21773,N_21721);
nand U21815 (N_21815,N_21626,N_21740);
nor U21816 (N_21816,N_21794,N_21659);
xnor U21817 (N_21817,N_21767,N_21718);
nor U21818 (N_21818,N_21602,N_21654);
or U21819 (N_21819,N_21693,N_21774);
and U21820 (N_21820,N_21667,N_21708);
and U21821 (N_21821,N_21636,N_21676);
or U21822 (N_21822,N_21666,N_21712);
or U21823 (N_21823,N_21786,N_21732);
nand U21824 (N_21824,N_21675,N_21799);
xor U21825 (N_21825,N_21634,N_21742);
nand U21826 (N_21826,N_21772,N_21785);
xnor U21827 (N_21827,N_21600,N_21699);
and U21828 (N_21828,N_21746,N_21630);
nor U21829 (N_21829,N_21758,N_21698);
nor U21830 (N_21830,N_21750,N_21606);
nand U21831 (N_21831,N_21789,N_21720);
or U21832 (N_21832,N_21747,N_21700);
or U21833 (N_21833,N_21629,N_21777);
nand U21834 (N_21834,N_21696,N_21797);
or U21835 (N_21835,N_21795,N_21670);
nor U21836 (N_21836,N_21605,N_21788);
or U21837 (N_21837,N_21735,N_21658);
or U21838 (N_21838,N_21682,N_21728);
xnor U21839 (N_21839,N_21624,N_21781);
nand U21840 (N_21840,N_21669,N_21779);
nand U21841 (N_21841,N_21617,N_21762);
xnor U21842 (N_21842,N_21757,N_21714);
or U21843 (N_21843,N_21715,N_21753);
nand U21844 (N_21844,N_21655,N_21619);
xnor U21845 (N_21845,N_21775,N_21625);
nor U21846 (N_21846,N_21652,N_21719);
nor U21847 (N_21847,N_21628,N_21607);
and U21848 (N_21848,N_21646,N_21725);
or U21849 (N_21849,N_21620,N_21662);
and U21850 (N_21850,N_21685,N_21660);
xor U21851 (N_21851,N_21731,N_21739);
nor U21852 (N_21852,N_21653,N_21734);
or U21853 (N_21853,N_21752,N_21778);
and U21854 (N_21854,N_21691,N_21694);
nor U21855 (N_21855,N_21637,N_21627);
nor U21856 (N_21856,N_21702,N_21640);
and U21857 (N_21857,N_21631,N_21695);
or U21858 (N_21858,N_21621,N_21770);
nor U21859 (N_21859,N_21665,N_21771);
nand U21860 (N_21860,N_21759,N_21679);
or U21861 (N_21861,N_21639,N_21729);
nor U21862 (N_21862,N_21678,N_21713);
xor U21863 (N_21863,N_21790,N_21683);
nand U21864 (N_21864,N_21689,N_21763);
xor U21865 (N_21865,N_21741,N_21798);
or U21866 (N_21866,N_21743,N_21650);
and U21867 (N_21867,N_21632,N_21730);
and U21868 (N_21868,N_21641,N_21663);
and U21869 (N_21869,N_21673,N_21610);
xor U21870 (N_21870,N_21792,N_21761);
xnor U21871 (N_21871,N_21706,N_21768);
nand U21872 (N_21872,N_21751,N_21766);
or U21873 (N_21873,N_21656,N_21647);
nand U21874 (N_21874,N_21614,N_21623);
nand U21875 (N_21875,N_21687,N_21733);
and U21876 (N_21876,N_21622,N_21784);
nand U21877 (N_21877,N_21791,N_21651);
nor U21878 (N_21878,N_21744,N_21765);
or U21879 (N_21879,N_21615,N_21608);
nor U21880 (N_21880,N_21710,N_21674);
and U21881 (N_21881,N_21644,N_21724);
xnor U21882 (N_21882,N_21760,N_21649);
and U21883 (N_21883,N_21709,N_21711);
nand U21884 (N_21884,N_21703,N_21722);
nand U21885 (N_21885,N_21780,N_21684);
xnor U21886 (N_21886,N_21612,N_21704);
xnor U21887 (N_21887,N_21748,N_21723);
nor U21888 (N_21888,N_21737,N_21633);
nand U21889 (N_21889,N_21738,N_21717);
xor U21890 (N_21890,N_21677,N_21635);
xor U21891 (N_21891,N_21793,N_21648);
nand U21892 (N_21892,N_21782,N_21642);
nand U21893 (N_21893,N_21603,N_21681);
nand U21894 (N_21894,N_21716,N_21787);
nand U21895 (N_21895,N_21745,N_21609);
or U21896 (N_21896,N_21657,N_21690);
and U21897 (N_21897,N_21618,N_21736);
or U21898 (N_21898,N_21701,N_21668);
nor U21899 (N_21899,N_21726,N_21611);
nand U21900 (N_21900,N_21659,N_21758);
nor U21901 (N_21901,N_21600,N_21730);
xor U21902 (N_21902,N_21640,N_21729);
and U21903 (N_21903,N_21631,N_21696);
nand U21904 (N_21904,N_21700,N_21717);
xor U21905 (N_21905,N_21729,N_21610);
nand U21906 (N_21906,N_21685,N_21680);
xor U21907 (N_21907,N_21778,N_21704);
nand U21908 (N_21908,N_21738,N_21683);
and U21909 (N_21909,N_21730,N_21630);
nor U21910 (N_21910,N_21746,N_21724);
nand U21911 (N_21911,N_21791,N_21710);
or U21912 (N_21912,N_21619,N_21675);
or U21913 (N_21913,N_21759,N_21790);
xnor U21914 (N_21914,N_21785,N_21776);
or U21915 (N_21915,N_21694,N_21711);
and U21916 (N_21916,N_21705,N_21770);
nand U21917 (N_21917,N_21723,N_21765);
or U21918 (N_21918,N_21656,N_21645);
and U21919 (N_21919,N_21681,N_21653);
nor U21920 (N_21920,N_21690,N_21765);
nor U21921 (N_21921,N_21766,N_21705);
nor U21922 (N_21922,N_21633,N_21705);
xor U21923 (N_21923,N_21638,N_21645);
or U21924 (N_21924,N_21727,N_21772);
and U21925 (N_21925,N_21646,N_21703);
nor U21926 (N_21926,N_21775,N_21743);
nor U21927 (N_21927,N_21792,N_21776);
and U21928 (N_21928,N_21663,N_21795);
xnor U21929 (N_21929,N_21699,N_21780);
and U21930 (N_21930,N_21749,N_21756);
and U21931 (N_21931,N_21761,N_21722);
or U21932 (N_21932,N_21702,N_21655);
or U21933 (N_21933,N_21788,N_21622);
nand U21934 (N_21934,N_21774,N_21785);
and U21935 (N_21935,N_21651,N_21605);
nand U21936 (N_21936,N_21639,N_21792);
or U21937 (N_21937,N_21754,N_21701);
nand U21938 (N_21938,N_21617,N_21787);
nor U21939 (N_21939,N_21700,N_21750);
or U21940 (N_21940,N_21660,N_21774);
and U21941 (N_21941,N_21744,N_21784);
and U21942 (N_21942,N_21708,N_21630);
nand U21943 (N_21943,N_21632,N_21783);
and U21944 (N_21944,N_21780,N_21625);
xnor U21945 (N_21945,N_21752,N_21711);
nor U21946 (N_21946,N_21757,N_21738);
or U21947 (N_21947,N_21634,N_21685);
xnor U21948 (N_21948,N_21690,N_21635);
or U21949 (N_21949,N_21786,N_21686);
or U21950 (N_21950,N_21656,N_21731);
nand U21951 (N_21951,N_21685,N_21726);
or U21952 (N_21952,N_21630,N_21717);
nor U21953 (N_21953,N_21795,N_21766);
or U21954 (N_21954,N_21648,N_21788);
xor U21955 (N_21955,N_21632,N_21723);
xnor U21956 (N_21956,N_21613,N_21747);
or U21957 (N_21957,N_21712,N_21651);
and U21958 (N_21958,N_21720,N_21719);
or U21959 (N_21959,N_21666,N_21730);
and U21960 (N_21960,N_21736,N_21697);
xnor U21961 (N_21961,N_21639,N_21613);
or U21962 (N_21962,N_21664,N_21744);
xnor U21963 (N_21963,N_21761,N_21798);
nand U21964 (N_21964,N_21702,N_21777);
nand U21965 (N_21965,N_21615,N_21768);
xnor U21966 (N_21966,N_21738,N_21760);
or U21967 (N_21967,N_21600,N_21656);
and U21968 (N_21968,N_21633,N_21618);
xnor U21969 (N_21969,N_21738,N_21699);
nor U21970 (N_21970,N_21695,N_21715);
and U21971 (N_21971,N_21606,N_21648);
nor U21972 (N_21972,N_21747,N_21659);
nor U21973 (N_21973,N_21614,N_21705);
or U21974 (N_21974,N_21701,N_21797);
and U21975 (N_21975,N_21639,N_21628);
nor U21976 (N_21976,N_21753,N_21744);
xnor U21977 (N_21977,N_21738,N_21746);
and U21978 (N_21978,N_21787,N_21610);
xor U21979 (N_21979,N_21758,N_21783);
xor U21980 (N_21980,N_21792,N_21677);
and U21981 (N_21981,N_21628,N_21714);
or U21982 (N_21982,N_21715,N_21772);
nand U21983 (N_21983,N_21684,N_21761);
nor U21984 (N_21984,N_21667,N_21798);
xnor U21985 (N_21985,N_21602,N_21738);
nor U21986 (N_21986,N_21789,N_21606);
and U21987 (N_21987,N_21775,N_21612);
nand U21988 (N_21988,N_21714,N_21703);
or U21989 (N_21989,N_21759,N_21657);
xnor U21990 (N_21990,N_21797,N_21662);
and U21991 (N_21991,N_21675,N_21674);
nor U21992 (N_21992,N_21663,N_21717);
and U21993 (N_21993,N_21654,N_21777);
nand U21994 (N_21994,N_21791,N_21742);
or U21995 (N_21995,N_21600,N_21774);
nor U21996 (N_21996,N_21654,N_21736);
and U21997 (N_21997,N_21716,N_21708);
xnor U21998 (N_21998,N_21616,N_21696);
nand U21999 (N_21999,N_21702,N_21784);
nor U22000 (N_22000,N_21916,N_21899);
nor U22001 (N_22001,N_21930,N_21929);
and U22002 (N_22002,N_21874,N_21820);
xnor U22003 (N_22003,N_21984,N_21831);
and U22004 (N_22004,N_21979,N_21876);
and U22005 (N_22005,N_21849,N_21810);
nor U22006 (N_22006,N_21924,N_21974);
or U22007 (N_22007,N_21942,N_21871);
xnor U22008 (N_22008,N_21903,N_21808);
xnor U22009 (N_22009,N_21980,N_21915);
nand U22010 (N_22010,N_21801,N_21837);
xnor U22011 (N_22011,N_21817,N_21989);
nor U22012 (N_22012,N_21813,N_21948);
xnor U22013 (N_22013,N_21986,N_21839);
nand U22014 (N_22014,N_21838,N_21856);
and U22015 (N_22015,N_21873,N_21882);
nand U22016 (N_22016,N_21997,N_21946);
nand U22017 (N_22017,N_21821,N_21963);
nor U22018 (N_22018,N_21823,N_21996);
nand U22019 (N_22019,N_21976,N_21975);
or U22020 (N_22020,N_21834,N_21912);
nor U22021 (N_22021,N_21988,N_21983);
nor U22022 (N_22022,N_21895,N_21847);
nand U22023 (N_22023,N_21933,N_21973);
nor U22024 (N_22024,N_21884,N_21832);
or U22025 (N_22025,N_21990,N_21928);
and U22026 (N_22026,N_21805,N_21978);
xnor U22027 (N_22027,N_21852,N_21841);
xor U22028 (N_22028,N_21936,N_21807);
xnor U22029 (N_22029,N_21938,N_21862);
and U22030 (N_22030,N_21944,N_21968);
and U22031 (N_22031,N_21966,N_21865);
or U22032 (N_22032,N_21888,N_21875);
nand U22033 (N_22033,N_21864,N_21926);
nor U22034 (N_22034,N_21935,N_21998);
nor U22035 (N_22035,N_21962,N_21870);
or U22036 (N_22036,N_21981,N_21812);
and U22037 (N_22037,N_21894,N_21958);
xor U22038 (N_22038,N_21851,N_21957);
or U22039 (N_22039,N_21896,N_21919);
or U22040 (N_22040,N_21941,N_21897);
nand U22041 (N_22041,N_21908,N_21858);
and U22042 (N_22042,N_21891,N_21954);
or U22043 (N_22043,N_21907,N_21932);
and U22044 (N_22044,N_21955,N_21971);
nand U22045 (N_22045,N_21911,N_21972);
xnor U22046 (N_22046,N_21993,N_21866);
nor U22047 (N_22047,N_21861,N_21960);
nand U22048 (N_22048,N_21868,N_21804);
nor U22049 (N_22049,N_21910,N_21854);
xor U22050 (N_22050,N_21937,N_21803);
and U22051 (N_22051,N_21991,N_21898);
nand U22052 (N_22052,N_21999,N_21889);
xor U22053 (N_22053,N_21835,N_21877);
nor U22054 (N_22054,N_21927,N_21800);
nand U22055 (N_22055,N_21920,N_21819);
or U22056 (N_22056,N_21947,N_21822);
and U22057 (N_22057,N_21853,N_21863);
or U22058 (N_22058,N_21995,N_21977);
nand U22059 (N_22059,N_21814,N_21860);
or U22060 (N_22060,N_21901,N_21917);
xor U22061 (N_22061,N_21982,N_21833);
nand U22062 (N_22062,N_21902,N_21952);
nor U22063 (N_22063,N_21830,N_21890);
nand U22064 (N_22064,N_21878,N_21816);
and U22065 (N_22065,N_21893,N_21953);
nand U22066 (N_22066,N_21818,N_21961);
or U22067 (N_22067,N_21943,N_21869);
and U22068 (N_22068,N_21950,N_21940);
nand U22069 (N_22069,N_21827,N_21922);
or U22070 (N_22070,N_21987,N_21811);
xnor U22071 (N_22071,N_21857,N_21836);
nand U22072 (N_22072,N_21842,N_21845);
and U22073 (N_22073,N_21918,N_21825);
nand U22074 (N_22074,N_21906,N_21850);
xor U22075 (N_22075,N_21959,N_21885);
nand U22076 (N_22076,N_21828,N_21887);
nand U22077 (N_22077,N_21809,N_21855);
nor U22078 (N_22078,N_21905,N_21969);
nand U22079 (N_22079,N_21892,N_21824);
nand U22080 (N_22080,N_21881,N_21872);
nand U22081 (N_22081,N_21909,N_21925);
or U22082 (N_22082,N_21992,N_21844);
xnor U22083 (N_22083,N_21843,N_21956);
xnor U22084 (N_22084,N_21815,N_21914);
xnor U22085 (N_22085,N_21923,N_21904);
nor U22086 (N_22086,N_21913,N_21945);
or U22087 (N_22087,N_21967,N_21921);
xor U22088 (N_22088,N_21840,N_21970);
xnor U22089 (N_22089,N_21939,N_21829);
xor U22090 (N_22090,N_21867,N_21802);
nand U22091 (N_22091,N_21859,N_21934);
xor U22092 (N_22092,N_21806,N_21951);
nor U22093 (N_22093,N_21965,N_21886);
nor U22094 (N_22094,N_21826,N_21931);
nor U22095 (N_22095,N_21883,N_21846);
nand U22096 (N_22096,N_21994,N_21880);
xor U22097 (N_22097,N_21985,N_21964);
nor U22098 (N_22098,N_21949,N_21879);
xor U22099 (N_22099,N_21848,N_21900);
nor U22100 (N_22100,N_21888,N_21867);
nor U22101 (N_22101,N_21990,N_21803);
nand U22102 (N_22102,N_21814,N_21839);
nand U22103 (N_22103,N_21804,N_21911);
and U22104 (N_22104,N_21938,N_21926);
xnor U22105 (N_22105,N_21962,N_21979);
or U22106 (N_22106,N_21818,N_21840);
xor U22107 (N_22107,N_21811,N_21835);
or U22108 (N_22108,N_21977,N_21997);
nor U22109 (N_22109,N_21934,N_21819);
and U22110 (N_22110,N_21809,N_21930);
nand U22111 (N_22111,N_21860,N_21872);
xor U22112 (N_22112,N_21813,N_21931);
nor U22113 (N_22113,N_21832,N_21915);
or U22114 (N_22114,N_21827,N_21867);
nand U22115 (N_22115,N_21940,N_21973);
and U22116 (N_22116,N_21832,N_21887);
nor U22117 (N_22117,N_21987,N_21834);
and U22118 (N_22118,N_21808,N_21931);
or U22119 (N_22119,N_21993,N_21919);
nand U22120 (N_22120,N_21964,N_21920);
or U22121 (N_22121,N_21954,N_21874);
nand U22122 (N_22122,N_21814,N_21845);
or U22123 (N_22123,N_21842,N_21948);
and U22124 (N_22124,N_21986,N_21930);
nor U22125 (N_22125,N_21878,N_21959);
or U22126 (N_22126,N_21895,N_21862);
nand U22127 (N_22127,N_21867,N_21850);
or U22128 (N_22128,N_21920,N_21827);
nand U22129 (N_22129,N_21950,N_21843);
xor U22130 (N_22130,N_21859,N_21972);
or U22131 (N_22131,N_21880,N_21986);
xnor U22132 (N_22132,N_21855,N_21868);
nor U22133 (N_22133,N_21925,N_21848);
nor U22134 (N_22134,N_21997,N_21993);
or U22135 (N_22135,N_21926,N_21879);
nor U22136 (N_22136,N_21983,N_21969);
nand U22137 (N_22137,N_21981,N_21953);
nor U22138 (N_22138,N_21846,N_21991);
nand U22139 (N_22139,N_21949,N_21829);
or U22140 (N_22140,N_21887,N_21829);
and U22141 (N_22141,N_21834,N_21921);
nand U22142 (N_22142,N_21941,N_21997);
nor U22143 (N_22143,N_21863,N_21937);
nand U22144 (N_22144,N_21983,N_21938);
and U22145 (N_22145,N_21831,N_21916);
nor U22146 (N_22146,N_21843,N_21942);
or U22147 (N_22147,N_21942,N_21917);
xor U22148 (N_22148,N_21871,N_21984);
or U22149 (N_22149,N_21992,N_21836);
xor U22150 (N_22150,N_21925,N_21877);
nand U22151 (N_22151,N_21842,N_21978);
and U22152 (N_22152,N_21993,N_21830);
nand U22153 (N_22153,N_21954,N_21943);
nand U22154 (N_22154,N_21905,N_21854);
xnor U22155 (N_22155,N_21840,N_21820);
nand U22156 (N_22156,N_21817,N_21986);
and U22157 (N_22157,N_21912,N_21816);
and U22158 (N_22158,N_21847,N_21848);
and U22159 (N_22159,N_21985,N_21826);
or U22160 (N_22160,N_21986,N_21816);
nor U22161 (N_22161,N_21981,N_21826);
xnor U22162 (N_22162,N_21868,N_21885);
xnor U22163 (N_22163,N_21854,N_21978);
xnor U22164 (N_22164,N_21839,N_21871);
nor U22165 (N_22165,N_21826,N_21873);
xnor U22166 (N_22166,N_21950,N_21901);
xor U22167 (N_22167,N_21951,N_21880);
xnor U22168 (N_22168,N_21913,N_21905);
and U22169 (N_22169,N_21877,N_21819);
and U22170 (N_22170,N_21816,N_21818);
xnor U22171 (N_22171,N_21925,N_21888);
nand U22172 (N_22172,N_21853,N_21909);
xor U22173 (N_22173,N_21876,N_21998);
or U22174 (N_22174,N_21961,N_21911);
nand U22175 (N_22175,N_21919,N_21931);
xor U22176 (N_22176,N_21964,N_21889);
nor U22177 (N_22177,N_21828,N_21910);
nor U22178 (N_22178,N_21854,N_21829);
nand U22179 (N_22179,N_21847,N_21898);
xnor U22180 (N_22180,N_21872,N_21800);
or U22181 (N_22181,N_21938,N_21824);
nand U22182 (N_22182,N_21863,N_21997);
xnor U22183 (N_22183,N_21883,N_21962);
nor U22184 (N_22184,N_21908,N_21842);
xor U22185 (N_22185,N_21939,N_21965);
nor U22186 (N_22186,N_21868,N_21850);
and U22187 (N_22187,N_21859,N_21874);
xnor U22188 (N_22188,N_21993,N_21979);
or U22189 (N_22189,N_21925,N_21894);
xnor U22190 (N_22190,N_21929,N_21946);
nor U22191 (N_22191,N_21829,N_21817);
nor U22192 (N_22192,N_21889,N_21996);
nor U22193 (N_22193,N_21820,N_21822);
nor U22194 (N_22194,N_21887,N_21972);
or U22195 (N_22195,N_21988,N_21990);
and U22196 (N_22196,N_21925,N_21962);
and U22197 (N_22197,N_21813,N_21855);
and U22198 (N_22198,N_21845,N_21910);
nand U22199 (N_22199,N_21973,N_21873);
nor U22200 (N_22200,N_22075,N_22030);
nor U22201 (N_22201,N_22032,N_22077);
nor U22202 (N_22202,N_22116,N_22037);
or U22203 (N_22203,N_22010,N_22029);
nor U22204 (N_22204,N_22117,N_22151);
nor U22205 (N_22205,N_22155,N_22174);
nor U22206 (N_22206,N_22104,N_22042);
nand U22207 (N_22207,N_22101,N_22018);
and U22208 (N_22208,N_22127,N_22109);
nor U22209 (N_22209,N_22064,N_22196);
nand U22210 (N_22210,N_22001,N_22097);
nor U22211 (N_22211,N_22192,N_22186);
nor U22212 (N_22212,N_22184,N_22195);
xor U22213 (N_22213,N_22039,N_22090);
nor U22214 (N_22214,N_22167,N_22121);
nand U22215 (N_22215,N_22180,N_22133);
and U22216 (N_22216,N_22038,N_22181);
or U22217 (N_22217,N_22126,N_22136);
nand U22218 (N_22218,N_22093,N_22140);
nand U22219 (N_22219,N_22106,N_22158);
nand U22220 (N_22220,N_22153,N_22049);
xnor U22221 (N_22221,N_22026,N_22144);
or U22222 (N_22222,N_22147,N_22150);
xor U22223 (N_22223,N_22040,N_22099);
nor U22224 (N_22224,N_22008,N_22103);
and U22225 (N_22225,N_22041,N_22028);
nand U22226 (N_22226,N_22080,N_22044);
nand U22227 (N_22227,N_22185,N_22115);
or U22228 (N_22228,N_22189,N_22123);
nand U22229 (N_22229,N_22194,N_22073);
xor U22230 (N_22230,N_22164,N_22062);
nor U22231 (N_22231,N_22013,N_22047);
nand U22232 (N_22232,N_22031,N_22059);
nand U22233 (N_22233,N_22119,N_22173);
or U22234 (N_22234,N_22125,N_22048);
xor U22235 (N_22235,N_22129,N_22182);
xor U22236 (N_22236,N_22162,N_22149);
nor U22237 (N_22237,N_22172,N_22091);
nor U22238 (N_22238,N_22120,N_22014);
or U22239 (N_22239,N_22095,N_22055);
nand U22240 (N_22240,N_22022,N_22067);
and U22241 (N_22241,N_22015,N_22003);
nand U22242 (N_22242,N_22060,N_22135);
or U22243 (N_22243,N_22154,N_22112);
nand U22244 (N_22244,N_22046,N_22083);
or U22245 (N_22245,N_22058,N_22124);
or U22246 (N_22246,N_22183,N_22110);
and U22247 (N_22247,N_22105,N_22078);
xnor U22248 (N_22248,N_22074,N_22171);
and U22249 (N_22249,N_22025,N_22139);
nor U22250 (N_22250,N_22156,N_22131);
nand U22251 (N_22251,N_22016,N_22056);
nand U22252 (N_22252,N_22193,N_22079);
and U22253 (N_22253,N_22069,N_22011);
or U22254 (N_22254,N_22066,N_22163);
nor U22255 (N_22255,N_22111,N_22197);
nor U22256 (N_22256,N_22088,N_22188);
nor U22257 (N_22257,N_22166,N_22034);
and U22258 (N_22258,N_22002,N_22084);
or U22259 (N_22259,N_22072,N_22145);
xnor U22260 (N_22260,N_22102,N_22085);
or U22261 (N_22261,N_22087,N_22024);
or U22262 (N_22262,N_22053,N_22138);
nor U22263 (N_22263,N_22000,N_22179);
and U22264 (N_22264,N_22178,N_22092);
and U22265 (N_22265,N_22198,N_22082);
nand U22266 (N_22266,N_22006,N_22177);
xnor U22267 (N_22267,N_22142,N_22033);
nand U22268 (N_22268,N_22023,N_22128);
nor U22269 (N_22269,N_22137,N_22020);
xnor U22270 (N_22270,N_22052,N_22118);
nor U22271 (N_22271,N_22130,N_22036);
or U22272 (N_22272,N_22021,N_22065);
nand U22273 (N_22273,N_22134,N_22165);
and U22274 (N_22274,N_22012,N_22094);
and U22275 (N_22275,N_22143,N_22170);
and U22276 (N_22276,N_22190,N_22176);
nor U22277 (N_22277,N_22199,N_22051);
and U22278 (N_22278,N_22152,N_22108);
nor U22279 (N_22279,N_22160,N_22045);
and U22280 (N_22280,N_22050,N_22063);
nand U22281 (N_22281,N_22043,N_22132);
xor U22282 (N_22282,N_22122,N_22175);
and U22283 (N_22283,N_22057,N_22146);
nand U22284 (N_22284,N_22004,N_22007);
nor U22285 (N_22285,N_22141,N_22068);
or U22286 (N_22286,N_22114,N_22070);
nor U22287 (N_22287,N_22161,N_22061);
or U22288 (N_22288,N_22009,N_22054);
nand U22289 (N_22289,N_22071,N_22113);
nand U22290 (N_22290,N_22168,N_22107);
nand U22291 (N_22291,N_22017,N_22089);
or U22292 (N_22292,N_22081,N_22148);
nand U22293 (N_22293,N_22005,N_22076);
and U22294 (N_22294,N_22098,N_22191);
xor U22295 (N_22295,N_22100,N_22035);
or U22296 (N_22296,N_22096,N_22159);
nor U22297 (N_22297,N_22157,N_22019);
or U22298 (N_22298,N_22169,N_22086);
or U22299 (N_22299,N_22027,N_22187);
xor U22300 (N_22300,N_22074,N_22044);
xnor U22301 (N_22301,N_22183,N_22150);
or U22302 (N_22302,N_22047,N_22196);
or U22303 (N_22303,N_22051,N_22078);
or U22304 (N_22304,N_22126,N_22105);
nor U22305 (N_22305,N_22189,N_22068);
nor U22306 (N_22306,N_22188,N_22107);
nand U22307 (N_22307,N_22121,N_22024);
xor U22308 (N_22308,N_22140,N_22034);
nor U22309 (N_22309,N_22161,N_22173);
xnor U22310 (N_22310,N_22081,N_22049);
xnor U22311 (N_22311,N_22190,N_22168);
and U22312 (N_22312,N_22082,N_22178);
and U22313 (N_22313,N_22025,N_22035);
xor U22314 (N_22314,N_22036,N_22115);
and U22315 (N_22315,N_22152,N_22021);
and U22316 (N_22316,N_22119,N_22100);
xor U22317 (N_22317,N_22007,N_22094);
nor U22318 (N_22318,N_22090,N_22029);
xnor U22319 (N_22319,N_22023,N_22187);
nor U22320 (N_22320,N_22122,N_22174);
xor U22321 (N_22321,N_22129,N_22199);
and U22322 (N_22322,N_22057,N_22094);
nand U22323 (N_22323,N_22094,N_22042);
or U22324 (N_22324,N_22172,N_22097);
and U22325 (N_22325,N_22127,N_22013);
xnor U22326 (N_22326,N_22173,N_22159);
and U22327 (N_22327,N_22024,N_22049);
xnor U22328 (N_22328,N_22131,N_22122);
and U22329 (N_22329,N_22166,N_22071);
xor U22330 (N_22330,N_22046,N_22054);
and U22331 (N_22331,N_22104,N_22069);
nor U22332 (N_22332,N_22002,N_22076);
and U22333 (N_22333,N_22157,N_22163);
nor U22334 (N_22334,N_22131,N_22121);
nand U22335 (N_22335,N_22113,N_22053);
and U22336 (N_22336,N_22078,N_22144);
nand U22337 (N_22337,N_22107,N_22172);
or U22338 (N_22338,N_22101,N_22120);
nand U22339 (N_22339,N_22120,N_22164);
nand U22340 (N_22340,N_22043,N_22014);
and U22341 (N_22341,N_22065,N_22013);
nor U22342 (N_22342,N_22104,N_22173);
and U22343 (N_22343,N_22123,N_22091);
xnor U22344 (N_22344,N_22002,N_22001);
nor U22345 (N_22345,N_22074,N_22045);
nor U22346 (N_22346,N_22072,N_22146);
nor U22347 (N_22347,N_22140,N_22177);
nand U22348 (N_22348,N_22120,N_22139);
or U22349 (N_22349,N_22175,N_22019);
nor U22350 (N_22350,N_22094,N_22167);
xnor U22351 (N_22351,N_22081,N_22149);
xor U22352 (N_22352,N_22017,N_22176);
or U22353 (N_22353,N_22060,N_22078);
xor U22354 (N_22354,N_22158,N_22073);
and U22355 (N_22355,N_22192,N_22019);
nand U22356 (N_22356,N_22034,N_22175);
nand U22357 (N_22357,N_22088,N_22185);
or U22358 (N_22358,N_22181,N_22092);
nand U22359 (N_22359,N_22031,N_22030);
nor U22360 (N_22360,N_22166,N_22010);
nand U22361 (N_22361,N_22195,N_22169);
and U22362 (N_22362,N_22118,N_22111);
xor U22363 (N_22363,N_22140,N_22170);
xnor U22364 (N_22364,N_22059,N_22074);
or U22365 (N_22365,N_22158,N_22144);
nand U22366 (N_22366,N_22163,N_22142);
nor U22367 (N_22367,N_22126,N_22110);
nor U22368 (N_22368,N_22092,N_22091);
or U22369 (N_22369,N_22110,N_22135);
and U22370 (N_22370,N_22004,N_22152);
and U22371 (N_22371,N_22159,N_22122);
and U22372 (N_22372,N_22197,N_22061);
xnor U22373 (N_22373,N_22165,N_22132);
nand U22374 (N_22374,N_22197,N_22170);
nand U22375 (N_22375,N_22158,N_22009);
xnor U22376 (N_22376,N_22119,N_22142);
or U22377 (N_22377,N_22078,N_22063);
or U22378 (N_22378,N_22128,N_22048);
or U22379 (N_22379,N_22044,N_22127);
or U22380 (N_22380,N_22118,N_22080);
nor U22381 (N_22381,N_22019,N_22064);
nor U22382 (N_22382,N_22094,N_22118);
or U22383 (N_22383,N_22073,N_22014);
xnor U22384 (N_22384,N_22187,N_22033);
nor U22385 (N_22385,N_22095,N_22140);
nand U22386 (N_22386,N_22140,N_22014);
nand U22387 (N_22387,N_22060,N_22051);
xor U22388 (N_22388,N_22182,N_22038);
xor U22389 (N_22389,N_22071,N_22055);
nor U22390 (N_22390,N_22108,N_22062);
nand U22391 (N_22391,N_22142,N_22064);
xor U22392 (N_22392,N_22083,N_22102);
xnor U22393 (N_22393,N_22175,N_22174);
xnor U22394 (N_22394,N_22158,N_22192);
nand U22395 (N_22395,N_22027,N_22087);
nand U22396 (N_22396,N_22078,N_22141);
nor U22397 (N_22397,N_22155,N_22085);
nor U22398 (N_22398,N_22162,N_22190);
xnor U22399 (N_22399,N_22194,N_22115);
or U22400 (N_22400,N_22261,N_22225);
nand U22401 (N_22401,N_22256,N_22378);
and U22402 (N_22402,N_22343,N_22339);
or U22403 (N_22403,N_22300,N_22203);
nand U22404 (N_22404,N_22220,N_22395);
and U22405 (N_22405,N_22307,N_22253);
xor U22406 (N_22406,N_22335,N_22348);
nor U22407 (N_22407,N_22292,N_22270);
or U22408 (N_22408,N_22340,N_22237);
or U22409 (N_22409,N_22252,N_22322);
nand U22410 (N_22410,N_22315,N_22217);
nand U22411 (N_22411,N_22254,N_22281);
nor U22412 (N_22412,N_22301,N_22357);
and U22413 (N_22413,N_22226,N_22235);
or U22414 (N_22414,N_22297,N_22334);
and U22415 (N_22415,N_22214,N_22286);
nand U22416 (N_22416,N_22383,N_22243);
or U22417 (N_22417,N_22313,N_22345);
nand U22418 (N_22418,N_22224,N_22371);
xor U22419 (N_22419,N_22287,N_22207);
xnor U22420 (N_22420,N_22306,N_22376);
xnor U22421 (N_22421,N_22344,N_22283);
xor U22422 (N_22422,N_22249,N_22304);
and U22423 (N_22423,N_22278,N_22316);
xor U22424 (N_22424,N_22231,N_22366);
nor U22425 (N_22425,N_22327,N_22245);
nand U22426 (N_22426,N_22389,N_22341);
nand U22427 (N_22427,N_22377,N_22309);
nand U22428 (N_22428,N_22265,N_22353);
xor U22429 (N_22429,N_22333,N_22317);
or U22430 (N_22430,N_22223,N_22330);
and U22431 (N_22431,N_22200,N_22209);
nor U22432 (N_22432,N_22387,N_22386);
nor U22433 (N_22433,N_22251,N_22221);
xnor U22434 (N_22434,N_22367,N_22218);
nand U22435 (N_22435,N_22296,N_22314);
nand U22436 (N_22436,N_22294,N_22241);
or U22437 (N_22437,N_22205,N_22234);
nand U22438 (N_22438,N_22239,N_22392);
nor U22439 (N_22439,N_22240,N_22321);
xnor U22440 (N_22440,N_22288,N_22215);
xor U22441 (N_22441,N_22364,N_22312);
nor U22442 (N_22442,N_22355,N_22279);
xor U22443 (N_22443,N_22238,N_22393);
xor U22444 (N_22444,N_22227,N_22388);
nand U22445 (N_22445,N_22338,N_22285);
nand U22446 (N_22446,N_22248,N_22271);
and U22447 (N_22447,N_22368,N_22291);
nor U22448 (N_22448,N_22267,N_22246);
and U22449 (N_22449,N_22391,N_22266);
nor U22450 (N_22450,N_22274,N_22210);
nor U22451 (N_22451,N_22381,N_22275);
and U22452 (N_22452,N_22396,N_22359);
and U22453 (N_22453,N_22372,N_22259);
nor U22454 (N_22454,N_22373,N_22332);
nand U22455 (N_22455,N_22276,N_22324);
nand U22456 (N_22456,N_22262,N_22349);
xor U22457 (N_22457,N_22318,N_22204);
xor U22458 (N_22458,N_22236,N_22384);
or U22459 (N_22459,N_22272,N_22212);
nor U22460 (N_22460,N_22289,N_22299);
and U22461 (N_22461,N_22319,N_22358);
nand U22462 (N_22462,N_22269,N_22208);
xor U22463 (N_22463,N_22303,N_22277);
or U22464 (N_22464,N_22255,N_22268);
nand U22465 (N_22465,N_22390,N_22382);
nand U22466 (N_22466,N_22201,N_22379);
or U22467 (N_22467,N_22228,N_22229);
or U22468 (N_22468,N_22244,N_22342);
xnor U22469 (N_22469,N_22305,N_22385);
nor U22470 (N_22470,N_22375,N_22351);
nand U22471 (N_22471,N_22350,N_22360);
or U22472 (N_22472,N_22399,N_22311);
or U22473 (N_22473,N_22216,N_22302);
or U22474 (N_22474,N_22346,N_22352);
nand U22475 (N_22475,N_22222,N_22284);
xnor U22476 (N_22476,N_22290,N_22337);
xor U22477 (N_22477,N_22250,N_22363);
and U22478 (N_22478,N_22325,N_22397);
xor U22479 (N_22479,N_22347,N_22369);
and U22480 (N_22480,N_22242,N_22320);
xor U22481 (N_22481,N_22329,N_22394);
xor U22482 (N_22482,N_22354,N_22247);
nand U22483 (N_22483,N_22213,N_22380);
or U22484 (N_22484,N_22398,N_22362);
nand U22485 (N_22485,N_22310,N_22331);
and U22486 (N_22486,N_22361,N_22260);
nand U22487 (N_22487,N_22233,N_22202);
nand U22488 (N_22488,N_22295,N_22230);
nand U22489 (N_22489,N_22326,N_22308);
nor U22490 (N_22490,N_22219,N_22206);
xor U22491 (N_22491,N_22211,N_22374);
nand U22492 (N_22492,N_22280,N_22328);
nand U22493 (N_22493,N_22282,N_22336);
nand U22494 (N_22494,N_22273,N_22232);
nor U22495 (N_22495,N_22258,N_22298);
or U22496 (N_22496,N_22356,N_22263);
xor U22497 (N_22497,N_22264,N_22323);
or U22498 (N_22498,N_22365,N_22370);
and U22499 (N_22499,N_22293,N_22257);
xnor U22500 (N_22500,N_22242,N_22358);
or U22501 (N_22501,N_22381,N_22380);
and U22502 (N_22502,N_22254,N_22313);
nand U22503 (N_22503,N_22359,N_22360);
or U22504 (N_22504,N_22220,N_22335);
nor U22505 (N_22505,N_22221,N_22374);
nand U22506 (N_22506,N_22213,N_22296);
and U22507 (N_22507,N_22250,N_22319);
xnor U22508 (N_22508,N_22371,N_22381);
nand U22509 (N_22509,N_22378,N_22302);
nor U22510 (N_22510,N_22272,N_22232);
or U22511 (N_22511,N_22300,N_22228);
xor U22512 (N_22512,N_22243,N_22241);
and U22513 (N_22513,N_22200,N_22346);
nor U22514 (N_22514,N_22236,N_22318);
and U22515 (N_22515,N_22338,N_22221);
xnor U22516 (N_22516,N_22279,N_22271);
or U22517 (N_22517,N_22261,N_22366);
and U22518 (N_22518,N_22242,N_22220);
and U22519 (N_22519,N_22300,N_22207);
xor U22520 (N_22520,N_22390,N_22347);
and U22521 (N_22521,N_22320,N_22391);
and U22522 (N_22522,N_22238,N_22240);
xnor U22523 (N_22523,N_22358,N_22388);
or U22524 (N_22524,N_22376,N_22389);
and U22525 (N_22525,N_22253,N_22279);
xor U22526 (N_22526,N_22272,N_22372);
and U22527 (N_22527,N_22250,N_22334);
xor U22528 (N_22528,N_22322,N_22311);
and U22529 (N_22529,N_22359,N_22298);
xor U22530 (N_22530,N_22267,N_22300);
and U22531 (N_22531,N_22387,N_22326);
or U22532 (N_22532,N_22331,N_22399);
and U22533 (N_22533,N_22249,N_22212);
nand U22534 (N_22534,N_22325,N_22232);
and U22535 (N_22535,N_22274,N_22338);
or U22536 (N_22536,N_22329,N_22231);
nand U22537 (N_22537,N_22364,N_22256);
and U22538 (N_22538,N_22383,N_22242);
nor U22539 (N_22539,N_22294,N_22309);
xnor U22540 (N_22540,N_22345,N_22308);
nand U22541 (N_22541,N_22349,N_22350);
nor U22542 (N_22542,N_22339,N_22391);
xor U22543 (N_22543,N_22251,N_22292);
and U22544 (N_22544,N_22200,N_22341);
or U22545 (N_22545,N_22386,N_22338);
xnor U22546 (N_22546,N_22309,N_22342);
xor U22547 (N_22547,N_22291,N_22217);
nand U22548 (N_22548,N_22235,N_22361);
or U22549 (N_22549,N_22390,N_22276);
or U22550 (N_22550,N_22324,N_22290);
or U22551 (N_22551,N_22329,N_22395);
nor U22552 (N_22552,N_22338,N_22365);
or U22553 (N_22553,N_22313,N_22361);
nor U22554 (N_22554,N_22296,N_22256);
nor U22555 (N_22555,N_22361,N_22249);
xor U22556 (N_22556,N_22354,N_22386);
nand U22557 (N_22557,N_22302,N_22396);
or U22558 (N_22558,N_22319,N_22210);
nand U22559 (N_22559,N_22258,N_22289);
or U22560 (N_22560,N_22210,N_22211);
and U22561 (N_22561,N_22320,N_22386);
or U22562 (N_22562,N_22367,N_22369);
and U22563 (N_22563,N_22326,N_22270);
xnor U22564 (N_22564,N_22236,N_22366);
nand U22565 (N_22565,N_22271,N_22299);
nor U22566 (N_22566,N_22388,N_22229);
and U22567 (N_22567,N_22374,N_22297);
and U22568 (N_22568,N_22249,N_22300);
xnor U22569 (N_22569,N_22350,N_22285);
and U22570 (N_22570,N_22292,N_22366);
nor U22571 (N_22571,N_22347,N_22356);
nand U22572 (N_22572,N_22361,N_22350);
and U22573 (N_22573,N_22272,N_22201);
xnor U22574 (N_22574,N_22211,N_22396);
nand U22575 (N_22575,N_22389,N_22318);
or U22576 (N_22576,N_22236,N_22324);
nand U22577 (N_22577,N_22241,N_22372);
nor U22578 (N_22578,N_22389,N_22327);
or U22579 (N_22579,N_22305,N_22358);
and U22580 (N_22580,N_22216,N_22241);
nor U22581 (N_22581,N_22348,N_22272);
nor U22582 (N_22582,N_22213,N_22348);
nand U22583 (N_22583,N_22348,N_22311);
nor U22584 (N_22584,N_22319,N_22344);
nor U22585 (N_22585,N_22329,N_22348);
nand U22586 (N_22586,N_22257,N_22398);
nand U22587 (N_22587,N_22335,N_22251);
nand U22588 (N_22588,N_22326,N_22393);
nor U22589 (N_22589,N_22270,N_22236);
nor U22590 (N_22590,N_22345,N_22352);
nor U22591 (N_22591,N_22392,N_22211);
xnor U22592 (N_22592,N_22244,N_22341);
xnor U22593 (N_22593,N_22387,N_22298);
and U22594 (N_22594,N_22274,N_22350);
nand U22595 (N_22595,N_22359,N_22261);
nor U22596 (N_22596,N_22340,N_22282);
and U22597 (N_22597,N_22337,N_22370);
and U22598 (N_22598,N_22212,N_22219);
nand U22599 (N_22599,N_22309,N_22307);
and U22600 (N_22600,N_22550,N_22553);
nor U22601 (N_22601,N_22425,N_22431);
or U22602 (N_22602,N_22445,N_22403);
or U22603 (N_22603,N_22551,N_22429);
or U22604 (N_22604,N_22498,N_22490);
nand U22605 (N_22605,N_22497,N_22510);
or U22606 (N_22606,N_22557,N_22484);
nand U22607 (N_22607,N_22458,N_22471);
nor U22608 (N_22608,N_22548,N_22584);
and U22609 (N_22609,N_22528,N_22437);
nor U22610 (N_22610,N_22424,N_22447);
or U22611 (N_22611,N_22442,N_22569);
and U22612 (N_22612,N_22438,N_22520);
xor U22613 (N_22613,N_22493,N_22521);
nor U22614 (N_22614,N_22596,N_22478);
nor U22615 (N_22615,N_22467,N_22430);
and U22616 (N_22616,N_22573,N_22441);
and U22617 (N_22617,N_22549,N_22411);
nand U22618 (N_22618,N_22558,N_22465);
or U22619 (N_22619,N_22402,N_22541);
xnor U22620 (N_22620,N_22422,N_22433);
and U22621 (N_22621,N_22470,N_22540);
and U22622 (N_22622,N_22439,N_22426);
nor U22623 (N_22623,N_22546,N_22462);
and U22624 (N_22624,N_22556,N_22542);
and U22625 (N_22625,N_22466,N_22476);
nor U22626 (N_22626,N_22531,N_22539);
xnor U22627 (N_22627,N_22468,N_22446);
nand U22628 (N_22628,N_22566,N_22544);
nor U22629 (N_22629,N_22489,N_22527);
or U22630 (N_22630,N_22545,N_22481);
or U22631 (N_22631,N_22502,N_22524);
or U22632 (N_22632,N_22513,N_22416);
or U22633 (N_22633,N_22496,N_22554);
or U22634 (N_22634,N_22451,N_22434);
nor U22635 (N_22635,N_22594,N_22579);
or U22636 (N_22636,N_22575,N_22555);
or U22637 (N_22637,N_22488,N_22483);
or U22638 (N_22638,N_22494,N_22583);
nand U22639 (N_22639,N_22532,N_22459);
nand U22640 (N_22640,N_22518,N_22537);
and U22641 (N_22641,N_22512,N_22593);
nor U22642 (N_22642,N_22595,N_22576);
or U22643 (N_22643,N_22519,N_22508);
nand U22644 (N_22644,N_22577,N_22535);
or U22645 (N_22645,N_22410,N_22506);
or U22646 (N_22646,N_22589,N_22412);
xor U22647 (N_22647,N_22507,N_22464);
xnor U22648 (N_22648,N_22563,N_22485);
and U22649 (N_22649,N_22590,N_22454);
nor U22650 (N_22650,N_22449,N_22534);
nor U22651 (N_22651,N_22533,N_22444);
xor U22652 (N_22652,N_22565,N_22413);
and U22653 (N_22653,N_22404,N_22419);
nor U22654 (N_22654,N_22516,N_22479);
or U22655 (N_22655,N_22503,N_22591);
nand U22656 (N_22656,N_22456,N_22435);
xor U22657 (N_22657,N_22529,N_22480);
xnor U22658 (N_22658,N_22486,N_22517);
nor U22659 (N_22659,N_22580,N_22515);
nor U22660 (N_22660,N_22559,N_22564);
or U22661 (N_22661,N_22582,N_22574);
nor U22662 (N_22662,N_22504,N_22585);
nand U22663 (N_22663,N_22436,N_22588);
or U22664 (N_22664,N_22423,N_22561);
xnor U22665 (N_22665,N_22409,N_22572);
nand U22666 (N_22666,N_22450,N_22511);
nand U22667 (N_22667,N_22432,N_22567);
nand U22668 (N_22668,N_22514,N_22405);
and U22669 (N_22669,N_22455,N_22525);
nand U22670 (N_22670,N_22536,N_22509);
xnor U22671 (N_22671,N_22560,N_22453);
or U22672 (N_22672,N_22420,N_22501);
xor U22673 (N_22673,N_22400,N_22407);
or U22674 (N_22674,N_22530,N_22408);
nand U22675 (N_22675,N_22587,N_22473);
xnor U22676 (N_22676,N_22570,N_22568);
nor U22677 (N_22677,N_22461,N_22562);
nand U22678 (N_22678,N_22463,N_22597);
and U22679 (N_22679,N_22469,N_22415);
nand U22680 (N_22680,N_22571,N_22475);
xnor U22681 (N_22681,N_22523,N_22505);
and U22682 (N_22682,N_22428,N_22452);
nand U22683 (N_22683,N_22586,N_22443);
and U22684 (N_22684,N_22460,N_22492);
or U22685 (N_22685,N_22500,N_22547);
or U22686 (N_22686,N_22522,N_22538);
or U22687 (N_22687,N_22418,N_22487);
nand U22688 (N_22688,N_22499,N_22491);
nor U22689 (N_22689,N_22526,N_22457);
nor U22690 (N_22690,N_22414,N_22440);
nor U22691 (N_22691,N_22482,N_22417);
or U22692 (N_22692,N_22474,N_22448);
xor U22693 (N_22693,N_22598,N_22472);
or U22694 (N_22694,N_22581,N_22592);
nor U22695 (N_22695,N_22543,N_22427);
and U22696 (N_22696,N_22578,N_22477);
nand U22697 (N_22697,N_22599,N_22406);
and U22698 (N_22698,N_22552,N_22495);
xnor U22699 (N_22699,N_22401,N_22421);
xor U22700 (N_22700,N_22484,N_22512);
nor U22701 (N_22701,N_22534,N_22590);
and U22702 (N_22702,N_22447,N_22488);
xor U22703 (N_22703,N_22414,N_22489);
and U22704 (N_22704,N_22564,N_22587);
nor U22705 (N_22705,N_22497,N_22490);
xnor U22706 (N_22706,N_22416,N_22581);
or U22707 (N_22707,N_22467,N_22531);
or U22708 (N_22708,N_22513,N_22406);
or U22709 (N_22709,N_22556,N_22575);
nor U22710 (N_22710,N_22457,N_22471);
xnor U22711 (N_22711,N_22544,N_22509);
xnor U22712 (N_22712,N_22470,N_22418);
and U22713 (N_22713,N_22530,N_22552);
nor U22714 (N_22714,N_22570,N_22439);
xor U22715 (N_22715,N_22445,N_22585);
or U22716 (N_22716,N_22513,N_22555);
xor U22717 (N_22717,N_22502,N_22499);
and U22718 (N_22718,N_22448,N_22491);
and U22719 (N_22719,N_22570,N_22581);
or U22720 (N_22720,N_22583,N_22477);
and U22721 (N_22721,N_22528,N_22537);
or U22722 (N_22722,N_22587,N_22502);
xnor U22723 (N_22723,N_22415,N_22575);
nor U22724 (N_22724,N_22551,N_22434);
and U22725 (N_22725,N_22405,N_22556);
xnor U22726 (N_22726,N_22477,N_22558);
and U22727 (N_22727,N_22444,N_22555);
nor U22728 (N_22728,N_22571,N_22507);
and U22729 (N_22729,N_22429,N_22421);
nor U22730 (N_22730,N_22583,N_22567);
nor U22731 (N_22731,N_22480,N_22509);
nand U22732 (N_22732,N_22557,N_22496);
xnor U22733 (N_22733,N_22470,N_22410);
nor U22734 (N_22734,N_22592,N_22463);
and U22735 (N_22735,N_22464,N_22409);
and U22736 (N_22736,N_22466,N_22555);
or U22737 (N_22737,N_22458,N_22588);
or U22738 (N_22738,N_22461,N_22445);
and U22739 (N_22739,N_22498,N_22569);
nor U22740 (N_22740,N_22519,N_22562);
xnor U22741 (N_22741,N_22589,N_22563);
and U22742 (N_22742,N_22478,N_22554);
and U22743 (N_22743,N_22476,N_22506);
or U22744 (N_22744,N_22542,N_22585);
or U22745 (N_22745,N_22488,N_22573);
nand U22746 (N_22746,N_22477,N_22432);
nor U22747 (N_22747,N_22466,N_22425);
xnor U22748 (N_22748,N_22533,N_22502);
or U22749 (N_22749,N_22450,N_22420);
nor U22750 (N_22750,N_22581,N_22573);
xnor U22751 (N_22751,N_22478,N_22529);
and U22752 (N_22752,N_22468,N_22536);
and U22753 (N_22753,N_22453,N_22577);
or U22754 (N_22754,N_22477,N_22408);
xnor U22755 (N_22755,N_22542,N_22521);
and U22756 (N_22756,N_22439,N_22524);
and U22757 (N_22757,N_22576,N_22525);
nor U22758 (N_22758,N_22528,N_22538);
nor U22759 (N_22759,N_22570,N_22497);
or U22760 (N_22760,N_22496,N_22402);
xnor U22761 (N_22761,N_22552,N_22443);
nand U22762 (N_22762,N_22432,N_22550);
nand U22763 (N_22763,N_22547,N_22573);
nor U22764 (N_22764,N_22489,N_22554);
or U22765 (N_22765,N_22492,N_22450);
xor U22766 (N_22766,N_22572,N_22486);
and U22767 (N_22767,N_22542,N_22449);
nor U22768 (N_22768,N_22553,N_22406);
nor U22769 (N_22769,N_22563,N_22584);
nor U22770 (N_22770,N_22449,N_22588);
or U22771 (N_22771,N_22481,N_22598);
or U22772 (N_22772,N_22474,N_22531);
and U22773 (N_22773,N_22422,N_22402);
or U22774 (N_22774,N_22445,N_22416);
xnor U22775 (N_22775,N_22599,N_22438);
nand U22776 (N_22776,N_22491,N_22435);
nor U22777 (N_22777,N_22407,N_22417);
or U22778 (N_22778,N_22527,N_22447);
or U22779 (N_22779,N_22538,N_22500);
nand U22780 (N_22780,N_22421,N_22481);
or U22781 (N_22781,N_22544,N_22416);
or U22782 (N_22782,N_22455,N_22462);
and U22783 (N_22783,N_22469,N_22540);
or U22784 (N_22784,N_22460,N_22582);
xor U22785 (N_22785,N_22598,N_22525);
xor U22786 (N_22786,N_22467,N_22449);
nand U22787 (N_22787,N_22473,N_22575);
nand U22788 (N_22788,N_22504,N_22437);
and U22789 (N_22789,N_22447,N_22588);
and U22790 (N_22790,N_22439,N_22461);
and U22791 (N_22791,N_22413,N_22541);
or U22792 (N_22792,N_22480,N_22468);
or U22793 (N_22793,N_22456,N_22551);
xnor U22794 (N_22794,N_22557,N_22410);
xor U22795 (N_22795,N_22581,N_22442);
nor U22796 (N_22796,N_22450,N_22537);
nor U22797 (N_22797,N_22407,N_22522);
nor U22798 (N_22798,N_22450,N_22436);
xnor U22799 (N_22799,N_22496,N_22542);
and U22800 (N_22800,N_22689,N_22747);
and U22801 (N_22801,N_22608,N_22642);
nor U22802 (N_22802,N_22783,N_22764);
or U22803 (N_22803,N_22659,N_22750);
nor U22804 (N_22804,N_22640,N_22768);
nor U22805 (N_22805,N_22675,N_22778);
xnor U22806 (N_22806,N_22795,N_22719);
xor U22807 (N_22807,N_22792,N_22717);
nor U22808 (N_22808,N_22767,N_22601);
and U22809 (N_22809,N_22623,N_22604);
nor U22810 (N_22810,N_22603,N_22761);
nor U22811 (N_22811,N_22686,N_22683);
nand U22812 (N_22812,N_22711,N_22721);
and U22813 (N_22813,N_22753,N_22724);
nor U22814 (N_22814,N_22664,N_22631);
nand U22815 (N_22815,N_22618,N_22799);
nand U22816 (N_22816,N_22648,N_22622);
nand U22817 (N_22817,N_22720,N_22661);
and U22818 (N_22818,N_22674,N_22679);
nand U22819 (N_22819,N_22716,N_22709);
nor U22820 (N_22820,N_22692,N_22676);
and U22821 (N_22821,N_22744,N_22673);
and U22822 (N_22822,N_22762,N_22777);
nor U22823 (N_22823,N_22649,N_22699);
nand U22824 (N_22824,N_22639,N_22791);
and U22825 (N_22825,N_22616,N_22663);
xnor U22826 (N_22826,N_22670,N_22650);
xor U22827 (N_22827,N_22694,N_22737);
or U22828 (N_22828,N_22605,N_22630);
nand U22829 (N_22829,N_22656,N_22684);
or U22830 (N_22830,N_22714,N_22697);
and U22831 (N_22831,N_22621,N_22730);
nor U22832 (N_22832,N_22669,N_22624);
or U22833 (N_22833,N_22695,N_22627);
xor U22834 (N_22834,N_22797,N_22609);
and U22835 (N_22835,N_22757,N_22781);
xor U22836 (N_22836,N_22643,N_22731);
and U22837 (N_22837,N_22790,N_22789);
xor U22838 (N_22838,N_22776,N_22617);
nor U22839 (N_22839,N_22668,N_22759);
and U22840 (N_22840,N_22615,N_22718);
and U22841 (N_22841,N_22633,N_22771);
and U22842 (N_22842,N_22727,N_22749);
or U22843 (N_22843,N_22612,N_22600);
xor U22844 (N_22844,N_22691,N_22681);
xnor U22845 (N_22845,N_22728,N_22652);
and U22846 (N_22846,N_22688,N_22754);
and U22847 (N_22847,N_22707,N_22715);
nand U22848 (N_22848,N_22756,N_22666);
or U22849 (N_22849,N_22613,N_22602);
or U22850 (N_22850,N_22638,N_22636);
nor U22851 (N_22851,N_22736,N_22770);
xor U22852 (N_22852,N_22745,N_22786);
and U22853 (N_22853,N_22733,N_22732);
and U22854 (N_22854,N_22634,N_22632);
nor U22855 (N_22855,N_22637,N_22712);
nor U22856 (N_22856,N_22700,N_22742);
or U22857 (N_22857,N_22769,N_22766);
xnor U22858 (N_22858,N_22620,N_22667);
xnor U22859 (N_22859,N_22782,N_22779);
xor U22860 (N_22860,N_22662,N_22738);
or U22861 (N_22861,N_22774,N_22696);
nor U22862 (N_22862,N_22748,N_22743);
xor U22863 (N_22863,N_22722,N_22657);
nor U22864 (N_22864,N_22693,N_22654);
and U22865 (N_22865,N_22784,N_22690);
or U22866 (N_22866,N_22702,N_22734);
and U22867 (N_22867,N_22785,N_22705);
xor U22868 (N_22868,N_22653,N_22625);
nand U22869 (N_22869,N_22704,N_22672);
nor U22870 (N_22870,N_22723,N_22796);
nor U22871 (N_22871,N_22698,N_22788);
and U22872 (N_22872,N_22687,N_22641);
nor U22873 (N_22873,N_22628,N_22752);
nor U22874 (N_22874,N_22701,N_22614);
nand U22875 (N_22875,N_22606,N_22725);
or U22876 (N_22876,N_22645,N_22706);
nand U22877 (N_22877,N_22787,N_22772);
nor U22878 (N_22878,N_22703,N_22793);
and U22879 (N_22879,N_22629,N_22610);
or U22880 (N_22880,N_22647,N_22677);
nor U22881 (N_22881,N_22798,N_22729);
nor U22882 (N_22882,N_22710,N_22611);
or U22883 (N_22883,N_22735,N_22760);
and U22884 (N_22884,N_22665,N_22671);
nand U22885 (N_22885,N_22682,N_22739);
nand U22886 (N_22886,N_22607,N_22619);
or U22887 (N_22887,N_22635,N_22773);
nand U22888 (N_22888,N_22746,N_22655);
or U22889 (N_22889,N_22646,N_22685);
nand U22890 (N_22890,N_22780,N_22626);
and U22891 (N_22891,N_22755,N_22713);
and U22892 (N_22892,N_22651,N_22726);
and U22893 (N_22893,N_22660,N_22678);
nor U22894 (N_22894,N_22741,N_22680);
nor U22895 (N_22895,N_22758,N_22644);
and U22896 (N_22896,N_22751,N_22708);
and U22897 (N_22897,N_22765,N_22794);
xnor U22898 (N_22898,N_22740,N_22763);
nand U22899 (N_22899,N_22775,N_22658);
and U22900 (N_22900,N_22683,N_22743);
nand U22901 (N_22901,N_22735,N_22782);
xnor U22902 (N_22902,N_22775,N_22652);
nor U22903 (N_22903,N_22773,N_22797);
nor U22904 (N_22904,N_22710,N_22689);
and U22905 (N_22905,N_22793,N_22600);
and U22906 (N_22906,N_22619,N_22747);
nor U22907 (N_22907,N_22706,N_22618);
or U22908 (N_22908,N_22727,N_22766);
and U22909 (N_22909,N_22764,N_22654);
nor U22910 (N_22910,N_22766,N_22701);
or U22911 (N_22911,N_22609,N_22779);
nor U22912 (N_22912,N_22606,N_22646);
nand U22913 (N_22913,N_22732,N_22711);
nand U22914 (N_22914,N_22737,N_22623);
xor U22915 (N_22915,N_22660,N_22628);
nand U22916 (N_22916,N_22659,N_22779);
nand U22917 (N_22917,N_22787,N_22676);
xor U22918 (N_22918,N_22682,N_22673);
nor U22919 (N_22919,N_22685,N_22707);
xnor U22920 (N_22920,N_22676,N_22721);
and U22921 (N_22921,N_22730,N_22743);
and U22922 (N_22922,N_22704,N_22669);
nand U22923 (N_22923,N_22793,N_22743);
or U22924 (N_22924,N_22792,N_22636);
xor U22925 (N_22925,N_22622,N_22756);
nor U22926 (N_22926,N_22619,N_22794);
nor U22927 (N_22927,N_22766,N_22742);
and U22928 (N_22928,N_22771,N_22749);
or U22929 (N_22929,N_22680,N_22665);
and U22930 (N_22930,N_22688,N_22781);
and U22931 (N_22931,N_22632,N_22775);
nor U22932 (N_22932,N_22655,N_22606);
xnor U22933 (N_22933,N_22674,N_22617);
xor U22934 (N_22934,N_22628,N_22770);
xnor U22935 (N_22935,N_22709,N_22659);
and U22936 (N_22936,N_22679,N_22755);
or U22937 (N_22937,N_22769,N_22623);
nor U22938 (N_22938,N_22796,N_22766);
xor U22939 (N_22939,N_22764,N_22741);
xnor U22940 (N_22940,N_22693,N_22757);
nor U22941 (N_22941,N_22681,N_22624);
and U22942 (N_22942,N_22669,N_22782);
nand U22943 (N_22943,N_22690,N_22675);
and U22944 (N_22944,N_22798,N_22727);
nand U22945 (N_22945,N_22654,N_22738);
nand U22946 (N_22946,N_22696,N_22727);
nand U22947 (N_22947,N_22691,N_22651);
xnor U22948 (N_22948,N_22705,N_22624);
xor U22949 (N_22949,N_22626,N_22636);
nand U22950 (N_22950,N_22766,N_22605);
nor U22951 (N_22951,N_22774,N_22760);
nand U22952 (N_22952,N_22678,N_22670);
and U22953 (N_22953,N_22761,N_22775);
or U22954 (N_22954,N_22772,N_22717);
or U22955 (N_22955,N_22669,N_22724);
nand U22956 (N_22956,N_22778,N_22722);
and U22957 (N_22957,N_22691,N_22791);
nand U22958 (N_22958,N_22767,N_22647);
or U22959 (N_22959,N_22665,N_22615);
and U22960 (N_22960,N_22670,N_22686);
nand U22961 (N_22961,N_22687,N_22625);
nor U22962 (N_22962,N_22797,N_22656);
nand U22963 (N_22963,N_22795,N_22709);
xor U22964 (N_22964,N_22724,N_22614);
xor U22965 (N_22965,N_22680,N_22789);
and U22966 (N_22966,N_22678,N_22695);
or U22967 (N_22967,N_22613,N_22793);
nand U22968 (N_22968,N_22799,N_22764);
or U22969 (N_22969,N_22664,N_22632);
nand U22970 (N_22970,N_22641,N_22700);
or U22971 (N_22971,N_22767,N_22726);
and U22972 (N_22972,N_22613,N_22794);
nor U22973 (N_22973,N_22720,N_22748);
or U22974 (N_22974,N_22667,N_22668);
and U22975 (N_22975,N_22674,N_22684);
or U22976 (N_22976,N_22741,N_22656);
xor U22977 (N_22977,N_22748,N_22719);
nor U22978 (N_22978,N_22647,N_22764);
nor U22979 (N_22979,N_22716,N_22705);
xnor U22980 (N_22980,N_22683,N_22604);
or U22981 (N_22981,N_22647,N_22778);
xor U22982 (N_22982,N_22657,N_22761);
nor U22983 (N_22983,N_22699,N_22689);
nor U22984 (N_22984,N_22662,N_22772);
xor U22985 (N_22985,N_22763,N_22772);
nand U22986 (N_22986,N_22657,N_22762);
or U22987 (N_22987,N_22784,N_22737);
nor U22988 (N_22988,N_22617,N_22793);
or U22989 (N_22989,N_22717,N_22766);
or U22990 (N_22990,N_22697,N_22660);
xnor U22991 (N_22991,N_22752,N_22621);
or U22992 (N_22992,N_22614,N_22711);
xnor U22993 (N_22993,N_22663,N_22639);
nor U22994 (N_22994,N_22792,N_22731);
and U22995 (N_22995,N_22643,N_22769);
and U22996 (N_22996,N_22622,N_22708);
nor U22997 (N_22997,N_22659,N_22743);
or U22998 (N_22998,N_22739,N_22792);
or U22999 (N_22999,N_22659,N_22781);
nand U23000 (N_23000,N_22821,N_22979);
nand U23001 (N_23001,N_22983,N_22814);
nand U23002 (N_23002,N_22966,N_22980);
or U23003 (N_23003,N_22865,N_22887);
nor U23004 (N_23004,N_22806,N_22815);
nand U23005 (N_23005,N_22990,N_22879);
or U23006 (N_23006,N_22803,N_22846);
or U23007 (N_23007,N_22858,N_22992);
nand U23008 (N_23008,N_22809,N_22948);
and U23009 (N_23009,N_22859,N_22964);
xnor U23010 (N_23010,N_22951,N_22974);
xnor U23011 (N_23011,N_22949,N_22971);
nand U23012 (N_23012,N_22837,N_22968);
xor U23013 (N_23013,N_22952,N_22900);
or U23014 (N_23014,N_22923,N_22993);
nand U23015 (N_23015,N_22870,N_22902);
nor U23016 (N_23016,N_22832,N_22978);
nand U23017 (N_23017,N_22824,N_22826);
and U23018 (N_23018,N_22972,N_22945);
or U23019 (N_23019,N_22893,N_22875);
and U23020 (N_23020,N_22871,N_22955);
and U23021 (N_23021,N_22867,N_22903);
nor U23022 (N_23022,N_22907,N_22954);
nor U23023 (N_23023,N_22982,N_22933);
and U23024 (N_23024,N_22841,N_22856);
or U23025 (N_23025,N_22901,N_22881);
or U23026 (N_23026,N_22931,N_22928);
nor U23027 (N_23027,N_22854,N_22976);
or U23028 (N_23028,N_22857,N_22929);
or U23029 (N_23029,N_22946,N_22831);
nand U23030 (N_23030,N_22950,N_22941);
nand U23031 (N_23031,N_22862,N_22812);
and U23032 (N_23032,N_22801,N_22961);
and U23033 (N_23033,N_22957,N_22996);
xnor U23034 (N_23034,N_22890,N_22849);
xor U23035 (N_23035,N_22823,N_22882);
or U23036 (N_23036,N_22943,N_22953);
nor U23037 (N_23037,N_22818,N_22899);
xor U23038 (N_23038,N_22851,N_22959);
or U23039 (N_23039,N_22868,N_22994);
nor U23040 (N_23040,N_22995,N_22883);
or U23041 (N_23041,N_22921,N_22897);
and U23042 (N_23042,N_22938,N_22805);
or U23043 (N_23043,N_22960,N_22936);
nor U23044 (N_23044,N_22986,N_22829);
nor U23045 (N_23045,N_22969,N_22984);
and U23046 (N_23046,N_22917,N_22885);
and U23047 (N_23047,N_22838,N_22888);
nor U23048 (N_23048,N_22898,N_22935);
nor U23049 (N_23049,N_22816,N_22991);
and U23050 (N_23050,N_22800,N_22911);
and U23051 (N_23051,N_22958,N_22834);
or U23052 (N_23052,N_22830,N_22817);
nand U23053 (N_23053,N_22988,N_22869);
xor U23054 (N_23054,N_22930,N_22910);
nand U23055 (N_23055,N_22916,N_22810);
or U23056 (N_23056,N_22934,N_22860);
and U23057 (N_23057,N_22909,N_22908);
and U23058 (N_23058,N_22915,N_22863);
xor U23059 (N_23059,N_22884,N_22876);
xnor U23060 (N_23060,N_22906,N_22820);
nand U23061 (N_23061,N_22914,N_22896);
xnor U23062 (N_23062,N_22813,N_22981);
and U23063 (N_23063,N_22874,N_22873);
nor U23064 (N_23064,N_22866,N_22963);
or U23065 (N_23065,N_22827,N_22927);
or U23066 (N_23066,N_22891,N_22872);
nand U23067 (N_23067,N_22877,N_22842);
and U23068 (N_23068,N_22926,N_22956);
nor U23069 (N_23069,N_22845,N_22836);
and U23070 (N_23070,N_22942,N_22895);
and U23071 (N_23071,N_22847,N_22886);
and U23072 (N_23072,N_22878,N_22999);
xnor U23073 (N_23073,N_22807,N_22989);
and U23074 (N_23074,N_22918,N_22844);
xnor U23075 (N_23075,N_22987,N_22973);
xor U23076 (N_23076,N_22802,N_22985);
nand U23077 (N_23077,N_22894,N_22839);
or U23078 (N_23078,N_22843,N_22925);
or U23079 (N_23079,N_22825,N_22905);
nand U23080 (N_23080,N_22904,N_22913);
xnor U23081 (N_23081,N_22944,N_22922);
nor U23082 (N_23082,N_22912,N_22819);
nor U23083 (N_23083,N_22939,N_22848);
nor U23084 (N_23084,N_22892,N_22970);
nand U23085 (N_23085,N_22822,N_22804);
and U23086 (N_23086,N_22975,N_22833);
and U23087 (N_23087,N_22962,N_22977);
nand U23088 (N_23088,N_22937,N_22840);
and U23089 (N_23089,N_22880,N_22997);
or U23090 (N_23090,N_22850,N_22853);
nor U23091 (N_23091,N_22919,N_22855);
xnor U23092 (N_23092,N_22932,N_22920);
nor U23093 (N_23093,N_22924,N_22835);
nand U23094 (N_23094,N_22828,N_22889);
xor U23095 (N_23095,N_22940,N_22947);
or U23096 (N_23096,N_22852,N_22998);
nand U23097 (N_23097,N_22811,N_22861);
or U23098 (N_23098,N_22808,N_22967);
xnor U23099 (N_23099,N_22864,N_22965);
xnor U23100 (N_23100,N_22943,N_22809);
nand U23101 (N_23101,N_22816,N_22899);
nand U23102 (N_23102,N_22924,N_22811);
and U23103 (N_23103,N_22903,N_22990);
nand U23104 (N_23104,N_22823,N_22997);
nand U23105 (N_23105,N_22987,N_22884);
nand U23106 (N_23106,N_22945,N_22854);
or U23107 (N_23107,N_22867,N_22918);
xor U23108 (N_23108,N_22855,N_22969);
or U23109 (N_23109,N_22994,N_22915);
nand U23110 (N_23110,N_22918,N_22968);
and U23111 (N_23111,N_22874,N_22803);
xor U23112 (N_23112,N_22828,N_22812);
nand U23113 (N_23113,N_22831,N_22809);
or U23114 (N_23114,N_22911,N_22858);
or U23115 (N_23115,N_22981,N_22875);
or U23116 (N_23116,N_22930,N_22981);
nand U23117 (N_23117,N_22819,N_22851);
xnor U23118 (N_23118,N_22840,N_22936);
xor U23119 (N_23119,N_22916,N_22898);
xor U23120 (N_23120,N_22811,N_22927);
xnor U23121 (N_23121,N_22859,N_22993);
xnor U23122 (N_23122,N_22859,N_22818);
or U23123 (N_23123,N_22887,N_22874);
or U23124 (N_23124,N_22822,N_22831);
and U23125 (N_23125,N_22968,N_22902);
nand U23126 (N_23126,N_22881,N_22921);
or U23127 (N_23127,N_22825,N_22887);
and U23128 (N_23128,N_22811,N_22954);
xnor U23129 (N_23129,N_22837,N_22956);
or U23130 (N_23130,N_22865,N_22880);
nand U23131 (N_23131,N_22835,N_22876);
or U23132 (N_23132,N_22854,N_22839);
or U23133 (N_23133,N_22960,N_22918);
xor U23134 (N_23134,N_22898,N_22939);
and U23135 (N_23135,N_22882,N_22907);
xor U23136 (N_23136,N_22914,N_22880);
or U23137 (N_23137,N_22964,N_22867);
nand U23138 (N_23138,N_22872,N_22925);
nor U23139 (N_23139,N_22968,N_22923);
nor U23140 (N_23140,N_22913,N_22946);
nor U23141 (N_23141,N_22866,N_22977);
and U23142 (N_23142,N_22929,N_22942);
or U23143 (N_23143,N_22985,N_22890);
nor U23144 (N_23144,N_22808,N_22911);
nand U23145 (N_23145,N_22809,N_22980);
xor U23146 (N_23146,N_22870,N_22839);
nand U23147 (N_23147,N_22849,N_22919);
or U23148 (N_23148,N_22839,N_22886);
and U23149 (N_23149,N_22828,N_22887);
nand U23150 (N_23150,N_22948,N_22985);
and U23151 (N_23151,N_22952,N_22998);
or U23152 (N_23152,N_22864,N_22929);
nand U23153 (N_23153,N_22933,N_22895);
and U23154 (N_23154,N_22837,N_22894);
or U23155 (N_23155,N_22831,N_22948);
or U23156 (N_23156,N_22913,N_22866);
and U23157 (N_23157,N_22863,N_22843);
nand U23158 (N_23158,N_22987,N_22811);
xor U23159 (N_23159,N_22872,N_22815);
xor U23160 (N_23160,N_22927,N_22840);
nand U23161 (N_23161,N_22831,N_22985);
or U23162 (N_23162,N_22902,N_22885);
and U23163 (N_23163,N_22935,N_22836);
and U23164 (N_23164,N_22859,N_22851);
xnor U23165 (N_23165,N_22941,N_22911);
and U23166 (N_23166,N_22810,N_22813);
nand U23167 (N_23167,N_22981,N_22956);
or U23168 (N_23168,N_22856,N_22863);
nor U23169 (N_23169,N_22875,N_22866);
nor U23170 (N_23170,N_22871,N_22891);
nand U23171 (N_23171,N_22909,N_22964);
nand U23172 (N_23172,N_22851,N_22911);
nor U23173 (N_23173,N_22999,N_22838);
nand U23174 (N_23174,N_22974,N_22818);
or U23175 (N_23175,N_22879,N_22994);
nand U23176 (N_23176,N_22862,N_22831);
and U23177 (N_23177,N_22848,N_22800);
nand U23178 (N_23178,N_22910,N_22911);
or U23179 (N_23179,N_22883,N_22868);
and U23180 (N_23180,N_22812,N_22858);
xor U23181 (N_23181,N_22864,N_22861);
and U23182 (N_23182,N_22958,N_22952);
nand U23183 (N_23183,N_22940,N_22803);
or U23184 (N_23184,N_22996,N_22953);
and U23185 (N_23185,N_22930,N_22813);
xnor U23186 (N_23186,N_22822,N_22930);
and U23187 (N_23187,N_22898,N_22856);
xor U23188 (N_23188,N_22967,N_22959);
xnor U23189 (N_23189,N_22805,N_22999);
nor U23190 (N_23190,N_22841,N_22864);
nand U23191 (N_23191,N_22959,N_22947);
and U23192 (N_23192,N_22961,N_22941);
or U23193 (N_23193,N_22852,N_22945);
xnor U23194 (N_23194,N_22967,N_22934);
nor U23195 (N_23195,N_22966,N_22961);
nand U23196 (N_23196,N_22815,N_22889);
or U23197 (N_23197,N_22919,N_22811);
nor U23198 (N_23198,N_22841,N_22928);
xnor U23199 (N_23199,N_22978,N_22895);
nand U23200 (N_23200,N_23176,N_23072);
nand U23201 (N_23201,N_23155,N_23062);
xnor U23202 (N_23202,N_23174,N_23011);
nand U23203 (N_23203,N_23066,N_23178);
or U23204 (N_23204,N_23167,N_23180);
or U23205 (N_23205,N_23032,N_23019);
or U23206 (N_23206,N_23024,N_23076);
and U23207 (N_23207,N_23004,N_23027);
xnor U23208 (N_23208,N_23035,N_23050);
nand U23209 (N_23209,N_23195,N_23103);
xor U23210 (N_23210,N_23157,N_23041);
and U23211 (N_23211,N_23048,N_23122);
xnor U23212 (N_23212,N_23012,N_23144);
or U23213 (N_23213,N_23057,N_23166);
nor U23214 (N_23214,N_23042,N_23110);
or U23215 (N_23215,N_23085,N_23160);
nand U23216 (N_23216,N_23086,N_23074);
nand U23217 (N_23217,N_23187,N_23156);
and U23218 (N_23218,N_23094,N_23138);
nand U23219 (N_23219,N_23111,N_23198);
xnor U23220 (N_23220,N_23083,N_23123);
nand U23221 (N_23221,N_23071,N_23133);
and U23222 (N_23222,N_23001,N_23149);
xnor U23223 (N_23223,N_23130,N_23113);
or U23224 (N_23224,N_23116,N_23164);
or U23225 (N_23225,N_23124,N_23018);
and U23226 (N_23226,N_23020,N_23080);
xnor U23227 (N_23227,N_23148,N_23095);
nand U23228 (N_23228,N_23179,N_23040);
xnor U23229 (N_23229,N_23135,N_23112);
nor U23230 (N_23230,N_23169,N_23096);
or U23231 (N_23231,N_23127,N_23092);
or U23232 (N_23232,N_23059,N_23049);
xor U23233 (N_23233,N_23044,N_23090);
nand U23234 (N_23234,N_23115,N_23191);
nand U23235 (N_23235,N_23053,N_23196);
nor U23236 (N_23236,N_23182,N_23104);
xor U23237 (N_23237,N_23039,N_23177);
nor U23238 (N_23238,N_23163,N_23189);
nand U23239 (N_23239,N_23052,N_23075);
or U23240 (N_23240,N_23109,N_23030);
and U23241 (N_23241,N_23036,N_23014);
nor U23242 (N_23242,N_23098,N_23134);
nand U23243 (N_23243,N_23100,N_23153);
or U23244 (N_23244,N_23046,N_23089);
and U23245 (N_23245,N_23070,N_23126);
nor U23246 (N_23246,N_23031,N_23136);
and U23247 (N_23247,N_23151,N_23033);
nor U23248 (N_23248,N_23114,N_23025);
xnor U23249 (N_23249,N_23056,N_23121);
nor U23250 (N_23250,N_23101,N_23088);
and U23251 (N_23251,N_23063,N_23184);
nor U23252 (N_23252,N_23162,N_23125);
and U23253 (N_23253,N_23007,N_23165);
xor U23254 (N_23254,N_23181,N_23051);
xor U23255 (N_23255,N_23108,N_23009);
or U23256 (N_23256,N_23190,N_23161);
and U23257 (N_23257,N_23168,N_23064);
nand U23258 (N_23258,N_23137,N_23026);
and U23259 (N_23259,N_23159,N_23006);
nand U23260 (N_23260,N_23139,N_23060);
nand U23261 (N_23261,N_23141,N_23034);
and U23262 (N_23262,N_23084,N_23154);
and U23263 (N_23263,N_23175,N_23017);
nor U23264 (N_23264,N_23147,N_23188);
or U23265 (N_23265,N_23091,N_23058);
nor U23266 (N_23266,N_23037,N_23023);
or U23267 (N_23267,N_23128,N_23077);
and U23268 (N_23268,N_23069,N_23106);
nor U23269 (N_23269,N_23003,N_23183);
xor U23270 (N_23270,N_23118,N_23132);
or U23271 (N_23271,N_23073,N_23005);
xor U23272 (N_23272,N_23172,N_23068);
xor U23273 (N_23273,N_23061,N_23143);
xor U23274 (N_23274,N_23199,N_23140);
nor U23275 (N_23275,N_23105,N_23120);
nand U23276 (N_23276,N_23185,N_23170);
nand U23277 (N_23277,N_23158,N_23081);
and U23278 (N_23278,N_23093,N_23067);
or U23279 (N_23279,N_23119,N_23099);
or U23280 (N_23280,N_23002,N_23150);
nand U23281 (N_23281,N_23008,N_23079);
and U23282 (N_23282,N_23029,N_23192);
nand U23283 (N_23283,N_23145,N_23047);
nand U23284 (N_23284,N_23054,N_23013);
or U23285 (N_23285,N_23193,N_23117);
nand U23286 (N_23286,N_23107,N_23065);
nor U23287 (N_23287,N_23082,N_23010);
xor U23288 (N_23288,N_23087,N_23173);
or U23289 (N_23289,N_23038,N_23021);
nand U23290 (N_23290,N_23055,N_23078);
and U23291 (N_23291,N_23022,N_23186);
nand U23292 (N_23292,N_23015,N_23146);
or U23293 (N_23293,N_23197,N_23097);
xnor U23294 (N_23294,N_23043,N_23016);
nor U23295 (N_23295,N_23102,N_23194);
or U23296 (N_23296,N_23000,N_23142);
nand U23297 (N_23297,N_23152,N_23171);
or U23298 (N_23298,N_23129,N_23045);
xnor U23299 (N_23299,N_23028,N_23131);
and U23300 (N_23300,N_23062,N_23071);
nand U23301 (N_23301,N_23139,N_23115);
or U23302 (N_23302,N_23078,N_23113);
and U23303 (N_23303,N_23143,N_23010);
and U23304 (N_23304,N_23178,N_23126);
nand U23305 (N_23305,N_23127,N_23002);
or U23306 (N_23306,N_23177,N_23185);
xnor U23307 (N_23307,N_23154,N_23147);
nand U23308 (N_23308,N_23073,N_23058);
nand U23309 (N_23309,N_23006,N_23053);
and U23310 (N_23310,N_23090,N_23125);
and U23311 (N_23311,N_23133,N_23011);
nor U23312 (N_23312,N_23095,N_23142);
and U23313 (N_23313,N_23179,N_23016);
and U23314 (N_23314,N_23007,N_23156);
nand U23315 (N_23315,N_23163,N_23078);
or U23316 (N_23316,N_23065,N_23036);
nand U23317 (N_23317,N_23066,N_23143);
nor U23318 (N_23318,N_23036,N_23140);
nand U23319 (N_23319,N_23028,N_23081);
nor U23320 (N_23320,N_23045,N_23168);
xor U23321 (N_23321,N_23096,N_23151);
nor U23322 (N_23322,N_23095,N_23145);
xnor U23323 (N_23323,N_23087,N_23081);
nor U23324 (N_23324,N_23007,N_23080);
nor U23325 (N_23325,N_23166,N_23199);
or U23326 (N_23326,N_23142,N_23160);
and U23327 (N_23327,N_23187,N_23064);
and U23328 (N_23328,N_23032,N_23002);
nand U23329 (N_23329,N_23026,N_23122);
nor U23330 (N_23330,N_23183,N_23187);
and U23331 (N_23331,N_23026,N_23090);
nor U23332 (N_23332,N_23133,N_23156);
nor U23333 (N_23333,N_23187,N_23005);
nor U23334 (N_23334,N_23023,N_23121);
or U23335 (N_23335,N_23101,N_23080);
nand U23336 (N_23336,N_23137,N_23107);
or U23337 (N_23337,N_23053,N_23125);
nand U23338 (N_23338,N_23082,N_23178);
nor U23339 (N_23339,N_23049,N_23121);
or U23340 (N_23340,N_23198,N_23007);
nand U23341 (N_23341,N_23154,N_23128);
or U23342 (N_23342,N_23164,N_23158);
nor U23343 (N_23343,N_23144,N_23157);
or U23344 (N_23344,N_23072,N_23198);
and U23345 (N_23345,N_23179,N_23114);
xor U23346 (N_23346,N_23139,N_23158);
and U23347 (N_23347,N_23025,N_23044);
and U23348 (N_23348,N_23149,N_23137);
or U23349 (N_23349,N_23003,N_23190);
and U23350 (N_23350,N_23117,N_23141);
or U23351 (N_23351,N_23015,N_23118);
or U23352 (N_23352,N_23011,N_23005);
and U23353 (N_23353,N_23170,N_23020);
or U23354 (N_23354,N_23052,N_23181);
nor U23355 (N_23355,N_23060,N_23063);
xnor U23356 (N_23356,N_23197,N_23053);
nor U23357 (N_23357,N_23037,N_23076);
or U23358 (N_23358,N_23025,N_23115);
xnor U23359 (N_23359,N_23009,N_23134);
and U23360 (N_23360,N_23066,N_23116);
nand U23361 (N_23361,N_23166,N_23055);
or U23362 (N_23362,N_23171,N_23044);
or U23363 (N_23363,N_23117,N_23066);
or U23364 (N_23364,N_23162,N_23122);
or U23365 (N_23365,N_23085,N_23026);
nor U23366 (N_23366,N_23023,N_23154);
nor U23367 (N_23367,N_23079,N_23067);
nor U23368 (N_23368,N_23102,N_23061);
xor U23369 (N_23369,N_23068,N_23098);
xnor U23370 (N_23370,N_23014,N_23049);
nor U23371 (N_23371,N_23046,N_23194);
nand U23372 (N_23372,N_23037,N_23102);
and U23373 (N_23373,N_23129,N_23105);
or U23374 (N_23374,N_23089,N_23075);
xor U23375 (N_23375,N_23022,N_23091);
and U23376 (N_23376,N_23192,N_23003);
nor U23377 (N_23377,N_23189,N_23063);
and U23378 (N_23378,N_23127,N_23034);
nor U23379 (N_23379,N_23149,N_23156);
nand U23380 (N_23380,N_23191,N_23061);
and U23381 (N_23381,N_23033,N_23188);
xor U23382 (N_23382,N_23099,N_23135);
nor U23383 (N_23383,N_23190,N_23100);
xnor U23384 (N_23384,N_23182,N_23070);
nand U23385 (N_23385,N_23146,N_23160);
nand U23386 (N_23386,N_23187,N_23124);
xnor U23387 (N_23387,N_23009,N_23187);
nor U23388 (N_23388,N_23041,N_23060);
nor U23389 (N_23389,N_23156,N_23120);
or U23390 (N_23390,N_23191,N_23113);
xor U23391 (N_23391,N_23179,N_23087);
nand U23392 (N_23392,N_23195,N_23118);
nand U23393 (N_23393,N_23153,N_23077);
or U23394 (N_23394,N_23108,N_23006);
nand U23395 (N_23395,N_23101,N_23028);
nand U23396 (N_23396,N_23122,N_23168);
xnor U23397 (N_23397,N_23070,N_23190);
nand U23398 (N_23398,N_23064,N_23034);
or U23399 (N_23399,N_23005,N_23003);
nor U23400 (N_23400,N_23242,N_23306);
xor U23401 (N_23401,N_23334,N_23340);
xnor U23402 (N_23402,N_23330,N_23368);
or U23403 (N_23403,N_23275,N_23345);
xor U23404 (N_23404,N_23256,N_23392);
nand U23405 (N_23405,N_23269,N_23273);
nor U23406 (N_23406,N_23315,N_23372);
nor U23407 (N_23407,N_23290,N_23332);
or U23408 (N_23408,N_23227,N_23270);
nand U23409 (N_23409,N_23311,N_23224);
xor U23410 (N_23410,N_23339,N_23376);
and U23411 (N_23411,N_23329,N_23302);
nand U23412 (N_23412,N_23327,N_23338);
nor U23413 (N_23413,N_23324,N_23211);
nor U23414 (N_23414,N_23346,N_23397);
nand U23415 (N_23415,N_23336,N_23285);
and U23416 (N_23416,N_23305,N_23284);
nor U23417 (N_23417,N_23205,N_23279);
xnor U23418 (N_23418,N_23248,N_23221);
nand U23419 (N_23419,N_23264,N_23274);
xnor U23420 (N_23420,N_23231,N_23283);
xnor U23421 (N_23421,N_23257,N_23241);
nand U23422 (N_23422,N_23371,N_23260);
nand U23423 (N_23423,N_23277,N_23355);
nand U23424 (N_23424,N_23230,N_23281);
or U23425 (N_23425,N_23347,N_23328);
nor U23426 (N_23426,N_23391,N_23249);
or U23427 (N_23427,N_23232,N_23208);
xor U23428 (N_23428,N_23335,N_23363);
nor U23429 (N_23429,N_23310,N_23389);
and U23430 (N_23430,N_23250,N_23353);
and U23431 (N_23431,N_23237,N_23265);
and U23432 (N_23432,N_23351,N_23243);
or U23433 (N_23433,N_23331,N_23276);
nor U23434 (N_23434,N_23268,N_23223);
nor U23435 (N_23435,N_23225,N_23254);
nand U23436 (N_23436,N_23228,N_23359);
nor U23437 (N_23437,N_23398,N_23291);
xnor U23438 (N_23438,N_23271,N_23222);
nor U23439 (N_23439,N_23364,N_23350);
nor U23440 (N_23440,N_23362,N_23356);
nand U23441 (N_23441,N_23213,N_23282);
nand U23442 (N_23442,N_23263,N_23344);
or U23443 (N_23443,N_23220,N_23236);
and U23444 (N_23444,N_23233,N_23289);
nor U23445 (N_23445,N_23394,N_23320);
and U23446 (N_23446,N_23323,N_23301);
and U23447 (N_23447,N_23349,N_23367);
nand U23448 (N_23448,N_23258,N_23203);
nor U23449 (N_23449,N_23385,N_23293);
or U23450 (N_23450,N_23202,N_23206);
nor U23451 (N_23451,N_23369,N_23292);
nor U23452 (N_23452,N_23266,N_23370);
or U23453 (N_23453,N_23382,N_23218);
nor U23454 (N_23454,N_23209,N_23316);
xor U23455 (N_23455,N_23314,N_23337);
nand U23456 (N_23456,N_23333,N_23272);
nand U23457 (N_23457,N_23381,N_23267);
xnor U23458 (N_23458,N_23318,N_23212);
and U23459 (N_23459,N_23360,N_23380);
nor U23460 (N_23460,N_23321,N_23378);
and U23461 (N_23461,N_23298,N_23294);
xor U23462 (N_23462,N_23200,N_23247);
xnor U23463 (N_23463,N_23280,N_23251);
nand U23464 (N_23464,N_23245,N_23357);
or U23465 (N_23465,N_23325,N_23217);
xor U23466 (N_23466,N_23216,N_23393);
and U23467 (N_23467,N_23375,N_23384);
nor U23468 (N_23468,N_23296,N_23210);
nor U23469 (N_23469,N_23322,N_23383);
and U23470 (N_23470,N_23244,N_23354);
or U23471 (N_23471,N_23259,N_23309);
nand U23472 (N_23472,N_23238,N_23304);
and U23473 (N_23473,N_23229,N_23255);
and U23474 (N_23474,N_23343,N_23240);
nor U23475 (N_23475,N_23379,N_23361);
and U23476 (N_23476,N_23396,N_23313);
and U23477 (N_23477,N_23286,N_23317);
nor U23478 (N_23478,N_23300,N_23307);
nor U23479 (N_23479,N_23219,N_23308);
nand U23480 (N_23480,N_23365,N_23295);
nor U23481 (N_23481,N_23377,N_23387);
xnor U23482 (N_23482,N_23246,N_23366);
xor U23483 (N_23483,N_23261,N_23395);
nor U23484 (N_23484,N_23374,N_23342);
nand U23485 (N_23485,N_23390,N_23201);
xnor U23486 (N_23486,N_23303,N_23288);
nor U23487 (N_23487,N_23253,N_23252);
nand U23488 (N_23488,N_23399,N_23341);
xor U23489 (N_23489,N_23348,N_23299);
nor U23490 (N_23490,N_23262,N_23239);
xnor U23491 (N_23491,N_23278,N_23207);
nor U23492 (N_23492,N_23358,N_23386);
nand U23493 (N_23493,N_23388,N_23204);
xnor U23494 (N_23494,N_23326,N_23226);
nand U23495 (N_23495,N_23234,N_23319);
and U23496 (N_23496,N_23214,N_23287);
or U23497 (N_23497,N_23352,N_23373);
or U23498 (N_23498,N_23235,N_23297);
nor U23499 (N_23499,N_23312,N_23215);
nor U23500 (N_23500,N_23269,N_23203);
nand U23501 (N_23501,N_23321,N_23296);
nor U23502 (N_23502,N_23288,N_23381);
or U23503 (N_23503,N_23326,N_23245);
or U23504 (N_23504,N_23300,N_23379);
and U23505 (N_23505,N_23322,N_23321);
nor U23506 (N_23506,N_23326,N_23319);
and U23507 (N_23507,N_23222,N_23395);
nand U23508 (N_23508,N_23216,N_23355);
nand U23509 (N_23509,N_23372,N_23324);
nand U23510 (N_23510,N_23313,N_23325);
or U23511 (N_23511,N_23218,N_23261);
and U23512 (N_23512,N_23395,N_23208);
or U23513 (N_23513,N_23373,N_23243);
xor U23514 (N_23514,N_23223,N_23396);
xnor U23515 (N_23515,N_23226,N_23330);
or U23516 (N_23516,N_23209,N_23387);
nand U23517 (N_23517,N_23219,N_23261);
or U23518 (N_23518,N_23344,N_23343);
xor U23519 (N_23519,N_23393,N_23357);
xnor U23520 (N_23520,N_23214,N_23273);
nand U23521 (N_23521,N_23254,N_23216);
or U23522 (N_23522,N_23347,N_23204);
or U23523 (N_23523,N_23250,N_23272);
xor U23524 (N_23524,N_23231,N_23343);
or U23525 (N_23525,N_23290,N_23342);
nor U23526 (N_23526,N_23243,N_23317);
nand U23527 (N_23527,N_23384,N_23219);
and U23528 (N_23528,N_23224,N_23231);
or U23529 (N_23529,N_23282,N_23369);
nor U23530 (N_23530,N_23356,N_23307);
and U23531 (N_23531,N_23279,N_23355);
and U23532 (N_23532,N_23310,N_23304);
xnor U23533 (N_23533,N_23342,N_23242);
or U23534 (N_23534,N_23352,N_23268);
or U23535 (N_23535,N_23231,N_23238);
nand U23536 (N_23536,N_23212,N_23364);
nand U23537 (N_23537,N_23337,N_23357);
nand U23538 (N_23538,N_23340,N_23217);
and U23539 (N_23539,N_23212,N_23251);
xnor U23540 (N_23540,N_23242,N_23246);
xnor U23541 (N_23541,N_23278,N_23367);
nand U23542 (N_23542,N_23391,N_23340);
or U23543 (N_23543,N_23235,N_23207);
nand U23544 (N_23544,N_23304,N_23201);
or U23545 (N_23545,N_23309,N_23356);
or U23546 (N_23546,N_23361,N_23231);
nor U23547 (N_23547,N_23332,N_23279);
or U23548 (N_23548,N_23211,N_23275);
nor U23549 (N_23549,N_23281,N_23267);
xor U23550 (N_23550,N_23272,N_23234);
nand U23551 (N_23551,N_23235,N_23208);
nand U23552 (N_23552,N_23371,N_23392);
and U23553 (N_23553,N_23392,N_23300);
xnor U23554 (N_23554,N_23262,N_23294);
and U23555 (N_23555,N_23224,N_23248);
nor U23556 (N_23556,N_23229,N_23297);
xor U23557 (N_23557,N_23331,N_23239);
nand U23558 (N_23558,N_23391,N_23267);
nand U23559 (N_23559,N_23376,N_23281);
nand U23560 (N_23560,N_23391,N_23392);
xnor U23561 (N_23561,N_23347,N_23315);
nor U23562 (N_23562,N_23250,N_23234);
or U23563 (N_23563,N_23276,N_23350);
nand U23564 (N_23564,N_23319,N_23207);
nor U23565 (N_23565,N_23399,N_23217);
and U23566 (N_23566,N_23234,N_23329);
or U23567 (N_23567,N_23211,N_23267);
xor U23568 (N_23568,N_23395,N_23213);
or U23569 (N_23569,N_23356,N_23237);
nand U23570 (N_23570,N_23264,N_23279);
and U23571 (N_23571,N_23272,N_23313);
or U23572 (N_23572,N_23316,N_23235);
nor U23573 (N_23573,N_23244,N_23298);
or U23574 (N_23574,N_23222,N_23263);
or U23575 (N_23575,N_23392,N_23304);
nor U23576 (N_23576,N_23276,N_23377);
or U23577 (N_23577,N_23248,N_23205);
nand U23578 (N_23578,N_23354,N_23284);
nand U23579 (N_23579,N_23208,N_23264);
or U23580 (N_23580,N_23227,N_23204);
nand U23581 (N_23581,N_23352,N_23323);
nor U23582 (N_23582,N_23288,N_23234);
nand U23583 (N_23583,N_23290,N_23398);
or U23584 (N_23584,N_23354,N_23253);
or U23585 (N_23585,N_23218,N_23281);
and U23586 (N_23586,N_23382,N_23352);
xor U23587 (N_23587,N_23242,N_23346);
and U23588 (N_23588,N_23293,N_23320);
nor U23589 (N_23589,N_23352,N_23357);
or U23590 (N_23590,N_23300,N_23327);
nand U23591 (N_23591,N_23293,N_23372);
and U23592 (N_23592,N_23222,N_23324);
nor U23593 (N_23593,N_23236,N_23395);
xor U23594 (N_23594,N_23386,N_23242);
and U23595 (N_23595,N_23362,N_23329);
or U23596 (N_23596,N_23248,N_23312);
or U23597 (N_23597,N_23356,N_23282);
or U23598 (N_23598,N_23370,N_23354);
or U23599 (N_23599,N_23311,N_23214);
nor U23600 (N_23600,N_23588,N_23501);
nor U23601 (N_23601,N_23579,N_23544);
or U23602 (N_23602,N_23516,N_23446);
or U23603 (N_23603,N_23570,N_23481);
and U23604 (N_23604,N_23448,N_23453);
or U23605 (N_23605,N_23592,N_23580);
or U23606 (N_23606,N_23495,N_23542);
or U23607 (N_23607,N_23566,N_23488);
and U23608 (N_23608,N_23530,N_23547);
and U23609 (N_23609,N_23513,N_23480);
and U23610 (N_23610,N_23593,N_23478);
nand U23611 (N_23611,N_23454,N_23496);
or U23612 (N_23612,N_23499,N_23461);
xnor U23613 (N_23613,N_23440,N_23597);
and U23614 (N_23614,N_23503,N_23517);
xnor U23615 (N_23615,N_23436,N_23466);
nor U23616 (N_23616,N_23443,N_23538);
xnor U23617 (N_23617,N_23489,N_23549);
nor U23618 (N_23618,N_23582,N_23458);
xor U23619 (N_23619,N_23433,N_23557);
nor U23620 (N_23620,N_23432,N_23509);
nor U23621 (N_23621,N_23518,N_23474);
nand U23622 (N_23622,N_23569,N_23519);
and U23623 (N_23623,N_23528,N_23429);
xnor U23624 (N_23624,N_23449,N_23545);
or U23625 (N_23625,N_23546,N_23423);
or U23626 (N_23626,N_23486,N_23533);
or U23627 (N_23627,N_23548,N_23527);
and U23628 (N_23628,N_23400,N_23441);
nor U23629 (N_23629,N_23438,N_23491);
nor U23630 (N_23630,N_23490,N_23583);
nand U23631 (N_23631,N_23596,N_23437);
nor U23632 (N_23632,N_23598,N_23444);
nand U23633 (N_23633,N_23567,N_23554);
xnor U23634 (N_23634,N_23418,N_23417);
nand U23635 (N_23635,N_23502,N_23492);
xnor U23636 (N_23636,N_23416,N_23479);
nor U23637 (N_23637,N_23578,N_23531);
nor U23638 (N_23638,N_23590,N_23473);
nor U23639 (N_23639,N_23435,N_23410);
nand U23640 (N_23640,N_23422,N_23482);
nand U23641 (N_23641,N_23556,N_23412);
nand U23642 (N_23642,N_23535,N_23575);
xor U23643 (N_23643,N_23468,N_23536);
nand U23644 (N_23644,N_23493,N_23512);
nor U23645 (N_23645,N_23576,N_23581);
nand U23646 (N_23646,N_23599,N_23430);
nor U23647 (N_23647,N_23476,N_23534);
nor U23648 (N_23648,N_23460,N_23463);
nand U23649 (N_23649,N_23451,N_23529);
nand U23650 (N_23650,N_23522,N_23484);
and U23651 (N_23651,N_23426,N_23439);
nor U23652 (N_23652,N_23550,N_23477);
nor U23653 (N_23653,N_23472,N_23427);
nand U23654 (N_23654,N_23541,N_23552);
and U23655 (N_23655,N_23524,N_23498);
or U23656 (N_23656,N_23521,N_23467);
nor U23657 (N_23657,N_23555,N_23471);
nand U23658 (N_23658,N_23523,N_23564);
nand U23659 (N_23659,N_23424,N_23562);
or U23660 (N_23660,N_23539,N_23526);
nand U23661 (N_23661,N_23514,N_23497);
xor U23662 (N_23662,N_23560,N_23589);
xor U23663 (N_23663,N_23540,N_23586);
or U23664 (N_23664,N_23457,N_23543);
nand U23665 (N_23665,N_23450,N_23431);
nand U23666 (N_23666,N_23500,N_23594);
and U23667 (N_23667,N_23507,N_23465);
and U23668 (N_23668,N_23574,N_23506);
or U23669 (N_23669,N_23403,N_23591);
and U23670 (N_23670,N_23456,N_23462);
or U23671 (N_23671,N_23572,N_23537);
xor U23672 (N_23672,N_23577,N_23563);
or U23673 (N_23673,N_23551,N_23464);
nor U23674 (N_23674,N_23428,N_23455);
nand U23675 (N_23675,N_23420,N_23510);
and U23676 (N_23676,N_23553,N_23413);
nor U23677 (N_23677,N_23505,N_23559);
or U23678 (N_23678,N_23402,N_23415);
nor U23679 (N_23679,N_23571,N_23404);
nand U23680 (N_23680,N_23584,N_23573);
or U23681 (N_23681,N_23520,N_23595);
nor U23682 (N_23682,N_23494,N_23504);
or U23683 (N_23683,N_23568,N_23469);
xor U23684 (N_23684,N_23452,N_23532);
xnor U23685 (N_23685,N_23447,N_23487);
nand U23686 (N_23686,N_23419,N_23442);
nor U23687 (N_23687,N_23421,N_23445);
nor U23688 (N_23688,N_23587,N_23409);
nor U23689 (N_23689,N_23459,N_23414);
xnor U23690 (N_23690,N_23425,N_23558);
or U23691 (N_23691,N_23485,N_23585);
nor U23692 (N_23692,N_23561,N_23470);
or U23693 (N_23693,N_23565,N_23434);
nand U23694 (N_23694,N_23405,N_23406);
or U23695 (N_23695,N_23408,N_23475);
xor U23696 (N_23696,N_23508,N_23411);
or U23697 (N_23697,N_23515,N_23525);
or U23698 (N_23698,N_23407,N_23511);
nor U23699 (N_23699,N_23483,N_23401);
or U23700 (N_23700,N_23458,N_23502);
nor U23701 (N_23701,N_23523,N_23487);
or U23702 (N_23702,N_23532,N_23472);
and U23703 (N_23703,N_23408,N_23500);
or U23704 (N_23704,N_23493,N_23525);
xnor U23705 (N_23705,N_23513,N_23582);
xnor U23706 (N_23706,N_23536,N_23487);
or U23707 (N_23707,N_23416,N_23419);
or U23708 (N_23708,N_23592,N_23453);
nand U23709 (N_23709,N_23430,N_23563);
nand U23710 (N_23710,N_23561,N_23415);
nand U23711 (N_23711,N_23527,N_23444);
xnor U23712 (N_23712,N_23599,N_23481);
nand U23713 (N_23713,N_23432,N_23536);
nand U23714 (N_23714,N_23471,N_23499);
xnor U23715 (N_23715,N_23512,N_23421);
nor U23716 (N_23716,N_23508,N_23494);
nand U23717 (N_23717,N_23562,N_23474);
and U23718 (N_23718,N_23531,N_23596);
or U23719 (N_23719,N_23504,N_23463);
xnor U23720 (N_23720,N_23438,N_23507);
and U23721 (N_23721,N_23506,N_23585);
and U23722 (N_23722,N_23461,N_23498);
and U23723 (N_23723,N_23561,N_23473);
or U23724 (N_23724,N_23449,N_23459);
or U23725 (N_23725,N_23407,N_23509);
and U23726 (N_23726,N_23562,N_23481);
and U23727 (N_23727,N_23468,N_23518);
or U23728 (N_23728,N_23458,N_23573);
xor U23729 (N_23729,N_23557,N_23503);
and U23730 (N_23730,N_23469,N_23501);
nand U23731 (N_23731,N_23502,N_23404);
or U23732 (N_23732,N_23584,N_23413);
or U23733 (N_23733,N_23522,N_23450);
or U23734 (N_23734,N_23563,N_23581);
xor U23735 (N_23735,N_23494,N_23460);
nand U23736 (N_23736,N_23585,N_23591);
xor U23737 (N_23737,N_23420,N_23508);
and U23738 (N_23738,N_23454,N_23522);
or U23739 (N_23739,N_23405,N_23574);
xnor U23740 (N_23740,N_23455,N_23465);
xor U23741 (N_23741,N_23562,N_23459);
or U23742 (N_23742,N_23595,N_23492);
nor U23743 (N_23743,N_23442,N_23476);
nand U23744 (N_23744,N_23440,N_23449);
nor U23745 (N_23745,N_23457,N_23517);
and U23746 (N_23746,N_23431,N_23536);
or U23747 (N_23747,N_23435,N_23415);
or U23748 (N_23748,N_23478,N_23596);
xnor U23749 (N_23749,N_23449,N_23469);
nor U23750 (N_23750,N_23416,N_23402);
and U23751 (N_23751,N_23546,N_23474);
or U23752 (N_23752,N_23481,N_23574);
nor U23753 (N_23753,N_23571,N_23455);
or U23754 (N_23754,N_23559,N_23510);
and U23755 (N_23755,N_23580,N_23455);
and U23756 (N_23756,N_23500,N_23474);
and U23757 (N_23757,N_23507,N_23517);
nand U23758 (N_23758,N_23403,N_23595);
nor U23759 (N_23759,N_23468,N_23497);
or U23760 (N_23760,N_23489,N_23514);
nand U23761 (N_23761,N_23465,N_23521);
nor U23762 (N_23762,N_23409,N_23415);
or U23763 (N_23763,N_23477,N_23421);
or U23764 (N_23764,N_23415,N_23440);
and U23765 (N_23765,N_23548,N_23546);
nor U23766 (N_23766,N_23473,N_23518);
xor U23767 (N_23767,N_23509,N_23538);
or U23768 (N_23768,N_23521,N_23502);
xor U23769 (N_23769,N_23475,N_23474);
or U23770 (N_23770,N_23433,N_23507);
or U23771 (N_23771,N_23522,N_23585);
nand U23772 (N_23772,N_23447,N_23410);
or U23773 (N_23773,N_23583,N_23404);
nor U23774 (N_23774,N_23515,N_23443);
and U23775 (N_23775,N_23517,N_23583);
nand U23776 (N_23776,N_23521,N_23472);
or U23777 (N_23777,N_23513,N_23470);
or U23778 (N_23778,N_23532,N_23502);
and U23779 (N_23779,N_23558,N_23422);
and U23780 (N_23780,N_23574,N_23596);
and U23781 (N_23781,N_23536,N_23403);
and U23782 (N_23782,N_23454,N_23502);
and U23783 (N_23783,N_23407,N_23584);
or U23784 (N_23784,N_23521,N_23515);
xnor U23785 (N_23785,N_23423,N_23545);
or U23786 (N_23786,N_23495,N_23476);
nor U23787 (N_23787,N_23590,N_23455);
xnor U23788 (N_23788,N_23537,N_23483);
or U23789 (N_23789,N_23477,N_23422);
nand U23790 (N_23790,N_23417,N_23552);
nor U23791 (N_23791,N_23417,N_23528);
nor U23792 (N_23792,N_23447,N_23552);
xnor U23793 (N_23793,N_23585,N_23477);
xnor U23794 (N_23794,N_23524,N_23517);
or U23795 (N_23795,N_23417,N_23430);
nor U23796 (N_23796,N_23500,N_23569);
or U23797 (N_23797,N_23462,N_23406);
xnor U23798 (N_23798,N_23414,N_23489);
or U23799 (N_23799,N_23515,N_23453);
nor U23800 (N_23800,N_23676,N_23702);
xnor U23801 (N_23801,N_23635,N_23709);
nand U23802 (N_23802,N_23721,N_23694);
xor U23803 (N_23803,N_23613,N_23615);
or U23804 (N_23804,N_23762,N_23682);
xnor U23805 (N_23805,N_23739,N_23792);
nor U23806 (N_23806,N_23628,N_23691);
xnor U23807 (N_23807,N_23750,N_23748);
nand U23808 (N_23808,N_23677,N_23690);
xnor U23809 (N_23809,N_23715,N_23793);
and U23810 (N_23810,N_23610,N_23678);
nand U23811 (N_23811,N_23617,N_23602);
nand U23812 (N_23812,N_23761,N_23772);
nor U23813 (N_23813,N_23708,N_23660);
nand U23814 (N_23814,N_23706,N_23714);
or U23815 (N_23815,N_23738,N_23783);
or U23816 (N_23816,N_23666,N_23695);
xnor U23817 (N_23817,N_23763,N_23625);
nor U23818 (N_23818,N_23747,N_23697);
and U23819 (N_23819,N_23681,N_23655);
and U23820 (N_23820,N_23674,N_23716);
nor U23821 (N_23821,N_23657,N_23670);
xor U23822 (N_23822,N_23760,N_23769);
nand U23823 (N_23823,N_23664,N_23774);
xnor U23824 (N_23824,N_23661,N_23600);
nand U23825 (N_23825,N_23742,N_23773);
or U23826 (N_23826,N_23645,N_23781);
or U23827 (N_23827,N_23603,N_23797);
or U23828 (N_23828,N_23638,N_23719);
nor U23829 (N_23829,N_23633,N_23786);
and U23830 (N_23830,N_23765,N_23705);
nor U23831 (N_23831,N_23731,N_23623);
or U23832 (N_23832,N_23746,N_23725);
and U23833 (N_23833,N_23640,N_23611);
or U23834 (N_23834,N_23679,N_23730);
xnor U23835 (N_23835,N_23777,N_23673);
nor U23836 (N_23836,N_23632,N_23629);
or U23837 (N_23837,N_23642,N_23794);
nor U23838 (N_23838,N_23790,N_23620);
or U23839 (N_23839,N_23624,N_23647);
xor U23840 (N_23840,N_23759,N_23718);
or U23841 (N_23841,N_23696,N_23758);
nor U23842 (N_23842,N_23771,N_23729);
nor U23843 (N_23843,N_23658,N_23728);
xor U23844 (N_23844,N_23733,N_23789);
and U23845 (N_23845,N_23631,N_23668);
nor U23846 (N_23846,N_23757,N_23654);
nor U23847 (N_23847,N_23675,N_23767);
nand U23848 (N_23848,N_23601,N_23780);
xnor U23849 (N_23849,N_23636,N_23752);
xor U23850 (N_23850,N_23639,N_23651);
nor U23851 (N_23851,N_23779,N_23604);
xnor U23852 (N_23852,N_23689,N_23768);
and U23853 (N_23853,N_23707,N_23724);
xor U23854 (N_23854,N_23699,N_23698);
or U23855 (N_23855,N_23643,N_23704);
and U23856 (N_23856,N_23741,N_23795);
or U23857 (N_23857,N_23656,N_23683);
and U23858 (N_23858,N_23778,N_23798);
nand U23859 (N_23859,N_23637,N_23693);
and U23860 (N_23860,N_23634,N_23665);
xnor U23861 (N_23861,N_23745,N_23700);
nand U23862 (N_23862,N_23616,N_23671);
xor U23863 (N_23863,N_23712,N_23717);
and U23864 (N_23864,N_23641,N_23653);
nand U23865 (N_23865,N_23650,N_23787);
nor U23866 (N_23866,N_23680,N_23764);
and U23867 (N_23867,N_23753,N_23776);
nand U23868 (N_23868,N_23732,N_23607);
or U23869 (N_23869,N_23740,N_23608);
nand U23870 (N_23870,N_23788,N_23692);
or U23871 (N_23871,N_23605,N_23737);
nor U23872 (N_23872,N_23703,N_23751);
xor U23873 (N_23873,N_23723,N_23614);
or U23874 (N_23874,N_23659,N_23722);
and U23875 (N_23875,N_23791,N_23622);
and U23876 (N_23876,N_23648,N_23685);
or U23877 (N_23877,N_23796,N_23736);
nand U23878 (N_23878,N_23652,N_23669);
nor U23879 (N_23879,N_23662,N_23619);
or U23880 (N_23880,N_23646,N_23701);
and U23881 (N_23881,N_23621,N_23687);
xnor U23882 (N_23882,N_23766,N_23756);
nor U23883 (N_23883,N_23684,N_23713);
and U23884 (N_23884,N_23784,N_23720);
nor U23885 (N_23885,N_23618,N_23606);
nand U23886 (N_23886,N_23744,N_23609);
and U23887 (N_23887,N_23710,N_23770);
xor U23888 (N_23888,N_23630,N_23749);
and U23889 (N_23889,N_23782,N_23785);
or U23890 (N_23890,N_23775,N_23755);
nand U23891 (N_23891,N_23627,N_23799);
or U23892 (N_23892,N_23711,N_23743);
xnor U23893 (N_23893,N_23644,N_23626);
nor U23894 (N_23894,N_23672,N_23734);
nor U23895 (N_23895,N_23726,N_23688);
nor U23896 (N_23896,N_23686,N_23735);
nor U23897 (N_23897,N_23727,N_23612);
nor U23898 (N_23898,N_23667,N_23663);
nor U23899 (N_23899,N_23754,N_23649);
and U23900 (N_23900,N_23721,N_23765);
nor U23901 (N_23901,N_23711,N_23669);
xnor U23902 (N_23902,N_23690,N_23641);
or U23903 (N_23903,N_23612,N_23730);
nor U23904 (N_23904,N_23724,N_23678);
nor U23905 (N_23905,N_23632,N_23635);
nor U23906 (N_23906,N_23788,N_23699);
nand U23907 (N_23907,N_23653,N_23609);
or U23908 (N_23908,N_23692,N_23781);
nand U23909 (N_23909,N_23764,N_23665);
xnor U23910 (N_23910,N_23734,N_23657);
and U23911 (N_23911,N_23775,N_23697);
xnor U23912 (N_23912,N_23624,N_23630);
or U23913 (N_23913,N_23661,N_23671);
or U23914 (N_23914,N_23793,N_23708);
and U23915 (N_23915,N_23703,N_23675);
xor U23916 (N_23916,N_23758,N_23701);
nor U23917 (N_23917,N_23647,N_23605);
and U23918 (N_23918,N_23764,N_23616);
nor U23919 (N_23919,N_23787,N_23654);
nand U23920 (N_23920,N_23713,N_23615);
and U23921 (N_23921,N_23684,N_23611);
and U23922 (N_23922,N_23797,N_23638);
xnor U23923 (N_23923,N_23623,N_23724);
xor U23924 (N_23924,N_23752,N_23782);
nand U23925 (N_23925,N_23688,N_23724);
nand U23926 (N_23926,N_23747,N_23694);
xnor U23927 (N_23927,N_23750,N_23775);
or U23928 (N_23928,N_23636,N_23622);
nor U23929 (N_23929,N_23652,N_23790);
xnor U23930 (N_23930,N_23743,N_23792);
and U23931 (N_23931,N_23752,N_23647);
xor U23932 (N_23932,N_23667,N_23717);
or U23933 (N_23933,N_23738,N_23705);
xnor U23934 (N_23934,N_23646,N_23601);
xnor U23935 (N_23935,N_23630,N_23602);
nand U23936 (N_23936,N_23610,N_23603);
or U23937 (N_23937,N_23620,N_23712);
nor U23938 (N_23938,N_23644,N_23622);
nor U23939 (N_23939,N_23731,N_23760);
nand U23940 (N_23940,N_23691,N_23664);
and U23941 (N_23941,N_23684,N_23772);
and U23942 (N_23942,N_23628,N_23748);
and U23943 (N_23943,N_23645,N_23666);
or U23944 (N_23944,N_23711,N_23744);
nand U23945 (N_23945,N_23678,N_23708);
xor U23946 (N_23946,N_23609,N_23724);
xnor U23947 (N_23947,N_23778,N_23632);
nor U23948 (N_23948,N_23687,N_23703);
and U23949 (N_23949,N_23711,N_23627);
nand U23950 (N_23950,N_23794,N_23682);
and U23951 (N_23951,N_23645,N_23725);
xnor U23952 (N_23952,N_23764,N_23600);
nand U23953 (N_23953,N_23733,N_23719);
nand U23954 (N_23954,N_23774,N_23656);
nand U23955 (N_23955,N_23640,N_23786);
xnor U23956 (N_23956,N_23707,N_23732);
or U23957 (N_23957,N_23734,N_23663);
nor U23958 (N_23958,N_23797,N_23627);
xor U23959 (N_23959,N_23718,N_23684);
nand U23960 (N_23960,N_23756,N_23691);
nand U23961 (N_23961,N_23675,N_23616);
nor U23962 (N_23962,N_23785,N_23753);
or U23963 (N_23963,N_23689,N_23646);
or U23964 (N_23964,N_23748,N_23667);
xnor U23965 (N_23965,N_23787,N_23625);
nand U23966 (N_23966,N_23750,N_23708);
nor U23967 (N_23967,N_23648,N_23725);
and U23968 (N_23968,N_23650,N_23734);
and U23969 (N_23969,N_23745,N_23730);
xor U23970 (N_23970,N_23697,N_23607);
nand U23971 (N_23971,N_23799,N_23698);
and U23972 (N_23972,N_23636,N_23641);
or U23973 (N_23973,N_23773,N_23753);
or U23974 (N_23974,N_23601,N_23710);
nand U23975 (N_23975,N_23752,N_23732);
and U23976 (N_23976,N_23713,N_23604);
nor U23977 (N_23977,N_23663,N_23732);
or U23978 (N_23978,N_23797,N_23769);
and U23979 (N_23979,N_23712,N_23638);
nor U23980 (N_23980,N_23799,N_23719);
nand U23981 (N_23981,N_23791,N_23741);
or U23982 (N_23982,N_23665,N_23635);
or U23983 (N_23983,N_23605,N_23700);
xnor U23984 (N_23984,N_23718,N_23626);
xnor U23985 (N_23985,N_23700,N_23735);
nor U23986 (N_23986,N_23605,N_23774);
nand U23987 (N_23987,N_23670,N_23764);
nand U23988 (N_23988,N_23721,N_23727);
nand U23989 (N_23989,N_23725,N_23674);
nand U23990 (N_23990,N_23724,N_23761);
or U23991 (N_23991,N_23627,N_23612);
and U23992 (N_23992,N_23776,N_23662);
nor U23993 (N_23993,N_23649,N_23753);
and U23994 (N_23994,N_23715,N_23603);
xor U23995 (N_23995,N_23706,N_23727);
xnor U23996 (N_23996,N_23734,N_23618);
and U23997 (N_23997,N_23645,N_23634);
xnor U23998 (N_23998,N_23739,N_23794);
nand U23999 (N_23999,N_23730,N_23689);
nor U24000 (N_24000,N_23933,N_23834);
and U24001 (N_24001,N_23996,N_23955);
or U24002 (N_24002,N_23942,N_23991);
nor U24003 (N_24003,N_23852,N_23995);
xnor U24004 (N_24004,N_23850,N_23838);
nand U24005 (N_24005,N_23874,N_23962);
and U24006 (N_24006,N_23988,N_23987);
or U24007 (N_24007,N_23811,N_23823);
nand U24008 (N_24008,N_23817,N_23935);
xnor U24009 (N_24009,N_23983,N_23913);
and U24010 (N_24010,N_23889,N_23865);
or U24011 (N_24011,N_23853,N_23894);
and U24012 (N_24012,N_23846,N_23974);
and U24013 (N_24013,N_23820,N_23978);
or U24014 (N_24014,N_23989,N_23867);
or U24015 (N_24015,N_23808,N_23914);
nand U24016 (N_24016,N_23931,N_23885);
or U24017 (N_24017,N_23806,N_23927);
nor U24018 (N_24018,N_23905,N_23875);
or U24019 (N_24019,N_23873,N_23814);
nand U24020 (N_24020,N_23948,N_23922);
and U24021 (N_24021,N_23803,N_23906);
and U24022 (N_24022,N_23804,N_23923);
or U24023 (N_24023,N_23925,N_23890);
or U24024 (N_24024,N_23899,N_23876);
xor U24025 (N_24025,N_23976,N_23959);
and U24026 (N_24026,N_23878,N_23815);
nand U24027 (N_24027,N_23807,N_23950);
or U24028 (N_24028,N_23810,N_23982);
xnor U24029 (N_24029,N_23980,N_23936);
and U24030 (N_24030,N_23902,N_23828);
nand U24031 (N_24031,N_23984,N_23877);
and U24032 (N_24032,N_23892,N_23891);
and U24033 (N_24033,N_23830,N_23930);
or U24034 (N_24034,N_23824,N_23845);
xor U24035 (N_24035,N_23926,N_23977);
nand U24036 (N_24036,N_23861,N_23829);
nand U24037 (N_24037,N_23896,N_23816);
nor U24038 (N_24038,N_23886,N_23985);
and U24039 (N_24039,N_23843,N_23919);
nor U24040 (N_24040,N_23941,N_23920);
nor U24041 (N_24041,N_23970,N_23897);
and U24042 (N_24042,N_23975,N_23882);
or U24043 (N_24043,N_23858,N_23837);
or U24044 (N_24044,N_23960,N_23818);
nand U24045 (N_24045,N_23871,N_23921);
nor U24046 (N_24046,N_23992,N_23822);
or U24047 (N_24047,N_23869,N_23964);
or U24048 (N_24048,N_23802,N_23883);
or U24049 (N_24049,N_23809,N_23957);
nand U24050 (N_24050,N_23842,N_23986);
and U24051 (N_24051,N_23958,N_23943);
xnor U24052 (N_24052,N_23827,N_23844);
or U24053 (N_24053,N_23847,N_23812);
nor U24054 (N_24054,N_23954,N_23893);
xnor U24055 (N_24055,N_23870,N_23934);
xnor U24056 (N_24056,N_23821,N_23912);
nor U24057 (N_24057,N_23915,N_23999);
or U24058 (N_24058,N_23813,N_23836);
nor U24059 (N_24059,N_23990,N_23872);
and U24060 (N_24060,N_23900,N_23805);
or U24061 (N_24061,N_23880,N_23833);
or U24062 (N_24062,N_23966,N_23835);
or U24063 (N_24063,N_23945,N_23911);
or U24064 (N_24064,N_23851,N_23981);
and U24065 (N_24065,N_23898,N_23916);
or U24066 (N_24066,N_23855,N_23917);
nor U24067 (N_24067,N_23863,N_23854);
or U24068 (N_24068,N_23903,N_23859);
and U24069 (N_24069,N_23961,N_23994);
or U24070 (N_24070,N_23857,N_23860);
or U24071 (N_24071,N_23848,N_23832);
and U24072 (N_24072,N_23862,N_23910);
xnor U24073 (N_24073,N_23884,N_23953);
or U24074 (N_24074,N_23952,N_23967);
nand U24075 (N_24075,N_23819,N_23826);
nand U24076 (N_24076,N_23831,N_23972);
or U24077 (N_24077,N_23868,N_23993);
and U24078 (N_24078,N_23968,N_23904);
xor U24079 (N_24079,N_23800,N_23971);
xor U24080 (N_24080,N_23888,N_23895);
nor U24081 (N_24081,N_23940,N_23944);
xnor U24082 (N_24082,N_23881,N_23998);
or U24083 (N_24083,N_23929,N_23946);
xor U24084 (N_24084,N_23928,N_23963);
xnor U24085 (N_24085,N_23973,N_23825);
nand U24086 (N_24086,N_23932,N_23887);
nor U24087 (N_24087,N_23918,N_23951);
nand U24088 (N_24088,N_23839,N_23947);
or U24089 (N_24089,N_23879,N_23938);
or U24090 (N_24090,N_23969,N_23849);
and U24091 (N_24091,N_23866,N_23939);
nand U24092 (N_24092,N_23864,N_23909);
or U24093 (N_24093,N_23840,N_23949);
nor U24094 (N_24094,N_23841,N_23979);
nand U24095 (N_24095,N_23907,N_23956);
and U24096 (N_24096,N_23801,N_23856);
nor U24097 (N_24097,N_23908,N_23901);
nor U24098 (N_24098,N_23965,N_23997);
nand U24099 (N_24099,N_23924,N_23937);
or U24100 (N_24100,N_23962,N_23998);
xnor U24101 (N_24101,N_23932,N_23897);
nor U24102 (N_24102,N_23863,N_23973);
and U24103 (N_24103,N_23966,N_23931);
nand U24104 (N_24104,N_23847,N_23915);
nand U24105 (N_24105,N_23981,N_23840);
nor U24106 (N_24106,N_23844,N_23803);
or U24107 (N_24107,N_23825,N_23996);
xor U24108 (N_24108,N_23870,N_23930);
and U24109 (N_24109,N_23816,N_23989);
nor U24110 (N_24110,N_23928,N_23887);
nand U24111 (N_24111,N_23832,N_23952);
or U24112 (N_24112,N_23895,N_23981);
nand U24113 (N_24113,N_23904,N_23914);
or U24114 (N_24114,N_23951,N_23941);
and U24115 (N_24115,N_23871,N_23812);
nor U24116 (N_24116,N_23869,N_23940);
xnor U24117 (N_24117,N_23994,N_23978);
nand U24118 (N_24118,N_23834,N_23838);
xor U24119 (N_24119,N_23806,N_23983);
xor U24120 (N_24120,N_23851,N_23943);
nand U24121 (N_24121,N_23909,N_23933);
xor U24122 (N_24122,N_23844,N_23840);
and U24123 (N_24123,N_23870,N_23885);
xnor U24124 (N_24124,N_23943,N_23875);
nand U24125 (N_24125,N_23996,N_23917);
and U24126 (N_24126,N_23882,N_23927);
or U24127 (N_24127,N_23823,N_23979);
and U24128 (N_24128,N_23849,N_23954);
or U24129 (N_24129,N_23892,N_23905);
and U24130 (N_24130,N_23875,N_23852);
and U24131 (N_24131,N_23833,N_23892);
nor U24132 (N_24132,N_23855,N_23818);
nor U24133 (N_24133,N_23977,N_23914);
and U24134 (N_24134,N_23820,N_23825);
nand U24135 (N_24135,N_23800,N_23893);
nand U24136 (N_24136,N_23982,N_23933);
nor U24137 (N_24137,N_23879,N_23802);
or U24138 (N_24138,N_23936,N_23961);
or U24139 (N_24139,N_23965,N_23951);
nand U24140 (N_24140,N_23999,N_23987);
or U24141 (N_24141,N_23825,N_23956);
nor U24142 (N_24142,N_23902,N_23873);
nand U24143 (N_24143,N_23931,N_23900);
xor U24144 (N_24144,N_23933,N_23879);
nor U24145 (N_24145,N_23818,N_23850);
nand U24146 (N_24146,N_23972,N_23905);
nand U24147 (N_24147,N_23846,N_23883);
and U24148 (N_24148,N_23841,N_23945);
nand U24149 (N_24149,N_23914,N_23953);
nor U24150 (N_24150,N_23847,N_23950);
nand U24151 (N_24151,N_23911,N_23894);
nor U24152 (N_24152,N_23907,N_23838);
or U24153 (N_24153,N_23967,N_23977);
nor U24154 (N_24154,N_23878,N_23959);
or U24155 (N_24155,N_23893,N_23880);
or U24156 (N_24156,N_23820,N_23870);
or U24157 (N_24157,N_23837,N_23937);
or U24158 (N_24158,N_23999,N_23924);
xnor U24159 (N_24159,N_23876,N_23862);
nor U24160 (N_24160,N_23935,N_23915);
nor U24161 (N_24161,N_23861,N_23827);
and U24162 (N_24162,N_23801,N_23892);
nor U24163 (N_24163,N_23861,N_23826);
nor U24164 (N_24164,N_23976,N_23992);
xor U24165 (N_24165,N_23987,N_23911);
and U24166 (N_24166,N_23991,N_23983);
xor U24167 (N_24167,N_23966,N_23909);
and U24168 (N_24168,N_23820,N_23894);
nand U24169 (N_24169,N_23899,N_23823);
or U24170 (N_24170,N_23864,N_23935);
or U24171 (N_24171,N_23997,N_23807);
or U24172 (N_24172,N_23871,N_23941);
and U24173 (N_24173,N_23857,N_23970);
xnor U24174 (N_24174,N_23849,N_23996);
or U24175 (N_24175,N_23940,N_23854);
nand U24176 (N_24176,N_23865,N_23826);
xnor U24177 (N_24177,N_23807,N_23825);
nand U24178 (N_24178,N_23861,N_23974);
xor U24179 (N_24179,N_23911,N_23895);
xnor U24180 (N_24180,N_23827,N_23862);
nor U24181 (N_24181,N_23939,N_23850);
nor U24182 (N_24182,N_23992,N_23843);
xnor U24183 (N_24183,N_23990,N_23873);
xor U24184 (N_24184,N_23802,N_23904);
nand U24185 (N_24185,N_23879,N_23881);
nor U24186 (N_24186,N_23883,N_23851);
xnor U24187 (N_24187,N_23889,N_23871);
nand U24188 (N_24188,N_23825,N_23919);
or U24189 (N_24189,N_23881,N_23988);
and U24190 (N_24190,N_23843,N_23977);
or U24191 (N_24191,N_23816,N_23873);
and U24192 (N_24192,N_23876,N_23955);
nand U24193 (N_24193,N_23959,N_23897);
and U24194 (N_24194,N_23841,N_23934);
nor U24195 (N_24195,N_23832,N_23973);
nand U24196 (N_24196,N_23921,N_23904);
or U24197 (N_24197,N_23887,N_23869);
nor U24198 (N_24198,N_23874,N_23865);
xor U24199 (N_24199,N_23933,N_23907);
nor U24200 (N_24200,N_24002,N_24136);
nor U24201 (N_24201,N_24022,N_24067);
nor U24202 (N_24202,N_24196,N_24047);
xor U24203 (N_24203,N_24194,N_24033);
xnor U24204 (N_24204,N_24100,N_24173);
xor U24205 (N_24205,N_24098,N_24017);
or U24206 (N_24206,N_24094,N_24040);
xor U24207 (N_24207,N_24110,N_24075);
xnor U24208 (N_24208,N_24108,N_24093);
nand U24209 (N_24209,N_24160,N_24074);
nand U24210 (N_24210,N_24113,N_24114);
xor U24211 (N_24211,N_24176,N_24054);
xor U24212 (N_24212,N_24050,N_24046);
and U24213 (N_24213,N_24123,N_24133);
nand U24214 (N_24214,N_24130,N_24115);
nor U24215 (N_24215,N_24101,N_24069);
nor U24216 (N_24216,N_24072,N_24184);
nor U24217 (N_24217,N_24161,N_24041);
nand U24218 (N_24218,N_24165,N_24052);
nand U24219 (N_24219,N_24006,N_24019);
or U24220 (N_24220,N_24013,N_24009);
xor U24221 (N_24221,N_24137,N_24150);
xnor U24222 (N_24222,N_24086,N_24018);
or U24223 (N_24223,N_24030,N_24151);
xor U24224 (N_24224,N_24039,N_24023);
nor U24225 (N_24225,N_24015,N_24126);
or U24226 (N_24226,N_24190,N_24037);
nor U24227 (N_24227,N_24059,N_24003);
nand U24228 (N_24228,N_24170,N_24167);
nand U24229 (N_24229,N_24099,N_24025);
xor U24230 (N_24230,N_24119,N_24053);
or U24231 (N_24231,N_24182,N_24042);
and U24232 (N_24232,N_24065,N_24080);
nor U24233 (N_24233,N_24112,N_24038);
or U24234 (N_24234,N_24177,N_24128);
nor U24235 (N_24235,N_24032,N_24021);
nand U24236 (N_24236,N_24149,N_24140);
nand U24237 (N_24237,N_24172,N_24031);
xor U24238 (N_24238,N_24084,N_24166);
and U24239 (N_24239,N_24058,N_24076);
or U24240 (N_24240,N_24091,N_24153);
nor U24241 (N_24241,N_24005,N_24174);
xor U24242 (N_24242,N_24066,N_24055);
nand U24243 (N_24243,N_24001,N_24044);
nand U24244 (N_24244,N_24043,N_24147);
nor U24245 (N_24245,N_24051,N_24168);
and U24246 (N_24246,N_24008,N_24068);
nand U24247 (N_24247,N_24121,N_24131);
or U24248 (N_24248,N_24198,N_24155);
or U24249 (N_24249,N_24132,N_24048);
and U24250 (N_24250,N_24000,N_24088);
xnor U24251 (N_24251,N_24197,N_24107);
and U24252 (N_24252,N_24135,N_24082);
nand U24253 (N_24253,N_24078,N_24189);
nor U24254 (N_24254,N_24192,N_24016);
and U24255 (N_24255,N_24122,N_24011);
nor U24256 (N_24256,N_24024,N_24036);
xor U24257 (N_24257,N_24143,N_24028);
or U24258 (N_24258,N_24109,N_24186);
nand U24259 (N_24259,N_24180,N_24061);
xnor U24260 (N_24260,N_24012,N_24146);
nor U24261 (N_24261,N_24105,N_24163);
or U24262 (N_24262,N_24027,N_24034);
xnor U24263 (N_24263,N_24079,N_24045);
or U24264 (N_24264,N_24129,N_24120);
and U24265 (N_24265,N_24157,N_24060);
nand U24266 (N_24266,N_24096,N_24199);
or U24267 (N_24267,N_24125,N_24158);
xnor U24268 (N_24268,N_24116,N_24090);
nor U24269 (N_24269,N_24144,N_24152);
xnor U24270 (N_24270,N_24178,N_24010);
xor U24271 (N_24271,N_24071,N_24141);
xor U24272 (N_24272,N_24077,N_24083);
nand U24273 (N_24273,N_24191,N_24164);
xnor U24274 (N_24274,N_24117,N_24162);
xnor U24275 (N_24275,N_24111,N_24118);
nor U24276 (N_24276,N_24188,N_24193);
and U24277 (N_24277,N_24092,N_24064);
and U24278 (N_24278,N_24156,N_24035);
and U24279 (N_24279,N_24049,N_24148);
xor U24280 (N_24280,N_24187,N_24159);
or U24281 (N_24281,N_24154,N_24139);
nor U24282 (N_24282,N_24062,N_24195);
nand U24283 (N_24283,N_24085,N_24095);
nand U24284 (N_24284,N_24087,N_24007);
or U24285 (N_24285,N_24104,N_24183);
xor U24286 (N_24286,N_24185,N_24004);
and U24287 (N_24287,N_24089,N_24020);
and U24288 (N_24288,N_24057,N_24056);
or U24289 (N_24289,N_24179,N_24134);
nand U24290 (N_24290,N_24026,N_24169);
and U24291 (N_24291,N_24124,N_24106);
and U24292 (N_24292,N_24073,N_24142);
nand U24293 (N_24293,N_24181,N_24014);
xor U24294 (N_24294,N_24127,N_24102);
nand U24295 (N_24295,N_24103,N_24081);
nand U24296 (N_24296,N_24029,N_24138);
and U24297 (N_24297,N_24063,N_24145);
xor U24298 (N_24298,N_24175,N_24070);
or U24299 (N_24299,N_24097,N_24171);
nor U24300 (N_24300,N_24140,N_24192);
nand U24301 (N_24301,N_24135,N_24101);
or U24302 (N_24302,N_24163,N_24173);
xor U24303 (N_24303,N_24161,N_24037);
or U24304 (N_24304,N_24074,N_24100);
xor U24305 (N_24305,N_24166,N_24183);
or U24306 (N_24306,N_24069,N_24168);
nor U24307 (N_24307,N_24189,N_24071);
nor U24308 (N_24308,N_24170,N_24065);
and U24309 (N_24309,N_24188,N_24106);
and U24310 (N_24310,N_24070,N_24101);
nor U24311 (N_24311,N_24118,N_24057);
xnor U24312 (N_24312,N_24095,N_24056);
nand U24313 (N_24313,N_24029,N_24160);
or U24314 (N_24314,N_24141,N_24152);
nor U24315 (N_24315,N_24049,N_24004);
nor U24316 (N_24316,N_24151,N_24128);
xnor U24317 (N_24317,N_24196,N_24154);
and U24318 (N_24318,N_24133,N_24062);
nor U24319 (N_24319,N_24181,N_24170);
xnor U24320 (N_24320,N_24024,N_24125);
xnor U24321 (N_24321,N_24159,N_24080);
and U24322 (N_24322,N_24136,N_24093);
or U24323 (N_24323,N_24147,N_24100);
and U24324 (N_24324,N_24167,N_24161);
or U24325 (N_24325,N_24046,N_24011);
xor U24326 (N_24326,N_24066,N_24112);
nand U24327 (N_24327,N_24193,N_24096);
and U24328 (N_24328,N_24142,N_24159);
nand U24329 (N_24329,N_24177,N_24007);
and U24330 (N_24330,N_24153,N_24130);
and U24331 (N_24331,N_24198,N_24115);
nor U24332 (N_24332,N_24137,N_24039);
xor U24333 (N_24333,N_24129,N_24109);
xor U24334 (N_24334,N_24121,N_24047);
nand U24335 (N_24335,N_24047,N_24146);
and U24336 (N_24336,N_24023,N_24034);
and U24337 (N_24337,N_24095,N_24130);
nor U24338 (N_24338,N_24042,N_24100);
nor U24339 (N_24339,N_24071,N_24183);
xnor U24340 (N_24340,N_24140,N_24045);
nand U24341 (N_24341,N_24139,N_24097);
nand U24342 (N_24342,N_24070,N_24050);
nand U24343 (N_24343,N_24041,N_24032);
or U24344 (N_24344,N_24165,N_24136);
nand U24345 (N_24345,N_24035,N_24053);
and U24346 (N_24346,N_24052,N_24011);
and U24347 (N_24347,N_24187,N_24175);
and U24348 (N_24348,N_24135,N_24054);
nor U24349 (N_24349,N_24041,N_24007);
nor U24350 (N_24350,N_24191,N_24153);
xor U24351 (N_24351,N_24168,N_24106);
xor U24352 (N_24352,N_24067,N_24152);
or U24353 (N_24353,N_24161,N_24040);
or U24354 (N_24354,N_24115,N_24171);
nor U24355 (N_24355,N_24159,N_24034);
nand U24356 (N_24356,N_24109,N_24138);
xor U24357 (N_24357,N_24082,N_24110);
and U24358 (N_24358,N_24171,N_24100);
or U24359 (N_24359,N_24046,N_24103);
and U24360 (N_24360,N_24099,N_24191);
or U24361 (N_24361,N_24101,N_24177);
nand U24362 (N_24362,N_24097,N_24136);
nand U24363 (N_24363,N_24191,N_24166);
or U24364 (N_24364,N_24002,N_24164);
and U24365 (N_24365,N_24092,N_24137);
nor U24366 (N_24366,N_24158,N_24023);
nor U24367 (N_24367,N_24161,N_24092);
nand U24368 (N_24368,N_24192,N_24085);
nor U24369 (N_24369,N_24172,N_24132);
xor U24370 (N_24370,N_24073,N_24199);
or U24371 (N_24371,N_24038,N_24075);
and U24372 (N_24372,N_24165,N_24135);
nand U24373 (N_24373,N_24098,N_24162);
nand U24374 (N_24374,N_24033,N_24030);
xnor U24375 (N_24375,N_24143,N_24179);
nand U24376 (N_24376,N_24172,N_24106);
and U24377 (N_24377,N_24049,N_24187);
nor U24378 (N_24378,N_24055,N_24037);
xnor U24379 (N_24379,N_24198,N_24062);
xor U24380 (N_24380,N_24188,N_24113);
nand U24381 (N_24381,N_24027,N_24112);
and U24382 (N_24382,N_24133,N_24081);
nor U24383 (N_24383,N_24080,N_24096);
or U24384 (N_24384,N_24008,N_24132);
and U24385 (N_24385,N_24168,N_24152);
or U24386 (N_24386,N_24193,N_24008);
xnor U24387 (N_24387,N_24027,N_24086);
nor U24388 (N_24388,N_24015,N_24117);
xor U24389 (N_24389,N_24140,N_24087);
and U24390 (N_24390,N_24128,N_24013);
nand U24391 (N_24391,N_24186,N_24194);
xor U24392 (N_24392,N_24025,N_24039);
xnor U24393 (N_24393,N_24091,N_24175);
xnor U24394 (N_24394,N_24166,N_24160);
nand U24395 (N_24395,N_24129,N_24054);
or U24396 (N_24396,N_24111,N_24034);
xor U24397 (N_24397,N_24061,N_24136);
and U24398 (N_24398,N_24109,N_24009);
nor U24399 (N_24399,N_24012,N_24088);
nand U24400 (N_24400,N_24281,N_24268);
or U24401 (N_24401,N_24362,N_24360);
and U24402 (N_24402,N_24265,N_24358);
and U24403 (N_24403,N_24361,N_24305);
and U24404 (N_24404,N_24391,N_24393);
and U24405 (N_24405,N_24229,N_24380);
nor U24406 (N_24406,N_24234,N_24346);
nand U24407 (N_24407,N_24215,N_24261);
nor U24408 (N_24408,N_24321,N_24343);
nor U24409 (N_24409,N_24236,N_24264);
nor U24410 (N_24410,N_24375,N_24308);
nand U24411 (N_24411,N_24299,N_24239);
or U24412 (N_24412,N_24385,N_24224);
nor U24413 (N_24413,N_24318,N_24206);
or U24414 (N_24414,N_24316,N_24230);
nand U24415 (N_24415,N_24392,N_24396);
nor U24416 (N_24416,N_24359,N_24306);
nor U24417 (N_24417,N_24214,N_24296);
or U24418 (N_24418,N_24325,N_24398);
and U24419 (N_24419,N_24347,N_24275);
nand U24420 (N_24420,N_24246,N_24207);
nor U24421 (N_24421,N_24201,N_24363);
nand U24422 (N_24422,N_24231,N_24217);
or U24423 (N_24423,N_24338,N_24319);
nor U24424 (N_24424,N_24288,N_24263);
and U24425 (N_24425,N_24381,N_24209);
nor U24426 (N_24426,N_24337,N_24252);
nor U24427 (N_24427,N_24241,N_24303);
nor U24428 (N_24428,N_24287,N_24249);
nor U24429 (N_24429,N_24386,N_24314);
xor U24430 (N_24430,N_24254,N_24378);
or U24431 (N_24431,N_24295,N_24341);
nor U24432 (N_24432,N_24245,N_24262);
nor U24433 (N_24433,N_24352,N_24388);
nor U24434 (N_24434,N_24307,N_24369);
nand U24435 (N_24435,N_24284,N_24350);
and U24436 (N_24436,N_24335,N_24267);
or U24437 (N_24437,N_24286,N_24329);
xnor U24438 (N_24438,N_24331,N_24202);
or U24439 (N_24439,N_24302,N_24317);
xor U24440 (N_24440,N_24205,N_24294);
xor U24441 (N_24441,N_24340,N_24367);
or U24442 (N_24442,N_24292,N_24270);
nand U24443 (N_24443,N_24237,N_24353);
xor U24444 (N_24444,N_24310,N_24372);
and U24445 (N_24445,N_24390,N_24300);
and U24446 (N_24446,N_24282,N_24330);
xor U24447 (N_24447,N_24216,N_24371);
or U24448 (N_24448,N_24218,N_24223);
nand U24449 (N_24449,N_24210,N_24212);
nor U24450 (N_24450,N_24211,N_24255);
or U24451 (N_24451,N_24271,N_24344);
or U24452 (N_24452,N_24221,N_24200);
nand U24453 (N_24453,N_24397,N_24357);
xnor U24454 (N_24454,N_24309,N_24289);
nand U24455 (N_24455,N_24290,N_24235);
xnor U24456 (N_24456,N_24356,N_24238);
or U24457 (N_24457,N_24315,N_24279);
xnor U24458 (N_24458,N_24313,N_24311);
and U24459 (N_24459,N_24364,N_24277);
nand U24460 (N_24460,N_24273,N_24333);
or U24461 (N_24461,N_24274,N_24213);
or U24462 (N_24462,N_24203,N_24240);
or U24463 (N_24463,N_24243,N_24228);
or U24464 (N_24464,N_24365,N_24373);
nor U24465 (N_24465,N_24354,N_24258);
or U24466 (N_24466,N_24253,N_24328);
xor U24467 (N_24467,N_24257,N_24382);
nand U24468 (N_24468,N_24349,N_24272);
xor U24469 (N_24469,N_24220,N_24280);
and U24470 (N_24470,N_24323,N_24204);
or U24471 (N_24471,N_24232,N_24374);
or U24472 (N_24472,N_24334,N_24285);
nor U24473 (N_24473,N_24379,N_24291);
or U24474 (N_24474,N_24348,N_24389);
and U24475 (N_24475,N_24377,N_24222);
nand U24476 (N_24476,N_24304,N_24225);
nand U24477 (N_24477,N_24250,N_24326);
nand U24478 (N_24478,N_24293,N_24312);
or U24479 (N_24479,N_24278,N_24242);
nand U24480 (N_24480,N_24283,N_24324);
xor U24481 (N_24481,N_24248,N_24336);
or U24482 (N_24482,N_24208,N_24301);
nor U24483 (N_24483,N_24355,N_24342);
nor U24484 (N_24484,N_24251,N_24320);
nor U24485 (N_24485,N_24339,N_24247);
xnor U24486 (N_24486,N_24276,N_24259);
or U24487 (N_24487,N_24256,N_24266);
xor U24488 (N_24488,N_24219,N_24370);
or U24489 (N_24489,N_24332,N_24384);
and U24490 (N_24490,N_24298,N_24394);
and U24491 (N_24491,N_24244,N_24226);
and U24492 (N_24492,N_24399,N_24345);
or U24493 (N_24493,N_24376,N_24322);
nand U24494 (N_24494,N_24383,N_24260);
or U24495 (N_24495,N_24327,N_24297);
xnor U24496 (N_24496,N_24395,N_24269);
nand U24497 (N_24497,N_24227,N_24366);
nand U24498 (N_24498,N_24351,N_24387);
nand U24499 (N_24499,N_24233,N_24368);
or U24500 (N_24500,N_24387,N_24383);
xor U24501 (N_24501,N_24206,N_24282);
nand U24502 (N_24502,N_24333,N_24396);
nand U24503 (N_24503,N_24288,N_24234);
nor U24504 (N_24504,N_24329,N_24251);
xor U24505 (N_24505,N_24330,N_24254);
nor U24506 (N_24506,N_24308,N_24259);
and U24507 (N_24507,N_24290,N_24278);
and U24508 (N_24508,N_24240,N_24358);
or U24509 (N_24509,N_24395,N_24246);
and U24510 (N_24510,N_24271,N_24357);
nor U24511 (N_24511,N_24299,N_24295);
or U24512 (N_24512,N_24218,N_24285);
or U24513 (N_24513,N_24250,N_24388);
nand U24514 (N_24514,N_24350,N_24223);
or U24515 (N_24515,N_24291,N_24355);
nand U24516 (N_24516,N_24290,N_24244);
nor U24517 (N_24517,N_24389,N_24279);
nor U24518 (N_24518,N_24210,N_24233);
nor U24519 (N_24519,N_24207,N_24327);
nand U24520 (N_24520,N_24235,N_24203);
and U24521 (N_24521,N_24286,N_24300);
xor U24522 (N_24522,N_24230,N_24337);
nand U24523 (N_24523,N_24315,N_24251);
nor U24524 (N_24524,N_24233,N_24375);
xor U24525 (N_24525,N_24339,N_24224);
or U24526 (N_24526,N_24341,N_24274);
nand U24527 (N_24527,N_24344,N_24277);
xnor U24528 (N_24528,N_24268,N_24317);
or U24529 (N_24529,N_24298,N_24340);
or U24530 (N_24530,N_24376,N_24272);
nor U24531 (N_24531,N_24237,N_24247);
xnor U24532 (N_24532,N_24361,N_24240);
nand U24533 (N_24533,N_24381,N_24205);
xor U24534 (N_24534,N_24288,N_24255);
or U24535 (N_24535,N_24321,N_24329);
xor U24536 (N_24536,N_24305,N_24375);
xor U24537 (N_24537,N_24327,N_24326);
or U24538 (N_24538,N_24369,N_24360);
nand U24539 (N_24539,N_24392,N_24324);
nor U24540 (N_24540,N_24382,N_24216);
nor U24541 (N_24541,N_24360,N_24202);
nor U24542 (N_24542,N_24227,N_24268);
or U24543 (N_24543,N_24399,N_24216);
xnor U24544 (N_24544,N_24349,N_24275);
xor U24545 (N_24545,N_24358,N_24372);
and U24546 (N_24546,N_24227,N_24393);
nand U24547 (N_24547,N_24307,N_24337);
xnor U24548 (N_24548,N_24270,N_24384);
and U24549 (N_24549,N_24381,N_24320);
nor U24550 (N_24550,N_24329,N_24250);
xor U24551 (N_24551,N_24289,N_24359);
or U24552 (N_24552,N_24284,N_24278);
and U24553 (N_24553,N_24362,N_24283);
nand U24554 (N_24554,N_24315,N_24235);
xor U24555 (N_24555,N_24327,N_24330);
or U24556 (N_24556,N_24335,N_24239);
xor U24557 (N_24557,N_24231,N_24355);
nor U24558 (N_24558,N_24381,N_24256);
xor U24559 (N_24559,N_24283,N_24248);
nand U24560 (N_24560,N_24349,N_24387);
nor U24561 (N_24561,N_24307,N_24241);
nand U24562 (N_24562,N_24314,N_24268);
xor U24563 (N_24563,N_24339,N_24284);
nand U24564 (N_24564,N_24225,N_24218);
and U24565 (N_24565,N_24208,N_24312);
or U24566 (N_24566,N_24383,N_24340);
xnor U24567 (N_24567,N_24241,N_24296);
xor U24568 (N_24568,N_24327,N_24335);
and U24569 (N_24569,N_24247,N_24337);
or U24570 (N_24570,N_24398,N_24244);
nand U24571 (N_24571,N_24286,N_24399);
nor U24572 (N_24572,N_24223,N_24361);
or U24573 (N_24573,N_24365,N_24315);
xor U24574 (N_24574,N_24263,N_24344);
nor U24575 (N_24575,N_24373,N_24239);
or U24576 (N_24576,N_24300,N_24263);
and U24577 (N_24577,N_24276,N_24354);
xor U24578 (N_24578,N_24335,N_24266);
xor U24579 (N_24579,N_24225,N_24316);
nor U24580 (N_24580,N_24214,N_24336);
or U24581 (N_24581,N_24390,N_24268);
xnor U24582 (N_24582,N_24246,N_24334);
nor U24583 (N_24583,N_24343,N_24277);
nand U24584 (N_24584,N_24307,N_24305);
and U24585 (N_24585,N_24362,N_24258);
nand U24586 (N_24586,N_24278,N_24283);
or U24587 (N_24587,N_24229,N_24328);
xnor U24588 (N_24588,N_24323,N_24392);
xor U24589 (N_24589,N_24266,N_24347);
xor U24590 (N_24590,N_24399,N_24217);
nand U24591 (N_24591,N_24303,N_24296);
nor U24592 (N_24592,N_24220,N_24245);
or U24593 (N_24593,N_24312,N_24321);
xor U24594 (N_24594,N_24297,N_24231);
nand U24595 (N_24595,N_24305,N_24313);
and U24596 (N_24596,N_24251,N_24396);
xnor U24597 (N_24597,N_24282,N_24312);
xor U24598 (N_24598,N_24334,N_24267);
xnor U24599 (N_24599,N_24209,N_24301);
nor U24600 (N_24600,N_24568,N_24435);
and U24601 (N_24601,N_24416,N_24409);
xor U24602 (N_24602,N_24547,N_24470);
nor U24603 (N_24603,N_24574,N_24509);
nand U24604 (N_24604,N_24408,N_24584);
nand U24605 (N_24605,N_24418,N_24407);
nand U24606 (N_24606,N_24592,N_24591);
xnor U24607 (N_24607,N_24532,N_24539);
or U24608 (N_24608,N_24537,N_24400);
xnor U24609 (N_24609,N_24410,N_24544);
and U24610 (N_24610,N_24546,N_24579);
and U24611 (N_24611,N_24458,N_24556);
nor U24612 (N_24612,N_24441,N_24548);
and U24613 (N_24613,N_24456,N_24545);
and U24614 (N_24614,N_24426,N_24535);
nand U24615 (N_24615,N_24413,N_24451);
and U24616 (N_24616,N_24436,N_24577);
nor U24617 (N_24617,N_24566,N_24484);
nor U24618 (N_24618,N_24581,N_24536);
nor U24619 (N_24619,N_24473,N_24583);
nor U24620 (N_24620,N_24538,N_24589);
xnor U24621 (N_24621,N_24524,N_24553);
nand U24622 (N_24622,N_24463,N_24464);
nor U24623 (N_24623,N_24531,N_24431);
nor U24624 (N_24624,N_24455,N_24467);
nand U24625 (N_24625,N_24576,N_24514);
or U24626 (N_24626,N_24453,N_24498);
nor U24627 (N_24627,N_24412,N_24502);
nand U24628 (N_24628,N_24447,N_24450);
nor U24629 (N_24629,N_24554,N_24454);
or U24630 (N_24630,N_24586,N_24555);
xnor U24631 (N_24631,N_24444,N_24421);
xor U24632 (N_24632,N_24445,N_24430);
nand U24633 (N_24633,N_24428,N_24575);
or U24634 (N_24634,N_24597,N_24533);
and U24635 (N_24635,N_24507,N_24442);
nand U24636 (N_24636,N_24596,N_24432);
or U24637 (N_24637,N_24540,N_24563);
or U24638 (N_24638,N_24526,N_24406);
xor U24639 (N_24639,N_24474,N_24560);
or U24640 (N_24640,N_24508,N_24465);
nand U24641 (N_24641,N_24452,N_24551);
nand U24642 (N_24642,N_24501,N_24529);
nand U24643 (N_24643,N_24469,N_24414);
and U24644 (N_24644,N_24521,N_24593);
xor U24645 (N_24645,N_24468,N_24565);
nand U24646 (N_24646,N_24588,N_24437);
or U24647 (N_24647,N_24482,N_24419);
xor U24648 (N_24648,N_24401,N_24481);
nor U24649 (N_24649,N_24585,N_24578);
and U24650 (N_24650,N_24534,N_24519);
and U24651 (N_24651,N_24487,N_24486);
nor U24652 (N_24652,N_24490,N_24512);
or U24653 (N_24653,N_24552,N_24569);
and U24654 (N_24654,N_24557,N_24423);
or U24655 (N_24655,N_24564,N_24530);
nand U24656 (N_24656,N_24504,N_24567);
and U24657 (N_24657,N_24523,N_24457);
or U24658 (N_24658,N_24477,N_24594);
and U24659 (N_24659,N_24562,N_24446);
and U24660 (N_24660,N_24479,N_24528);
nor U24661 (N_24661,N_24402,N_24494);
and U24662 (N_24662,N_24550,N_24422);
nand U24663 (N_24663,N_24438,N_24543);
xor U24664 (N_24664,N_24449,N_24522);
nand U24665 (N_24665,N_24572,N_24542);
xor U24666 (N_24666,N_24466,N_24489);
nand U24667 (N_24667,N_24461,N_24580);
xor U24668 (N_24668,N_24516,N_24496);
or U24669 (N_24669,N_24493,N_24460);
xnor U24670 (N_24670,N_24520,N_24478);
or U24671 (N_24671,N_24443,N_24515);
nand U24672 (N_24672,N_24510,N_24518);
nor U24673 (N_24673,N_24499,N_24415);
or U24674 (N_24674,N_24527,N_24483);
or U24675 (N_24675,N_24492,N_24513);
nand U24676 (N_24676,N_24573,N_24439);
or U24677 (N_24677,N_24459,N_24429);
and U24678 (N_24678,N_24411,N_24505);
and U24679 (N_24679,N_24558,N_24485);
nand U24680 (N_24680,N_24525,N_24403);
nand U24681 (N_24681,N_24595,N_24517);
nor U24682 (N_24682,N_24404,N_24424);
nand U24683 (N_24683,N_24549,N_24476);
or U24684 (N_24684,N_24497,N_24480);
xnor U24685 (N_24685,N_24587,N_24434);
xnor U24686 (N_24686,N_24433,N_24590);
xor U24687 (N_24687,N_24503,N_24427);
or U24688 (N_24688,N_24471,N_24448);
and U24689 (N_24689,N_24559,N_24500);
nand U24690 (N_24690,N_24598,N_24440);
nor U24691 (N_24691,N_24472,N_24570);
and U24692 (N_24692,N_24462,N_24541);
and U24693 (N_24693,N_24506,N_24420);
xnor U24694 (N_24694,N_24582,N_24417);
nand U24695 (N_24695,N_24571,N_24405);
xor U24696 (N_24696,N_24475,N_24561);
nor U24697 (N_24697,N_24425,N_24599);
nor U24698 (N_24698,N_24491,N_24495);
and U24699 (N_24699,N_24488,N_24511);
or U24700 (N_24700,N_24596,N_24498);
nand U24701 (N_24701,N_24498,N_24457);
and U24702 (N_24702,N_24568,N_24430);
nor U24703 (N_24703,N_24414,N_24482);
xnor U24704 (N_24704,N_24461,N_24545);
and U24705 (N_24705,N_24455,N_24418);
or U24706 (N_24706,N_24476,N_24532);
or U24707 (N_24707,N_24588,N_24491);
nor U24708 (N_24708,N_24468,N_24432);
and U24709 (N_24709,N_24512,N_24433);
xnor U24710 (N_24710,N_24556,N_24435);
nand U24711 (N_24711,N_24471,N_24422);
and U24712 (N_24712,N_24590,N_24580);
nand U24713 (N_24713,N_24583,N_24529);
and U24714 (N_24714,N_24420,N_24558);
xnor U24715 (N_24715,N_24478,N_24419);
nand U24716 (N_24716,N_24407,N_24442);
nand U24717 (N_24717,N_24509,N_24592);
or U24718 (N_24718,N_24545,N_24453);
nand U24719 (N_24719,N_24567,N_24493);
nand U24720 (N_24720,N_24478,N_24451);
and U24721 (N_24721,N_24474,N_24551);
xnor U24722 (N_24722,N_24593,N_24478);
and U24723 (N_24723,N_24497,N_24511);
and U24724 (N_24724,N_24568,N_24439);
and U24725 (N_24725,N_24460,N_24406);
and U24726 (N_24726,N_24568,N_24552);
and U24727 (N_24727,N_24542,N_24497);
or U24728 (N_24728,N_24469,N_24404);
xor U24729 (N_24729,N_24440,N_24446);
or U24730 (N_24730,N_24459,N_24567);
xnor U24731 (N_24731,N_24443,N_24428);
and U24732 (N_24732,N_24583,N_24410);
nand U24733 (N_24733,N_24452,N_24450);
and U24734 (N_24734,N_24558,N_24537);
xnor U24735 (N_24735,N_24488,N_24549);
or U24736 (N_24736,N_24455,N_24473);
nor U24737 (N_24737,N_24532,N_24596);
nand U24738 (N_24738,N_24486,N_24457);
and U24739 (N_24739,N_24542,N_24460);
or U24740 (N_24740,N_24509,N_24500);
nand U24741 (N_24741,N_24412,N_24448);
xnor U24742 (N_24742,N_24488,N_24407);
or U24743 (N_24743,N_24454,N_24563);
and U24744 (N_24744,N_24506,N_24552);
or U24745 (N_24745,N_24420,N_24571);
nor U24746 (N_24746,N_24448,N_24580);
and U24747 (N_24747,N_24511,N_24538);
or U24748 (N_24748,N_24426,N_24451);
or U24749 (N_24749,N_24423,N_24494);
xor U24750 (N_24750,N_24483,N_24512);
or U24751 (N_24751,N_24438,N_24556);
nand U24752 (N_24752,N_24567,N_24584);
nor U24753 (N_24753,N_24576,N_24431);
or U24754 (N_24754,N_24432,N_24528);
or U24755 (N_24755,N_24452,N_24502);
xnor U24756 (N_24756,N_24501,N_24559);
and U24757 (N_24757,N_24427,N_24439);
nor U24758 (N_24758,N_24409,N_24506);
and U24759 (N_24759,N_24437,N_24485);
and U24760 (N_24760,N_24506,N_24493);
xnor U24761 (N_24761,N_24494,N_24527);
xnor U24762 (N_24762,N_24465,N_24513);
nand U24763 (N_24763,N_24446,N_24415);
and U24764 (N_24764,N_24410,N_24423);
or U24765 (N_24765,N_24511,N_24461);
xnor U24766 (N_24766,N_24433,N_24491);
or U24767 (N_24767,N_24440,N_24536);
or U24768 (N_24768,N_24476,N_24436);
xor U24769 (N_24769,N_24550,N_24548);
or U24770 (N_24770,N_24482,N_24578);
and U24771 (N_24771,N_24470,N_24410);
xnor U24772 (N_24772,N_24557,N_24545);
or U24773 (N_24773,N_24520,N_24491);
or U24774 (N_24774,N_24544,N_24568);
xnor U24775 (N_24775,N_24579,N_24412);
or U24776 (N_24776,N_24571,N_24438);
xor U24777 (N_24777,N_24416,N_24448);
or U24778 (N_24778,N_24464,N_24588);
or U24779 (N_24779,N_24571,N_24598);
or U24780 (N_24780,N_24414,N_24523);
or U24781 (N_24781,N_24525,N_24541);
nand U24782 (N_24782,N_24597,N_24448);
nand U24783 (N_24783,N_24435,N_24548);
xnor U24784 (N_24784,N_24581,N_24580);
nand U24785 (N_24785,N_24464,N_24467);
or U24786 (N_24786,N_24564,N_24541);
nor U24787 (N_24787,N_24495,N_24420);
nor U24788 (N_24788,N_24595,N_24422);
nor U24789 (N_24789,N_24500,N_24489);
xnor U24790 (N_24790,N_24432,N_24531);
nor U24791 (N_24791,N_24428,N_24450);
or U24792 (N_24792,N_24586,N_24596);
and U24793 (N_24793,N_24404,N_24435);
and U24794 (N_24794,N_24540,N_24543);
nand U24795 (N_24795,N_24453,N_24590);
xnor U24796 (N_24796,N_24521,N_24468);
nand U24797 (N_24797,N_24532,N_24418);
or U24798 (N_24798,N_24547,N_24586);
xnor U24799 (N_24799,N_24527,N_24532);
and U24800 (N_24800,N_24644,N_24692);
xnor U24801 (N_24801,N_24756,N_24605);
nor U24802 (N_24802,N_24714,N_24722);
and U24803 (N_24803,N_24728,N_24705);
nand U24804 (N_24804,N_24740,N_24764);
xnor U24805 (N_24805,N_24752,N_24733);
xnor U24806 (N_24806,N_24769,N_24698);
or U24807 (N_24807,N_24782,N_24663);
nor U24808 (N_24808,N_24646,N_24638);
nand U24809 (N_24809,N_24632,N_24795);
nand U24810 (N_24810,N_24647,N_24741);
xnor U24811 (N_24811,N_24763,N_24745);
xor U24812 (N_24812,N_24772,N_24676);
xnor U24813 (N_24813,N_24630,N_24721);
xor U24814 (N_24814,N_24717,N_24601);
or U24815 (N_24815,N_24732,N_24729);
or U24816 (N_24816,N_24662,N_24648);
and U24817 (N_24817,N_24688,N_24703);
nor U24818 (N_24818,N_24642,N_24734);
nor U24819 (N_24819,N_24726,N_24725);
or U24820 (N_24820,N_24679,N_24742);
xnor U24821 (N_24821,N_24727,N_24607);
nor U24822 (N_24822,N_24671,N_24609);
or U24823 (N_24823,N_24748,N_24779);
and U24824 (N_24824,N_24751,N_24767);
xor U24825 (N_24825,N_24694,N_24738);
nand U24826 (N_24826,N_24656,N_24700);
xnor U24827 (N_24827,N_24696,N_24716);
nand U24828 (N_24828,N_24675,N_24623);
and U24829 (N_24829,N_24672,N_24634);
or U24830 (N_24830,N_24786,N_24602);
xor U24831 (N_24831,N_24793,N_24617);
nand U24832 (N_24832,N_24674,N_24689);
nand U24833 (N_24833,N_24753,N_24655);
or U24834 (N_24834,N_24669,N_24754);
nand U24835 (N_24835,N_24771,N_24693);
and U24836 (N_24836,N_24710,N_24720);
and U24837 (N_24837,N_24673,N_24766);
nor U24838 (N_24838,N_24666,N_24610);
or U24839 (N_24839,N_24639,N_24724);
and U24840 (N_24840,N_24780,N_24788);
and U24841 (N_24841,N_24690,N_24635);
nand U24842 (N_24842,N_24627,N_24667);
xor U24843 (N_24843,N_24701,N_24785);
nor U24844 (N_24844,N_24774,N_24650);
and U24845 (N_24845,N_24739,N_24744);
nand U24846 (N_24846,N_24678,N_24747);
xnor U24847 (N_24847,N_24783,N_24711);
nor U24848 (N_24848,N_24677,N_24730);
xnor U24849 (N_24849,N_24704,N_24787);
xnor U24850 (N_24850,N_24640,N_24612);
nor U24851 (N_24851,N_24737,N_24723);
and U24852 (N_24852,N_24684,N_24791);
or U24853 (N_24853,N_24658,N_24629);
nor U24854 (N_24854,N_24637,N_24759);
xnor U24855 (N_24855,N_24603,N_24636);
nor U24856 (N_24856,N_24781,N_24622);
and U24857 (N_24857,N_24633,N_24682);
nand U24858 (N_24858,N_24695,N_24628);
or U24859 (N_24859,N_24765,N_24613);
nand U24860 (N_24860,N_24743,N_24621);
or U24861 (N_24861,N_24625,N_24624);
or U24862 (N_24862,N_24615,N_24652);
and U24863 (N_24863,N_24794,N_24768);
or U24864 (N_24864,N_24608,N_24718);
nor U24865 (N_24865,N_24683,N_24619);
xnor U24866 (N_24866,N_24657,N_24626);
or U24867 (N_24867,N_24604,N_24736);
or U24868 (N_24868,N_24702,N_24762);
nand U24869 (N_24869,N_24776,N_24707);
and U24870 (N_24870,N_24775,N_24749);
nand U24871 (N_24871,N_24686,N_24755);
and U24872 (N_24872,N_24691,N_24661);
nand U24873 (N_24873,N_24699,N_24761);
and U24874 (N_24874,N_24643,N_24653);
and U24875 (N_24875,N_24697,N_24790);
nand U24876 (N_24876,N_24799,N_24777);
nor U24877 (N_24877,N_24758,N_24789);
xnor U24878 (N_24878,N_24735,N_24746);
or U24879 (N_24879,N_24778,N_24645);
or U24880 (N_24880,N_24600,N_24792);
nand U24881 (N_24881,N_24798,N_24680);
nand U24882 (N_24882,N_24709,N_24654);
or U24883 (N_24883,N_24606,N_24620);
and U24884 (N_24884,N_24668,N_24651);
nor U24885 (N_24885,N_24784,N_24713);
or U24886 (N_24886,N_24750,N_24681);
and U24887 (N_24887,N_24641,N_24708);
nor U24888 (N_24888,N_24670,N_24660);
and U24889 (N_24889,N_24614,N_24760);
and U24890 (N_24890,N_24611,N_24659);
nand U24891 (N_24891,N_24618,N_24719);
nor U24892 (N_24892,N_24649,N_24796);
nand U24893 (N_24893,N_24665,N_24712);
nand U24894 (N_24894,N_24731,N_24770);
or U24895 (N_24895,N_24773,N_24631);
or U24896 (N_24896,N_24664,N_24685);
or U24897 (N_24897,N_24687,N_24757);
nor U24898 (N_24898,N_24715,N_24797);
or U24899 (N_24899,N_24706,N_24616);
nor U24900 (N_24900,N_24725,N_24748);
xor U24901 (N_24901,N_24746,N_24627);
or U24902 (N_24902,N_24701,N_24732);
nor U24903 (N_24903,N_24669,N_24784);
nand U24904 (N_24904,N_24688,N_24758);
nor U24905 (N_24905,N_24763,N_24747);
and U24906 (N_24906,N_24778,N_24663);
nor U24907 (N_24907,N_24647,N_24760);
xor U24908 (N_24908,N_24754,N_24635);
nor U24909 (N_24909,N_24709,N_24688);
nor U24910 (N_24910,N_24774,N_24642);
nor U24911 (N_24911,N_24655,N_24632);
nor U24912 (N_24912,N_24717,N_24624);
nand U24913 (N_24913,N_24683,N_24718);
xnor U24914 (N_24914,N_24625,N_24636);
and U24915 (N_24915,N_24780,N_24688);
nand U24916 (N_24916,N_24618,N_24680);
xor U24917 (N_24917,N_24604,N_24655);
xor U24918 (N_24918,N_24790,N_24724);
or U24919 (N_24919,N_24793,N_24668);
xnor U24920 (N_24920,N_24625,N_24703);
or U24921 (N_24921,N_24625,N_24691);
nand U24922 (N_24922,N_24620,N_24676);
nor U24923 (N_24923,N_24713,N_24764);
nand U24924 (N_24924,N_24634,N_24643);
nand U24925 (N_24925,N_24763,N_24777);
and U24926 (N_24926,N_24771,N_24764);
xor U24927 (N_24927,N_24611,N_24646);
nor U24928 (N_24928,N_24653,N_24763);
or U24929 (N_24929,N_24706,N_24695);
and U24930 (N_24930,N_24675,N_24644);
nor U24931 (N_24931,N_24701,N_24781);
nand U24932 (N_24932,N_24779,N_24656);
xor U24933 (N_24933,N_24662,N_24790);
nor U24934 (N_24934,N_24794,N_24612);
and U24935 (N_24935,N_24620,N_24751);
or U24936 (N_24936,N_24789,N_24779);
xnor U24937 (N_24937,N_24656,N_24755);
or U24938 (N_24938,N_24780,N_24652);
xnor U24939 (N_24939,N_24699,N_24789);
nand U24940 (N_24940,N_24700,N_24777);
xnor U24941 (N_24941,N_24761,N_24785);
nor U24942 (N_24942,N_24762,N_24632);
nor U24943 (N_24943,N_24655,N_24614);
and U24944 (N_24944,N_24727,N_24611);
or U24945 (N_24945,N_24704,N_24643);
or U24946 (N_24946,N_24757,N_24688);
nor U24947 (N_24947,N_24630,N_24775);
nand U24948 (N_24948,N_24769,N_24755);
xor U24949 (N_24949,N_24604,N_24795);
and U24950 (N_24950,N_24715,N_24736);
nor U24951 (N_24951,N_24706,N_24699);
nand U24952 (N_24952,N_24774,N_24743);
xor U24953 (N_24953,N_24714,N_24790);
or U24954 (N_24954,N_24790,N_24780);
nor U24955 (N_24955,N_24712,N_24779);
and U24956 (N_24956,N_24637,N_24752);
nand U24957 (N_24957,N_24675,N_24744);
xnor U24958 (N_24958,N_24664,N_24647);
nor U24959 (N_24959,N_24768,N_24723);
nor U24960 (N_24960,N_24669,N_24642);
and U24961 (N_24961,N_24711,N_24737);
and U24962 (N_24962,N_24713,N_24641);
nor U24963 (N_24963,N_24767,N_24705);
nand U24964 (N_24964,N_24677,N_24627);
nor U24965 (N_24965,N_24682,N_24754);
nor U24966 (N_24966,N_24619,N_24768);
nand U24967 (N_24967,N_24705,N_24674);
nor U24968 (N_24968,N_24637,N_24765);
xnor U24969 (N_24969,N_24731,N_24787);
xor U24970 (N_24970,N_24796,N_24626);
and U24971 (N_24971,N_24730,N_24688);
nor U24972 (N_24972,N_24601,N_24764);
and U24973 (N_24973,N_24607,N_24665);
or U24974 (N_24974,N_24745,N_24631);
nand U24975 (N_24975,N_24707,N_24730);
xnor U24976 (N_24976,N_24787,N_24705);
xnor U24977 (N_24977,N_24789,N_24619);
xnor U24978 (N_24978,N_24653,N_24629);
nor U24979 (N_24979,N_24690,N_24606);
or U24980 (N_24980,N_24727,N_24650);
xor U24981 (N_24981,N_24715,N_24640);
nor U24982 (N_24982,N_24735,N_24751);
nand U24983 (N_24983,N_24769,N_24673);
nor U24984 (N_24984,N_24623,N_24710);
nand U24985 (N_24985,N_24695,N_24745);
or U24986 (N_24986,N_24671,N_24734);
or U24987 (N_24987,N_24750,N_24677);
xor U24988 (N_24988,N_24757,N_24736);
xor U24989 (N_24989,N_24745,N_24785);
xnor U24990 (N_24990,N_24686,N_24685);
and U24991 (N_24991,N_24774,N_24747);
or U24992 (N_24992,N_24705,N_24716);
nor U24993 (N_24993,N_24675,N_24692);
nand U24994 (N_24994,N_24694,N_24696);
or U24995 (N_24995,N_24612,N_24708);
nor U24996 (N_24996,N_24754,N_24740);
xnor U24997 (N_24997,N_24706,N_24713);
xor U24998 (N_24998,N_24719,N_24708);
or U24999 (N_24999,N_24639,N_24669);
or U25000 (N_25000,N_24973,N_24839);
xor U25001 (N_25001,N_24933,N_24834);
nand U25002 (N_25002,N_24959,N_24838);
xnor U25003 (N_25003,N_24999,N_24945);
and U25004 (N_25004,N_24910,N_24829);
and U25005 (N_25005,N_24966,N_24887);
nand U25006 (N_25006,N_24875,N_24872);
nand U25007 (N_25007,N_24918,N_24901);
or U25008 (N_25008,N_24821,N_24914);
nor U25009 (N_25009,N_24857,N_24814);
xnor U25010 (N_25010,N_24979,N_24915);
nor U25011 (N_25011,N_24936,N_24950);
and U25012 (N_25012,N_24801,N_24853);
or U25013 (N_25013,N_24997,N_24967);
and U25014 (N_25014,N_24826,N_24990);
xor U25015 (N_25015,N_24837,N_24934);
and U25016 (N_25016,N_24965,N_24948);
and U25017 (N_25017,N_24820,N_24920);
xnor U25018 (N_25018,N_24895,N_24974);
nor U25019 (N_25019,N_24893,N_24816);
and U25020 (N_25020,N_24832,N_24806);
nor U25021 (N_25021,N_24874,N_24971);
or U25022 (N_25022,N_24984,N_24902);
or U25023 (N_25023,N_24946,N_24908);
or U25024 (N_25024,N_24889,N_24835);
xnor U25025 (N_25025,N_24843,N_24937);
nand U25026 (N_25026,N_24878,N_24928);
and U25027 (N_25027,N_24852,N_24962);
or U25028 (N_25028,N_24953,N_24909);
nor U25029 (N_25029,N_24932,N_24939);
nor U25030 (N_25030,N_24951,N_24811);
and U25031 (N_25031,N_24830,N_24960);
xnor U25032 (N_25032,N_24970,N_24961);
nand U25033 (N_25033,N_24880,N_24803);
and U25034 (N_25034,N_24942,N_24916);
nor U25035 (N_25035,N_24868,N_24822);
xor U25036 (N_25036,N_24849,N_24804);
and U25037 (N_25037,N_24963,N_24956);
and U25038 (N_25038,N_24841,N_24993);
xor U25039 (N_25039,N_24957,N_24988);
nand U25040 (N_25040,N_24989,N_24846);
nand U25041 (N_25041,N_24969,N_24975);
xnor U25042 (N_25042,N_24824,N_24845);
and U25043 (N_25043,N_24877,N_24917);
nor U25044 (N_25044,N_24972,N_24850);
xor U25045 (N_25045,N_24919,N_24865);
xor U25046 (N_25046,N_24848,N_24888);
nor U25047 (N_25047,N_24983,N_24952);
nor U25048 (N_25048,N_24827,N_24949);
or U25049 (N_25049,N_24858,N_24860);
or U25050 (N_25050,N_24886,N_24922);
nor U25051 (N_25051,N_24815,N_24964);
nor U25052 (N_25052,N_24905,N_24879);
nand U25053 (N_25053,N_24925,N_24998);
xnor U25054 (N_25054,N_24991,N_24996);
and U25055 (N_25055,N_24900,N_24883);
xnor U25056 (N_25056,N_24992,N_24987);
nor U25057 (N_25057,N_24958,N_24851);
nand U25058 (N_25058,N_24930,N_24885);
nand U25059 (N_25059,N_24861,N_24844);
xor U25060 (N_25060,N_24947,N_24955);
and U25061 (N_25061,N_24819,N_24809);
or U25062 (N_25062,N_24840,N_24935);
xnor U25063 (N_25063,N_24944,N_24929);
nand U25064 (N_25064,N_24856,N_24892);
xor U25065 (N_25065,N_24876,N_24923);
and U25066 (N_25066,N_24982,N_24800);
xnor U25067 (N_25067,N_24904,N_24926);
or U25068 (N_25068,N_24940,N_24985);
nand U25069 (N_25069,N_24943,N_24825);
nand U25070 (N_25070,N_24976,N_24995);
or U25071 (N_25071,N_24882,N_24981);
and U25072 (N_25072,N_24911,N_24899);
or U25073 (N_25073,N_24836,N_24831);
and U25074 (N_25074,N_24906,N_24828);
and U25075 (N_25075,N_24833,N_24818);
nor U25076 (N_25076,N_24896,N_24808);
xnor U25077 (N_25077,N_24881,N_24907);
or U25078 (N_25078,N_24807,N_24912);
xnor U25079 (N_25079,N_24859,N_24898);
nor U25080 (N_25080,N_24894,N_24986);
nand U25081 (N_25081,N_24873,N_24871);
xor U25082 (N_25082,N_24862,N_24931);
and U25083 (N_25083,N_24810,N_24842);
nor U25084 (N_25084,N_24897,N_24847);
or U25085 (N_25085,N_24927,N_24805);
nor U25086 (N_25086,N_24890,N_24941);
nor U25087 (N_25087,N_24921,N_24891);
or U25088 (N_25088,N_24913,N_24813);
nor U25089 (N_25089,N_24802,N_24812);
or U25090 (N_25090,N_24968,N_24869);
xor U25091 (N_25091,N_24854,N_24903);
nand U25092 (N_25092,N_24870,N_24817);
xnor U25093 (N_25093,N_24978,N_24924);
and U25094 (N_25094,N_24938,N_24866);
or U25095 (N_25095,N_24994,N_24980);
xor U25096 (N_25096,N_24977,N_24867);
nand U25097 (N_25097,N_24863,N_24954);
xor U25098 (N_25098,N_24855,N_24864);
and U25099 (N_25099,N_24884,N_24823);
and U25100 (N_25100,N_24918,N_24963);
and U25101 (N_25101,N_24977,N_24849);
and U25102 (N_25102,N_24819,N_24852);
nor U25103 (N_25103,N_24948,N_24908);
and U25104 (N_25104,N_24987,N_24934);
nand U25105 (N_25105,N_24808,N_24883);
and U25106 (N_25106,N_24877,N_24846);
xor U25107 (N_25107,N_24804,N_24855);
nand U25108 (N_25108,N_24990,N_24978);
or U25109 (N_25109,N_24830,N_24992);
nand U25110 (N_25110,N_24855,N_24930);
nor U25111 (N_25111,N_24926,N_24955);
xnor U25112 (N_25112,N_24959,N_24979);
or U25113 (N_25113,N_24891,N_24951);
nor U25114 (N_25114,N_24920,N_24918);
and U25115 (N_25115,N_24816,N_24968);
or U25116 (N_25116,N_24944,N_24934);
or U25117 (N_25117,N_24810,N_24900);
xor U25118 (N_25118,N_24956,N_24826);
xor U25119 (N_25119,N_24816,N_24828);
nor U25120 (N_25120,N_24913,N_24807);
or U25121 (N_25121,N_24841,N_24869);
nand U25122 (N_25122,N_24928,N_24914);
and U25123 (N_25123,N_24878,N_24879);
and U25124 (N_25124,N_24874,N_24856);
xnor U25125 (N_25125,N_24890,N_24864);
nand U25126 (N_25126,N_24911,N_24810);
or U25127 (N_25127,N_24833,N_24888);
nor U25128 (N_25128,N_24926,N_24833);
xnor U25129 (N_25129,N_24930,N_24912);
and U25130 (N_25130,N_24969,N_24965);
xor U25131 (N_25131,N_24997,N_24818);
nand U25132 (N_25132,N_24901,N_24982);
nor U25133 (N_25133,N_24841,N_24910);
and U25134 (N_25134,N_24858,N_24856);
nor U25135 (N_25135,N_24914,N_24870);
nand U25136 (N_25136,N_24859,N_24802);
and U25137 (N_25137,N_24818,N_24913);
and U25138 (N_25138,N_24984,N_24817);
or U25139 (N_25139,N_24803,N_24929);
or U25140 (N_25140,N_24900,N_24947);
xor U25141 (N_25141,N_24985,N_24909);
and U25142 (N_25142,N_24916,N_24875);
xor U25143 (N_25143,N_24892,N_24977);
and U25144 (N_25144,N_24889,N_24971);
or U25145 (N_25145,N_24950,N_24934);
or U25146 (N_25146,N_24835,N_24960);
or U25147 (N_25147,N_24916,N_24931);
and U25148 (N_25148,N_24982,N_24959);
nor U25149 (N_25149,N_24905,N_24817);
and U25150 (N_25150,N_24959,N_24898);
xor U25151 (N_25151,N_24809,N_24964);
xor U25152 (N_25152,N_24802,N_24878);
and U25153 (N_25153,N_24888,N_24907);
xor U25154 (N_25154,N_24832,N_24974);
nand U25155 (N_25155,N_24851,N_24820);
and U25156 (N_25156,N_24856,N_24977);
nor U25157 (N_25157,N_24869,N_24817);
nand U25158 (N_25158,N_24801,N_24877);
and U25159 (N_25159,N_24944,N_24991);
xor U25160 (N_25160,N_24926,N_24843);
xor U25161 (N_25161,N_24981,N_24977);
nand U25162 (N_25162,N_24957,N_24925);
nor U25163 (N_25163,N_24891,N_24963);
or U25164 (N_25164,N_24881,N_24944);
or U25165 (N_25165,N_24936,N_24800);
or U25166 (N_25166,N_24952,N_24874);
xnor U25167 (N_25167,N_24846,N_24813);
xor U25168 (N_25168,N_24859,N_24838);
and U25169 (N_25169,N_24864,N_24857);
nand U25170 (N_25170,N_24977,N_24966);
and U25171 (N_25171,N_24802,N_24804);
nor U25172 (N_25172,N_24969,N_24924);
and U25173 (N_25173,N_24805,N_24981);
xnor U25174 (N_25174,N_24927,N_24937);
nor U25175 (N_25175,N_24950,N_24882);
and U25176 (N_25176,N_24921,N_24810);
or U25177 (N_25177,N_24950,N_24825);
or U25178 (N_25178,N_24926,N_24887);
nor U25179 (N_25179,N_24822,N_24812);
or U25180 (N_25180,N_24853,N_24985);
nor U25181 (N_25181,N_24879,N_24971);
nor U25182 (N_25182,N_24951,N_24802);
or U25183 (N_25183,N_24852,N_24844);
nand U25184 (N_25184,N_24985,N_24861);
nor U25185 (N_25185,N_24870,N_24935);
nor U25186 (N_25186,N_24815,N_24873);
nor U25187 (N_25187,N_24920,N_24928);
nand U25188 (N_25188,N_24865,N_24875);
or U25189 (N_25189,N_24878,N_24938);
xor U25190 (N_25190,N_24955,N_24887);
xor U25191 (N_25191,N_24839,N_24941);
nand U25192 (N_25192,N_24950,N_24818);
nor U25193 (N_25193,N_24820,N_24983);
and U25194 (N_25194,N_24806,N_24837);
and U25195 (N_25195,N_24892,N_24893);
nor U25196 (N_25196,N_24960,N_24965);
nor U25197 (N_25197,N_24887,N_24842);
nand U25198 (N_25198,N_24943,N_24858);
xnor U25199 (N_25199,N_24813,N_24984);
and U25200 (N_25200,N_25103,N_25172);
and U25201 (N_25201,N_25059,N_25142);
xnor U25202 (N_25202,N_25073,N_25149);
nor U25203 (N_25203,N_25091,N_25062);
nor U25204 (N_25204,N_25116,N_25079);
nor U25205 (N_25205,N_25027,N_25184);
nor U25206 (N_25206,N_25072,N_25085);
or U25207 (N_25207,N_25055,N_25045);
and U25208 (N_25208,N_25113,N_25191);
nand U25209 (N_25209,N_25030,N_25012);
nand U25210 (N_25210,N_25100,N_25003);
and U25211 (N_25211,N_25040,N_25178);
xor U25212 (N_25212,N_25174,N_25037);
and U25213 (N_25213,N_25197,N_25154);
and U25214 (N_25214,N_25041,N_25068);
and U25215 (N_25215,N_25161,N_25133);
nor U25216 (N_25216,N_25118,N_25104);
nor U25217 (N_25217,N_25028,N_25084);
or U25218 (N_25218,N_25060,N_25175);
nand U25219 (N_25219,N_25156,N_25016);
nor U25220 (N_25220,N_25014,N_25135);
nor U25221 (N_25221,N_25017,N_25098);
or U25222 (N_25222,N_25058,N_25026);
and U25223 (N_25223,N_25078,N_25173);
and U25224 (N_25224,N_25129,N_25034);
and U25225 (N_25225,N_25164,N_25095);
xor U25226 (N_25226,N_25155,N_25150);
and U25227 (N_25227,N_25198,N_25018);
and U25228 (N_25228,N_25131,N_25046);
or U25229 (N_25229,N_25199,N_25127);
nand U25230 (N_25230,N_25130,N_25106);
and U25231 (N_25231,N_25109,N_25057);
nand U25232 (N_25232,N_25020,N_25089);
nand U25233 (N_25233,N_25061,N_25176);
or U25234 (N_25234,N_25092,N_25010);
xor U25235 (N_25235,N_25013,N_25187);
and U25236 (N_25236,N_25140,N_25080);
xor U25237 (N_25237,N_25152,N_25067);
and U25238 (N_25238,N_25105,N_25157);
or U25239 (N_25239,N_25076,N_25169);
xnor U25240 (N_25240,N_25117,N_25033);
nor U25241 (N_25241,N_25075,N_25163);
or U25242 (N_25242,N_25185,N_25043);
nor U25243 (N_25243,N_25193,N_25086);
and U25244 (N_25244,N_25071,N_25053);
nand U25245 (N_25245,N_25036,N_25125);
nand U25246 (N_25246,N_25048,N_25151);
nand U25247 (N_25247,N_25143,N_25170);
nand U25248 (N_25248,N_25107,N_25194);
nor U25249 (N_25249,N_25179,N_25165);
nand U25250 (N_25250,N_25001,N_25132);
nor U25251 (N_25251,N_25141,N_25112);
nor U25252 (N_25252,N_25167,N_25035);
nor U25253 (N_25253,N_25019,N_25190);
or U25254 (N_25254,N_25038,N_25160);
nor U25255 (N_25255,N_25144,N_25094);
nand U25256 (N_25256,N_25052,N_25096);
or U25257 (N_25257,N_25015,N_25134);
nor U25258 (N_25258,N_25145,N_25128);
nand U25259 (N_25259,N_25002,N_25114);
or U25260 (N_25260,N_25093,N_25101);
and U25261 (N_25261,N_25147,N_25074);
and U25262 (N_25262,N_25121,N_25153);
xnor U25263 (N_25263,N_25021,N_25077);
or U25264 (N_25264,N_25166,N_25146);
and U25265 (N_25265,N_25087,N_25006);
nand U25266 (N_25266,N_25032,N_25183);
or U25267 (N_25267,N_25102,N_25024);
and U25268 (N_25268,N_25065,N_25063);
xor U25269 (N_25269,N_25124,N_25011);
nor U25270 (N_25270,N_25069,N_25186);
and U25271 (N_25271,N_25181,N_25050);
and U25272 (N_25272,N_25136,N_25042);
nor U25273 (N_25273,N_25138,N_25099);
nor U25274 (N_25274,N_25056,N_25188);
and U25275 (N_25275,N_25051,N_25159);
nand U25276 (N_25276,N_25039,N_25054);
nand U25277 (N_25277,N_25110,N_25044);
and U25278 (N_25278,N_25139,N_25090);
nand U25279 (N_25279,N_25049,N_25082);
and U25280 (N_25280,N_25023,N_25123);
nor U25281 (N_25281,N_25097,N_25171);
xor U25282 (N_25282,N_25088,N_25196);
nor U25283 (N_25283,N_25119,N_25158);
nor U25284 (N_25284,N_25031,N_25064);
xnor U25285 (N_25285,N_25000,N_25005);
and U25286 (N_25286,N_25189,N_25192);
nand U25287 (N_25287,N_25008,N_25126);
nor U25288 (N_25288,N_25111,N_25108);
nand U25289 (N_25289,N_25122,N_25029);
or U25290 (N_25290,N_25070,N_25182);
nand U25291 (N_25291,N_25047,N_25115);
nor U25292 (N_25292,N_25009,N_25137);
nor U25293 (N_25293,N_25022,N_25177);
nor U25294 (N_25294,N_25148,N_25081);
nand U25295 (N_25295,N_25066,N_25195);
or U25296 (N_25296,N_25004,N_25025);
nor U25297 (N_25297,N_25083,N_25162);
xor U25298 (N_25298,N_25007,N_25120);
nand U25299 (N_25299,N_25168,N_25180);
nand U25300 (N_25300,N_25156,N_25031);
xor U25301 (N_25301,N_25080,N_25112);
or U25302 (N_25302,N_25061,N_25187);
or U25303 (N_25303,N_25169,N_25116);
or U25304 (N_25304,N_25074,N_25089);
or U25305 (N_25305,N_25051,N_25064);
nand U25306 (N_25306,N_25150,N_25151);
xnor U25307 (N_25307,N_25089,N_25139);
nor U25308 (N_25308,N_25120,N_25012);
and U25309 (N_25309,N_25019,N_25076);
and U25310 (N_25310,N_25172,N_25111);
or U25311 (N_25311,N_25095,N_25170);
nand U25312 (N_25312,N_25052,N_25021);
and U25313 (N_25313,N_25014,N_25129);
or U25314 (N_25314,N_25076,N_25105);
or U25315 (N_25315,N_25165,N_25081);
xor U25316 (N_25316,N_25028,N_25147);
xor U25317 (N_25317,N_25099,N_25181);
xnor U25318 (N_25318,N_25172,N_25147);
or U25319 (N_25319,N_25181,N_25121);
xor U25320 (N_25320,N_25165,N_25014);
nor U25321 (N_25321,N_25120,N_25043);
nor U25322 (N_25322,N_25186,N_25101);
nor U25323 (N_25323,N_25182,N_25088);
and U25324 (N_25324,N_25168,N_25170);
or U25325 (N_25325,N_25089,N_25133);
nand U25326 (N_25326,N_25070,N_25004);
nand U25327 (N_25327,N_25064,N_25127);
nor U25328 (N_25328,N_25017,N_25085);
nor U25329 (N_25329,N_25138,N_25170);
or U25330 (N_25330,N_25145,N_25041);
xor U25331 (N_25331,N_25120,N_25116);
xor U25332 (N_25332,N_25099,N_25162);
xor U25333 (N_25333,N_25128,N_25028);
nand U25334 (N_25334,N_25139,N_25065);
nor U25335 (N_25335,N_25065,N_25060);
nand U25336 (N_25336,N_25061,N_25069);
nor U25337 (N_25337,N_25098,N_25033);
nand U25338 (N_25338,N_25025,N_25173);
or U25339 (N_25339,N_25020,N_25123);
nor U25340 (N_25340,N_25031,N_25008);
or U25341 (N_25341,N_25172,N_25014);
nor U25342 (N_25342,N_25021,N_25197);
nor U25343 (N_25343,N_25058,N_25123);
nor U25344 (N_25344,N_25098,N_25034);
nand U25345 (N_25345,N_25037,N_25195);
or U25346 (N_25346,N_25001,N_25057);
xnor U25347 (N_25347,N_25025,N_25160);
xnor U25348 (N_25348,N_25125,N_25132);
xnor U25349 (N_25349,N_25141,N_25038);
or U25350 (N_25350,N_25190,N_25125);
nor U25351 (N_25351,N_25184,N_25119);
xnor U25352 (N_25352,N_25002,N_25046);
xnor U25353 (N_25353,N_25030,N_25084);
or U25354 (N_25354,N_25097,N_25137);
nor U25355 (N_25355,N_25043,N_25004);
nor U25356 (N_25356,N_25186,N_25153);
or U25357 (N_25357,N_25050,N_25150);
nand U25358 (N_25358,N_25126,N_25065);
nand U25359 (N_25359,N_25008,N_25038);
nor U25360 (N_25360,N_25052,N_25079);
or U25361 (N_25361,N_25080,N_25088);
or U25362 (N_25362,N_25019,N_25066);
xor U25363 (N_25363,N_25031,N_25080);
nand U25364 (N_25364,N_25195,N_25119);
nor U25365 (N_25365,N_25165,N_25164);
nand U25366 (N_25366,N_25005,N_25128);
nand U25367 (N_25367,N_25148,N_25036);
nor U25368 (N_25368,N_25084,N_25049);
or U25369 (N_25369,N_25055,N_25061);
xnor U25370 (N_25370,N_25001,N_25026);
or U25371 (N_25371,N_25000,N_25081);
and U25372 (N_25372,N_25020,N_25096);
xor U25373 (N_25373,N_25119,N_25012);
or U25374 (N_25374,N_25152,N_25135);
nor U25375 (N_25375,N_25129,N_25103);
or U25376 (N_25376,N_25069,N_25199);
and U25377 (N_25377,N_25170,N_25008);
and U25378 (N_25378,N_25024,N_25132);
and U25379 (N_25379,N_25130,N_25045);
and U25380 (N_25380,N_25106,N_25073);
and U25381 (N_25381,N_25086,N_25029);
and U25382 (N_25382,N_25007,N_25100);
and U25383 (N_25383,N_25049,N_25061);
nand U25384 (N_25384,N_25112,N_25023);
or U25385 (N_25385,N_25188,N_25183);
nand U25386 (N_25386,N_25026,N_25119);
nand U25387 (N_25387,N_25079,N_25057);
nor U25388 (N_25388,N_25162,N_25114);
and U25389 (N_25389,N_25080,N_25183);
nor U25390 (N_25390,N_25021,N_25028);
nand U25391 (N_25391,N_25025,N_25108);
or U25392 (N_25392,N_25069,N_25109);
and U25393 (N_25393,N_25053,N_25036);
and U25394 (N_25394,N_25162,N_25110);
nor U25395 (N_25395,N_25083,N_25065);
and U25396 (N_25396,N_25052,N_25043);
and U25397 (N_25397,N_25198,N_25132);
and U25398 (N_25398,N_25164,N_25101);
or U25399 (N_25399,N_25190,N_25004);
or U25400 (N_25400,N_25291,N_25300);
nor U25401 (N_25401,N_25331,N_25380);
or U25402 (N_25402,N_25277,N_25249);
nand U25403 (N_25403,N_25242,N_25229);
and U25404 (N_25404,N_25353,N_25203);
and U25405 (N_25405,N_25234,N_25215);
nor U25406 (N_25406,N_25251,N_25317);
nand U25407 (N_25407,N_25263,N_25398);
and U25408 (N_25408,N_25364,N_25385);
nor U25409 (N_25409,N_25332,N_25301);
or U25410 (N_25410,N_25265,N_25395);
nand U25411 (N_25411,N_25318,N_25302);
or U25412 (N_25412,N_25220,N_25360);
nand U25413 (N_25413,N_25367,N_25206);
nand U25414 (N_25414,N_25337,N_25393);
xor U25415 (N_25415,N_25389,N_25376);
xnor U25416 (N_25416,N_25351,N_25270);
and U25417 (N_25417,N_25333,N_25328);
nand U25418 (N_25418,N_25289,N_25382);
and U25419 (N_25419,N_25299,N_25239);
or U25420 (N_25420,N_25285,N_25288);
and U25421 (N_25421,N_25325,N_25207);
nand U25422 (N_25422,N_25287,N_25227);
or U25423 (N_25423,N_25292,N_25322);
nor U25424 (N_25424,N_25261,N_25241);
and U25425 (N_25425,N_25238,N_25218);
and U25426 (N_25426,N_25280,N_25375);
and U25427 (N_25427,N_25230,N_25305);
or U25428 (N_25428,N_25272,N_25212);
nor U25429 (N_25429,N_25358,N_25345);
nor U25430 (N_25430,N_25315,N_25286);
nor U25431 (N_25431,N_25210,N_25250);
xor U25432 (N_25432,N_25293,N_25271);
nand U25433 (N_25433,N_25278,N_25245);
nor U25434 (N_25434,N_25372,N_25384);
xnor U25435 (N_25435,N_25254,N_25267);
nand U25436 (N_25436,N_25314,N_25205);
or U25437 (N_25437,N_25316,N_25379);
nand U25438 (N_25438,N_25269,N_25327);
nand U25439 (N_25439,N_25303,N_25296);
or U25440 (N_25440,N_25248,N_25324);
nand U25441 (N_25441,N_25223,N_25275);
nand U25442 (N_25442,N_25397,N_25244);
nor U25443 (N_25443,N_25386,N_25309);
and U25444 (N_25444,N_25281,N_25363);
nand U25445 (N_25445,N_25394,N_25214);
and U25446 (N_25446,N_25396,N_25335);
nand U25447 (N_25447,N_25326,N_25336);
nor U25448 (N_25448,N_25355,N_25243);
or U25449 (N_25449,N_25297,N_25264);
xor U25450 (N_25450,N_25334,N_25362);
nand U25451 (N_25451,N_25202,N_25259);
xor U25452 (N_25452,N_25330,N_25252);
nand U25453 (N_25453,N_25258,N_25217);
or U25454 (N_25454,N_25260,N_25295);
xnor U25455 (N_25455,N_25329,N_25356);
xor U25456 (N_25456,N_25304,N_25366);
or U25457 (N_25457,N_25361,N_25392);
and U25458 (N_25458,N_25221,N_25357);
xnor U25459 (N_25459,N_25354,N_25200);
xor U25460 (N_25460,N_25310,N_25344);
nor U25461 (N_25461,N_25348,N_25219);
nand U25462 (N_25462,N_25339,N_25388);
nand U25463 (N_25463,N_25308,N_25283);
and U25464 (N_25464,N_25222,N_25381);
or U25465 (N_25465,N_25232,N_25311);
nand U25466 (N_25466,N_25320,N_25266);
or U25467 (N_25467,N_25284,N_25323);
or U25468 (N_25468,N_25370,N_25236);
and U25469 (N_25469,N_25312,N_25383);
or U25470 (N_25470,N_25313,N_25262);
nand U25471 (N_25471,N_25274,N_25273);
and U25472 (N_25472,N_25365,N_25253);
xnor U25473 (N_25473,N_25225,N_25349);
xor U25474 (N_25474,N_25298,N_25359);
xnor U25475 (N_25475,N_25352,N_25231);
nor U25476 (N_25476,N_25342,N_25226);
nand U25477 (N_25477,N_25390,N_25340);
nand U25478 (N_25478,N_25247,N_25346);
and U25479 (N_25479,N_25368,N_25256);
nor U25480 (N_25480,N_25387,N_25378);
xor U25481 (N_25481,N_25240,N_25290);
nand U25482 (N_25482,N_25341,N_25319);
xor U25483 (N_25483,N_25237,N_25257);
nand U25484 (N_25484,N_25307,N_25228);
nand U25485 (N_25485,N_25369,N_25373);
xnor U25486 (N_25486,N_25201,N_25391);
nand U25487 (N_25487,N_25204,N_25338);
and U25488 (N_25488,N_25268,N_25235);
and U25489 (N_25489,N_25216,N_25347);
xor U25490 (N_25490,N_25374,N_25306);
and U25491 (N_25491,N_25371,N_25294);
nor U25492 (N_25492,N_25208,N_25377);
or U25493 (N_25493,N_25321,N_25276);
or U25494 (N_25494,N_25224,N_25399);
and U25495 (N_25495,N_25211,N_25213);
nand U25496 (N_25496,N_25282,N_25343);
nor U25497 (N_25497,N_25246,N_25255);
xor U25498 (N_25498,N_25279,N_25233);
xnor U25499 (N_25499,N_25209,N_25350);
or U25500 (N_25500,N_25364,N_25287);
or U25501 (N_25501,N_25358,N_25363);
nor U25502 (N_25502,N_25228,N_25229);
nor U25503 (N_25503,N_25225,N_25243);
or U25504 (N_25504,N_25263,N_25343);
nor U25505 (N_25505,N_25202,N_25328);
xor U25506 (N_25506,N_25213,N_25363);
and U25507 (N_25507,N_25274,N_25299);
or U25508 (N_25508,N_25393,N_25203);
nor U25509 (N_25509,N_25284,N_25324);
or U25510 (N_25510,N_25302,N_25323);
nor U25511 (N_25511,N_25239,N_25203);
nand U25512 (N_25512,N_25351,N_25232);
and U25513 (N_25513,N_25214,N_25249);
or U25514 (N_25514,N_25210,N_25311);
nor U25515 (N_25515,N_25349,N_25253);
nor U25516 (N_25516,N_25324,N_25239);
nor U25517 (N_25517,N_25320,N_25238);
or U25518 (N_25518,N_25275,N_25248);
or U25519 (N_25519,N_25315,N_25309);
nor U25520 (N_25520,N_25382,N_25234);
xnor U25521 (N_25521,N_25206,N_25256);
xor U25522 (N_25522,N_25387,N_25243);
nand U25523 (N_25523,N_25231,N_25314);
and U25524 (N_25524,N_25298,N_25356);
nor U25525 (N_25525,N_25279,N_25219);
xnor U25526 (N_25526,N_25313,N_25338);
nor U25527 (N_25527,N_25262,N_25306);
nand U25528 (N_25528,N_25312,N_25380);
and U25529 (N_25529,N_25311,N_25305);
nor U25530 (N_25530,N_25396,N_25345);
nand U25531 (N_25531,N_25277,N_25275);
and U25532 (N_25532,N_25312,N_25256);
nor U25533 (N_25533,N_25395,N_25387);
or U25534 (N_25534,N_25349,N_25297);
nand U25535 (N_25535,N_25362,N_25271);
nand U25536 (N_25536,N_25266,N_25317);
and U25537 (N_25537,N_25277,N_25238);
and U25538 (N_25538,N_25368,N_25275);
and U25539 (N_25539,N_25261,N_25391);
xor U25540 (N_25540,N_25285,N_25328);
xnor U25541 (N_25541,N_25213,N_25296);
nor U25542 (N_25542,N_25260,N_25223);
nand U25543 (N_25543,N_25351,N_25244);
nor U25544 (N_25544,N_25326,N_25253);
nor U25545 (N_25545,N_25303,N_25353);
nand U25546 (N_25546,N_25201,N_25380);
nor U25547 (N_25547,N_25319,N_25215);
and U25548 (N_25548,N_25318,N_25399);
nand U25549 (N_25549,N_25391,N_25326);
xnor U25550 (N_25550,N_25350,N_25279);
and U25551 (N_25551,N_25349,N_25389);
nand U25552 (N_25552,N_25300,N_25349);
or U25553 (N_25553,N_25219,N_25317);
or U25554 (N_25554,N_25330,N_25357);
and U25555 (N_25555,N_25352,N_25271);
xnor U25556 (N_25556,N_25261,N_25302);
or U25557 (N_25557,N_25240,N_25288);
and U25558 (N_25558,N_25321,N_25242);
or U25559 (N_25559,N_25235,N_25287);
xnor U25560 (N_25560,N_25307,N_25283);
nand U25561 (N_25561,N_25289,N_25293);
and U25562 (N_25562,N_25238,N_25367);
and U25563 (N_25563,N_25273,N_25344);
xor U25564 (N_25564,N_25393,N_25253);
xnor U25565 (N_25565,N_25309,N_25236);
or U25566 (N_25566,N_25325,N_25352);
and U25567 (N_25567,N_25290,N_25258);
xnor U25568 (N_25568,N_25219,N_25309);
nand U25569 (N_25569,N_25381,N_25212);
or U25570 (N_25570,N_25390,N_25302);
nor U25571 (N_25571,N_25380,N_25228);
nand U25572 (N_25572,N_25382,N_25282);
nor U25573 (N_25573,N_25298,N_25308);
nor U25574 (N_25574,N_25207,N_25338);
or U25575 (N_25575,N_25285,N_25381);
and U25576 (N_25576,N_25279,N_25356);
or U25577 (N_25577,N_25254,N_25303);
and U25578 (N_25578,N_25280,N_25288);
or U25579 (N_25579,N_25280,N_25212);
and U25580 (N_25580,N_25371,N_25335);
nand U25581 (N_25581,N_25384,N_25327);
nor U25582 (N_25582,N_25349,N_25344);
nand U25583 (N_25583,N_25376,N_25379);
nand U25584 (N_25584,N_25398,N_25333);
and U25585 (N_25585,N_25345,N_25297);
nand U25586 (N_25586,N_25335,N_25271);
nand U25587 (N_25587,N_25343,N_25243);
nor U25588 (N_25588,N_25272,N_25209);
nor U25589 (N_25589,N_25200,N_25323);
and U25590 (N_25590,N_25232,N_25341);
and U25591 (N_25591,N_25207,N_25258);
nand U25592 (N_25592,N_25377,N_25237);
and U25593 (N_25593,N_25265,N_25367);
or U25594 (N_25594,N_25392,N_25310);
and U25595 (N_25595,N_25280,N_25386);
or U25596 (N_25596,N_25288,N_25228);
and U25597 (N_25597,N_25348,N_25293);
or U25598 (N_25598,N_25288,N_25260);
xnor U25599 (N_25599,N_25312,N_25200);
xor U25600 (N_25600,N_25414,N_25523);
nor U25601 (N_25601,N_25453,N_25590);
or U25602 (N_25602,N_25576,N_25521);
xor U25603 (N_25603,N_25489,N_25456);
and U25604 (N_25604,N_25574,N_25567);
and U25605 (N_25605,N_25515,N_25497);
xor U25606 (N_25606,N_25470,N_25540);
nor U25607 (N_25607,N_25500,N_25455);
xnor U25608 (N_25608,N_25416,N_25427);
and U25609 (N_25609,N_25522,N_25437);
and U25610 (N_25610,N_25546,N_25492);
nand U25611 (N_25611,N_25424,N_25578);
and U25612 (N_25612,N_25401,N_25496);
and U25613 (N_25613,N_25431,N_25494);
nor U25614 (N_25614,N_25513,N_25573);
xnor U25615 (N_25615,N_25566,N_25507);
nand U25616 (N_25616,N_25538,N_25529);
xor U25617 (N_25617,N_25563,N_25429);
nand U25618 (N_25618,N_25584,N_25543);
and U25619 (N_25619,N_25545,N_25419);
nand U25620 (N_25620,N_25461,N_25595);
nand U25621 (N_25621,N_25498,N_25537);
nor U25622 (N_25622,N_25508,N_25493);
or U25623 (N_25623,N_25514,N_25482);
nor U25624 (N_25624,N_25555,N_25525);
xor U25625 (N_25625,N_25553,N_25598);
nor U25626 (N_25626,N_25516,N_25532);
xnor U25627 (N_25627,N_25594,N_25559);
xor U25628 (N_25628,N_25432,N_25568);
or U25629 (N_25629,N_25544,N_25491);
nor U25630 (N_25630,N_25487,N_25585);
xor U25631 (N_25631,N_25589,N_25588);
and U25632 (N_25632,N_25435,N_25531);
xor U25633 (N_25633,N_25418,N_25475);
and U25634 (N_25634,N_25448,N_25443);
nand U25635 (N_25635,N_25421,N_25481);
xor U25636 (N_25636,N_25577,N_25423);
or U25637 (N_25637,N_25518,N_25509);
and U25638 (N_25638,N_25548,N_25527);
or U25639 (N_25639,N_25557,N_25445);
xnor U25640 (N_25640,N_25503,N_25413);
nand U25641 (N_25641,N_25474,N_25466);
nand U25642 (N_25642,N_25486,N_25438);
or U25643 (N_25643,N_25417,N_25458);
nand U25644 (N_25644,N_25471,N_25571);
and U25645 (N_25645,N_25406,N_25404);
xnor U25646 (N_25646,N_25441,N_25450);
nand U25647 (N_25647,N_25551,N_25597);
xnor U25648 (N_25648,N_25436,N_25550);
or U25649 (N_25649,N_25463,N_25444);
nor U25650 (N_25650,N_25415,N_25407);
and U25651 (N_25651,N_25465,N_25517);
nand U25652 (N_25652,N_25593,N_25402);
and U25653 (N_25653,N_25542,N_25549);
nor U25654 (N_25654,N_25490,N_25459);
xor U25655 (N_25655,N_25468,N_25512);
and U25656 (N_25656,N_25579,N_25556);
or U25657 (N_25657,N_25575,N_25581);
or U25658 (N_25658,N_25425,N_25564);
and U25659 (N_25659,N_25484,N_25467);
xor U25660 (N_25660,N_25591,N_25505);
or U25661 (N_25661,N_25580,N_25539);
nand U25662 (N_25662,N_25485,N_25569);
and U25663 (N_25663,N_25442,N_25422);
and U25664 (N_25664,N_25510,N_25460);
or U25665 (N_25665,N_25535,N_25451);
or U25666 (N_25666,N_25477,N_25586);
xor U25667 (N_25667,N_25583,N_25526);
xor U25668 (N_25668,N_25530,N_25552);
nand U25669 (N_25669,N_25506,N_25558);
nor U25670 (N_25670,N_25408,N_25480);
nor U25671 (N_25671,N_25454,N_25428);
nor U25672 (N_25672,N_25528,N_25560);
nand U25673 (N_25673,N_25533,N_25504);
or U25674 (N_25674,N_25473,N_25501);
and U25675 (N_25675,N_25440,N_25439);
nor U25676 (N_25676,N_25434,N_25446);
and U25677 (N_25677,N_25405,N_25534);
nor U25678 (N_25678,N_25479,N_25476);
nand U25679 (N_25679,N_25472,N_25449);
nor U25680 (N_25680,N_25587,N_25499);
and U25681 (N_25681,N_25596,N_25547);
nand U25682 (N_25682,N_25478,N_25420);
or U25683 (N_25683,N_25452,N_25599);
nand U25684 (N_25684,N_25511,N_25541);
and U25685 (N_25685,N_25433,N_25412);
xnor U25686 (N_25686,N_25469,N_25536);
and U25687 (N_25687,N_25447,N_25561);
and U25688 (N_25688,N_25524,N_25411);
and U25689 (N_25689,N_25430,N_25554);
and U25690 (N_25690,N_25426,N_25570);
and U25691 (N_25691,N_25483,N_25592);
nand U25692 (N_25692,N_25457,N_25403);
or U25693 (N_25693,N_25410,N_25464);
or U25694 (N_25694,N_25562,N_25400);
xor U25695 (N_25695,N_25565,N_25519);
or U25696 (N_25696,N_25462,N_25495);
or U25697 (N_25697,N_25572,N_25409);
and U25698 (N_25698,N_25488,N_25582);
nand U25699 (N_25699,N_25520,N_25502);
xor U25700 (N_25700,N_25500,N_25582);
and U25701 (N_25701,N_25542,N_25555);
and U25702 (N_25702,N_25585,N_25504);
and U25703 (N_25703,N_25551,N_25425);
nand U25704 (N_25704,N_25543,N_25412);
nor U25705 (N_25705,N_25419,N_25538);
or U25706 (N_25706,N_25552,N_25484);
nand U25707 (N_25707,N_25541,N_25503);
nand U25708 (N_25708,N_25479,N_25403);
nor U25709 (N_25709,N_25488,N_25440);
nand U25710 (N_25710,N_25431,N_25511);
nor U25711 (N_25711,N_25528,N_25456);
or U25712 (N_25712,N_25419,N_25566);
nor U25713 (N_25713,N_25547,N_25454);
nand U25714 (N_25714,N_25592,N_25551);
nor U25715 (N_25715,N_25403,N_25592);
nand U25716 (N_25716,N_25452,N_25438);
xnor U25717 (N_25717,N_25425,N_25472);
nand U25718 (N_25718,N_25587,N_25494);
nor U25719 (N_25719,N_25591,N_25516);
nor U25720 (N_25720,N_25519,N_25466);
and U25721 (N_25721,N_25568,N_25476);
nand U25722 (N_25722,N_25448,N_25518);
nor U25723 (N_25723,N_25497,N_25430);
xnor U25724 (N_25724,N_25454,N_25509);
xnor U25725 (N_25725,N_25577,N_25513);
nand U25726 (N_25726,N_25574,N_25403);
nand U25727 (N_25727,N_25593,N_25523);
xnor U25728 (N_25728,N_25561,N_25551);
or U25729 (N_25729,N_25574,N_25543);
nor U25730 (N_25730,N_25425,N_25470);
or U25731 (N_25731,N_25504,N_25538);
or U25732 (N_25732,N_25561,N_25538);
nor U25733 (N_25733,N_25506,N_25426);
and U25734 (N_25734,N_25418,N_25561);
nor U25735 (N_25735,N_25490,N_25466);
or U25736 (N_25736,N_25499,N_25591);
nor U25737 (N_25737,N_25501,N_25553);
nand U25738 (N_25738,N_25590,N_25445);
xnor U25739 (N_25739,N_25461,N_25505);
nor U25740 (N_25740,N_25575,N_25508);
xor U25741 (N_25741,N_25403,N_25560);
and U25742 (N_25742,N_25462,N_25598);
nand U25743 (N_25743,N_25416,N_25595);
or U25744 (N_25744,N_25496,N_25464);
or U25745 (N_25745,N_25450,N_25434);
and U25746 (N_25746,N_25436,N_25561);
and U25747 (N_25747,N_25480,N_25599);
nor U25748 (N_25748,N_25424,N_25559);
and U25749 (N_25749,N_25481,N_25484);
or U25750 (N_25750,N_25400,N_25418);
and U25751 (N_25751,N_25585,N_25519);
nor U25752 (N_25752,N_25411,N_25417);
nand U25753 (N_25753,N_25591,N_25482);
xor U25754 (N_25754,N_25593,N_25493);
xnor U25755 (N_25755,N_25534,N_25552);
and U25756 (N_25756,N_25405,N_25450);
nand U25757 (N_25757,N_25457,N_25503);
or U25758 (N_25758,N_25591,N_25513);
xnor U25759 (N_25759,N_25519,N_25419);
or U25760 (N_25760,N_25488,N_25484);
nand U25761 (N_25761,N_25462,N_25571);
nor U25762 (N_25762,N_25436,N_25540);
and U25763 (N_25763,N_25462,N_25413);
nor U25764 (N_25764,N_25506,N_25452);
nor U25765 (N_25765,N_25432,N_25435);
nor U25766 (N_25766,N_25407,N_25483);
nor U25767 (N_25767,N_25498,N_25570);
nor U25768 (N_25768,N_25522,N_25574);
or U25769 (N_25769,N_25455,N_25420);
xnor U25770 (N_25770,N_25575,N_25457);
or U25771 (N_25771,N_25463,N_25465);
or U25772 (N_25772,N_25549,N_25584);
nor U25773 (N_25773,N_25598,N_25548);
or U25774 (N_25774,N_25460,N_25466);
nand U25775 (N_25775,N_25487,N_25498);
nor U25776 (N_25776,N_25570,N_25510);
or U25777 (N_25777,N_25499,N_25452);
xnor U25778 (N_25778,N_25511,N_25575);
nand U25779 (N_25779,N_25522,N_25555);
nand U25780 (N_25780,N_25514,N_25515);
and U25781 (N_25781,N_25449,N_25486);
or U25782 (N_25782,N_25524,N_25400);
or U25783 (N_25783,N_25555,N_25599);
nor U25784 (N_25784,N_25474,N_25528);
xor U25785 (N_25785,N_25576,N_25449);
nor U25786 (N_25786,N_25536,N_25448);
nand U25787 (N_25787,N_25473,N_25527);
nand U25788 (N_25788,N_25537,N_25459);
nand U25789 (N_25789,N_25562,N_25475);
nand U25790 (N_25790,N_25455,N_25501);
and U25791 (N_25791,N_25523,N_25522);
nor U25792 (N_25792,N_25534,N_25571);
and U25793 (N_25793,N_25556,N_25479);
nand U25794 (N_25794,N_25409,N_25402);
or U25795 (N_25795,N_25554,N_25466);
or U25796 (N_25796,N_25570,N_25505);
xnor U25797 (N_25797,N_25444,N_25436);
or U25798 (N_25798,N_25443,N_25508);
or U25799 (N_25799,N_25413,N_25488);
nor U25800 (N_25800,N_25757,N_25744);
nor U25801 (N_25801,N_25669,N_25722);
and U25802 (N_25802,N_25738,N_25629);
or U25803 (N_25803,N_25699,N_25636);
or U25804 (N_25804,N_25655,N_25729);
and U25805 (N_25805,N_25670,N_25718);
xor U25806 (N_25806,N_25614,N_25685);
nor U25807 (N_25807,N_25740,N_25657);
nor U25808 (N_25808,N_25688,N_25733);
or U25809 (N_25809,N_25761,N_25696);
and U25810 (N_25810,N_25640,N_25634);
xnor U25811 (N_25811,N_25664,N_25773);
nand U25812 (N_25812,N_25695,N_25608);
nand U25813 (N_25813,N_25754,N_25734);
and U25814 (N_25814,N_25626,N_25735);
nor U25815 (N_25815,N_25790,N_25766);
or U25816 (N_25816,N_25706,N_25715);
or U25817 (N_25817,N_25653,N_25713);
xnor U25818 (N_25818,N_25776,N_25794);
xor U25819 (N_25819,N_25788,N_25707);
nand U25820 (N_25820,N_25753,N_25749);
nor U25821 (N_25821,N_25624,N_25795);
and U25822 (N_25822,N_25779,N_25726);
or U25823 (N_25823,N_25770,N_25642);
or U25824 (N_25824,N_25789,N_25651);
xor U25825 (N_25825,N_25680,N_25625);
nor U25826 (N_25826,N_25727,N_25768);
xor U25827 (N_25827,N_25676,N_25648);
and U25828 (N_25828,N_25792,N_25787);
xor U25829 (N_25829,N_25622,N_25697);
xnor U25830 (N_25830,N_25662,N_25742);
nand U25831 (N_25831,N_25633,N_25791);
and U25832 (N_25832,N_25755,N_25705);
nor U25833 (N_25833,N_25691,N_25674);
nor U25834 (N_25834,N_25668,N_25708);
xnor U25835 (N_25835,N_25635,N_25687);
or U25836 (N_25836,N_25678,N_25796);
and U25837 (N_25837,N_25739,N_25743);
or U25838 (N_25838,N_25702,N_25728);
nor U25839 (N_25839,N_25745,N_25602);
nor U25840 (N_25840,N_25782,N_25660);
nand U25841 (N_25841,N_25617,N_25641);
and U25842 (N_25842,N_25772,N_25725);
nor U25843 (N_25843,N_25701,N_25665);
nand U25844 (N_25844,N_25737,N_25724);
nand U25845 (N_25845,N_25709,N_25760);
nor U25846 (N_25846,N_25656,N_25628);
and U25847 (N_25847,N_25717,N_25777);
nand U25848 (N_25848,N_25730,N_25606);
and U25849 (N_25849,N_25661,N_25767);
nor U25850 (N_25850,N_25667,N_25630);
and U25851 (N_25851,N_25654,N_25682);
or U25852 (N_25852,N_25639,N_25644);
or U25853 (N_25853,N_25720,N_25683);
nand U25854 (N_25854,N_25632,N_25751);
nor U25855 (N_25855,N_25611,N_25603);
or U25856 (N_25856,N_25741,N_25612);
and U25857 (N_25857,N_25693,N_25650);
or U25858 (N_25858,N_25620,N_25769);
xnor U25859 (N_25859,N_25649,N_25659);
xor U25860 (N_25860,N_25619,N_25600);
xor U25861 (N_25861,N_25797,N_25690);
nor U25862 (N_25862,N_25675,N_25613);
nand U25863 (N_25863,N_25646,N_25780);
nor U25864 (N_25864,N_25618,N_25736);
nand U25865 (N_25865,N_25771,N_25643);
xnor U25866 (N_25866,N_25746,N_25694);
nor U25867 (N_25867,N_25714,N_25673);
or U25868 (N_25868,N_25679,N_25627);
nor U25869 (N_25869,N_25677,N_25704);
nor U25870 (N_25870,N_25700,N_25623);
or U25871 (N_25871,N_25616,N_25672);
nor U25872 (N_25872,N_25793,N_25681);
and U25873 (N_25873,N_25658,N_25692);
or U25874 (N_25874,N_25610,N_25703);
or U25875 (N_25875,N_25689,N_25719);
nand U25876 (N_25876,N_25615,N_25786);
or U25877 (N_25877,N_25638,N_25647);
nand U25878 (N_25878,N_25621,N_25710);
nand U25879 (N_25879,N_25775,N_25732);
or U25880 (N_25880,N_25750,N_25604);
and U25881 (N_25881,N_25631,N_25764);
nor U25882 (N_25882,N_25723,N_25609);
xnor U25883 (N_25883,N_25731,N_25686);
nand U25884 (N_25884,N_25663,N_25712);
nand U25885 (N_25885,N_25785,N_25684);
or U25886 (N_25886,N_25666,N_25671);
xnor U25887 (N_25887,N_25765,N_25756);
or U25888 (N_25888,N_25759,N_25652);
xor U25889 (N_25889,N_25778,N_25698);
or U25890 (N_25890,N_25774,N_25601);
nor U25891 (N_25891,N_25763,N_25748);
nand U25892 (N_25892,N_25637,N_25758);
xnor U25893 (N_25893,N_25607,N_25752);
nand U25894 (N_25894,N_25747,N_25711);
nand U25895 (N_25895,N_25783,N_25798);
nor U25896 (N_25896,N_25645,N_25781);
or U25897 (N_25897,N_25762,N_25716);
and U25898 (N_25898,N_25605,N_25721);
nor U25899 (N_25899,N_25799,N_25784);
and U25900 (N_25900,N_25795,N_25676);
and U25901 (N_25901,N_25632,N_25675);
nand U25902 (N_25902,N_25717,N_25723);
and U25903 (N_25903,N_25618,N_25751);
xor U25904 (N_25904,N_25634,N_25715);
nand U25905 (N_25905,N_25618,N_25638);
or U25906 (N_25906,N_25683,N_25692);
xnor U25907 (N_25907,N_25686,N_25792);
xor U25908 (N_25908,N_25793,N_25631);
nand U25909 (N_25909,N_25607,N_25619);
nor U25910 (N_25910,N_25611,N_25769);
nand U25911 (N_25911,N_25740,N_25642);
nor U25912 (N_25912,N_25774,N_25653);
xnor U25913 (N_25913,N_25635,N_25726);
and U25914 (N_25914,N_25738,N_25606);
xor U25915 (N_25915,N_25793,N_25613);
nand U25916 (N_25916,N_25647,N_25729);
nor U25917 (N_25917,N_25741,N_25754);
nand U25918 (N_25918,N_25698,N_25682);
and U25919 (N_25919,N_25623,N_25796);
nor U25920 (N_25920,N_25680,N_25754);
xnor U25921 (N_25921,N_25661,N_25658);
and U25922 (N_25922,N_25770,N_25692);
or U25923 (N_25923,N_25610,N_25712);
and U25924 (N_25924,N_25712,N_25757);
and U25925 (N_25925,N_25699,N_25767);
and U25926 (N_25926,N_25751,N_25774);
or U25927 (N_25927,N_25649,N_25686);
nand U25928 (N_25928,N_25788,N_25779);
xor U25929 (N_25929,N_25757,N_25617);
nand U25930 (N_25930,N_25723,N_25682);
and U25931 (N_25931,N_25769,N_25729);
or U25932 (N_25932,N_25639,N_25665);
nor U25933 (N_25933,N_25673,N_25719);
and U25934 (N_25934,N_25763,N_25670);
nor U25935 (N_25935,N_25621,N_25602);
xor U25936 (N_25936,N_25780,N_25710);
xor U25937 (N_25937,N_25798,N_25746);
nor U25938 (N_25938,N_25787,N_25735);
and U25939 (N_25939,N_25664,N_25785);
nor U25940 (N_25940,N_25654,N_25607);
xor U25941 (N_25941,N_25762,N_25789);
or U25942 (N_25942,N_25649,N_25769);
xnor U25943 (N_25943,N_25602,N_25750);
nand U25944 (N_25944,N_25783,N_25624);
and U25945 (N_25945,N_25726,N_25680);
nand U25946 (N_25946,N_25751,N_25711);
xnor U25947 (N_25947,N_25697,N_25706);
or U25948 (N_25948,N_25639,N_25722);
and U25949 (N_25949,N_25738,N_25697);
xnor U25950 (N_25950,N_25630,N_25750);
nor U25951 (N_25951,N_25692,N_25616);
and U25952 (N_25952,N_25746,N_25714);
or U25953 (N_25953,N_25607,N_25702);
nor U25954 (N_25954,N_25609,N_25710);
and U25955 (N_25955,N_25694,N_25625);
nand U25956 (N_25956,N_25766,N_25723);
xnor U25957 (N_25957,N_25763,N_25673);
nor U25958 (N_25958,N_25727,N_25741);
and U25959 (N_25959,N_25718,N_25782);
and U25960 (N_25960,N_25775,N_25731);
and U25961 (N_25961,N_25619,N_25659);
and U25962 (N_25962,N_25627,N_25674);
or U25963 (N_25963,N_25650,N_25768);
xnor U25964 (N_25964,N_25761,N_25659);
xor U25965 (N_25965,N_25679,N_25696);
nor U25966 (N_25966,N_25711,N_25754);
nand U25967 (N_25967,N_25656,N_25604);
and U25968 (N_25968,N_25690,N_25764);
and U25969 (N_25969,N_25621,N_25760);
xnor U25970 (N_25970,N_25768,N_25773);
nand U25971 (N_25971,N_25742,N_25661);
nor U25972 (N_25972,N_25707,N_25709);
nor U25973 (N_25973,N_25735,N_25767);
or U25974 (N_25974,N_25697,N_25790);
or U25975 (N_25975,N_25797,N_25612);
nand U25976 (N_25976,N_25641,N_25691);
nor U25977 (N_25977,N_25624,N_25727);
and U25978 (N_25978,N_25621,N_25626);
xnor U25979 (N_25979,N_25695,N_25625);
nand U25980 (N_25980,N_25700,N_25784);
and U25981 (N_25981,N_25655,N_25716);
nand U25982 (N_25982,N_25735,N_25667);
xnor U25983 (N_25983,N_25626,N_25761);
nor U25984 (N_25984,N_25672,N_25613);
and U25985 (N_25985,N_25659,N_25747);
and U25986 (N_25986,N_25658,N_25789);
nor U25987 (N_25987,N_25709,N_25677);
or U25988 (N_25988,N_25647,N_25764);
and U25989 (N_25989,N_25712,N_25793);
or U25990 (N_25990,N_25659,N_25671);
xor U25991 (N_25991,N_25678,N_25649);
nand U25992 (N_25992,N_25796,N_25765);
nor U25993 (N_25993,N_25722,N_25603);
nand U25994 (N_25994,N_25701,N_25661);
or U25995 (N_25995,N_25627,N_25790);
or U25996 (N_25996,N_25730,N_25649);
nor U25997 (N_25997,N_25665,N_25728);
and U25998 (N_25998,N_25731,N_25745);
and U25999 (N_25999,N_25664,N_25757);
and U26000 (N_26000,N_25983,N_25823);
or U26001 (N_26001,N_25954,N_25842);
xnor U26002 (N_26002,N_25966,N_25905);
nand U26003 (N_26003,N_25888,N_25994);
xnor U26004 (N_26004,N_25865,N_25924);
nand U26005 (N_26005,N_25858,N_25897);
xor U26006 (N_26006,N_25876,N_25894);
or U26007 (N_26007,N_25805,N_25998);
nand U26008 (N_26008,N_25863,N_25943);
nand U26009 (N_26009,N_25811,N_25980);
and U26010 (N_26010,N_25871,N_25856);
or U26011 (N_26011,N_25893,N_25997);
xnor U26012 (N_26012,N_25907,N_25984);
or U26013 (N_26013,N_25806,N_25898);
and U26014 (N_26014,N_25908,N_25970);
or U26015 (N_26015,N_25890,N_25835);
nor U26016 (N_26016,N_25962,N_25839);
and U26017 (N_26017,N_25985,N_25853);
nand U26018 (N_26018,N_25800,N_25855);
nand U26019 (N_26019,N_25934,N_25827);
xnor U26020 (N_26020,N_25838,N_25901);
nor U26021 (N_26021,N_25953,N_25830);
or U26022 (N_26022,N_25967,N_25957);
nand U26023 (N_26023,N_25919,N_25882);
or U26024 (N_26024,N_25933,N_25891);
or U26025 (N_26025,N_25921,N_25955);
and U26026 (N_26026,N_25875,N_25964);
nor U26027 (N_26027,N_25836,N_25889);
xor U26028 (N_26028,N_25941,N_25944);
or U26029 (N_26029,N_25996,N_25850);
and U26030 (N_26030,N_25990,N_25815);
nand U26031 (N_26031,N_25832,N_25900);
and U26032 (N_26032,N_25961,N_25834);
nand U26033 (N_26033,N_25862,N_25860);
or U26034 (N_26034,N_25988,N_25932);
or U26035 (N_26035,N_25959,N_25958);
xnor U26036 (N_26036,N_25975,N_25825);
or U26037 (N_26037,N_25820,N_25952);
nor U26038 (N_26038,N_25948,N_25803);
and U26039 (N_26039,N_25982,N_25885);
and U26040 (N_26040,N_25881,N_25991);
and U26041 (N_26041,N_25945,N_25937);
nor U26042 (N_26042,N_25971,N_25965);
or U26043 (N_26043,N_25981,N_25930);
and U26044 (N_26044,N_25931,N_25849);
xor U26045 (N_26045,N_25939,N_25845);
and U26046 (N_26046,N_25977,N_25883);
nor U26047 (N_26047,N_25804,N_25826);
and U26048 (N_26048,N_25949,N_25868);
nand U26049 (N_26049,N_25851,N_25950);
nand U26050 (N_26050,N_25879,N_25947);
or U26051 (N_26051,N_25816,N_25940);
and U26052 (N_26052,N_25963,N_25916);
nor U26053 (N_26053,N_25837,N_25802);
xnor U26054 (N_26054,N_25911,N_25843);
nor U26055 (N_26055,N_25809,N_25848);
nand U26056 (N_26056,N_25818,N_25925);
and U26057 (N_26057,N_25833,N_25844);
and U26058 (N_26058,N_25903,N_25841);
or U26059 (N_26059,N_25928,N_25866);
nor U26060 (N_26060,N_25920,N_25935);
and U26061 (N_26061,N_25895,N_25810);
nor U26062 (N_26062,N_25912,N_25979);
nor U26063 (N_26063,N_25884,N_25859);
nand U26064 (N_26064,N_25847,N_25951);
or U26065 (N_26065,N_25887,N_25880);
xor U26066 (N_26066,N_25929,N_25918);
or U26067 (N_26067,N_25993,N_25814);
and U26068 (N_26068,N_25813,N_25995);
xor U26069 (N_26069,N_25822,N_25909);
and U26070 (N_26070,N_25854,N_25904);
nor U26071 (N_26071,N_25999,N_25978);
or U26072 (N_26072,N_25892,N_25956);
or U26073 (N_26073,N_25828,N_25913);
nor U26074 (N_26074,N_25922,N_25886);
xnor U26075 (N_26075,N_25872,N_25992);
and U26076 (N_26076,N_25829,N_25869);
nor U26077 (N_26077,N_25846,N_25986);
or U26078 (N_26078,N_25821,N_25972);
nand U26079 (N_26079,N_25852,N_25867);
xor U26080 (N_26080,N_25808,N_25927);
or U26081 (N_26081,N_25974,N_25969);
xor U26082 (N_26082,N_25917,N_25936);
nor U26083 (N_26083,N_25812,N_25801);
or U26084 (N_26084,N_25899,N_25861);
nor U26085 (N_26085,N_25926,N_25878);
nor U26086 (N_26086,N_25914,N_25938);
and U26087 (N_26087,N_25864,N_25923);
xnor U26088 (N_26088,N_25946,N_25968);
and U26089 (N_26089,N_25831,N_25989);
or U26090 (N_26090,N_25874,N_25915);
nand U26091 (N_26091,N_25906,N_25910);
nor U26092 (N_26092,N_25987,N_25873);
nor U26093 (N_26093,N_25960,N_25896);
xor U26094 (N_26094,N_25817,N_25870);
nor U26095 (N_26095,N_25819,N_25840);
or U26096 (N_26096,N_25976,N_25877);
nor U26097 (N_26097,N_25902,N_25942);
nand U26098 (N_26098,N_25824,N_25857);
nor U26099 (N_26099,N_25973,N_25807);
nor U26100 (N_26100,N_25852,N_25908);
xor U26101 (N_26101,N_25846,N_25981);
or U26102 (N_26102,N_25894,N_25803);
xor U26103 (N_26103,N_25837,N_25929);
xor U26104 (N_26104,N_25836,N_25834);
and U26105 (N_26105,N_25815,N_25962);
nand U26106 (N_26106,N_25874,N_25809);
and U26107 (N_26107,N_25916,N_25848);
xnor U26108 (N_26108,N_25913,N_25811);
xnor U26109 (N_26109,N_25945,N_25840);
nand U26110 (N_26110,N_25801,N_25810);
and U26111 (N_26111,N_25932,N_25881);
nand U26112 (N_26112,N_25933,N_25955);
and U26113 (N_26113,N_25996,N_25972);
and U26114 (N_26114,N_25968,N_25835);
nand U26115 (N_26115,N_25970,N_25822);
and U26116 (N_26116,N_25845,N_25865);
or U26117 (N_26117,N_25826,N_25835);
or U26118 (N_26118,N_25868,N_25900);
nand U26119 (N_26119,N_25892,N_25906);
or U26120 (N_26120,N_25909,N_25929);
nand U26121 (N_26121,N_25881,N_25983);
and U26122 (N_26122,N_25988,N_25930);
nand U26123 (N_26123,N_25957,N_25945);
and U26124 (N_26124,N_25856,N_25807);
or U26125 (N_26125,N_25979,N_25929);
or U26126 (N_26126,N_25867,N_25938);
nor U26127 (N_26127,N_25935,N_25994);
nand U26128 (N_26128,N_25988,N_25964);
nor U26129 (N_26129,N_25856,N_25924);
nor U26130 (N_26130,N_25932,N_25964);
nor U26131 (N_26131,N_25854,N_25884);
nor U26132 (N_26132,N_25943,N_25966);
nor U26133 (N_26133,N_25803,N_25853);
xor U26134 (N_26134,N_25828,N_25809);
nand U26135 (N_26135,N_25957,N_25845);
xnor U26136 (N_26136,N_25974,N_25978);
or U26137 (N_26137,N_25823,N_25953);
or U26138 (N_26138,N_25927,N_25843);
xor U26139 (N_26139,N_25943,N_25969);
and U26140 (N_26140,N_25934,N_25971);
or U26141 (N_26141,N_25957,N_25937);
and U26142 (N_26142,N_25813,N_25949);
or U26143 (N_26143,N_25857,N_25897);
xnor U26144 (N_26144,N_25989,N_25865);
or U26145 (N_26145,N_25998,N_25869);
nand U26146 (N_26146,N_25922,N_25806);
xor U26147 (N_26147,N_25998,N_25930);
or U26148 (N_26148,N_25941,N_25931);
xor U26149 (N_26149,N_25988,N_25920);
nor U26150 (N_26150,N_25956,N_25937);
nor U26151 (N_26151,N_25894,N_25847);
nand U26152 (N_26152,N_25851,N_25864);
nand U26153 (N_26153,N_25992,N_25991);
nand U26154 (N_26154,N_25977,N_25967);
and U26155 (N_26155,N_25945,N_25904);
or U26156 (N_26156,N_25989,N_25923);
nor U26157 (N_26157,N_25804,N_25939);
xnor U26158 (N_26158,N_25966,N_25861);
nand U26159 (N_26159,N_25870,N_25998);
and U26160 (N_26160,N_25815,N_25853);
nor U26161 (N_26161,N_25928,N_25932);
or U26162 (N_26162,N_25877,N_25904);
and U26163 (N_26163,N_25987,N_25841);
nand U26164 (N_26164,N_25950,N_25814);
and U26165 (N_26165,N_25832,N_25951);
nand U26166 (N_26166,N_25806,N_25918);
or U26167 (N_26167,N_25907,N_25833);
and U26168 (N_26168,N_25952,N_25840);
xnor U26169 (N_26169,N_25885,N_25858);
nor U26170 (N_26170,N_25989,N_25880);
or U26171 (N_26171,N_25828,N_25946);
nor U26172 (N_26172,N_25815,N_25827);
nor U26173 (N_26173,N_25878,N_25948);
nand U26174 (N_26174,N_25990,N_25818);
and U26175 (N_26175,N_25900,N_25856);
nor U26176 (N_26176,N_25809,N_25807);
nor U26177 (N_26177,N_25948,N_25810);
xnor U26178 (N_26178,N_25892,N_25813);
nor U26179 (N_26179,N_25860,N_25953);
or U26180 (N_26180,N_25932,N_25971);
or U26181 (N_26181,N_25825,N_25947);
nand U26182 (N_26182,N_25976,N_25950);
nor U26183 (N_26183,N_25897,N_25983);
and U26184 (N_26184,N_25910,N_25891);
and U26185 (N_26185,N_25965,N_25822);
or U26186 (N_26186,N_25875,N_25834);
and U26187 (N_26187,N_25819,N_25938);
nor U26188 (N_26188,N_25896,N_25889);
nor U26189 (N_26189,N_25871,N_25995);
and U26190 (N_26190,N_25867,N_25861);
or U26191 (N_26191,N_25899,N_25858);
or U26192 (N_26192,N_25998,N_25893);
nor U26193 (N_26193,N_25902,N_25929);
and U26194 (N_26194,N_25985,N_25937);
and U26195 (N_26195,N_25908,N_25828);
xor U26196 (N_26196,N_25802,N_25809);
and U26197 (N_26197,N_25935,N_25865);
or U26198 (N_26198,N_25879,N_25852);
or U26199 (N_26199,N_25913,N_25960);
xor U26200 (N_26200,N_26061,N_26005);
and U26201 (N_26201,N_26027,N_26145);
nor U26202 (N_26202,N_26163,N_26065);
nand U26203 (N_26203,N_26055,N_26081);
and U26204 (N_26204,N_26096,N_26199);
and U26205 (N_26205,N_26113,N_26095);
or U26206 (N_26206,N_26020,N_26013);
or U26207 (N_26207,N_26181,N_26058);
and U26208 (N_26208,N_26141,N_26149);
nand U26209 (N_26209,N_26067,N_26093);
nand U26210 (N_26210,N_26080,N_26110);
nand U26211 (N_26211,N_26084,N_26085);
xnor U26212 (N_26212,N_26125,N_26073);
xnor U26213 (N_26213,N_26015,N_26017);
nor U26214 (N_26214,N_26046,N_26071);
or U26215 (N_26215,N_26038,N_26120);
nand U26216 (N_26216,N_26083,N_26197);
xnor U26217 (N_26217,N_26025,N_26063);
xnor U26218 (N_26218,N_26036,N_26170);
or U26219 (N_26219,N_26030,N_26042);
or U26220 (N_26220,N_26147,N_26186);
nor U26221 (N_26221,N_26105,N_26010);
nor U26222 (N_26222,N_26131,N_26161);
and U26223 (N_26223,N_26012,N_26086);
and U26224 (N_26224,N_26182,N_26164);
nand U26225 (N_26225,N_26040,N_26000);
and U26226 (N_26226,N_26088,N_26158);
xor U26227 (N_26227,N_26142,N_26069);
nor U26228 (N_26228,N_26139,N_26099);
nand U26229 (N_26229,N_26014,N_26137);
nor U26230 (N_26230,N_26072,N_26003);
and U26231 (N_26231,N_26074,N_26165);
or U26232 (N_26232,N_26190,N_26053);
nor U26233 (N_26233,N_26060,N_26172);
or U26234 (N_26234,N_26196,N_26114);
xnor U26235 (N_26235,N_26009,N_26091);
nor U26236 (N_26236,N_26117,N_26011);
nor U26237 (N_26237,N_26127,N_26001);
nand U26238 (N_26238,N_26188,N_26126);
nor U26239 (N_26239,N_26066,N_26050);
nor U26240 (N_26240,N_26097,N_26191);
nand U26241 (N_26241,N_26189,N_26129);
nand U26242 (N_26242,N_26123,N_26180);
and U26243 (N_26243,N_26037,N_26192);
and U26244 (N_26244,N_26168,N_26174);
or U26245 (N_26245,N_26140,N_26079);
and U26246 (N_26246,N_26023,N_26008);
or U26247 (N_26247,N_26116,N_26106);
nor U26248 (N_26248,N_26185,N_26184);
nor U26249 (N_26249,N_26135,N_26103);
and U26250 (N_26250,N_26193,N_26018);
xnor U26251 (N_26251,N_26183,N_26049);
nor U26252 (N_26252,N_26100,N_26138);
nand U26253 (N_26253,N_26162,N_26173);
xor U26254 (N_26254,N_26104,N_26102);
and U26255 (N_26255,N_26016,N_26143);
or U26256 (N_26256,N_26068,N_26152);
xor U26257 (N_26257,N_26178,N_26035);
or U26258 (N_26258,N_26052,N_26054);
and U26259 (N_26259,N_26156,N_26087);
nor U26260 (N_26260,N_26109,N_26177);
nor U26261 (N_26261,N_26124,N_26128);
or U26262 (N_26262,N_26176,N_26033);
nand U26263 (N_26263,N_26167,N_26146);
nand U26264 (N_26264,N_26078,N_26032);
and U26265 (N_26265,N_26029,N_26090);
xor U26266 (N_26266,N_26155,N_26059);
or U26267 (N_26267,N_26175,N_26019);
nor U26268 (N_26268,N_26169,N_26151);
nand U26269 (N_26269,N_26062,N_26198);
xor U26270 (N_26270,N_26118,N_26107);
or U26271 (N_26271,N_26021,N_26166);
or U26272 (N_26272,N_26121,N_26101);
or U26273 (N_26273,N_26075,N_26187);
xnor U26274 (N_26274,N_26006,N_26108);
xnor U26275 (N_26275,N_26115,N_26026);
or U26276 (N_26276,N_26039,N_26092);
and U26277 (N_26277,N_26041,N_26195);
nand U26278 (N_26278,N_26004,N_26130);
or U26279 (N_26279,N_26076,N_26007);
and U26280 (N_26280,N_26070,N_26150);
xnor U26281 (N_26281,N_26144,N_26194);
or U26282 (N_26282,N_26134,N_26044);
or U26283 (N_26283,N_26119,N_26034);
nand U26284 (N_26284,N_26064,N_26002);
or U26285 (N_26285,N_26094,N_26122);
and U26286 (N_26286,N_26153,N_26132);
nand U26287 (N_26287,N_26159,N_26077);
and U26288 (N_26288,N_26112,N_26024);
xnor U26289 (N_26289,N_26171,N_26048);
or U26290 (N_26290,N_26056,N_26057);
nor U26291 (N_26291,N_26148,N_26045);
or U26292 (N_26292,N_26179,N_26022);
xor U26293 (N_26293,N_26157,N_26111);
or U26294 (N_26294,N_26082,N_26154);
nand U26295 (N_26295,N_26136,N_26089);
or U26296 (N_26296,N_26043,N_26031);
nand U26297 (N_26297,N_26028,N_26098);
and U26298 (N_26298,N_26133,N_26047);
nand U26299 (N_26299,N_26051,N_26160);
and U26300 (N_26300,N_26109,N_26070);
nor U26301 (N_26301,N_26069,N_26092);
nor U26302 (N_26302,N_26182,N_26090);
nand U26303 (N_26303,N_26062,N_26089);
or U26304 (N_26304,N_26140,N_26053);
and U26305 (N_26305,N_26185,N_26038);
nor U26306 (N_26306,N_26168,N_26059);
xor U26307 (N_26307,N_26190,N_26032);
and U26308 (N_26308,N_26051,N_26140);
nand U26309 (N_26309,N_26182,N_26038);
xnor U26310 (N_26310,N_26025,N_26159);
nand U26311 (N_26311,N_26177,N_26097);
nand U26312 (N_26312,N_26062,N_26179);
nand U26313 (N_26313,N_26097,N_26099);
or U26314 (N_26314,N_26118,N_26199);
xor U26315 (N_26315,N_26121,N_26180);
xor U26316 (N_26316,N_26035,N_26112);
nor U26317 (N_26317,N_26158,N_26185);
nor U26318 (N_26318,N_26178,N_26111);
nand U26319 (N_26319,N_26084,N_26190);
xor U26320 (N_26320,N_26154,N_26110);
and U26321 (N_26321,N_26139,N_26013);
nand U26322 (N_26322,N_26194,N_26177);
xor U26323 (N_26323,N_26185,N_26075);
and U26324 (N_26324,N_26123,N_26112);
or U26325 (N_26325,N_26171,N_26107);
nor U26326 (N_26326,N_26183,N_26142);
nor U26327 (N_26327,N_26133,N_26072);
and U26328 (N_26328,N_26194,N_26063);
and U26329 (N_26329,N_26059,N_26128);
or U26330 (N_26330,N_26100,N_26065);
or U26331 (N_26331,N_26102,N_26155);
nor U26332 (N_26332,N_26006,N_26058);
and U26333 (N_26333,N_26140,N_26065);
xnor U26334 (N_26334,N_26140,N_26197);
nand U26335 (N_26335,N_26096,N_26101);
and U26336 (N_26336,N_26045,N_26147);
or U26337 (N_26337,N_26195,N_26001);
nand U26338 (N_26338,N_26089,N_26146);
nor U26339 (N_26339,N_26183,N_26148);
xnor U26340 (N_26340,N_26108,N_26061);
and U26341 (N_26341,N_26094,N_26044);
or U26342 (N_26342,N_26084,N_26033);
nor U26343 (N_26343,N_26193,N_26127);
nor U26344 (N_26344,N_26062,N_26186);
and U26345 (N_26345,N_26018,N_26033);
nand U26346 (N_26346,N_26061,N_26017);
nand U26347 (N_26347,N_26047,N_26142);
xor U26348 (N_26348,N_26092,N_26191);
xnor U26349 (N_26349,N_26175,N_26073);
and U26350 (N_26350,N_26020,N_26111);
xnor U26351 (N_26351,N_26142,N_26106);
xor U26352 (N_26352,N_26091,N_26163);
or U26353 (N_26353,N_26032,N_26126);
or U26354 (N_26354,N_26011,N_26070);
nand U26355 (N_26355,N_26187,N_26190);
and U26356 (N_26356,N_26120,N_26113);
and U26357 (N_26357,N_26152,N_26168);
or U26358 (N_26358,N_26106,N_26035);
nand U26359 (N_26359,N_26163,N_26052);
nand U26360 (N_26360,N_26073,N_26019);
and U26361 (N_26361,N_26145,N_26068);
or U26362 (N_26362,N_26058,N_26119);
nand U26363 (N_26363,N_26014,N_26062);
nand U26364 (N_26364,N_26144,N_26183);
and U26365 (N_26365,N_26154,N_26096);
nand U26366 (N_26366,N_26074,N_26142);
nand U26367 (N_26367,N_26015,N_26153);
or U26368 (N_26368,N_26081,N_26085);
nor U26369 (N_26369,N_26065,N_26133);
nand U26370 (N_26370,N_26035,N_26060);
nor U26371 (N_26371,N_26105,N_26085);
or U26372 (N_26372,N_26010,N_26029);
and U26373 (N_26373,N_26000,N_26181);
and U26374 (N_26374,N_26006,N_26174);
nor U26375 (N_26375,N_26011,N_26089);
or U26376 (N_26376,N_26089,N_26109);
and U26377 (N_26377,N_26005,N_26000);
xnor U26378 (N_26378,N_26021,N_26182);
nand U26379 (N_26379,N_26064,N_26140);
xnor U26380 (N_26380,N_26133,N_26045);
and U26381 (N_26381,N_26061,N_26125);
nor U26382 (N_26382,N_26020,N_26007);
nor U26383 (N_26383,N_26118,N_26187);
and U26384 (N_26384,N_26094,N_26164);
nor U26385 (N_26385,N_26181,N_26007);
xor U26386 (N_26386,N_26116,N_26082);
xnor U26387 (N_26387,N_26061,N_26016);
or U26388 (N_26388,N_26170,N_26031);
nand U26389 (N_26389,N_26107,N_26054);
xor U26390 (N_26390,N_26167,N_26115);
nand U26391 (N_26391,N_26016,N_26069);
or U26392 (N_26392,N_26144,N_26198);
or U26393 (N_26393,N_26169,N_26152);
or U26394 (N_26394,N_26190,N_26050);
and U26395 (N_26395,N_26104,N_26148);
and U26396 (N_26396,N_26091,N_26177);
nor U26397 (N_26397,N_26090,N_26129);
xor U26398 (N_26398,N_26143,N_26181);
nand U26399 (N_26399,N_26183,N_26083);
or U26400 (N_26400,N_26241,N_26211);
xnor U26401 (N_26401,N_26365,N_26351);
nand U26402 (N_26402,N_26218,N_26399);
and U26403 (N_26403,N_26254,N_26301);
nor U26404 (N_26404,N_26347,N_26208);
xor U26405 (N_26405,N_26333,N_26345);
nand U26406 (N_26406,N_26242,N_26348);
or U26407 (N_26407,N_26258,N_26205);
and U26408 (N_26408,N_26277,N_26363);
nor U26409 (N_26409,N_26248,N_26369);
nand U26410 (N_26410,N_26366,N_26284);
or U26411 (N_26411,N_26316,N_26393);
nand U26412 (N_26412,N_26278,N_26377);
or U26413 (N_26413,N_26265,N_26297);
xnor U26414 (N_26414,N_26331,N_26384);
or U26415 (N_26415,N_26302,N_26370);
or U26416 (N_26416,N_26314,N_26246);
nor U26417 (N_26417,N_26274,N_26255);
nor U26418 (N_26418,N_26360,N_26334);
and U26419 (N_26419,N_26210,N_26263);
or U26420 (N_26420,N_26381,N_26332);
and U26421 (N_26421,N_26359,N_26286);
and U26422 (N_26422,N_26323,N_26256);
and U26423 (N_26423,N_26391,N_26388);
nor U26424 (N_26424,N_26229,N_26321);
nand U26425 (N_26425,N_26244,N_26367);
nor U26426 (N_26426,N_26220,N_26392);
or U26427 (N_26427,N_26230,N_26235);
xor U26428 (N_26428,N_26298,N_26260);
xnor U26429 (N_26429,N_26259,N_26398);
nor U26430 (N_26430,N_26269,N_26342);
nand U26431 (N_26431,N_26335,N_26231);
xor U26432 (N_26432,N_26293,N_26253);
nor U26433 (N_26433,N_26315,N_26380);
xnor U26434 (N_26434,N_26313,N_26336);
nor U26435 (N_26435,N_26238,N_26202);
nand U26436 (N_26436,N_26320,N_26225);
nand U26437 (N_26437,N_26206,N_26352);
nor U26438 (N_26438,N_26326,N_26328);
nor U26439 (N_26439,N_26249,N_26362);
nor U26440 (N_26440,N_26330,N_26361);
or U26441 (N_26441,N_26243,N_26350);
nor U26442 (N_26442,N_26287,N_26329);
or U26443 (N_26443,N_26250,N_26295);
nor U26444 (N_26444,N_26273,N_26291);
and U26445 (N_26445,N_26397,N_26276);
and U26446 (N_26446,N_26378,N_26324);
and U26447 (N_26447,N_26288,N_26371);
and U26448 (N_26448,N_26309,N_26306);
nor U26449 (N_26449,N_26312,N_26212);
nor U26450 (N_26450,N_26261,N_26354);
xor U26451 (N_26451,N_26376,N_26307);
nor U26452 (N_26452,N_26214,N_26358);
and U26453 (N_26453,N_26386,N_26394);
and U26454 (N_26454,N_26383,N_26264);
xor U26455 (N_26455,N_26285,N_26389);
or U26456 (N_26456,N_26234,N_26237);
nand U26457 (N_26457,N_26281,N_26222);
nor U26458 (N_26458,N_26353,N_26305);
xnor U26459 (N_26459,N_26340,N_26279);
nor U26460 (N_26460,N_26357,N_26201);
or U26461 (N_26461,N_26387,N_26343);
nand U26462 (N_26462,N_26251,N_26325);
or U26463 (N_26463,N_26200,N_26346);
and U26464 (N_26464,N_26204,N_26322);
or U26465 (N_26465,N_26339,N_26247);
and U26466 (N_26466,N_26266,N_26221);
and U26467 (N_26467,N_26318,N_26268);
or U26468 (N_26468,N_26310,N_26395);
or U26469 (N_26469,N_26292,N_26217);
nor U26470 (N_26470,N_26213,N_26344);
nor U26471 (N_26471,N_26304,N_26372);
or U26472 (N_26472,N_26319,N_26207);
nor U26473 (N_26473,N_26368,N_26272);
xnor U26474 (N_26474,N_26396,N_26233);
nand U26475 (N_26475,N_26262,N_26209);
or U26476 (N_26476,N_26223,N_26215);
or U26477 (N_26477,N_26390,N_26338);
and U26478 (N_26478,N_26252,N_26240);
nand U26479 (N_26479,N_26349,N_26228);
or U26480 (N_26480,N_26232,N_26300);
or U26481 (N_26481,N_26373,N_26303);
nand U26482 (N_26482,N_26337,N_26270);
or U26483 (N_26483,N_26267,N_26226);
nor U26484 (N_26484,N_26282,N_26374);
nand U26485 (N_26485,N_26271,N_26382);
nand U26486 (N_26486,N_26216,N_26245);
or U26487 (N_26487,N_26239,N_26275);
nor U26488 (N_26488,N_26385,N_26224);
and U26489 (N_26489,N_26289,N_26379);
nand U26490 (N_26490,N_26294,N_26283);
and U26491 (N_26491,N_26375,N_26296);
nand U26492 (N_26492,N_26299,N_26355);
xor U26493 (N_26493,N_26219,N_26308);
nand U26494 (N_26494,N_26203,N_26227);
nand U26495 (N_26495,N_26311,N_26341);
xnor U26496 (N_26496,N_26280,N_26290);
xnor U26497 (N_26497,N_26257,N_26364);
and U26498 (N_26498,N_26356,N_26317);
or U26499 (N_26499,N_26236,N_26327);
and U26500 (N_26500,N_26347,N_26286);
and U26501 (N_26501,N_26324,N_26317);
and U26502 (N_26502,N_26298,N_26385);
nand U26503 (N_26503,N_26215,N_26380);
nand U26504 (N_26504,N_26397,N_26278);
nand U26505 (N_26505,N_26342,N_26261);
and U26506 (N_26506,N_26276,N_26333);
and U26507 (N_26507,N_26230,N_26252);
nor U26508 (N_26508,N_26263,N_26274);
nor U26509 (N_26509,N_26359,N_26358);
and U26510 (N_26510,N_26261,N_26252);
and U26511 (N_26511,N_26308,N_26320);
or U26512 (N_26512,N_26303,N_26272);
nor U26513 (N_26513,N_26210,N_26318);
nand U26514 (N_26514,N_26334,N_26252);
or U26515 (N_26515,N_26340,N_26222);
and U26516 (N_26516,N_26397,N_26353);
nor U26517 (N_26517,N_26226,N_26225);
and U26518 (N_26518,N_26365,N_26388);
nand U26519 (N_26519,N_26363,N_26341);
or U26520 (N_26520,N_26288,N_26369);
or U26521 (N_26521,N_26280,N_26388);
or U26522 (N_26522,N_26297,N_26388);
nand U26523 (N_26523,N_26357,N_26265);
or U26524 (N_26524,N_26280,N_26332);
and U26525 (N_26525,N_26369,N_26250);
or U26526 (N_26526,N_26298,N_26397);
nand U26527 (N_26527,N_26231,N_26396);
or U26528 (N_26528,N_26332,N_26207);
xnor U26529 (N_26529,N_26313,N_26398);
and U26530 (N_26530,N_26347,N_26389);
nor U26531 (N_26531,N_26379,N_26254);
nor U26532 (N_26532,N_26228,N_26252);
nor U26533 (N_26533,N_26242,N_26376);
and U26534 (N_26534,N_26316,N_26315);
or U26535 (N_26535,N_26301,N_26327);
nor U26536 (N_26536,N_26207,N_26381);
xor U26537 (N_26537,N_26361,N_26277);
or U26538 (N_26538,N_26384,N_26377);
or U26539 (N_26539,N_26287,N_26223);
or U26540 (N_26540,N_26282,N_26395);
xor U26541 (N_26541,N_26359,N_26287);
nand U26542 (N_26542,N_26312,N_26260);
nor U26543 (N_26543,N_26247,N_26212);
or U26544 (N_26544,N_26319,N_26313);
and U26545 (N_26545,N_26254,N_26296);
and U26546 (N_26546,N_26253,N_26393);
or U26547 (N_26547,N_26281,N_26382);
and U26548 (N_26548,N_26330,N_26275);
or U26549 (N_26549,N_26398,N_26280);
or U26550 (N_26550,N_26333,N_26351);
nand U26551 (N_26551,N_26235,N_26339);
nand U26552 (N_26552,N_26358,N_26206);
xnor U26553 (N_26553,N_26263,N_26244);
or U26554 (N_26554,N_26270,N_26268);
and U26555 (N_26555,N_26304,N_26320);
nor U26556 (N_26556,N_26361,N_26356);
xnor U26557 (N_26557,N_26255,N_26290);
nand U26558 (N_26558,N_26379,N_26318);
and U26559 (N_26559,N_26383,N_26292);
nor U26560 (N_26560,N_26208,N_26355);
and U26561 (N_26561,N_26350,N_26229);
and U26562 (N_26562,N_26341,N_26297);
nand U26563 (N_26563,N_26358,N_26223);
nor U26564 (N_26564,N_26373,N_26377);
nor U26565 (N_26565,N_26270,N_26242);
or U26566 (N_26566,N_26231,N_26225);
or U26567 (N_26567,N_26385,N_26356);
nor U26568 (N_26568,N_26396,N_26228);
and U26569 (N_26569,N_26337,N_26342);
or U26570 (N_26570,N_26354,N_26284);
nand U26571 (N_26571,N_26287,N_26347);
nand U26572 (N_26572,N_26237,N_26310);
nand U26573 (N_26573,N_26339,N_26284);
or U26574 (N_26574,N_26298,N_26395);
or U26575 (N_26575,N_26243,N_26217);
nand U26576 (N_26576,N_26318,N_26249);
nor U26577 (N_26577,N_26324,N_26345);
xnor U26578 (N_26578,N_26212,N_26206);
nor U26579 (N_26579,N_26371,N_26265);
xnor U26580 (N_26580,N_26390,N_26251);
and U26581 (N_26581,N_26306,N_26235);
xor U26582 (N_26582,N_26228,N_26243);
or U26583 (N_26583,N_26263,N_26284);
and U26584 (N_26584,N_26305,N_26255);
nor U26585 (N_26585,N_26214,N_26241);
nor U26586 (N_26586,N_26369,N_26299);
nand U26587 (N_26587,N_26396,N_26282);
or U26588 (N_26588,N_26227,N_26390);
nand U26589 (N_26589,N_26241,N_26335);
nand U26590 (N_26590,N_26396,N_26257);
and U26591 (N_26591,N_26216,N_26248);
or U26592 (N_26592,N_26253,N_26269);
nor U26593 (N_26593,N_26330,N_26295);
or U26594 (N_26594,N_26230,N_26277);
nand U26595 (N_26595,N_26285,N_26362);
xnor U26596 (N_26596,N_26391,N_26364);
and U26597 (N_26597,N_26294,N_26371);
and U26598 (N_26598,N_26343,N_26204);
and U26599 (N_26599,N_26247,N_26276);
or U26600 (N_26600,N_26462,N_26487);
or U26601 (N_26601,N_26498,N_26473);
and U26602 (N_26602,N_26412,N_26468);
nand U26603 (N_26603,N_26515,N_26556);
and U26604 (N_26604,N_26507,N_26585);
nor U26605 (N_26605,N_26534,N_26416);
xnor U26606 (N_26606,N_26547,N_26566);
or U26607 (N_26607,N_26550,N_26489);
nand U26608 (N_26608,N_26434,N_26400);
nor U26609 (N_26609,N_26413,N_26436);
and U26610 (N_26610,N_26432,N_26450);
xor U26611 (N_26611,N_26441,N_26465);
nand U26612 (N_26612,N_26483,N_26414);
nand U26613 (N_26613,N_26578,N_26563);
nand U26614 (N_26614,N_26418,N_26423);
or U26615 (N_26615,N_26417,N_26580);
nand U26616 (N_26616,N_26577,N_26594);
xor U26617 (N_26617,N_26530,N_26470);
nor U26618 (N_26618,N_26497,N_26519);
or U26619 (N_26619,N_26479,N_26404);
or U26620 (N_26620,N_26491,N_26539);
or U26621 (N_26621,N_26407,N_26512);
nor U26622 (N_26622,N_26527,N_26456);
nor U26623 (N_26623,N_26503,N_26453);
and U26624 (N_26624,N_26542,N_26435);
nand U26625 (N_26625,N_26583,N_26559);
xor U26626 (N_26626,N_26537,N_26403);
nor U26627 (N_26627,N_26447,N_26525);
xnor U26628 (N_26628,N_26562,N_26558);
and U26629 (N_26629,N_26457,N_26471);
xor U26630 (N_26630,N_26523,N_26579);
and U26631 (N_26631,N_26484,N_26406);
and U26632 (N_26632,N_26409,N_26575);
and U26633 (N_26633,N_26474,N_26415);
or U26634 (N_26634,N_26442,N_26514);
nor U26635 (N_26635,N_26561,N_26596);
nor U26636 (N_26636,N_26463,N_26564);
nor U26637 (N_26637,N_26475,N_26521);
nor U26638 (N_26638,N_26439,N_26428);
nor U26639 (N_26639,N_26421,N_26531);
nand U26640 (N_26640,N_26524,N_26422);
nand U26641 (N_26641,N_26482,N_26501);
and U26642 (N_26642,N_26509,N_26528);
and U26643 (N_26643,N_26576,N_26591);
and U26644 (N_26644,N_26593,N_26598);
xnor U26645 (N_26645,N_26536,N_26533);
or U26646 (N_26646,N_26466,N_26455);
nor U26647 (N_26647,N_26557,N_26540);
and U26648 (N_26648,N_26546,N_26518);
or U26649 (N_26649,N_26590,N_26448);
nor U26650 (N_26650,N_26568,N_26516);
nor U26651 (N_26651,N_26510,N_26460);
xor U26652 (N_26652,N_26438,N_26597);
and U26653 (N_26653,N_26488,N_26410);
and U26654 (N_26654,N_26437,N_26419);
xor U26655 (N_26655,N_26451,N_26567);
nand U26656 (N_26656,N_26425,N_26467);
or U26657 (N_26657,N_26511,N_26552);
or U26658 (N_26658,N_26469,N_26493);
nor U26659 (N_26659,N_26582,N_26459);
or U26660 (N_26660,N_26508,N_26573);
or U26661 (N_26661,N_26526,N_26443);
nor U26662 (N_26662,N_26545,N_26586);
or U26663 (N_26663,N_26553,N_26560);
or U26664 (N_26664,N_26420,N_26587);
and U26665 (N_26665,N_26569,N_26485);
nand U26666 (N_26666,N_26431,N_26541);
and U26667 (N_26667,N_26506,N_26424);
and U26668 (N_26668,N_26500,N_26520);
or U26669 (N_26669,N_26571,N_26551);
or U26670 (N_26670,N_26529,N_26490);
nand U26671 (N_26671,N_26555,N_26408);
nor U26672 (N_26672,N_26445,N_26532);
nor U26673 (N_26673,N_26472,N_26427);
nor U26674 (N_26674,N_26452,N_26599);
nor U26675 (N_26675,N_26495,N_26574);
xor U26676 (N_26676,N_26589,N_26544);
nand U26677 (N_26677,N_26581,N_26543);
and U26678 (N_26678,N_26478,N_26461);
and U26679 (N_26679,N_26446,N_26405);
and U26680 (N_26680,N_26538,N_26458);
or U26681 (N_26681,N_26480,N_26426);
nor U26682 (N_26682,N_26433,N_26595);
xnor U26683 (N_26683,N_26588,N_26499);
or U26684 (N_26684,N_26496,N_26505);
and U26685 (N_26685,N_26411,N_26584);
nand U26686 (N_26686,N_26430,N_26522);
nor U26687 (N_26687,N_26401,N_26570);
nand U26688 (N_26688,N_26502,N_26449);
and U26689 (N_26689,N_26494,N_26492);
or U26690 (N_26690,N_26592,N_26554);
nor U26691 (N_26691,N_26464,N_26486);
and U26692 (N_26692,N_26477,N_26444);
xnor U26693 (N_26693,N_26440,N_26549);
xor U26694 (N_26694,N_26535,N_26517);
and U26695 (N_26695,N_26565,N_26454);
and U26696 (N_26696,N_26481,N_26429);
nand U26697 (N_26697,N_26402,N_26572);
nand U26698 (N_26698,N_26504,N_26476);
xnor U26699 (N_26699,N_26513,N_26548);
nand U26700 (N_26700,N_26434,N_26446);
or U26701 (N_26701,N_26528,N_26597);
nand U26702 (N_26702,N_26511,N_26506);
xnor U26703 (N_26703,N_26579,N_26581);
or U26704 (N_26704,N_26500,N_26421);
or U26705 (N_26705,N_26515,N_26579);
nand U26706 (N_26706,N_26448,N_26477);
nand U26707 (N_26707,N_26426,N_26546);
xor U26708 (N_26708,N_26403,N_26418);
nand U26709 (N_26709,N_26533,N_26430);
or U26710 (N_26710,N_26427,N_26421);
and U26711 (N_26711,N_26440,N_26508);
and U26712 (N_26712,N_26504,N_26474);
nor U26713 (N_26713,N_26491,N_26513);
or U26714 (N_26714,N_26412,N_26453);
or U26715 (N_26715,N_26472,N_26585);
and U26716 (N_26716,N_26415,N_26572);
xnor U26717 (N_26717,N_26475,N_26510);
or U26718 (N_26718,N_26439,N_26467);
nor U26719 (N_26719,N_26416,N_26424);
xnor U26720 (N_26720,N_26552,N_26477);
or U26721 (N_26721,N_26451,N_26555);
nand U26722 (N_26722,N_26413,N_26553);
xor U26723 (N_26723,N_26440,N_26497);
xnor U26724 (N_26724,N_26491,N_26510);
and U26725 (N_26725,N_26405,N_26550);
nor U26726 (N_26726,N_26439,N_26406);
and U26727 (N_26727,N_26424,N_26533);
nor U26728 (N_26728,N_26403,N_26471);
nand U26729 (N_26729,N_26419,N_26569);
nand U26730 (N_26730,N_26540,N_26526);
nand U26731 (N_26731,N_26467,N_26562);
or U26732 (N_26732,N_26543,N_26532);
or U26733 (N_26733,N_26539,N_26564);
nor U26734 (N_26734,N_26580,N_26472);
xnor U26735 (N_26735,N_26547,N_26578);
nor U26736 (N_26736,N_26502,N_26539);
nand U26737 (N_26737,N_26521,N_26552);
nor U26738 (N_26738,N_26532,N_26437);
xor U26739 (N_26739,N_26417,N_26540);
nand U26740 (N_26740,N_26452,N_26445);
and U26741 (N_26741,N_26474,N_26499);
or U26742 (N_26742,N_26426,N_26403);
or U26743 (N_26743,N_26483,N_26552);
nand U26744 (N_26744,N_26534,N_26432);
and U26745 (N_26745,N_26570,N_26548);
nor U26746 (N_26746,N_26464,N_26460);
nand U26747 (N_26747,N_26557,N_26524);
or U26748 (N_26748,N_26478,N_26407);
and U26749 (N_26749,N_26469,N_26590);
xor U26750 (N_26750,N_26449,N_26496);
or U26751 (N_26751,N_26537,N_26567);
nand U26752 (N_26752,N_26546,N_26437);
xnor U26753 (N_26753,N_26415,N_26465);
nand U26754 (N_26754,N_26500,N_26514);
nand U26755 (N_26755,N_26557,N_26579);
nor U26756 (N_26756,N_26450,N_26510);
or U26757 (N_26757,N_26481,N_26525);
nor U26758 (N_26758,N_26408,N_26536);
and U26759 (N_26759,N_26402,N_26587);
nand U26760 (N_26760,N_26453,N_26537);
nand U26761 (N_26761,N_26495,N_26567);
nor U26762 (N_26762,N_26421,N_26450);
xor U26763 (N_26763,N_26512,N_26473);
nand U26764 (N_26764,N_26541,N_26565);
nand U26765 (N_26765,N_26555,N_26480);
and U26766 (N_26766,N_26488,N_26553);
or U26767 (N_26767,N_26508,N_26480);
and U26768 (N_26768,N_26508,N_26490);
or U26769 (N_26769,N_26501,N_26525);
xor U26770 (N_26770,N_26590,N_26453);
xnor U26771 (N_26771,N_26421,N_26550);
nor U26772 (N_26772,N_26423,N_26560);
and U26773 (N_26773,N_26420,N_26573);
xor U26774 (N_26774,N_26470,N_26407);
or U26775 (N_26775,N_26444,N_26580);
or U26776 (N_26776,N_26527,N_26458);
xnor U26777 (N_26777,N_26562,N_26570);
nor U26778 (N_26778,N_26533,N_26402);
or U26779 (N_26779,N_26420,N_26452);
and U26780 (N_26780,N_26420,N_26592);
nand U26781 (N_26781,N_26457,N_26452);
and U26782 (N_26782,N_26585,N_26480);
xor U26783 (N_26783,N_26559,N_26502);
or U26784 (N_26784,N_26576,N_26413);
xnor U26785 (N_26785,N_26538,N_26594);
nor U26786 (N_26786,N_26508,N_26598);
and U26787 (N_26787,N_26469,N_26548);
xnor U26788 (N_26788,N_26436,N_26468);
nor U26789 (N_26789,N_26435,N_26571);
nand U26790 (N_26790,N_26566,N_26440);
nor U26791 (N_26791,N_26419,N_26446);
and U26792 (N_26792,N_26489,N_26546);
nand U26793 (N_26793,N_26412,N_26580);
xor U26794 (N_26794,N_26411,N_26406);
or U26795 (N_26795,N_26475,N_26407);
nor U26796 (N_26796,N_26450,N_26438);
and U26797 (N_26797,N_26469,N_26506);
and U26798 (N_26798,N_26476,N_26563);
xor U26799 (N_26799,N_26422,N_26550);
xor U26800 (N_26800,N_26793,N_26792);
nor U26801 (N_26801,N_26611,N_26649);
and U26802 (N_26802,N_26702,N_26716);
and U26803 (N_26803,N_26652,N_26607);
nor U26804 (N_26804,N_26646,N_26747);
nand U26805 (N_26805,N_26633,N_26643);
or U26806 (N_26806,N_26679,N_26713);
and U26807 (N_26807,N_26710,N_26757);
or U26808 (N_26808,N_26615,N_26619);
nand U26809 (N_26809,N_26794,N_26778);
or U26810 (N_26810,N_26651,N_26623);
xnor U26811 (N_26811,N_26715,N_26630);
nand U26812 (N_26812,N_26682,N_26637);
xor U26813 (N_26813,N_26610,N_26684);
xor U26814 (N_26814,N_26670,N_26791);
or U26815 (N_26815,N_26730,N_26740);
and U26816 (N_26816,N_26654,N_26688);
and U26817 (N_26817,N_26663,N_26734);
and U26818 (N_26818,N_26746,N_26602);
nor U26819 (N_26819,N_26647,N_26711);
and U26820 (N_26820,N_26661,N_26770);
or U26821 (N_26821,N_26726,N_26681);
xnor U26822 (N_26822,N_26763,N_26600);
nand U26823 (N_26823,N_26714,N_26621);
and U26824 (N_26824,N_26634,N_26674);
nor U26825 (N_26825,N_26613,N_26790);
and U26826 (N_26826,N_26744,N_26699);
and U26827 (N_26827,N_26781,N_26616);
xnor U26828 (N_26828,N_26754,N_26627);
nand U26829 (N_26829,N_26690,N_26689);
nand U26830 (N_26830,N_26625,N_26709);
xnor U26831 (N_26831,N_26717,N_26776);
xnor U26832 (N_26832,N_26760,N_26631);
nand U26833 (N_26833,N_26641,N_26669);
nand U26834 (N_26834,N_26635,N_26788);
and U26835 (N_26835,N_26624,N_26782);
xor U26836 (N_26836,N_26737,N_26756);
nor U26837 (N_26837,N_26604,N_26609);
and U26838 (N_26838,N_26695,N_26777);
nand U26839 (N_26839,N_26771,N_26706);
and U26840 (N_26840,N_26729,N_26718);
nand U26841 (N_26841,N_26626,N_26755);
xnor U26842 (N_26842,N_26725,N_26666);
xor U26843 (N_26843,N_26759,N_26748);
and U26844 (N_26844,N_26766,N_26603);
nand U26845 (N_26845,N_26796,N_26692);
or U26846 (N_26846,N_26783,N_26799);
nor U26847 (N_26847,N_26798,N_26693);
nor U26848 (N_26848,N_26787,N_26617);
or U26849 (N_26849,N_26698,N_26638);
xor U26850 (N_26850,N_26780,N_26785);
nand U26851 (N_26851,N_26675,N_26753);
and U26852 (N_26852,N_26605,N_26705);
nor U26853 (N_26853,N_26697,N_26700);
nor U26854 (N_26854,N_26636,N_26752);
nand U26855 (N_26855,N_26696,N_26742);
or U26856 (N_26856,N_26601,N_26680);
xnor U26857 (N_26857,N_26648,N_26797);
or U26858 (N_26858,N_26673,N_26655);
or U26859 (N_26859,N_26677,N_26743);
or U26860 (N_26860,N_26614,N_26775);
and U26861 (N_26861,N_26704,N_26618);
or U26862 (N_26862,N_26632,N_26768);
or U26863 (N_26863,N_26741,N_26691);
and U26864 (N_26864,N_26694,N_26721);
nand U26865 (N_26865,N_26620,N_26733);
and U26866 (N_26866,N_26660,N_26749);
or U26867 (N_26867,N_26645,N_26758);
nor U26868 (N_26868,N_26779,N_26640);
xor U26869 (N_26869,N_26720,N_26685);
xor U26870 (N_26870,N_26750,N_26656);
nand U26871 (N_26871,N_26761,N_26658);
or U26872 (N_26872,N_26784,N_26774);
nor U26873 (N_26873,N_26629,N_26722);
and U26874 (N_26874,N_26606,N_26686);
xnor U26875 (N_26875,N_26664,N_26653);
nand U26876 (N_26876,N_26659,N_26765);
nand U26877 (N_26877,N_26767,N_26657);
xnor U26878 (N_26878,N_26642,N_26703);
nor U26879 (N_26879,N_26724,N_26732);
nor U26880 (N_26880,N_26665,N_26727);
or U26881 (N_26881,N_26751,N_26769);
nand U26882 (N_26882,N_26712,N_26683);
xnor U26883 (N_26883,N_26736,N_26668);
or U26884 (N_26884,N_26707,N_26676);
or U26885 (N_26885,N_26701,N_26719);
xnor U26886 (N_26886,N_26662,N_26687);
and U26887 (N_26887,N_26612,N_26639);
nor U26888 (N_26888,N_26795,N_26735);
nor U26889 (N_26889,N_26745,N_26731);
or U26890 (N_26890,N_26608,N_26678);
nor U26891 (N_26891,N_26628,N_26667);
nand U26892 (N_26892,N_26672,N_26764);
or U26893 (N_26893,N_26739,N_26738);
and U26894 (N_26894,N_26789,N_26773);
xnor U26895 (N_26895,N_26622,N_26723);
or U26896 (N_26896,N_26708,N_26762);
nand U26897 (N_26897,N_26728,N_26650);
and U26898 (N_26898,N_26786,N_26644);
nor U26899 (N_26899,N_26671,N_26772);
xnor U26900 (N_26900,N_26786,N_26789);
or U26901 (N_26901,N_26781,N_26700);
nor U26902 (N_26902,N_26652,N_26780);
nor U26903 (N_26903,N_26688,N_26774);
xor U26904 (N_26904,N_26730,N_26791);
and U26905 (N_26905,N_26644,N_26767);
nor U26906 (N_26906,N_26740,N_26648);
or U26907 (N_26907,N_26722,N_26632);
and U26908 (N_26908,N_26672,N_26663);
and U26909 (N_26909,N_26767,N_26791);
and U26910 (N_26910,N_26696,N_26714);
xor U26911 (N_26911,N_26605,N_26688);
and U26912 (N_26912,N_26682,N_26799);
or U26913 (N_26913,N_26754,N_26766);
xor U26914 (N_26914,N_26636,N_26634);
nor U26915 (N_26915,N_26728,N_26707);
or U26916 (N_26916,N_26728,N_26749);
and U26917 (N_26917,N_26657,N_26734);
xor U26918 (N_26918,N_26781,N_26629);
and U26919 (N_26919,N_26780,N_26690);
xor U26920 (N_26920,N_26696,N_26700);
nor U26921 (N_26921,N_26756,N_26705);
and U26922 (N_26922,N_26717,N_26759);
xor U26923 (N_26923,N_26781,N_26637);
and U26924 (N_26924,N_26798,N_26727);
and U26925 (N_26925,N_26700,N_26756);
nor U26926 (N_26926,N_26608,N_26702);
nand U26927 (N_26927,N_26605,N_26664);
and U26928 (N_26928,N_26679,N_26772);
nand U26929 (N_26929,N_26672,N_26773);
xor U26930 (N_26930,N_26768,N_26697);
nand U26931 (N_26931,N_26642,N_26686);
and U26932 (N_26932,N_26667,N_26713);
nand U26933 (N_26933,N_26669,N_26757);
and U26934 (N_26934,N_26771,N_26641);
nand U26935 (N_26935,N_26679,N_26761);
and U26936 (N_26936,N_26625,N_26675);
or U26937 (N_26937,N_26779,N_26736);
xor U26938 (N_26938,N_26627,N_26685);
xnor U26939 (N_26939,N_26677,N_26753);
xor U26940 (N_26940,N_26661,N_26797);
nand U26941 (N_26941,N_26727,N_26661);
xor U26942 (N_26942,N_26796,N_26762);
xnor U26943 (N_26943,N_26662,N_26673);
nand U26944 (N_26944,N_26799,N_26757);
or U26945 (N_26945,N_26782,N_26623);
nand U26946 (N_26946,N_26730,N_26690);
xor U26947 (N_26947,N_26797,N_26655);
xor U26948 (N_26948,N_26733,N_26713);
and U26949 (N_26949,N_26727,N_26745);
and U26950 (N_26950,N_26746,N_26727);
and U26951 (N_26951,N_26697,N_26670);
xor U26952 (N_26952,N_26736,N_26703);
nand U26953 (N_26953,N_26600,N_26753);
and U26954 (N_26954,N_26660,N_26733);
or U26955 (N_26955,N_26795,N_26646);
xnor U26956 (N_26956,N_26754,N_26663);
nand U26957 (N_26957,N_26690,N_26688);
xor U26958 (N_26958,N_26614,N_26617);
nor U26959 (N_26959,N_26727,N_26774);
nand U26960 (N_26960,N_26674,N_26658);
or U26961 (N_26961,N_26622,N_26691);
nand U26962 (N_26962,N_26737,N_26746);
xnor U26963 (N_26963,N_26625,N_26695);
or U26964 (N_26964,N_26717,N_26767);
and U26965 (N_26965,N_26609,N_26727);
or U26966 (N_26966,N_26710,N_26601);
xnor U26967 (N_26967,N_26691,N_26733);
xnor U26968 (N_26968,N_26788,N_26730);
nor U26969 (N_26969,N_26776,N_26713);
or U26970 (N_26970,N_26792,N_26653);
nand U26971 (N_26971,N_26661,N_26716);
xnor U26972 (N_26972,N_26698,N_26692);
and U26973 (N_26973,N_26658,N_26637);
nor U26974 (N_26974,N_26762,N_26675);
nand U26975 (N_26975,N_26753,N_26733);
and U26976 (N_26976,N_26765,N_26693);
nor U26977 (N_26977,N_26614,N_26678);
nand U26978 (N_26978,N_26752,N_26669);
nor U26979 (N_26979,N_26698,N_26642);
xor U26980 (N_26980,N_26649,N_26762);
nor U26981 (N_26981,N_26688,N_26616);
nor U26982 (N_26982,N_26753,N_26693);
nand U26983 (N_26983,N_26613,N_26638);
and U26984 (N_26984,N_26746,N_26642);
nand U26985 (N_26985,N_26773,N_26608);
and U26986 (N_26986,N_26676,N_26729);
nand U26987 (N_26987,N_26635,N_26701);
xor U26988 (N_26988,N_26669,N_26767);
nor U26989 (N_26989,N_26730,N_26670);
or U26990 (N_26990,N_26726,N_26740);
nand U26991 (N_26991,N_26750,N_26659);
xnor U26992 (N_26992,N_26656,N_26655);
xor U26993 (N_26993,N_26611,N_26740);
nor U26994 (N_26994,N_26708,N_26756);
xor U26995 (N_26995,N_26683,N_26611);
xor U26996 (N_26996,N_26745,N_26730);
or U26997 (N_26997,N_26711,N_26708);
and U26998 (N_26998,N_26757,N_26692);
and U26999 (N_26999,N_26636,N_26708);
xnor U27000 (N_27000,N_26850,N_26961);
nor U27001 (N_27001,N_26976,N_26889);
and U27002 (N_27002,N_26873,N_26855);
or U27003 (N_27003,N_26859,N_26864);
or U27004 (N_27004,N_26836,N_26970);
nand U27005 (N_27005,N_26877,N_26931);
nand U27006 (N_27006,N_26977,N_26974);
nor U27007 (N_27007,N_26915,N_26923);
nand U27008 (N_27008,N_26980,N_26929);
xor U27009 (N_27009,N_26806,N_26817);
and U27010 (N_27010,N_26904,N_26868);
xnor U27011 (N_27011,N_26853,N_26852);
nand U27012 (N_27012,N_26835,N_26825);
nand U27013 (N_27013,N_26919,N_26858);
nor U27014 (N_27014,N_26870,N_26813);
xnor U27015 (N_27015,N_26972,N_26905);
or U27016 (N_27016,N_26883,N_26869);
xor U27017 (N_27017,N_26935,N_26992);
xor U27018 (N_27018,N_26899,N_26914);
nor U27019 (N_27019,N_26936,N_26903);
xor U27020 (N_27020,N_26824,N_26885);
or U27021 (N_27021,N_26981,N_26998);
nand U27022 (N_27022,N_26909,N_26847);
or U27023 (N_27023,N_26930,N_26967);
and U27024 (N_27024,N_26938,N_26928);
xnor U27025 (N_27025,N_26900,N_26818);
nor U27026 (N_27026,N_26865,N_26962);
xor U27027 (N_27027,N_26990,N_26941);
nor U27028 (N_27028,N_26827,N_26879);
or U27029 (N_27029,N_26861,N_26902);
or U27030 (N_27030,N_26907,N_26964);
xnor U27031 (N_27031,N_26893,N_26839);
xor U27032 (N_27032,N_26815,N_26888);
nand U27033 (N_27033,N_26988,N_26921);
nor U27034 (N_27034,N_26840,N_26841);
and U27035 (N_27035,N_26978,N_26801);
or U27036 (N_27036,N_26809,N_26917);
xnor U27037 (N_27037,N_26922,N_26856);
xnor U27038 (N_27038,N_26854,N_26802);
or U27039 (N_27039,N_26830,N_26822);
and U27040 (N_27040,N_26881,N_26829);
and U27041 (N_27041,N_26804,N_26811);
and U27042 (N_27042,N_26983,N_26913);
or U27043 (N_27043,N_26860,N_26866);
nand U27044 (N_27044,N_26947,N_26969);
or U27045 (N_27045,N_26934,N_26956);
nand U27046 (N_27046,N_26901,N_26832);
and U27047 (N_27047,N_26871,N_26842);
or U27048 (N_27048,N_26987,N_26942);
nor U27049 (N_27049,N_26872,N_26966);
nand U27050 (N_27050,N_26918,N_26912);
or U27051 (N_27051,N_26939,N_26985);
and U27052 (N_27052,N_26882,N_26807);
nand U27053 (N_27053,N_26857,N_26989);
and U27054 (N_27054,N_26927,N_26810);
nand U27055 (N_27055,N_26991,N_26932);
nand U27056 (N_27056,N_26895,N_26803);
xnor U27057 (N_27057,N_26819,N_26958);
and U27058 (N_27058,N_26837,N_26875);
nand U27059 (N_27059,N_26826,N_26960);
nand U27060 (N_27060,N_26816,N_26876);
xor U27061 (N_27061,N_26880,N_26925);
xor U27062 (N_27062,N_26821,N_26805);
xor U27063 (N_27063,N_26954,N_26926);
or U27064 (N_27064,N_26812,N_26973);
xnor U27065 (N_27065,N_26995,N_26844);
nor U27066 (N_27066,N_26999,N_26924);
and U27067 (N_27067,N_26949,N_26823);
and U27068 (N_27068,N_26937,N_26982);
xnor U27069 (N_27069,N_26993,N_26948);
xor U27070 (N_27070,N_26996,N_26979);
xor U27071 (N_27071,N_26833,N_26968);
xor U27072 (N_27072,N_26952,N_26944);
nor U27073 (N_27073,N_26862,N_26814);
nand U27074 (N_27074,N_26984,N_26890);
nand U27075 (N_27075,N_26874,N_26846);
or U27076 (N_27076,N_26943,N_26955);
nand U27077 (N_27077,N_26911,N_26916);
or U27078 (N_27078,N_26878,N_26959);
xor U27079 (N_27079,N_26845,N_26994);
xor U27080 (N_27080,N_26886,N_26965);
xnor U27081 (N_27081,N_26891,N_26851);
nor U27082 (N_27082,N_26945,N_26953);
and U27083 (N_27083,N_26838,N_26892);
nor U27084 (N_27084,N_26951,N_26940);
nor U27085 (N_27085,N_26997,N_26828);
xor U27086 (N_27086,N_26887,N_26820);
xnor U27087 (N_27087,N_26946,N_26867);
nor U27088 (N_27088,N_26957,N_26975);
and U27089 (N_27089,N_26910,N_26986);
xor U27090 (N_27090,N_26808,N_26800);
nand U27091 (N_27091,N_26884,N_26896);
nand U27092 (N_27092,N_26834,N_26971);
and U27093 (N_27093,N_26863,N_26906);
nand U27094 (N_27094,N_26849,N_26933);
nor U27095 (N_27095,N_26848,N_26894);
nand U27096 (N_27096,N_26920,N_26908);
nand U27097 (N_27097,N_26897,N_26898);
nor U27098 (N_27098,N_26963,N_26843);
nor U27099 (N_27099,N_26950,N_26831);
xor U27100 (N_27100,N_26836,N_26957);
and U27101 (N_27101,N_26817,N_26914);
xor U27102 (N_27102,N_26922,N_26869);
xnor U27103 (N_27103,N_26868,N_26812);
nand U27104 (N_27104,N_26843,N_26999);
nand U27105 (N_27105,N_26894,N_26902);
nor U27106 (N_27106,N_26837,N_26901);
nand U27107 (N_27107,N_26818,N_26977);
or U27108 (N_27108,N_26934,N_26960);
nor U27109 (N_27109,N_26888,N_26960);
xnor U27110 (N_27110,N_26982,N_26927);
nor U27111 (N_27111,N_26965,N_26940);
or U27112 (N_27112,N_26866,N_26804);
xnor U27113 (N_27113,N_26955,N_26866);
xnor U27114 (N_27114,N_26875,N_26872);
nand U27115 (N_27115,N_26964,N_26982);
xor U27116 (N_27116,N_26974,N_26804);
nand U27117 (N_27117,N_26844,N_26936);
nand U27118 (N_27118,N_26829,N_26816);
nor U27119 (N_27119,N_26828,N_26867);
nor U27120 (N_27120,N_26990,N_26818);
nand U27121 (N_27121,N_26848,N_26919);
nand U27122 (N_27122,N_26934,N_26985);
nor U27123 (N_27123,N_26957,N_26902);
and U27124 (N_27124,N_26939,N_26894);
nand U27125 (N_27125,N_26869,N_26889);
or U27126 (N_27126,N_26981,N_26942);
xor U27127 (N_27127,N_26852,N_26941);
xnor U27128 (N_27128,N_26989,N_26944);
or U27129 (N_27129,N_26948,N_26891);
and U27130 (N_27130,N_26960,N_26900);
or U27131 (N_27131,N_26953,N_26904);
and U27132 (N_27132,N_26835,N_26848);
and U27133 (N_27133,N_26953,N_26829);
or U27134 (N_27134,N_26805,N_26818);
nand U27135 (N_27135,N_26906,N_26990);
xnor U27136 (N_27136,N_26984,N_26957);
nor U27137 (N_27137,N_26936,N_26901);
nand U27138 (N_27138,N_26820,N_26847);
and U27139 (N_27139,N_26960,N_26861);
and U27140 (N_27140,N_26913,N_26831);
nor U27141 (N_27141,N_26815,N_26852);
xnor U27142 (N_27142,N_26867,N_26971);
xor U27143 (N_27143,N_26828,N_26812);
xor U27144 (N_27144,N_26976,N_26972);
or U27145 (N_27145,N_26820,N_26917);
nand U27146 (N_27146,N_26833,N_26929);
or U27147 (N_27147,N_26916,N_26848);
nor U27148 (N_27148,N_26975,N_26825);
or U27149 (N_27149,N_26909,N_26940);
or U27150 (N_27150,N_26884,N_26963);
nand U27151 (N_27151,N_26923,N_26842);
nand U27152 (N_27152,N_26886,N_26824);
or U27153 (N_27153,N_26964,N_26804);
xnor U27154 (N_27154,N_26955,N_26935);
nor U27155 (N_27155,N_26957,N_26832);
nand U27156 (N_27156,N_26803,N_26836);
xnor U27157 (N_27157,N_26873,N_26899);
or U27158 (N_27158,N_26897,N_26995);
nor U27159 (N_27159,N_26954,N_26915);
or U27160 (N_27160,N_26876,N_26945);
or U27161 (N_27161,N_26889,N_26816);
or U27162 (N_27162,N_26874,N_26934);
and U27163 (N_27163,N_26939,N_26962);
and U27164 (N_27164,N_26909,N_26921);
or U27165 (N_27165,N_26823,N_26892);
or U27166 (N_27166,N_26864,N_26834);
or U27167 (N_27167,N_26896,N_26823);
nor U27168 (N_27168,N_26869,N_26945);
xor U27169 (N_27169,N_26995,N_26876);
nand U27170 (N_27170,N_26969,N_26884);
nand U27171 (N_27171,N_26970,N_26895);
xnor U27172 (N_27172,N_26983,N_26896);
nand U27173 (N_27173,N_26924,N_26848);
and U27174 (N_27174,N_26893,N_26900);
nor U27175 (N_27175,N_26926,N_26937);
and U27176 (N_27176,N_26849,N_26998);
or U27177 (N_27177,N_26823,N_26866);
and U27178 (N_27178,N_26856,N_26982);
xor U27179 (N_27179,N_26935,N_26946);
and U27180 (N_27180,N_26890,N_26987);
or U27181 (N_27181,N_26881,N_26917);
nand U27182 (N_27182,N_26971,N_26868);
xor U27183 (N_27183,N_26833,N_26921);
or U27184 (N_27184,N_26898,N_26831);
and U27185 (N_27185,N_26914,N_26951);
nand U27186 (N_27186,N_26843,N_26936);
nand U27187 (N_27187,N_26925,N_26814);
and U27188 (N_27188,N_26827,N_26945);
nand U27189 (N_27189,N_26887,N_26967);
and U27190 (N_27190,N_26875,N_26927);
and U27191 (N_27191,N_26837,N_26934);
xor U27192 (N_27192,N_26858,N_26996);
xnor U27193 (N_27193,N_26812,N_26830);
or U27194 (N_27194,N_26935,N_26862);
xor U27195 (N_27195,N_26939,N_26877);
nor U27196 (N_27196,N_26874,N_26902);
xor U27197 (N_27197,N_26891,N_26843);
xnor U27198 (N_27198,N_26882,N_26825);
nand U27199 (N_27199,N_26879,N_26993);
xnor U27200 (N_27200,N_27005,N_27086);
or U27201 (N_27201,N_27154,N_27021);
nor U27202 (N_27202,N_27111,N_27167);
xor U27203 (N_27203,N_27183,N_27031);
nor U27204 (N_27204,N_27185,N_27126);
nand U27205 (N_27205,N_27008,N_27056);
and U27206 (N_27206,N_27013,N_27047);
xor U27207 (N_27207,N_27182,N_27015);
nor U27208 (N_27208,N_27035,N_27022);
xnor U27209 (N_27209,N_27194,N_27083);
xor U27210 (N_27210,N_27124,N_27119);
or U27211 (N_27211,N_27026,N_27190);
xnor U27212 (N_27212,N_27001,N_27188);
nor U27213 (N_27213,N_27040,N_27156);
nor U27214 (N_27214,N_27048,N_27072);
and U27215 (N_27215,N_27071,N_27191);
nor U27216 (N_27216,N_27087,N_27020);
and U27217 (N_27217,N_27069,N_27060);
or U27218 (N_27218,N_27046,N_27024);
nand U27219 (N_27219,N_27019,N_27145);
and U27220 (N_27220,N_27062,N_27142);
or U27221 (N_27221,N_27042,N_27067);
xnor U27222 (N_27222,N_27058,N_27192);
nand U27223 (N_27223,N_27039,N_27178);
and U27224 (N_27224,N_27011,N_27152);
or U27225 (N_27225,N_27118,N_27163);
nand U27226 (N_27226,N_27112,N_27187);
xnor U27227 (N_27227,N_27085,N_27121);
xnor U27228 (N_27228,N_27010,N_27164);
xor U27229 (N_27229,N_27106,N_27171);
or U27230 (N_27230,N_27168,N_27029);
xor U27231 (N_27231,N_27033,N_27144);
and U27232 (N_27232,N_27094,N_27081);
and U27233 (N_27233,N_27147,N_27198);
nand U27234 (N_27234,N_27051,N_27055);
xor U27235 (N_27235,N_27115,N_27009);
nor U27236 (N_27236,N_27180,N_27075);
nand U27237 (N_27237,N_27107,N_27063);
and U27238 (N_27238,N_27113,N_27120);
or U27239 (N_27239,N_27128,N_27123);
or U27240 (N_27240,N_27172,N_27109);
and U27241 (N_27241,N_27018,N_27125);
and U27242 (N_27242,N_27199,N_27030);
nand U27243 (N_27243,N_27016,N_27155);
xnor U27244 (N_27244,N_27002,N_27140);
and U27245 (N_27245,N_27004,N_27050);
nor U27246 (N_27246,N_27057,N_27197);
xor U27247 (N_27247,N_27027,N_27161);
or U27248 (N_27248,N_27138,N_27162);
xnor U27249 (N_27249,N_27149,N_27132);
or U27250 (N_27250,N_27127,N_27089);
and U27251 (N_27251,N_27041,N_27000);
nand U27252 (N_27252,N_27014,N_27099);
xnor U27253 (N_27253,N_27076,N_27017);
xor U27254 (N_27254,N_27160,N_27176);
xor U27255 (N_27255,N_27007,N_27100);
nor U27256 (N_27256,N_27059,N_27157);
nor U27257 (N_27257,N_27037,N_27146);
nand U27258 (N_27258,N_27065,N_27052);
nand U27259 (N_27259,N_27032,N_27003);
nand U27260 (N_27260,N_27074,N_27139);
xor U27261 (N_27261,N_27064,N_27122);
xnor U27262 (N_27262,N_27023,N_27141);
and U27263 (N_27263,N_27151,N_27091);
or U27264 (N_27264,N_27102,N_27136);
nand U27265 (N_27265,N_27179,N_27038);
or U27266 (N_27266,N_27073,N_27165);
nor U27267 (N_27267,N_27070,N_27130);
nand U27268 (N_27268,N_27043,N_27170);
and U27269 (N_27269,N_27097,N_27082);
and U27270 (N_27270,N_27061,N_27135);
or U27271 (N_27271,N_27159,N_27079);
nand U27272 (N_27272,N_27054,N_27080);
xnor U27273 (N_27273,N_27095,N_27034);
nand U27274 (N_27274,N_27093,N_27193);
xnor U27275 (N_27275,N_27196,N_27066);
or U27276 (N_27276,N_27186,N_27114);
nor U27277 (N_27277,N_27006,N_27150);
nor U27278 (N_27278,N_27090,N_27134);
and U27279 (N_27279,N_27104,N_27110);
nand U27280 (N_27280,N_27049,N_27133);
xor U27281 (N_27281,N_27174,N_27195);
nor U27282 (N_27282,N_27158,N_27131);
or U27283 (N_27283,N_27096,N_27153);
and U27284 (N_27284,N_27053,N_27084);
xnor U27285 (N_27285,N_27044,N_27088);
nand U27286 (N_27286,N_27103,N_27078);
nand U27287 (N_27287,N_27173,N_27184);
xnor U27288 (N_27288,N_27068,N_27025);
or U27289 (N_27289,N_27148,N_27166);
nand U27290 (N_27290,N_27137,N_27177);
xnor U27291 (N_27291,N_27116,N_27028);
nor U27292 (N_27292,N_27092,N_27098);
and U27293 (N_27293,N_27045,N_27189);
xor U27294 (N_27294,N_27105,N_27012);
nand U27295 (N_27295,N_27117,N_27181);
xor U27296 (N_27296,N_27129,N_27101);
nor U27297 (N_27297,N_27169,N_27036);
or U27298 (N_27298,N_27143,N_27077);
nand U27299 (N_27299,N_27108,N_27175);
and U27300 (N_27300,N_27022,N_27004);
and U27301 (N_27301,N_27103,N_27066);
xnor U27302 (N_27302,N_27058,N_27074);
or U27303 (N_27303,N_27118,N_27151);
nor U27304 (N_27304,N_27162,N_27059);
and U27305 (N_27305,N_27115,N_27107);
or U27306 (N_27306,N_27186,N_27182);
nand U27307 (N_27307,N_27157,N_27181);
xor U27308 (N_27308,N_27093,N_27074);
and U27309 (N_27309,N_27156,N_27132);
or U27310 (N_27310,N_27174,N_27012);
or U27311 (N_27311,N_27002,N_27078);
or U27312 (N_27312,N_27157,N_27061);
nand U27313 (N_27313,N_27180,N_27099);
and U27314 (N_27314,N_27182,N_27157);
or U27315 (N_27315,N_27109,N_27094);
nor U27316 (N_27316,N_27012,N_27146);
xnor U27317 (N_27317,N_27114,N_27094);
nor U27318 (N_27318,N_27137,N_27053);
xnor U27319 (N_27319,N_27119,N_27055);
and U27320 (N_27320,N_27136,N_27035);
nand U27321 (N_27321,N_27150,N_27184);
xor U27322 (N_27322,N_27040,N_27006);
nor U27323 (N_27323,N_27087,N_27048);
xnor U27324 (N_27324,N_27179,N_27186);
nand U27325 (N_27325,N_27196,N_27199);
and U27326 (N_27326,N_27008,N_27117);
and U27327 (N_27327,N_27197,N_27039);
nor U27328 (N_27328,N_27130,N_27188);
or U27329 (N_27329,N_27117,N_27184);
or U27330 (N_27330,N_27192,N_27160);
or U27331 (N_27331,N_27141,N_27177);
and U27332 (N_27332,N_27183,N_27018);
nand U27333 (N_27333,N_27012,N_27091);
or U27334 (N_27334,N_27115,N_27046);
or U27335 (N_27335,N_27108,N_27069);
nand U27336 (N_27336,N_27136,N_27148);
nor U27337 (N_27337,N_27148,N_27142);
and U27338 (N_27338,N_27190,N_27063);
nor U27339 (N_27339,N_27029,N_27161);
nand U27340 (N_27340,N_27000,N_27019);
xor U27341 (N_27341,N_27130,N_27002);
nor U27342 (N_27342,N_27021,N_27137);
nor U27343 (N_27343,N_27047,N_27152);
nand U27344 (N_27344,N_27005,N_27002);
nor U27345 (N_27345,N_27182,N_27009);
and U27346 (N_27346,N_27066,N_27085);
nor U27347 (N_27347,N_27132,N_27102);
xnor U27348 (N_27348,N_27057,N_27048);
nand U27349 (N_27349,N_27172,N_27167);
xor U27350 (N_27350,N_27128,N_27097);
nor U27351 (N_27351,N_27007,N_27098);
nor U27352 (N_27352,N_27000,N_27009);
nand U27353 (N_27353,N_27022,N_27008);
nand U27354 (N_27354,N_27147,N_27003);
or U27355 (N_27355,N_27113,N_27063);
and U27356 (N_27356,N_27138,N_27160);
and U27357 (N_27357,N_27157,N_27197);
xnor U27358 (N_27358,N_27171,N_27078);
nor U27359 (N_27359,N_27006,N_27005);
xor U27360 (N_27360,N_27085,N_27124);
nand U27361 (N_27361,N_27118,N_27080);
or U27362 (N_27362,N_27063,N_27081);
or U27363 (N_27363,N_27066,N_27003);
nand U27364 (N_27364,N_27031,N_27155);
and U27365 (N_27365,N_27125,N_27025);
nand U27366 (N_27366,N_27154,N_27167);
xor U27367 (N_27367,N_27042,N_27009);
or U27368 (N_27368,N_27088,N_27042);
xnor U27369 (N_27369,N_27142,N_27057);
and U27370 (N_27370,N_27136,N_27163);
or U27371 (N_27371,N_27010,N_27029);
nor U27372 (N_27372,N_27153,N_27009);
or U27373 (N_27373,N_27135,N_27018);
or U27374 (N_27374,N_27021,N_27155);
and U27375 (N_27375,N_27198,N_27177);
or U27376 (N_27376,N_27076,N_27109);
and U27377 (N_27377,N_27082,N_27068);
or U27378 (N_27378,N_27137,N_27126);
nand U27379 (N_27379,N_27039,N_27087);
nor U27380 (N_27380,N_27182,N_27010);
and U27381 (N_27381,N_27087,N_27138);
or U27382 (N_27382,N_27053,N_27155);
nand U27383 (N_27383,N_27102,N_27040);
nor U27384 (N_27384,N_27161,N_27013);
nor U27385 (N_27385,N_27161,N_27160);
or U27386 (N_27386,N_27000,N_27109);
or U27387 (N_27387,N_27118,N_27189);
xor U27388 (N_27388,N_27098,N_27135);
or U27389 (N_27389,N_27066,N_27142);
nor U27390 (N_27390,N_27187,N_27014);
or U27391 (N_27391,N_27162,N_27030);
nand U27392 (N_27392,N_27123,N_27127);
and U27393 (N_27393,N_27163,N_27063);
and U27394 (N_27394,N_27179,N_27141);
xnor U27395 (N_27395,N_27123,N_27118);
and U27396 (N_27396,N_27148,N_27186);
nand U27397 (N_27397,N_27189,N_27181);
and U27398 (N_27398,N_27164,N_27133);
and U27399 (N_27399,N_27183,N_27101);
nor U27400 (N_27400,N_27283,N_27241);
or U27401 (N_27401,N_27232,N_27338);
and U27402 (N_27402,N_27367,N_27388);
nor U27403 (N_27403,N_27380,N_27213);
and U27404 (N_27404,N_27206,N_27219);
xor U27405 (N_27405,N_27242,N_27278);
xnor U27406 (N_27406,N_27256,N_27217);
xor U27407 (N_27407,N_27296,N_27318);
xor U27408 (N_27408,N_27287,N_27246);
xor U27409 (N_27409,N_27393,N_27286);
nor U27410 (N_27410,N_27260,N_27204);
or U27411 (N_27411,N_27366,N_27381);
nand U27412 (N_27412,N_27284,N_27292);
xnor U27413 (N_27413,N_27325,N_27382);
nor U27414 (N_27414,N_27220,N_27319);
and U27415 (N_27415,N_27379,N_27300);
nand U27416 (N_27416,N_27384,N_27394);
xor U27417 (N_27417,N_27279,N_27351);
nor U27418 (N_27418,N_27348,N_27343);
and U27419 (N_27419,N_27224,N_27275);
nor U27420 (N_27420,N_27259,N_27329);
or U27421 (N_27421,N_27211,N_27373);
or U27422 (N_27422,N_27282,N_27293);
xnor U27423 (N_27423,N_27386,N_27316);
nand U27424 (N_27424,N_27214,N_27363);
nand U27425 (N_27425,N_27266,N_27268);
nor U27426 (N_27426,N_27238,N_27299);
or U27427 (N_27427,N_27378,N_27265);
or U27428 (N_27428,N_27371,N_27372);
or U27429 (N_27429,N_27294,N_27333);
nand U27430 (N_27430,N_27236,N_27234);
and U27431 (N_27431,N_27389,N_27280);
nand U27432 (N_27432,N_27304,N_27326);
xnor U27433 (N_27433,N_27233,N_27344);
nor U27434 (N_27434,N_27311,N_27269);
and U27435 (N_27435,N_27322,N_27362);
nor U27436 (N_27436,N_27355,N_27261);
xor U27437 (N_27437,N_27387,N_27200);
and U27438 (N_27438,N_27276,N_27359);
nor U27439 (N_27439,N_27302,N_27267);
nand U27440 (N_27440,N_27291,N_27334);
nor U27441 (N_27441,N_27315,N_27353);
or U27442 (N_27442,N_27277,N_27215);
nor U27443 (N_27443,N_27222,N_27207);
and U27444 (N_27444,N_27339,N_27397);
or U27445 (N_27445,N_27229,N_27263);
or U27446 (N_27446,N_27203,N_27376);
or U27447 (N_27447,N_27210,N_27347);
or U27448 (N_27448,N_27264,N_27385);
nor U27449 (N_27449,N_27288,N_27226);
and U27450 (N_27450,N_27370,N_27395);
nand U27451 (N_27451,N_27336,N_27352);
nor U27452 (N_27452,N_27324,N_27340);
and U27453 (N_27453,N_27231,N_27240);
xnor U27454 (N_27454,N_27391,N_27361);
nand U27455 (N_27455,N_27308,N_27377);
nand U27456 (N_27456,N_27349,N_27369);
or U27457 (N_27457,N_27321,N_27335);
or U27458 (N_27458,N_27228,N_27201);
nand U27459 (N_27459,N_27356,N_27342);
nor U27460 (N_27460,N_27332,N_27247);
nand U27461 (N_27461,N_27255,N_27257);
and U27462 (N_27462,N_27297,N_27237);
or U27463 (N_27463,N_27274,N_27360);
and U27464 (N_27464,N_27227,N_27244);
xnor U27465 (N_27465,N_27248,N_27230);
nor U27466 (N_27466,N_27272,N_27253);
xor U27467 (N_27467,N_27309,N_27375);
and U27468 (N_27468,N_27209,N_27350);
nor U27469 (N_27469,N_27354,N_27305);
and U27470 (N_27470,N_27271,N_27368);
nand U27471 (N_27471,N_27320,N_27298);
nor U27472 (N_27472,N_27235,N_27313);
nand U27473 (N_27473,N_27251,N_27258);
nor U27474 (N_27474,N_27374,N_27383);
xnor U27475 (N_27475,N_27317,N_27285);
nor U27476 (N_27476,N_27323,N_27398);
or U27477 (N_27477,N_27212,N_27327);
xnor U27478 (N_27478,N_27307,N_27289);
nand U27479 (N_27479,N_27341,N_27358);
or U27480 (N_27480,N_27290,N_27310);
and U27481 (N_27481,N_27396,N_27202);
xor U27482 (N_27482,N_27314,N_27364);
xnor U27483 (N_27483,N_27223,N_27250);
xor U27484 (N_27484,N_27270,N_27249);
xnor U27485 (N_27485,N_27221,N_27254);
or U27486 (N_27486,N_27243,N_27239);
xor U27487 (N_27487,N_27301,N_27218);
and U27488 (N_27488,N_27357,N_27216);
or U27489 (N_27489,N_27295,N_27328);
and U27490 (N_27490,N_27205,N_27281);
nor U27491 (N_27491,N_27337,N_27330);
and U27492 (N_27492,N_27306,N_27245);
nand U27493 (N_27493,N_27345,N_27225);
xnor U27494 (N_27494,N_27392,N_27399);
xor U27495 (N_27495,N_27208,N_27252);
nor U27496 (N_27496,N_27303,N_27390);
nor U27497 (N_27497,N_27262,N_27365);
or U27498 (N_27498,N_27346,N_27331);
nor U27499 (N_27499,N_27273,N_27312);
nand U27500 (N_27500,N_27257,N_27277);
or U27501 (N_27501,N_27306,N_27375);
and U27502 (N_27502,N_27376,N_27270);
or U27503 (N_27503,N_27394,N_27374);
xnor U27504 (N_27504,N_27282,N_27275);
or U27505 (N_27505,N_27248,N_27372);
nor U27506 (N_27506,N_27279,N_27326);
nand U27507 (N_27507,N_27209,N_27274);
and U27508 (N_27508,N_27306,N_27244);
nand U27509 (N_27509,N_27358,N_27310);
or U27510 (N_27510,N_27341,N_27290);
nand U27511 (N_27511,N_27348,N_27269);
nor U27512 (N_27512,N_27244,N_27398);
and U27513 (N_27513,N_27396,N_27316);
nand U27514 (N_27514,N_27315,N_27344);
nand U27515 (N_27515,N_27230,N_27266);
and U27516 (N_27516,N_27364,N_27274);
nand U27517 (N_27517,N_27361,N_27324);
nand U27518 (N_27518,N_27236,N_27273);
and U27519 (N_27519,N_27293,N_27241);
and U27520 (N_27520,N_27391,N_27235);
nand U27521 (N_27521,N_27234,N_27349);
nand U27522 (N_27522,N_27324,N_27280);
or U27523 (N_27523,N_27227,N_27374);
nor U27524 (N_27524,N_27256,N_27238);
nor U27525 (N_27525,N_27323,N_27294);
or U27526 (N_27526,N_27364,N_27362);
xor U27527 (N_27527,N_27285,N_27379);
nand U27528 (N_27528,N_27266,N_27387);
and U27529 (N_27529,N_27280,N_27217);
nand U27530 (N_27530,N_27349,N_27215);
or U27531 (N_27531,N_27243,N_27333);
or U27532 (N_27532,N_27220,N_27248);
and U27533 (N_27533,N_27342,N_27308);
or U27534 (N_27534,N_27275,N_27287);
and U27535 (N_27535,N_27205,N_27261);
and U27536 (N_27536,N_27232,N_27213);
or U27537 (N_27537,N_27333,N_27210);
xor U27538 (N_27538,N_27313,N_27209);
xor U27539 (N_27539,N_27359,N_27221);
and U27540 (N_27540,N_27223,N_27210);
nor U27541 (N_27541,N_27393,N_27340);
nand U27542 (N_27542,N_27391,N_27334);
nand U27543 (N_27543,N_27311,N_27234);
nand U27544 (N_27544,N_27359,N_27390);
nor U27545 (N_27545,N_27244,N_27368);
or U27546 (N_27546,N_27268,N_27322);
nor U27547 (N_27547,N_27227,N_27294);
and U27548 (N_27548,N_27377,N_27260);
nand U27549 (N_27549,N_27339,N_27241);
nor U27550 (N_27550,N_27386,N_27207);
nor U27551 (N_27551,N_27274,N_27220);
nand U27552 (N_27552,N_27341,N_27376);
nand U27553 (N_27553,N_27346,N_27382);
nand U27554 (N_27554,N_27314,N_27272);
nor U27555 (N_27555,N_27210,N_27280);
xnor U27556 (N_27556,N_27210,N_27393);
and U27557 (N_27557,N_27292,N_27271);
xor U27558 (N_27558,N_27277,N_27332);
xor U27559 (N_27559,N_27279,N_27265);
nor U27560 (N_27560,N_27398,N_27222);
or U27561 (N_27561,N_27380,N_27360);
xor U27562 (N_27562,N_27311,N_27397);
nor U27563 (N_27563,N_27340,N_27334);
or U27564 (N_27564,N_27217,N_27380);
nor U27565 (N_27565,N_27255,N_27326);
nor U27566 (N_27566,N_27377,N_27252);
or U27567 (N_27567,N_27200,N_27201);
xnor U27568 (N_27568,N_27271,N_27321);
nor U27569 (N_27569,N_27229,N_27280);
nand U27570 (N_27570,N_27224,N_27360);
or U27571 (N_27571,N_27267,N_27276);
xnor U27572 (N_27572,N_27323,N_27272);
nand U27573 (N_27573,N_27380,N_27349);
nand U27574 (N_27574,N_27212,N_27233);
nand U27575 (N_27575,N_27345,N_27390);
nor U27576 (N_27576,N_27386,N_27378);
xor U27577 (N_27577,N_27269,N_27389);
nor U27578 (N_27578,N_27354,N_27376);
and U27579 (N_27579,N_27296,N_27389);
nand U27580 (N_27580,N_27363,N_27332);
nand U27581 (N_27581,N_27226,N_27304);
nor U27582 (N_27582,N_27207,N_27349);
and U27583 (N_27583,N_27371,N_27360);
nor U27584 (N_27584,N_27314,N_27294);
nand U27585 (N_27585,N_27230,N_27269);
nor U27586 (N_27586,N_27354,N_27364);
nand U27587 (N_27587,N_27373,N_27213);
or U27588 (N_27588,N_27317,N_27313);
xor U27589 (N_27589,N_27205,N_27243);
and U27590 (N_27590,N_27293,N_27307);
xnor U27591 (N_27591,N_27355,N_27286);
xnor U27592 (N_27592,N_27212,N_27364);
nor U27593 (N_27593,N_27286,N_27232);
nand U27594 (N_27594,N_27388,N_27230);
xnor U27595 (N_27595,N_27292,N_27253);
xnor U27596 (N_27596,N_27301,N_27374);
nand U27597 (N_27597,N_27367,N_27257);
xnor U27598 (N_27598,N_27333,N_27332);
xnor U27599 (N_27599,N_27387,N_27207);
xnor U27600 (N_27600,N_27499,N_27497);
xnor U27601 (N_27601,N_27508,N_27567);
and U27602 (N_27602,N_27477,N_27498);
and U27603 (N_27603,N_27436,N_27560);
xnor U27604 (N_27604,N_27543,N_27413);
nor U27605 (N_27605,N_27506,N_27561);
nor U27606 (N_27606,N_27553,N_27580);
nand U27607 (N_27607,N_27406,N_27472);
xor U27608 (N_27608,N_27599,N_27407);
nor U27609 (N_27609,N_27539,N_27434);
and U27610 (N_27610,N_27473,N_27431);
xor U27611 (N_27611,N_27405,N_27519);
nand U27612 (N_27612,N_27520,N_27596);
nand U27613 (N_27613,N_27556,N_27452);
or U27614 (N_27614,N_27540,N_27428);
xor U27615 (N_27615,N_27448,N_27447);
and U27616 (N_27616,N_27418,N_27583);
nor U27617 (N_27617,N_27491,N_27569);
and U27618 (N_27618,N_27527,N_27455);
nand U27619 (N_27619,N_27588,N_27492);
xor U27620 (N_27620,N_27458,N_27410);
nand U27621 (N_27621,N_27423,N_27579);
nor U27622 (N_27622,N_27409,N_27421);
or U27623 (N_27623,N_27595,N_27453);
or U27624 (N_27624,N_27403,N_27594);
nand U27625 (N_27625,N_27451,N_27441);
nor U27626 (N_27626,N_27416,N_27521);
nand U27627 (N_27627,N_27442,N_27440);
and U27628 (N_27628,N_27568,N_27545);
and U27629 (N_27629,N_27470,N_27511);
xnor U27630 (N_27630,N_27577,N_27534);
nand U27631 (N_27631,N_27515,N_27429);
nor U27632 (N_27632,N_27538,N_27495);
nor U27633 (N_27633,N_27463,N_27524);
nand U27634 (N_27634,N_27526,N_27541);
xor U27635 (N_27635,N_27479,N_27544);
and U27636 (N_27636,N_27536,N_27454);
nand U27637 (N_27637,N_27435,N_27562);
xnor U27638 (N_27638,N_27411,N_27427);
nand U27639 (N_27639,N_27507,N_27550);
nor U27640 (N_27640,N_27547,N_27500);
xnor U27641 (N_27641,N_27563,N_27484);
xor U27642 (N_27642,N_27485,N_27419);
nor U27643 (N_27643,N_27528,N_27462);
and U27644 (N_27644,N_27433,N_27518);
nand U27645 (N_27645,N_27586,N_27505);
or U27646 (N_27646,N_27408,N_27587);
xnor U27647 (N_27647,N_27558,N_27465);
nor U27648 (N_27648,N_27486,N_27517);
nand U27649 (N_27649,N_27482,N_27461);
nor U27650 (N_27650,N_27552,N_27555);
or U27651 (N_27651,N_27483,N_27474);
and U27652 (N_27652,N_27570,N_27457);
nor U27653 (N_27653,N_27529,N_27464);
or U27654 (N_27654,N_27468,N_27597);
and U27655 (N_27655,N_27488,N_27523);
nand U27656 (N_27656,N_27459,N_27489);
nand U27657 (N_27657,N_27422,N_27456);
or U27658 (N_27658,N_27578,N_27509);
nor U27659 (N_27659,N_27559,N_27471);
or U27660 (N_27660,N_27557,N_27549);
or U27661 (N_27661,N_27490,N_27487);
xnor U27662 (N_27662,N_27576,N_27513);
or U27663 (N_27663,N_27525,N_27400);
nand U27664 (N_27664,N_27478,N_27445);
nor U27665 (N_27665,N_27530,N_27466);
nand U27666 (N_27666,N_27446,N_27574);
and U27667 (N_27667,N_27516,N_27546);
nor U27668 (N_27668,N_27494,N_27598);
nand U27669 (N_27669,N_27417,N_27554);
nand U27670 (N_27670,N_27591,N_27480);
nor U27671 (N_27671,N_27532,N_27512);
or U27672 (N_27672,N_27493,N_27582);
and U27673 (N_27673,N_27592,N_27589);
nor U27674 (N_27674,N_27438,N_27402);
or U27675 (N_27675,N_27533,N_27496);
xor U27676 (N_27676,N_27432,N_27430);
or U27677 (N_27677,N_27412,N_27425);
nand U27678 (N_27678,N_27449,N_27575);
nor U27679 (N_27679,N_27503,N_27572);
and U27680 (N_27680,N_27537,N_27510);
or U27681 (N_27681,N_27450,N_27565);
nand U27682 (N_27682,N_27460,N_27593);
nor U27683 (N_27683,N_27585,N_27522);
and U27684 (N_27684,N_27426,N_27481);
nor U27685 (N_27685,N_27584,N_27548);
nand U27686 (N_27686,N_27551,N_27571);
and U27687 (N_27687,N_27476,N_27564);
xor U27688 (N_27688,N_27469,N_27531);
xnor U27689 (N_27689,N_27414,N_27514);
nor U27690 (N_27690,N_27535,N_27401);
xor U27691 (N_27691,N_27504,N_27467);
and U27692 (N_27692,N_27420,N_27444);
nand U27693 (N_27693,N_27475,N_27566);
or U27694 (N_27694,N_27443,N_27501);
nand U27695 (N_27695,N_27542,N_27573);
xor U27696 (N_27696,N_27404,N_27439);
nor U27697 (N_27697,N_27415,N_27424);
xor U27698 (N_27698,N_27437,N_27590);
nor U27699 (N_27699,N_27581,N_27502);
xor U27700 (N_27700,N_27513,N_27477);
xor U27701 (N_27701,N_27500,N_27574);
or U27702 (N_27702,N_27572,N_27588);
nor U27703 (N_27703,N_27437,N_27561);
xor U27704 (N_27704,N_27528,N_27472);
nand U27705 (N_27705,N_27542,N_27591);
nor U27706 (N_27706,N_27498,N_27402);
and U27707 (N_27707,N_27475,N_27528);
xor U27708 (N_27708,N_27519,N_27531);
and U27709 (N_27709,N_27508,N_27549);
nor U27710 (N_27710,N_27552,N_27444);
and U27711 (N_27711,N_27465,N_27575);
or U27712 (N_27712,N_27590,N_27436);
xnor U27713 (N_27713,N_27416,N_27431);
and U27714 (N_27714,N_27410,N_27580);
or U27715 (N_27715,N_27415,N_27454);
xnor U27716 (N_27716,N_27448,N_27464);
xnor U27717 (N_27717,N_27446,N_27461);
nand U27718 (N_27718,N_27518,N_27444);
xnor U27719 (N_27719,N_27523,N_27408);
nor U27720 (N_27720,N_27459,N_27475);
nand U27721 (N_27721,N_27475,N_27584);
nor U27722 (N_27722,N_27409,N_27407);
nand U27723 (N_27723,N_27553,N_27597);
and U27724 (N_27724,N_27416,N_27478);
nor U27725 (N_27725,N_27545,N_27493);
nand U27726 (N_27726,N_27462,N_27406);
xor U27727 (N_27727,N_27511,N_27566);
and U27728 (N_27728,N_27559,N_27424);
nor U27729 (N_27729,N_27592,N_27596);
and U27730 (N_27730,N_27529,N_27504);
and U27731 (N_27731,N_27543,N_27492);
nor U27732 (N_27732,N_27459,N_27425);
nor U27733 (N_27733,N_27413,N_27455);
nand U27734 (N_27734,N_27566,N_27407);
and U27735 (N_27735,N_27524,N_27428);
and U27736 (N_27736,N_27438,N_27566);
nor U27737 (N_27737,N_27479,N_27429);
or U27738 (N_27738,N_27590,N_27448);
or U27739 (N_27739,N_27552,N_27460);
and U27740 (N_27740,N_27459,N_27473);
xnor U27741 (N_27741,N_27418,N_27560);
nor U27742 (N_27742,N_27442,N_27475);
nor U27743 (N_27743,N_27437,N_27410);
or U27744 (N_27744,N_27448,N_27488);
xnor U27745 (N_27745,N_27497,N_27564);
and U27746 (N_27746,N_27485,N_27458);
and U27747 (N_27747,N_27537,N_27444);
xnor U27748 (N_27748,N_27505,N_27483);
and U27749 (N_27749,N_27461,N_27549);
nor U27750 (N_27750,N_27436,N_27412);
and U27751 (N_27751,N_27400,N_27452);
and U27752 (N_27752,N_27590,N_27446);
xor U27753 (N_27753,N_27574,N_27428);
xor U27754 (N_27754,N_27575,N_27526);
xnor U27755 (N_27755,N_27527,N_27428);
and U27756 (N_27756,N_27522,N_27491);
or U27757 (N_27757,N_27505,N_27420);
or U27758 (N_27758,N_27458,N_27571);
xnor U27759 (N_27759,N_27426,N_27493);
xnor U27760 (N_27760,N_27532,N_27475);
xnor U27761 (N_27761,N_27574,N_27523);
nand U27762 (N_27762,N_27472,N_27544);
or U27763 (N_27763,N_27543,N_27572);
or U27764 (N_27764,N_27441,N_27590);
xnor U27765 (N_27765,N_27544,N_27422);
and U27766 (N_27766,N_27524,N_27430);
or U27767 (N_27767,N_27510,N_27593);
and U27768 (N_27768,N_27515,N_27432);
nor U27769 (N_27769,N_27593,N_27555);
and U27770 (N_27770,N_27589,N_27498);
nor U27771 (N_27771,N_27471,N_27476);
and U27772 (N_27772,N_27541,N_27584);
nand U27773 (N_27773,N_27454,N_27519);
and U27774 (N_27774,N_27530,N_27501);
nor U27775 (N_27775,N_27483,N_27518);
xor U27776 (N_27776,N_27541,N_27463);
or U27777 (N_27777,N_27515,N_27542);
nand U27778 (N_27778,N_27554,N_27460);
nand U27779 (N_27779,N_27549,N_27472);
xnor U27780 (N_27780,N_27440,N_27530);
nand U27781 (N_27781,N_27461,N_27586);
xnor U27782 (N_27782,N_27463,N_27455);
nand U27783 (N_27783,N_27534,N_27581);
nand U27784 (N_27784,N_27445,N_27409);
nand U27785 (N_27785,N_27477,N_27570);
and U27786 (N_27786,N_27488,N_27588);
nor U27787 (N_27787,N_27450,N_27417);
and U27788 (N_27788,N_27596,N_27544);
and U27789 (N_27789,N_27484,N_27568);
nand U27790 (N_27790,N_27547,N_27478);
and U27791 (N_27791,N_27480,N_27541);
and U27792 (N_27792,N_27565,N_27558);
and U27793 (N_27793,N_27429,N_27448);
or U27794 (N_27794,N_27578,N_27515);
nor U27795 (N_27795,N_27517,N_27574);
nor U27796 (N_27796,N_27508,N_27412);
nor U27797 (N_27797,N_27540,N_27464);
or U27798 (N_27798,N_27423,N_27431);
or U27799 (N_27799,N_27419,N_27544);
and U27800 (N_27800,N_27661,N_27691);
or U27801 (N_27801,N_27767,N_27774);
nand U27802 (N_27802,N_27778,N_27716);
or U27803 (N_27803,N_27792,N_27710);
or U27804 (N_27804,N_27646,N_27742);
nor U27805 (N_27805,N_27754,N_27623);
nand U27806 (N_27806,N_27731,N_27604);
xor U27807 (N_27807,N_27748,N_27768);
nor U27808 (N_27808,N_27746,N_27682);
nand U27809 (N_27809,N_27672,N_27795);
nor U27810 (N_27810,N_27684,N_27689);
or U27811 (N_27811,N_27735,N_27685);
and U27812 (N_27812,N_27680,N_27793);
xnor U27813 (N_27813,N_27694,N_27780);
or U27814 (N_27814,N_27616,N_27743);
xor U27815 (N_27815,N_27787,N_27621);
or U27816 (N_27816,N_27772,N_27690);
and U27817 (N_27817,N_27622,N_27679);
and U27818 (N_27818,N_27618,N_27688);
xor U27819 (N_27819,N_27643,N_27744);
and U27820 (N_27820,N_27711,N_27714);
nand U27821 (N_27821,N_27655,N_27627);
xnor U27822 (N_27822,N_27602,N_27794);
nor U27823 (N_27823,N_27662,N_27739);
nand U27824 (N_27824,N_27649,N_27770);
nor U27825 (N_27825,N_27712,N_27611);
or U27826 (N_27826,N_27750,N_27784);
nand U27827 (N_27827,N_27773,N_27632);
nor U27828 (N_27828,N_27757,N_27600);
and U27829 (N_27829,N_27628,N_27747);
and U27830 (N_27830,N_27771,N_27633);
xnor U27831 (N_27831,N_27670,N_27658);
nor U27832 (N_27832,N_27620,N_27706);
nor U27833 (N_27833,N_27657,N_27740);
nor U27834 (N_27834,N_27652,N_27610);
nor U27835 (N_27835,N_27749,N_27631);
and U27836 (N_27836,N_27665,N_27736);
nand U27837 (N_27837,N_27613,N_27675);
and U27838 (N_27838,N_27727,N_27785);
or U27839 (N_27839,N_27713,N_27733);
nand U27840 (N_27840,N_27634,N_27698);
nor U27841 (N_27841,N_27734,N_27777);
and U27842 (N_27842,N_27697,N_27723);
nor U27843 (N_27843,N_27776,N_27607);
nand U27844 (N_27844,N_27717,N_27701);
and U27845 (N_27845,N_27700,N_27637);
nand U27846 (N_27846,N_27756,N_27696);
and U27847 (N_27847,N_27606,N_27603);
and U27848 (N_27848,N_27615,N_27671);
nand U27849 (N_27849,N_27751,N_27763);
nand U27850 (N_27850,N_27720,N_27612);
nand U27851 (N_27851,N_27715,N_27630);
nor U27852 (N_27852,N_27692,N_27636);
nand U27853 (N_27853,N_27726,N_27703);
or U27854 (N_27854,N_27766,N_27617);
nor U27855 (N_27855,N_27686,N_27759);
nand U27856 (N_27856,N_27608,N_27660);
nor U27857 (N_27857,N_27728,N_27641);
and U27858 (N_27858,N_27656,N_27666);
and U27859 (N_27859,N_27659,N_27753);
nor U27860 (N_27860,N_27640,N_27765);
xor U27861 (N_27861,N_27722,N_27648);
or U27862 (N_27862,N_27769,N_27729);
and U27863 (N_27863,N_27695,N_27687);
or U27864 (N_27864,N_27642,N_27725);
or U27865 (N_27865,N_27762,N_27668);
xor U27866 (N_27866,N_27718,N_27654);
nand U27867 (N_27867,N_27745,N_27699);
nor U27868 (N_27868,N_27798,N_27626);
and U27869 (N_27869,N_27799,N_27709);
or U27870 (N_27870,N_27605,N_27779);
and U27871 (N_27871,N_27719,N_27781);
and U27872 (N_27872,N_27619,N_27789);
and U27873 (N_27873,N_27667,N_27644);
xnor U27874 (N_27874,N_27760,N_27758);
nand U27875 (N_27875,N_27796,N_27786);
or U27876 (N_27876,N_27741,N_27663);
or U27877 (N_27877,N_27707,N_27752);
nor U27878 (N_27878,N_27782,N_27678);
nand U27879 (N_27879,N_27614,N_27635);
or U27880 (N_27880,N_27788,N_27764);
nand U27881 (N_27881,N_27704,N_27783);
nand U27882 (N_27882,N_27730,N_27693);
nand U27883 (N_27883,N_27677,N_27797);
xnor U27884 (N_27884,N_27647,N_27681);
nand U27885 (N_27885,N_27676,N_27653);
nand U27886 (N_27886,N_27683,N_27791);
and U27887 (N_27887,N_27702,N_27790);
nor U27888 (N_27888,N_27625,N_27639);
xor U27889 (N_27889,N_27624,N_27651);
or U27890 (N_27890,N_27738,N_27629);
xor U27891 (N_27891,N_27664,N_27673);
xnor U27892 (N_27892,N_27761,N_27732);
nand U27893 (N_27893,N_27737,N_27705);
or U27894 (N_27894,N_27674,N_27638);
xnor U27895 (N_27895,N_27721,N_27669);
nor U27896 (N_27896,N_27708,N_27650);
or U27897 (N_27897,N_27601,N_27755);
or U27898 (N_27898,N_27775,N_27724);
nor U27899 (N_27899,N_27609,N_27645);
nor U27900 (N_27900,N_27733,N_27693);
or U27901 (N_27901,N_27748,N_27756);
nand U27902 (N_27902,N_27790,N_27640);
xnor U27903 (N_27903,N_27712,N_27628);
and U27904 (N_27904,N_27677,N_27705);
nor U27905 (N_27905,N_27710,N_27782);
nand U27906 (N_27906,N_27670,N_27717);
nand U27907 (N_27907,N_27634,N_27799);
xnor U27908 (N_27908,N_27759,N_27657);
and U27909 (N_27909,N_27707,N_27631);
xnor U27910 (N_27910,N_27704,N_27651);
nand U27911 (N_27911,N_27789,N_27675);
or U27912 (N_27912,N_27737,N_27744);
or U27913 (N_27913,N_27799,N_27654);
nand U27914 (N_27914,N_27627,N_27635);
nand U27915 (N_27915,N_27756,N_27716);
or U27916 (N_27916,N_27619,N_27627);
xnor U27917 (N_27917,N_27645,N_27633);
and U27918 (N_27918,N_27751,N_27757);
nand U27919 (N_27919,N_27761,N_27707);
or U27920 (N_27920,N_27732,N_27788);
xor U27921 (N_27921,N_27658,N_27798);
xnor U27922 (N_27922,N_27606,N_27769);
nor U27923 (N_27923,N_27708,N_27712);
nor U27924 (N_27924,N_27787,N_27657);
xor U27925 (N_27925,N_27704,N_27770);
xor U27926 (N_27926,N_27615,N_27693);
nor U27927 (N_27927,N_27732,N_27638);
and U27928 (N_27928,N_27774,N_27795);
nor U27929 (N_27929,N_27730,N_27751);
nand U27930 (N_27930,N_27791,N_27799);
nand U27931 (N_27931,N_27766,N_27762);
nor U27932 (N_27932,N_27643,N_27651);
nor U27933 (N_27933,N_27643,N_27734);
and U27934 (N_27934,N_27774,N_27606);
nand U27935 (N_27935,N_27684,N_27657);
and U27936 (N_27936,N_27645,N_27739);
or U27937 (N_27937,N_27645,N_27744);
and U27938 (N_27938,N_27695,N_27655);
nor U27939 (N_27939,N_27679,N_27646);
nor U27940 (N_27940,N_27722,N_27612);
nand U27941 (N_27941,N_27787,N_27703);
or U27942 (N_27942,N_27712,N_27642);
nand U27943 (N_27943,N_27651,N_27698);
and U27944 (N_27944,N_27768,N_27786);
nor U27945 (N_27945,N_27656,N_27687);
or U27946 (N_27946,N_27638,N_27620);
nor U27947 (N_27947,N_27726,N_27741);
nand U27948 (N_27948,N_27724,N_27736);
or U27949 (N_27949,N_27731,N_27711);
or U27950 (N_27950,N_27623,N_27670);
nand U27951 (N_27951,N_27792,N_27653);
or U27952 (N_27952,N_27651,N_27731);
and U27953 (N_27953,N_27719,N_27647);
nand U27954 (N_27954,N_27711,N_27790);
or U27955 (N_27955,N_27664,N_27724);
or U27956 (N_27956,N_27696,N_27688);
nor U27957 (N_27957,N_27739,N_27791);
and U27958 (N_27958,N_27780,N_27603);
or U27959 (N_27959,N_27604,N_27634);
and U27960 (N_27960,N_27665,N_27715);
nor U27961 (N_27961,N_27647,N_27608);
nor U27962 (N_27962,N_27685,N_27792);
or U27963 (N_27963,N_27620,N_27690);
and U27964 (N_27964,N_27619,N_27702);
and U27965 (N_27965,N_27664,N_27726);
nor U27966 (N_27966,N_27606,N_27731);
nor U27967 (N_27967,N_27727,N_27775);
xor U27968 (N_27968,N_27712,N_27785);
and U27969 (N_27969,N_27702,N_27719);
and U27970 (N_27970,N_27650,N_27696);
and U27971 (N_27971,N_27760,N_27633);
and U27972 (N_27972,N_27743,N_27608);
or U27973 (N_27973,N_27753,N_27756);
or U27974 (N_27974,N_27759,N_27741);
nand U27975 (N_27975,N_27771,N_27787);
and U27976 (N_27976,N_27618,N_27748);
and U27977 (N_27977,N_27655,N_27700);
or U27978 (N_27978,N_27631,N_27712);
nor U27979 (N_27979,N_27744,N_27725);
nor U27980 (N_27980,N_27685,N_27704);
xnor U27981 (N_27981,N_27660,N_27754);
xnor U27982 (N_27982,N_27732,N_27735);
and U27983 (N_27983,N_27653,N_27709);
or U27984 (N_27984,N_27722,N_27773);
xnor U27985 (N_27985,N_27686,N_27623);
and U27986 (N_27986,N_27721,N_27674);
and U27987 (N_27987,N_27646,N_27608);
nor U27988 (N_27988,N_27718,N_27764);
nand U27989 (N_27989,N_27715,N_27645);
xor U27990 (N_27990,N_27780,N_27609);
and U27991 (N_27991,N_27689,N_27760);
nand U27992 (N_27992,N_27703,N_27729);
or U27993 (N_27993,N_27736,N_27650);
nand U27994 (N_27994,N_27729,N_27788);
xnor U27995 (N_27995,N_27678,N_27684);
nor U27996 (N_27996,N_27741,N_27779);
xor U27997 (N_27997,N_27687,N_27615);
or U27998 (N_27998,N_27790,N_27740);
nor U27999 (N_27999,N_27723,N_27799);
and U28000 (N_28000,N_27879,N_27918);
or U28001 (N_28001,N_27977,N_27835);
nand U28002 (N_28002,N_27899,N_27983);
xor U28003 (N_28003,N_27968,N_27829);
nor U28004 (N_28004,N_27851,N_27913);
or U28005 (N_28005,N_27874,N_27950);
or U28006 (N_28006,N_27807,N_27903);
xnor U28007 (N_28007,N_27854,N_27831);
and U28008 (N_28008,N_27900,N_27933);
nand U28009 (N_28009,N_27992,N_27883);
xnor U28010 (N_28010,N_27898,N_27914);
nand U28011 (N_28011,N_27974,N_27980);
nand U28012 (N_28012,N_27818,N_27975);
or U28013 (N_28013,N_27924,N_27940);
nand U28014 (N_28014,N_27902,N_27886);
nand U28015 (N_28015,N_27810,N_27931);
and U28016 (N_28016,N_27986,N_27912);
or U28017 (N_28017,N_27809,N_27866);
and U28018 (N_28018,N_27988,N_27859);
and U28019 (N_28019,N_27990,N_27885);
nand U28020 (N_28020,N_27826,N_27962);
and U28021 (N_28021,N_27836,N_27817);
nand U28022 (N_28022,N_27812,N_27932);
or U28023 (N_28023,N_27887,N_27845);
nor U28024 (N_28024,N_27981,N_27965);
and U28025 (N_28025,N_27890,N_27978);
or U28026 (N_28026,N_27844,N_27853);
xor U28027 (N_28027,N_27889,N_27856);
xnor U28028 (N_28028,N_27852,N_27953);
nor U28029 (N_28029,N_27848,N_27846);
and U28030 (N_28030,N_27919,N_27942);
nor U28031 (N_28031,N_27995,N_27934);
and U28032 (N_28032,N_27849,N_27880);
nand U28033 (N_28033,N_27909,N_27833);
nor U28034 (N_28034,N_27939,N_27935);
nor U28035 (N_28035,N_27927,N_27842);
xor U28036 (N_28036,N_27806,N_27905);
nand U28037 (N_28037,N_27923,N_27840);
nor U28038 (N_28038,N_27949,N_27930);
nand U28039 (N_28039,N_27827,N_27838);
nor U28040 (N_28040,N_27928,N_27922);
and U28041 (N_28041,N_27819,N_27999);
and U28042 (N_28042,N_27864,N_27982);
nand U28043 (N_28043,N_27834,N_27998);
nand U28044 (N_28044,N_27804,N_27989);
and U28045 (N_28045,N_27870,N_27910);
nand U28046 (N_28046,N_27901,N_27825);
nand U28047 (N_28047,N_27956,N_27882);
nand U28048 (N_28048,N_27997,N_27957);
and U28049 (N_28049,N_27802,N_27970);
nor U28050 (N_28050,N_27813,N_27821);
and U28051 (N_28051,N_27801,N_27803);
nand U28052 (N_28052,N_27987,N_27892);
xor U28053 (N_28053,N_27985,N_27960);
nor U28054 (N_28054,N_27943,N_27920);
and U28055 (N_28055,N_27959,N_27993);
xnor U28056 (N_28056,N_27839,N_27969);
or U28057 (N_28057,N_27863,N_27921);
xor U28058 (N_28058,N_27904,N_27830);
and U28059 (N_28059,N_27843,N_27808);
or U28060 (N_28060,N_27971,N_27929);
or U28061 (N_28061,N_27907,N_27891);
and U28062 (N_28062,N_27832,N_27966);
nand U28063 (N_28063,N_27868,N_27952);
nor U28064 (N_28064,N_27937,N_27822);
xor U28065 (N_28065,N_27936,N_27850);
or U28066 (N_28066,N_27915,N_27994);
or U28067 (N_28067,N_27893,N_27945);
nor U28068 (N_28068,N_27847,N_27955);
or U28069 (N_28069,N_27858,N_27961);
nor U28070 (N_28070,N_27973,N_27871);
or U28071 (N_28071,N_27823,N_27897);
nor U28072 (N_28072,N_27954,N_27861);
or U28073 (N_28073,N_27947,N_27869);
nor U28074 (N_28074,N_27878,N_27877);
xnor U28075 (N_28075,N_27805,N_27815);
nor U28076 (N_28076,N_27958,N_27925);
and U28077 (N_28077,N_27948,N_27991);
xor U28078 (N_28078,N_27916,N_27865);
or U28079 (N_28079,N_27814,N_27996);
or U28080 (N_28080,N_27875,N_27926);
and U28081 (N_28081,N_27896,N_27906);
nand U28082 (N_28082,N_27911,N_27976);
and U28083 (N_28083,N_27824,N_27938);
and U28084 (N_28084,N_27944,N_27855);
xnor U28085 (N_28085,N_27841,N_27837);
and U28086 (N_28086,N_27884,N_27967);
and U28087 (N_28087,N_27816,N_27964);
and U28088 (N_28088,N_27984,N_27895);
nand U28089 (N_28089,N_27820,N_27941);
nand U28090 (N_28090,N_27972,N_27881);
xnor U28091 (N_28091,N_27917,N_27862);
or U28092 (N_28092,N_27946,N_27888);
nor U28093 (N_28093,N_27894,N_27867);
or U28094 (N_28094,N_27908,N_27951);
or U28095 (N_28095,N_27860,N_27979);
nor U28096 (N_28096,N_27828,N_27811);
nor U28097 (N_28097,N_27963,N_27876);
nor U28098 (N_28098,N_27857,N_27873);
nand U28099 (N_28099,N_27872,N_27800);
nand U28100 (N_28100,N_27975,N_27990);
nand U28101 (N_28101,N_27839,N_27973);
nand U28102 (N_28102,N_27859,N_27914);
and U28103 (N_28103,N_27828,N_27966);
nand U28104 (N_28104,N_27890,N_27938);
or U28105 (N_28105,N_27837,N_27986);
or U28106 (N_28106,N_27967,N_27863);
nand U28107 (N_28107,N_27900,N_27864);
or U28108 (N_28108,N_27985,N_27872);
xnor U28109 (N_28109,N_27865,N_27927);
nor U28110 (N_28110,N_27872,N_27884);
and U28111 (N_28111,N_27990,N_27887);
or U28112 (N_28112,N_27851,N_27977);
or U28113 (N_28113,N_27958,N_27813);
nand U28114 (N_28114,N_27937,N_27883);
xor U28115 (N_28115,N_27926,N_27903);
or U28116 (N_28116,N_27977,N_27840);
or U28117 (N_28117,N_27880,N_27845);
nand U28118 (N_28118,N_27845,N_27825);
or U28119 (N_28119,N_27996,N_27884);
and U28120 (N_28120,N_27829,N_27987);
and U28121 (N_28121,N_27912,N_27958);
or U28122 (N_28122,N_27883,N_27976);
nand U28123 (N_28123,N_27805,N_27897);
xor U28124 (N_28124,N_27953,N_27956);
and U28125 (N_28125,N_27928,N_27858);
and U28126 (N_28126,N_27856,N_27903);
or U28127 (N_28127,N_27887,N_27927);
nand U28128 (N_28128,N_27948,N_27893);
and U28129 (N_28129,N_27877,N_27852);
nand U28130 (N_28130,N_27868,N_27824);
xnor U28131 (N_28131,N_27984,N_27947);
and U28132 (N_28132,N_27866,N_27980);
nor U28133 (N_28133,N_27978,N_27935);
xnor U28134 (N_28134,N_27943,N_27995);
xor U28135 (N_28135,N_27878,N_27801);
or U28136 (N_28136,N_27924,N_27979);
nor U28137 (N_28137,N_27840,N_27844);
xnor U28138 (N_28138,N_27944,N_27883);
xor U28139 (N_28139,N_27979,N_27926);
or U28140 (N_28140,N_27967,N_27800);
and U28141 (N_28141,N_27829,N_27818);
nor U28142 (N_28142,N_27865,N_27968);
or U28143 (N_28143,N_27957,N_27941);
or U28144 (N_28144,N_27873,N_27924);
xnor U28145 (N_28145,N_27956,N_27862);
xnor U28146 (N_28146,N_27886,N_27892);
nand U28147 (N_28147,N_27916,N_27978);
nand U28148 (N_28148,N_27863,N_27859);
xnor U28149 (N_28149,N_27882,N_27841);
xor U28150 (N_28150,N_27874,N_27803);
xor U28151 (N_28151,N_27999,N_27940);
xnor U28152 (N_28152,N_27874,N_27927);
and U28153 (N_28153,N_27876,N_27889);
or U28154 (N_28154,N_27809,N_27998);
nor U28155 (N_28155,N_27827,N_27966);
xor U28156 (N_28156,N_27801,N_27817);
or U28157 (N_28157,N_27844,N_27889);
or U28158 (N_28158,N_27860,N_27916);
and U28159 (N_28159,N_27956,N_27949);
and U28160 (N_28160,N_27903,N_27945);
and U28161 (N_28161,N_27844,N_27877);
or U28162 (N_28162,N_27836,N_27851);
nand U28163 (N_28163,N_27950,N_27940);
or U28164 (N_28164,N_27812,N_27854);
or U28165 (N_28165,N_27829,N_27888);
or U28166 (N_28166,N_27907,N_27910);
xor U28167 (N_28167,N_27978,N_27854);
nand U28168 (N_28168,N_27836,N_27959);
xor U28169 (N_28169,N_27950,N_27981);
nand U28170 (N_28170,N_27920,N_27862);
nand U28171 (N_28171,N_27989,N_27815);
and U28172 (N_28172,N_27995,N_27805);
or U28173 (N_28173,N_27883,N_27808);
and U28174 (N_28174,N_27915,N_27917);
and U28175 (N_28175,N_27962,N_27993);
or U28176 (N_28176,N_27835,N_27946);
nor U28177 (N_28177,N_27962,N_27903);
and U28178 (N_28178,N_27899,N_27975);
and U28179 (N_28179,N_27996,N_27861);
xnor U28180 (N_28180,N_27889,N_27833);
nand U28181 (N_28181,N_27849,N_27953);
and U28182 (N_28182,N_27989,N_27898);
xor U28183 (N_28183,N_27927,N_27895);
nor U28184 (N_28184,N_27922,N_27978);
xnor U28185 (N_28185,N_27852,N_27913);
xnor U28186 (N_28186,N_27813,N_27873);
nor U28187 (N_28187,N_27847,N_27863);
nand U28188 (N_28188,N_27906,N_27900);
nand U28189 (N_28189,N_27918,N_27835);
and U28190 (N_28190,N_27832,N_27843);
nor U28191 (N_28191,N_27825,N_27982);
or U28192 (N_28192,N_27857,N_27868);
nand U28193 (N_28193,N_27934,N_27937);
nand U28194 (N_28194,N_27996,N_27946);
xnor U28195 (N_28195,N_27998,N_27852);
or U28196 (N_28196,N_27981,N_27888);
nand U28197 (N_28197,N_27846,N_27833);
nand U28198 (N_28198,N_27924,N_27820);
and U28199 (N_28199,N_27853,N_27964);
nor U28200 (N_28200,N_28093,N_28095);
or U28201 (N_28201,N_28140,N_28187);
and U28202 (N_28202,N_28182,N_28133);
xor U28203 (N_28203,N_28045,N_28127);
xor U28204 (N_28204,N_28157,N_28101);
and U28205 (N_28205,N_28084,N_28022);
nand U28206 (N_28206,N_28145,N_28110);
and U28207 (N_28207,N_28158,N_28112);
nor U28208 (N_28208,N_28195,N_28180);
xnor U28209 (N_28209,N_28020,N_28085);
or U28210 (N_28210,N_28049,N_28164);
nor U28211 (N_28211,N_28094,N_28038);
xor U28212 (N_28212,N_28194,N_28011);
xor U28213 (N_28213,N_28114,N_28048);
xnor U28214 (N_28214,N_28014,N_28088);
nand U28215 (N_28215,N_28188,N_28021);
nor U28216 (N_28216,N_28016,N_28064);
nor U28217 (N_28217,N_28097,N_28081);
nor U28218 (N_28218,N_28120,N_28192);
nor U28219 (N_28219,N_28099,N_28154);
and U28220 (N_28220,N_28080,N_28092);
or U28221 (N_28221,N_28172,N_28159);
nand U28222 (N_28222,N_28148,N_28035);
nand U28223 (N_28223,N_28190,N_28034);
nor U28224 (N_28224,N_28000,N_28115);
xor U28225 (N_28225,N_28005,N_28065);
or U28226 (N_28226,N_28197,N_28130);
or U28227 (N_28227,N_28089,N_28044);
xor U28228 (N_28228,N_28067,N_28186);
xor U28229 (N_28229,N_28010,N_28036);
nand U28230 (N_28230,N_28123,N_28150);
or U28231 (N_28231,N_28052,N_28122);
or U28232 (N_28232,N_28050,N_28006);
and U28233 (N_28233,N_28073,N_28124);
or U28234 (N_28234,N_28129,N_28107);
nor U28235 (N_28235,N_28160,N_28071);
nand U28236 (N_28236,N_28030,N_28146);
nand U28237 (N_28237,N_28131,N_28165);
or U28238 (N_28238,N_28141,N_28032);
nor U28239 (N_28239,N_28104,N_28009);
nor U28240 (N_28240,N_28173,N_28075);
nor U28241 (N_28241,N_28024,N_28174);
and U28242 (N_28242,N_28139,N_28061);
nor U28243 (N_28243,N_28161,N_28128);
nand U28244 (N_28244,N_28198,N_28012);
nand U28245 (N_28245,N_28119,N_28117);
or U28246 (N_28246,N_28134,N_28070);
xnor U28247 (N_28247,N_28082,N_28111);
nand U28248 (N_28248,N_28175,N_28183);
or U28249 (N_28249,N_28166,N_28008);
nor U28250 (N_28250,N_28137,N_28057);
or U28251 (N_28251,N_28033,N_28185);
nand U28252 (N_28252,N_28152,N_28015);
nor U28253 (N_28253,N_28121,N_28037);
nand U28254 (N_28254,N_28191,N_28087);
or U28255 (N_28255,N_28149,N_28078);
or U28256 (N_28256,N_28076,N_28066);
and U28257 (N_28257,N_28068,N_28059);
and U28258 (N_28258,N_28125,N_28100);
nand U28259 (N_28259,N_28113,N_28156);
or U28260 (N_28260,N_28162,N_28151);
or U28261 (N_28261,N_28083,N_28102);
nand U28262 (N_28262,N_28108,N_28147);
nand U28263 (N_28263,N_28019,N_28105);
nand U28264 (N_28264,N_28039,N_28031);
or U28265 (N_28265,N_28136,N_28199);
or U28266 (N_28266,N_28060,N_28023);
nand U28267 (N_28267,N_28053,N_28002);
or U28268 (N_28268,N_28074,N_28153);
or U28269 (N_28269,N_28043,N_28013);
or U28270 (N_28270,N_28007,N_28062);
nand U28271 (N_28271,N_28069,N_28004);
or U28272 (N_28272,N_28106,N_28091);
xor U28273 (N_28273,N_28055,N_28118);
or U28274 (N_28274,N_28029,N_28193);
nor U28275 (N_28275,N_28063,N_28181);
nor U28276 (N_28276,N_28189,N_28135);
nor U28277 (N_28277,N_28026,N_28098);
xnor U28278 (N_28278,N_28058,N_28177);
nor U28279 (N_28279,N_28077,N_28178);
nand U28280 (N_28280,N_28126,N_28086);
or U28281 (N_28281,N_28116,N_28040);
or U28282 (N_28282,N_28167,N_28168);
xnor U28283 (N_28283,N_28003,N_28170);
or U28284 (N_28284,N_28001,N_28169);
or U28285 (N_28285,N_28176,N_28047);
nand U28286 (N_28286,N_28143,N_28142);
xor U28287 (N_28287,N_28171,N_28196);
nor U28288 (N_28288,N_28138,N_28051);
xnor U28289 (N_28289,N_28184,N_28072);
or U28290 (N_28290,N_28096,N_28090);
nor U28291 (N_28291,N_28079,N_28163);
and U28292 (N_28292,N_28017,N_28109);
or U28293 (N_28293,N_28042,N_28155);
or U28294 (N_28294,N_28132,N_28056);
nor U28295 (N_28295,N_28103,N_28179);
xor U28296 (N_28296,N_28144,N_28027);
or U28297 (N_28297,N_28018,N_28025);
xor U28298 (N_28298,N_28041,N_28028);
xnor U28299 (N_28299,N_28046,N_28054);
nor U28300 (N_28300,N_28086,N_28033);
nand U28301 (N_28301,N_28040,N_28123);
or U28302 (N_28302,N_28169,N_28111);
nand U28303 (N_28303,N_28154,N_28129);
xor U28304 (N_28304,N_28081,N_28114);
nand U28305 (N_28305,N_28011,N_28139);
nand U28306 (N_28306,N_28166,N_28159);
nor U28307 (N_28307,N_28140,N_28070);
nor U28308 (N_28308,N_28198,N_28083);
or U28309 (N_28309,N_28105,N_28161);
nor U28310 (N_28310,N_28142,N_28159);
nand U28311 (N_28311,N_28153,N_28073);
and U28312 (N_28312,N_28098,N_28068);
nor U28313 (N_28313,N_28135,N_28077);
nor U28314 (N_28314,N_28031,N_28092);
xor U28315 (N_28315,N_28130,N_28067);
or U28316 (N_28316,N_28034,N_28084);
xor U28317 (N_28317,N_28092,N_28141);
and U28318 (N_28318,N_28066,N_28043);
nand U28319 (N_28319,N_28035,N_28167);
xnor U28320 (N_28320,N_28135,N_28032);
nand U28321 (N_28321,N_28146,N_28188);
xor U28322 (N_28322,N_28054,N_28031);
nor U28323 (N_28323,N_28118,N_28031);
nand U28324 (N_28324,N_28016,N_28098);
nand U28325 (N_28325,N_28098,N_28088);
nand U28326 (N_28326,N_28117,N_28068);
and U28327 (N_28327,N_28056,N_28101);
and U28328 (N_28328,N_28115,N_28082);
or U28329 (N_28329,N_28188,N_28134);
nor U28330 (N_28330,N_28041,N_28017);
and U28331 (N_28331,N_28128,N_28158);
and U28332 (N_28332,N_28012,N_28106);
nor U28333 (N_28333,N_28069,N_28031);
or U28334 (N_28334,N_28103,N_28078);
xnor U28335 (N_28335,N_28015,N_28072);
nor U28336 (N_28336,N_28111,N_28028);
xor U28337 (N_28337,N_28043,N_28135);
or U28338 (N_28338,N_28076,N_28073);
nand U28339 (N_28339,N_28040,N_28010);
xor U28340 (N_28340,N_28058,N_28116);
and U28341 (N_28341,N_28060,N_28138);
nor U28342 (N_28342,N_28067,N_28123);
or U28343 (N_28343,N_28095,N_28180);
and U28344 (N_28344,N_28038,N_28054);
nor U28345 (N_28345,N_28076,N_28110);
or U28346 (N_28346,N_28052,N_28018);
xnor U28347 (N_28347,N_28098,N_28101);
xnor U28348 (N_28348,N_28005,N_28126);
and U28349 (N_28349,N_28097,N_28144);
or U28350 (N_28350,N_28075,N_28023);
nand U28351 (N_28351,N_28080,N_28015);
and U28352 (N_28352,N_28090,N_28005);
or U28353 (N_28353,N_28180,N_28183);
xnor U28354 (N_28354,N_28094,N_28176);
nand U28355 (N_28355,N_28100,N_28079);
xor U28356 (N_28356,N_28029,N_28073);
xor U28357 (N_28357,N_28191,N_28171);
and U28358 (N_28358,N_28075,N_28030);
nor U28359 (N_28359,N_28120,N_28039);
nand U28360 (N_28360,N_28091,N_28117);
nand U28361 (N_28361,N_28015,N_28151);
and U28362 (N_28362,N_28059,N_28178);
and U28363 (N_28363,N_28163,N_28175);
xor U28364 (N_28364,N_28191,N_28033);
and U28365 (N_28365,N_28111,N_28035);
and U28366 (N_28366,N_28175,N_28081);
or U28367 (N_28367,N_28124,N_28020);
or U28368 (N_28368,N_28004,N_28140);
nor U28369 (N_28369,N_28060,N_28119);
nand U28370 (N_28370,N_28112,N_28022);
or U28371 (N_28371,N_28034,N_28120);
or U28372 (N_28372,N_28096,N_28097);
nand U28373 (N_28373,N_28031,N_28111);
nor U28374 (N_28374,N_28194,N_28123);
and U28375 (N_28375,N_28038,N_28010);
or U28376 (N_28376,N_28172,N_28139);
and U28377 (N_28377,N_28082,N_28014);
nor U28378 (N_28378,N_28117,N_28010);
or U28379 (N_28379,N_28131,N_28052);
or U28380 (N_28380,N_28027,N_28055);
and U28381 (N_28381,N_28050,N_28191);
nor U28382 (N_28382,N_28053,N_28055);
or U28383 (N_28383,N_28165,N_28190);
xor U28384 (N_28384,N_28104,N_28168);
nor U28385 (N_28385,N_28191,N_28119);
and U28386 (N_28386,N_28020,N_28167);
nor U28387 (N_28387,N_28118,N_28048);
xor U28388 (N_28388,N_28143,N_28190);
xnor U28389 (N_28389,N_28180,N_28120);
xnor U28390 (N_28390,N_28060,N_28066);
and U28391 (N_28391,N_28054,N_28077);
or U28392 (N_28392,N_28038,N_28001);
and U28393 (N_28393,N_28098,N_28145);
nor U28394 (N_28394,N_28115,N_28176);
xnor U28395 (N_28395,N_28066,N_28061);
nand U28396 (N_28396,N_28163,N_28134);
xnor U28397 (N_28397,N_28100,N_28072);
and U28398 (N_28398,N_28166,N_28011);
or U28399 (N_28399,N_28162,N_28116);
nor U28400 (N_28400,N_28301,N_28267);
nor U28401 (N_28401,N_28296,N_28393);
nor U28402 (N_28402,N_28307,N_28209);
and U28403 (N_28403,N_28237,N_28367);
nand U28404 (N_28404,N_28366,N_28335);
or U28405 (N_28405,N_28349,N_28392);
or U28406 (N_28406,N_28266,N_28302);
or U28407 (N_28407,N_28255,N_28394);
nand U28408 (N_28408,N_28279,N_28397);
xor U28409 (N_28409,N_28399,N_28344);
and U28410 (N_28410,N_28239,N_28238);
nor U28411 (N_28411,N_28345,N_28231);
nand U28412 (N_28412,N_28329,N_28292);
xnor U28413 (N_28413,N_28351,N_28265);
and U28414 (N_28414,N_28340,N_28253);
xnor U28415 (N_28415,N_28378,N_28202);
nor U28416 (N_28416,N_28334,N_28306);
nor U28417 (N_28417,N_28230,N_28234);
and U28418 (N_28418,N_28374,N_28336);
or U28419 (N_28419,N_28208,N_28369);
or U28420 (N_28420,N_28201,N_28224);
xnor U28421 (N_28421,N_28368,N_28256);
or U28422 (N_28422,N_28298,N_28317);
xnor U28423 (N_28423,N_28246,N_28288);
or U28424 (N_28424,N_28229,N_28376);
nand U28425 (N_28425,N_28293,N_28385);
nand U28426 (N_28426,N_28278,N_28322);
or U28427 (N_28427,N_28291,N_28272);
and U28428 (N_28428,N_28299,N_28284);
or U28429 (N_28429,N_28373,N_28310);
nand U28430 (N_28430,N_28295,N_28371);
xor U28431 (N_28431,N_28361,N_28252);
xnor U28432 (N_28432,N_28262,N_28372);
and U28433 (N_28433,N_28219,N_28289);
or U28434 (N_28434,N_28270,N_28206);
nand U28435 (N_28435,N_28387,N_28247);
xnor U28436 (N_28436,N_28323,N_28314);
or U28437 (N_28437,N_28282,N_28381);
and U28438 (N_28438,N_28297,N_28382);
nand U28439 (N_28439,N_28386,N_28333);
xor U28440 (N_28440,N_28359,N_28241);
or U28441 (N_28441,N_28342,N_28330);
nor U28442 (N_28442,N_28218,N_28346);
xnor U28443 (N_28443,N_28365,N_28261);
or U28444 (N_28444,N_28204,N_28325);
xor U28445 (N_28445,N_28259,N_28287);
and U28446 (N_28446,N_28352,N_28347);
and U28447 (N_28447,N_28227,N_28271);
nor U28448 (N_28448,N_28380,N_28274);
xnor U28449 (N_28449,N_28254,N_28250);
nand U28450 (N_28450,N_28258,N_28205);
nor U28451 (N_28451,N_28236,N_28275);
and U28452 (N_28452,N_28348,N_28277);
xor U28453 (N_28453,N_28243,N_28364);
nand U28454 (N_28454,N_28300,N_28264);
nor U28455 (N_28455,N_28221,N_28309);
nand U28456 (N_28456,N_28211,N_28281);
nor U28457 (N_28457,N_28316,N_28244);
and U28458 (N_28458,N_28327,N_28290);
or U28459 (N_28459,N_28398,N_28356);
or U28460 (N_28460,N_28222,N_28226);
nand U28461 (N_28461,N_28280,N_28355);
nand U28462 (N_28462,N_28311,N_28269);
and U28463 (N_28463,N_28220,N_28248);
nor U28464 (N_28464,N_28212,N_28363);
or U28465 (N_28465,N_28326,N_28263);
or U28466 (N_28466,N_28388,N_28353);
xnor U28467 (N_28467,N_28232,N_28242);
and U28468 (N_28468,N_28315,N_28319);
nor U28469 (N_28469,N_28350,N_28228);
nor U28470 (N_28470,N_28313,N_28303);
nor U28471 (N_28471,N_28207,N_28338);
nand U28472 (N_28472,N_28249,N_28321);
and U28473 (N_28473,N_28260,N_28308);
or U28474 (N_28474,N_28215,N_28233);
nor U28475 (N_28475,N_28379,N_28268);
and U28476 (N_28476,N_28304,N_28390);
xnor U28477 (N_28477,N_28337,N_28273);
xnor U28478 (N_28478,N_28339,N_28245);
xor U28479 (N_28479,N_28203,N_28312);
xor U28480 (N_28480,N_28251,N_28391);
nand U28481 (N_28481,N_28370,N_28213);
xor U28482 (N_28482,N_28362,N_28384);
xor U28483 (N_28483,N_28360,N_28395);
xor U28484 (N_28484,N_28375,N_28354);
nor U28485 (N_28485,N_28389,N_28320);
and U28486 (N_28486,N_28216,N_28305);
nand U28487 (N_28487,N_28294,N_28324);
nor U28488 (N_28488,N_28318,N_28357);
nor U28489 (N_28489,N_28283,N_28225);
nor U28490 (N_28490,N_28286,N_28358);
nor U28491 (N_28491,N_28223,N_28210);
and U28492 (N_28492,N_28240,N_28383);
or U28493 (N_28493,N_28341,N_28257);
or U28494 (N_28494,N_28276,N_28285);
xor U28495 (N_28495,N_28343,N_28214);
xnor U28496 (N_28496,N_28396,N_28328);
or U28497 (N_28497,N_28377,N_28217);
xor U28498 (N_28498,N_28332,N_28331);
or U28499 (N_28499,N_28200,N_28235);
and U28500 (N_28500,N_28325,N_28245);
and U28501 (N_28501,N_28289,N_28313);
nor U28502 (N_28502,N_28383,N_28331);
and U28503 (N_28503,N_28386,N_28230);
nand U28504 (N_28504,N_28283,N_28361);
nor U28505 (N_28505,N_28380,N_28217);
or U28506 (N_28506,N_28369,N_28317);
or U28507 (N_28507,N_28229,N_28263);
nand U28508 (N_28508,N_28316,N_28334);
nor U28509 (N_28509,N_28255,N_28259);
xnor U28510 (N_28510,N_28361,N_28233);
or U28511 (N_28511,N_28286,N_28284);
and U28512 (N_28512,N_28355,N_28339);
nor U28513 (N_28513,N_28280,N_28392);
nand U28514 (N_28514,N_28350,N_28281);
or U28515 (N_28515,N_28302,N_28298);
nor U28516 (N_28516,N_28294,N_28253);
and U28517 (N_28517,N_28234,N_28295);
or U28518 (N_28518,N_28307,N_28353);
nor U28519 (N_28519,N_28238,N_28224);
or U28520 (N_28520,N_28349,N_28341);
nand U28521 (N_28521,N_28205,N_28347);
and U28522 (N_28522,N_28264,N_28388);
nand U28523 (N_28523,N_28311,N_28315);
or U28524 (N_28524,N_28383,N_28347);
and U28525 (N_28525,N_28392,N_28250);
nand U28526 (N_28526,N_28350,N_28200);
nor U28527 (N_28527,N_28297,N_28257);
xor U28528 (N_28528,N_28214,N_28246);
nor U28529 (N_28529,N_28359,N_28310);
or U28530 (N_28530,N_28332,N_28315);
xor U28531 (N_28531,N_28377,N_28281);
and U28532 (N_28532,N_28309,N_28274);
nand U28533 (N_28533,N_28312,N_28294);
xor U28534 (N_28534,N_28345,N_28331);
nand U28535 (N_28535,N_28285,N_28270);
xor U28536 (N_28536,N_28248,N_28298);
nand U28537 (N_28537,N_28302,N_28367);
nand U28538 (N_28538,N_28272,N_28213);
and U28539 (N_28539,N_28202,N_28291);
and U28540 (N_28540,N_28342,N_28239);
nor U28541 (N_28541,N_28280,N_28391);
or U28542 (N_28542,N_28263,N_28322);
and U28543 (N_28543,N_28311,N_28394);
and U28544 (N_28544,N_28347,N_28296);
or U28545 (N_28545,N_28326,N_28346);
or U28546 (N_28546,N_28247,N_28337);
or U28547 (N_28547,N_28234,N_28290);
xnor U28548 (N_28548,N_28380,N_28384);
nor U28549 (N_28549,N_28286,N_28274);
and U28550 (N_28550,N_28396,N_28289);
nor U28551 (N_28551,N_28241,N_28381);
nand U28552 (N_28552,N_28268,N_28212);
and U28553 (N_28553,N_28249,N_28366);
or U28554 (N_28554,N_28262,N_28359);
nand U28555 (N_28555,N_28323,N_28366);
and U28556 (N_28556,N_28209,N_28242);
nand U28557 (N_28557,N_28234,N_28338);
xor U28558 (N_28558,N_28289,N_28256);
or U28559 (N_28559,N_28246,N_28285);
and U28560 (N_28560,N_28264,N_28324);
or U28561 (N_28561,N_28315,N_28261);
or U28562 (N_28562,N_28255,N_28284);
nor U28563 (N_28563,N_28284,N_28230);
nand U28564 (N_28564,N_28314,N_28369);
and U28565 (N_28565,N_28265,N_28357);
and U28566 (N_28566,N_28269,N_28292);
nand U28567 (N_28567,N_28371,N_28284);
xor U28568 (N_28568,N_28294,N_28273);
and U28569 (N_28569,N_28269,N_28350);
and U28570 (N_28570,N_28374,N_28328);
or U28571 (N_28571,N_28393,N_28262);
xor U28572 (N_28572,N_28333,N_28201);
nand U28573 (N_28573,N_28340,N_28307);
xor U28574 (N_28574,N_28286,N_28239);
or U28575 (N_28575,N_28339,N_28269);
and U28576 (N_28576,N_28202,N_28301);
or U28577 (N_28577,N_28397,N_28233);
xnor U28578 (N_28578,N_28297,N_28324);
and U28579 (N_28579,N_28383,N_28349);
nand U28580 (N_28580,N_28384,N_28304);
nor U28581 (N_28581,N_28273,N_28282);
or U28582 (N_28582,N_28296,N_28390);
xnor U28583 (N_28583,N_28314,N_28330);
nand U28584 (N_28584,N_28228,N_28222);
xnor U28585 (N_28585,N_28340,N_28339);
nor U28586 (N_28586,N_28337,N_28373);
nor U28587 (N_28587,N_28254,N_28377);
xor U28588 (N_28588,N_28326,N_28267);
xnor U28589 (N_28589,N_28291,N_28258);
nor U28590 (N_28590,N_28255,N_28247);
nor U28591 (N_28591,N_28240,N_28349);
xor U28592 (N_28592,N_28372,N_28204);
xnor U28593 (N_28593,N_28295,N_28231);
and U28594 (N_28594,N_28313,N_28225);
or U28595 (N_28595,N_28334,N_28237);
nor U28596 (N_28596,N_28349,N_28235);
or U28597 (N_28597,N_28346,N_28311);
xor U28598 (N_28598,N_28274,N_28222);
nand U28599 (N_28599,N_28216,N_28359);
and U28600 (N_28600,N_28588,N_28404);
xnor U28601 (N_28601,N_28523,N_28538);
nor U28602 (N_28602,N_28505,N_28550);
and U28603 (N_28603,N_28443,N_28534);
and U28604 (N_28604,N_28420,N_28496);
or U28605 (N_28605,N_28484,N_28573);
nor U28606 (N_28606,N_28545,N_28528);
nor U28607 (N_28607,N_28515,N_28421);
nand U28608 (N_28608,N_28444,N_28530);
or U28609 (N_28609,N_28522,N_28463);
nand U28610 (N_28610,N_28467,N_28480);
or U28611 (N_28611,N_28596,N_28532);
nand U28612 (N_28612,N_28439,N_28424);
nand U28613 (N_28613,N_28524,N_28462);
xnor U28614 (N_28614,N_28442,N_28542);
nor U28615 (N_28615,N_28475,N_28431);
or U28616 (N_28616,N_28422,N_28509);
and U28617 (N_28617,N_28473,N_28437);
xor U28618 (N_28618,N_28568,N_28458);
or U28619 (N_28619,N_28429,N_28460);
nand U28620 (N_28620,N_28579,N_28586);
xnor U28621 (N_28621,N_28436,N_28500);
nand U28622 (N_28622,N_28518,N_28571);
or U28623 (N_28623,N_28565,N_28453);
xor U28624 (N_28624,N_28427,N_28526);
nand U28625 (N_28625,N_28445,N_28537);
nand U28626 (N_28626,N_28451,N_28447);
and U28627 (N_28627,N_28511,N_28557);
or U28628 (N_28628,N_28481,N_28470);
nor U28629 (N_28629,N_28591,N_28413);
or U28630 (N_28630,N_28501,N_28527);
nor U28631 (N_28631,N_28461,N_28455);
or U28632 (N_28632,N_28598,N_28589);
nand U28633 (N_28633,N_28578,N_28418);
xnor U28634 (N_28634,N_28508,N_28547);
and U28635 (N_28635,N_28465,N_28417);
nand U28636 (N_28636,N_28449,N_28407);
xnor U28637 (N_28637,N_28503,N_28432);
xor U28638 (N_28638,N_28502,N_28599);
nor U28639 (N_28639,N_28577,N_28492);
and U28640 (N_28640,N_28477,N_28519);
nor U28641 (N_28641,N_28574,N_28498);
xor U28642 (N_28642,N_28543,N_28561);
xnor U28643 (N_28643,N_28535,N_28454);
and U28644 (N_28644,N_28569,N_28540);
and U28645 (N_28645,N_28576,N_28552);
and U28646 (N_28646,N_28474,N_28488);
and U28647 (N_28647,N_28464,N_28411);
and U28648 (N_28648,N_28597,N_28580);
and U28649 (N_28649,N_28433,N_28582);
nor U28650 (N_28650,N_28567,N_28520);
xnor U28651 (N_28651,N_28416,N_28548);
and U28652 (N_28652,N_28494,N_28593);
or U28653 (N_28653,N_28479,N_28441);
nand U28654 (N_28654,N_28434,N_28452);
xor U28655 (N_28655,N_28403,N_28400);
xnor U28656 (N_28656,N_28435,N_28493);
nand U28657 (N_28657,N_28584,N_28525);
or U28658 (N_28658,N_28570,N_28562);
nor U28659 (N_28659,N_28560,N_28556);
and U28660 (N_28660,N_28476,N_28531);
nand U28661 (N_28661,N_28425,N_28456);
or U28662 (N_28662,N_28533,N_28472);
or U28663 (N_28663,N_28541,N_28595);
nand U28664 (N_28664,N_28536,N_28409);
nand U28665 (N_28665,N_28410,N_28405);
and U28666 (N_28666,N_28482,N_28551);
nand U28667 (N_28667,N_28521,N_28513);
xor U28668 (N_28668,N_28468,N_28558);
or U28669 (N_28669,N_28566,N_28544);
nand U28670 (N_28670,N_28450,N_28555);
xnor U28671 (N_28671,N_28485,N_28572);
nand U28672 (N_28672,N_28559,N_28415);
xor U28673 (N_28673,N_28510,N_28457);
xor U28674 (N_28674,N_28402,N_28554);
and U28675 (N_28675,N_28430,N_28512);
and U28676 (N_28676,N_28490,N_28448);
or U28677 (N_28677,N_28563,N_28497);
nor U28678 (N_28678,N_28592,N_28590);
and U28679 (N_28679,N_28419,N_28517);
and U28680 (N_28680,N_28471,N_28440);
nand U28681 (N_28681,N_28491,N_28529);
nor U28682 (N_28682,N_28478,N_28587);
xor U28683 (N_28683,N_28575,N_28553);
and U28684 (N_28684,N_28514,N_28585);
or U28685 (N_28685,N_28581,N_28483);
or U28686 (N_28686,N_28507,N_28487);
and U28687 (N_28687,N_28408,N_28539);
xor U28688 (N_28688,N_28406,N_28466);
nand U28689 (N_28689,N_28495,N_28516);
xnor U28690 (N_28690,N_28546,N_28549);
and U28691 (N_28691,N_28499,N_28564);
nand U28692 (N_28692,N_28401,N_28469);
xnor U28693 (N_28693,N_28414,N_28412);
and U28694 (N_28694,N_28506,N_28426);
and U28695 (N_28695,N_28594,N_28583);
xor U28696 (N_28696,N_28489,N_28438);
xnor U28697 (N_28697,N_28459,N_28486);
xnor U28698 (N_28698,N_28428,N_28423);
nand U28699 (N_28699,N_28504,N_28446);
or U28700 (N_28700,N_28406,N_28529);
or U28701 (N_28701,N_28403,N_28422);
or U28702 (N_28702,N_28564,N_28580);
nand U28703 (N_28703,N_28571,N_28548);
and U28704 (N_28704,N_28548,N_28592);
xnor U28705 (N_28705,N_28533,N_28411);
nand U28706 (N_28706,N_28454,N_28481);
or U28707 (N_28707,N_28414,N_28543);
or U28708 (N_28708,N_28425,N_28589);
nor U28709 (N_28709,N_28587,N_28569);
nand U28710 (N_28710,N_28442,N_28439);
and U28711 (N_28711,N_28477,N_28508);
nor U28712 (N_28712,N_28415,N_28518);
xor U28713 (N_28713,N_28504,N_28588);
xnor U28714 (N_28714,N_28578,N_28450);
or U28715 (N_28715,N_28447,N_28512);
nand U28716 (N_28716,N_28463,N_28422);
nor U28717 (N_28717,N_28597,N_28408);
nand U28718 (N_28718,N_28550,N_28410);
and U28719 (N_28719,N_28547,N_28444);
and U28720 (N_28720,N_28434,N_28407);
xnor U28721 (N_28721,N_28485,N_28429);
or U28722 (N_28722,N_28491,N_28501);
and U28723 (N_28723,N_28573,N_28571);
nand U28724 (N_28724,N_28439,N_28433);
xor U28725 (N_28725,N_28530,N_28569);
xor U28726 (N_28726,N_28544,N_28494);
nor U28727 (N_28727,N_28537,N_28418);
nand U28728 (N_28728,N_28417,N_28507);
nand U28729 (N_28729,N_28565,N_28436);
nor U28730 (N_28730,N_28558,N_28586);
nor U28731 (N_28731,N_28537,N_28426);
xnor U28732 (N_28732,N_28564,N_28597);
and U28733 (N_28733,N_28456,N_28564);
xnor U28734 (N_28734,N_28443,N_28565);
and U28735 (N_28735,N_28434,N_28531);
nand U28736 (N_28736,N_28461,N_28525);
or U28737 (N_28737,N_28581,N_28504);
or U28738 (N_28738,N_28416,N_28542);
and U28739 (N_28739,N_28593,N_28515);
or U28740 (N_28740,N_28460,N_28459);
nor U28741 (N_28741,N_28588,N_28532);
and U28742 (N_28742,N_28589,N_28412);
nor U28743 (N_28743,N_28457,N_28486);
and U28744 (N_28744,N_28497,N_28577);
xor U28745 (N_28745,N_28459,N_28409);
nand U28746 (N_28746,N_28489,N_28463);
or U28747 (N_28747,N_28556,N_28411);
and U28748 (N_28748,N_28472,N_28514);
or U28749 (N_28749,N_28597,N_28570);
nand U28750 (N_28750,N_28537,N_28505);
and U28751 (N_28751,N_28513,N_28440);
xnor U28752 (N_28752,N_28487,N_28455);
xor U28753 (N_28753,N_28593,N_28531);
nor U28754 (N_28754,N_28420,N_28470);
nor U28755 (N_28755,N_28458,N_28406);
nor U28756 (N_28756,N_28570,N_28505);
and U28757 (N_28757,N_28599,N_28579);
or U28758 (N_28758,N_28458,N_28475);
and U28759 (N_28759,N_28509,N_28421);
nand U28760 (N_28760,N_28560,N_28575);
xnor U28761 (N_28761,N_28452,N_28475);
xor U28762 (N_28762,N_28413,N_28550);
or U28763 (N_28763,N_28579,N_28499);
and U28764 (N_28764,N_28500,N_28532);
and U28765 (N_28765,N_28458,N_28592);
nand U28766 (N_28766,N_28482,N_28404);
and U28767 (N_28767,N_28421,N_28553);
nand U28768 (N_28768,N_28495,N_28510);
nand U28769 (N_28769,N_28480,N_28495);
and U28770 (N_28770,N_28597,N_28587);
nand U28771 (N_28771,N_28538,N_28484);
xnor U28772 (N_28772,N_28473,N_28455);
nor U28773 (N_28773,N_28445,N_28440);
xnor U28774 (N_28774,N_28544,N_28478);
and U28775 (N_28775,N_28420,N_28500);
or U28776 (N_28776,N_28582,N_28593);
nand U28777 (N_28777,N_28532,N_28479);
nand U28778 (N_28778,N_28554,N_28524);
nand U28779 (N_28779,N_28460,N_28564);
xor U28780 (N_28780,N_28498,N_28537);
xnor U28781 (N_28781,N_28446,N_28524);
xnor U28782 (N_28782,N_28429,N_28582);
or U28783 (N_28783,N_28413,N_28444);
nand U28784 (N_28784,N_28522,N_28479);
or U28785 (N_28785,N_28561,N_28402);
nor U28786 (N_28786,N_28490,N_28528);
nand U28787 (N_28787,N_28530,N_28594);
and U28788 (N_28788,N_28520,N_28467);
and U28789 (N_28789,N_28534,N_28500);
xnor U28790 (N_28790,N_28411,N_28438);
nor U28791 (N_28791,N_28444,N_28564);
xor U28792 (N_28792,N_28449,N_28590);
xor U28793 (N_28793,N_28435,N_28457);
nand U28794 (N_28794,N_28434,N_28559);
and U28795 (N_28795,N_28480,N_28464);
xor U28796 (N_28796,N_28498,N_28509);
and U28797 (N_28797,N_28443,N_28442);
and U28798 (N_28798,N_28452,N_28425);
and U28799 (N_28799,N_28466,N_28476);
nor U28800 (N_28800,N_28756,N_28649);
and U28801 (N_28801,N_28679,N_28769);
and U28802 (N_28802,N_28669,N_28779);
xor U28803 (N_28803,N_28621,N_28688);
xor U28804 (N_28804,N_28662,N_28623);
xor U28805 (N_28805,N_28765,N_28608);
or U28806 (N_28806,N_28778,N_28722);
and U28807 (N_28807,N_28788,N_28663);
or U28808 (N_28808,N_28785,N_28772);
and U28809 (N_28809,N_28696,N_28665);
xnor U28810 (N_28810,N_28745,N_28757);
nand U28811 (N_28811,N_28768,N_28796);
nor U28812 (N_28812,N_28707,N_28658);
and U28813 (N_28813,N_28750,N_28746);
nor U28814 (N_28814,N_28681,N_28701);
nand U28815 (N_28815,N_28791,N_28712);
and U28816 (N_28816,N_28790,N_28693);
xor U28817 (N_28817,N_28773,N_28715);
xnor U28818 (N_28818,N_28735,N_28651);
xor U28819 (N_28819,N_28683,N_28695);
or U28820 (N_28820,N_28781,N_28766);
nand U28821 (N_28821,N_28793,N_28603);
or U28822 (N_28822,N_28761,N_28748);
or U28823 (N_28823,N_28615,N_28640);
xor U28824 (N_28824,N_28638,N_28648);
xor U28825 (N_28825,N_28607,N_28720);
and U28826 (N_28826,N_28616,N_28789);
nor U28827 (N_28827,N_28653,N_28717);
and U28828 (N_28828,N_28786,N_28742);
nor U28829 (N_28829,N_28727,N_28784);
or U28830 (N_28830,N_28703,N_28776);
and U28831 (N_28831,N_28737,N_28689);
nor U28832 (N_28832,N_28645,N_28747);
or U28833 (N_28833,N_28646,N_28626);
xnor U28834 (N_28834,N_28628,N_28733);
xnor U28835 (N_28835,N_28754,N_28780);
nor U28836 (N_28836,N_28680,N_28667);
and U28837 (N_28837,N_28611,N_28619);
or U28838 (N_28838,N_28631,N_28726);
or U28839 (N_28839,N_28751,N_28674);
and U28840 (N_28840,N_28795,N_28633);
and U28841 (N_28841,N_28714,N_28601);
and U28842 (N_28842,N_28650,N_28702);
and U28843 (N_28843,N_28738,N_28659);
xor U28844 (N_28844,N_28661,N_28618);
nand U28845 (N_28845,N_28713,N_28610);
nand U28846 (N_28846,N_28764,N_28692);
or U28847 (N_28847,N_28760,N_28668);
and U28848 (N_28848,N_28632,N_28637);
and U28849 (N_28849,N_28798,N_28716);
xnor U28850 (N_28850,N_28752,N_28759);
or U28851 (N_28851,N_28787,N_28636);
nor U28852 (N_28852,N_28676,N_28670);
or U28853 (N_28853,N_28634,N_28725);
nand U28854 (N_28854,N_28777,N_28739);
xor U28855 (N_28855,N_28605,N_28771);
nand U28856 (N_28856,N_28691,N_28635);
or U28857 (N_28857,N_28654,N_28718);
and U28858 (N_28858,N_28673,N_28794);
or U28859 (N_28859,N_28684,N_28710);
nor U28860 (N_28860,N_28709,N_28723);
xor U28861 (N_28861,N_28644,N_28762);
nand U28862 (N_28862,N_28770,N_28629);
xnor U28863 (N_28863,N_28774,N_28617);
nor U28864 (N_28864,N_28706,N_28731);
xor U28865 (N_28865,N_28678,N_28763);
xor U28866 (N_28866,N_28767,N_28729);
nor U28867 (N_28867,N_28620,N_28698);
nor U28868 (N_28868,N_28606,N_28604);
nor U28869 (N_28869,N_28630,N_28799);
nor U28870 (N_28870,N_28749,N_28753);
nand U28871 (N_28871,N_28743,N_28721);
nand U28872 (N_28872,N_28677,N_28647);
and U28873 (N_28873,N_28700,N_28643);
or U28874 (N_28874,N_28666,N_28792);
or U28875 (N_28875,N_28622,N_28641);
nand U28876 (N_28876,N_28656,N_28600);
nand U28877 (N_28877,N_28655,N_28613);
xnor U28878 (N_28878,N_28734,N_28625);
nor U28879 (N_28879,N_28694,N_28657);
nor U28880 (N_28880,N_28612,N_28740);
or U28881 (N_28881,N_28782,N_28624);
nor U28882 (N_28882,N_28660,N_28705);
nor U28883 (N_28883,N_28736,N_28685);
nor U28884 (N_28884,N_28783,N_28652);
nand U28885 (N_28885,N_28744,N_28686);
nand U28886 (N_28886,N_28602,N_28728);
xor U28887 (N_28887,N_28609,N_28708);
nand U28888 (N_28888,N_28755,N_28724);
xnor U28889 (N_28889,N_28627,N_28687);
and U28890 (N_28890,N_28699,N_28697);
nor U28891 (N_28891,N_28642,N_28664);
and U28892 (N_28892,N_28741,N_28732);
xor U28893 (N_28893,N_28719,N_28675);
nand U28894 (N_28894,N_28690,N_28797);
and U28895 (N_28895,N_28730,N_28711);
xor U28896 (N_28896,N_28639,N_28672);
nand U28897 (N_28897,N_28671,N_28704);
and U28898 (N_28898,N_28614,N_28758);
nor U28899 (N_28899,N_28682,N_28775);
and U28900 (N_28900,N_28671,N_28795);
xor U28901 (N_28901,N_28667,N_28718);
nand U28902 (N_28902,N_28628,N_28672);
nand U28903 (N_28903,N_28779,N_28737);
or U28904 (N_28904,N_28782,N_28721);
and U28905 (N_28905,N_28630,N_28676);
or U28906 (N_28906,N_28602,N_28601);
nand U28907 (N_28907,N_28787,N_28694);
and U28908 (N_28908,N_28716,N_28738);
nand U28909 (N_28909,N_28758,N_28605);
and U28910 (N_28910,N_28775,N_28799);
nor U28911 (N_28911,N_28704,N_28603);
nand U28912 (N_28912,N_28693,N_28774);
or U28913 (N_28913,N_28603,N_28759);
nor U28914 (N_28914,N_28747,N_28662);
or U28915 (N_28915,N_28612,N_28789);
xor U28916 (N_28916,N_28623,N_28607);
nor U28917 (N_28917,N_28684,N_28687);
and U28918 (N_28918,N_28694,N_28631);
nor U28919 (N_28919,N_28764,N_28752);
nor U28920 (N_28920,N_28795,N_28765);
xor U28921 (N_28921,N_28775,N_28784);
or U28922 (N_28922,N_28763,N_28720);
nor U28923 (N_28923,N_28633,N_28768);
xnor U28924 (N_28924,N_28607,N_28631);
xor U28925 (N_28925,N_28753,N_28727);
nand U28926 (N_28926,N_28659,N_28769);
and U28927 (N_28927,N_28658,N_28721);
and U28928 (N_28928,N_28768,N_28737);
nand U28929 (N_28929,N_28620,N_28690);
or U28930 (N_28930,N_28738,N_28790);
nor U28931 (N_28931,N_28681,N_28612);
nor U28932 (N_28932,N_28784,N_28636);
and U28933 (N_28933,N_28623,N_28704);
nand U28934 (N_28934,N_28710,N_28673);
and U28935 (N_28935,N_28752,N_28728);
and U28936 (N_28936,N_28624,N_28608);
nand U28937 (N_28937,N_28714,N_28777);
nor U28938 (N_28938,N_28746,N_28630);
or U28939 (N_28939,N_28698,N_28739);
and U28940 (N_28940,N_28683,N_28603);
xor U28941 (N_28941,N_28666,N_28702);
nand U28942 (N_28942,N_28603,N_28786);
nand U28943 (N_28943,N_28747,N_28623);
nand U28944 (N_28944,N_28617,N_28635);
xor U28945 (N_28945,N_28641,N_28645);
or U28946 (N_28946,N_28795,N_28645);
and U28947 (N_28947,N_28612,N_28693);
xor U28948 (N_28948,N_28798,N_28763);
nor U28949 (N_28949,N_28605,N_28722);
or U28950 (N_28950,N_28720,N_28653);
and U28951 (N_28951,N_28691,N_28687);
nor U28952 (N_28952,N_28687,N_28672);
xnor U28953 (N_28953,N_28635,N_28636);
xor U28954 (N_28954,N_28709,N_28771);
or U28955 (N_28955,N_28640,N_28667);
nand U28956 (N_28956,N_28649,N_28635);
or U28957 (N_28957,N_28601,N_28623);
xor U28958 (N_28958,N_28795,N_28647);
or U28959 (N_28959,N_28767,N_28711);
nor U28960 (N_28960,N_28709,N_28694);
nor U28961 (N_28961,N_28747,N_28630);
xnor U28962 (N_28962,N_28706,N_28665);
or U28963 (N_28963,N_28644,N_28647);
and U28964 (N_28964,N_28688,N_28660);
nor U28965 (N_28965,N_28751,N_28727);
nor U28966 (N_28966,N_28724,N_28723);
nor U28967 (N_28967,N_28666,N_28683);
nor U28968 (N_28968,N_28789,N_28662);
and U28969 (N_28969,N_28758,N_28604);
or U28970 (N_28970,N_28609,N_28663);
and U28971 (N_28971,N_28733,N_28718);
xor U28972 (N_28972,N_28713,N_28743);
nor U28973 (N_28973,N_28751,N_28718);
nor U28974 (N_28974,N_28790,N_28773);
and U28975 (N_28975,N_28634,N_28757);
xnor U28976 (N_28976,N_28727,N_28729);
or U28977 (N_28977,N_28784,N_28709);
nor U28978 (N_28978,N_28787,N_28601);
or U28979 (N_28979,N_28783,N_28771);
nand U28980 (N_28980,N_28615,N_28691);
nand U28981 (N_28981,N_28789,N_28633);
or U28982 (N_28982,N_28621,N_28608);
and U28983 (N_28983,N_28724,N_28754);
nor U28984 (N_28984,N_28795,N_28700);
nand U28985 (N_28985,N_28757,N_28621);
xor U28986 (N_28986,N_28697,N_28667);
or U28987 (N_28987,N_28729,N_28639);
and U28988 (N_28988,N_28694,N_28730);
or U28989 (N_28989,N_28792,N_28605);
nand U28990 (N_28990,N_28768,N_28617);
xnor U28991 (N_28991,N_28793,N_28621);
or U28992 (N_28992,N_28611,N_28641);
and U28993 (N_28993,N_28718,N_28696);
and U28994 (N_28994,N_28792,N_28614);
or U28995 (N_28995,N_28786,N_28626);
or U28996 (N_28996,N_28764,N_28644);
or U28997 (N_28997,N_28633,N_28669);
xnor U28998 (N_28998,N_28727,N_28758);
and U28999 (N_28999,N_28636,N_28696);
nor U29000 (N_29000,N_28852,N_28895);
nand U29001 (N_29001,N_28841,N_28894);
or U29002 (N_29002,N_28840,N_28866);
xnor U29003 (N_29003,N_28872,N_28849);
nand U29004 (N_29004,N_28941,N_28805);
and U29005 (N_29005,N_28980,N_28951);
or U29006 (N_29006,N_28931,N_28915);
nor U29007 (N_29007,N_28820,N_28998);
and U29008 (N_29008,N_28833,N_28892);
nand U29009 (N_29009,N_28832,N_28873);
nor U29010 (N_29010,N_28933,N_28870);
or U29011 (N_29011,N_28878,N_28958);
nand U29012 (N_29012,N_28874,N_28854);
or U29013 (N_29013,N_28903,N_28896);
and U29014 (N_29014,N_28856,N_28992);
nor U29015 (N_29015,N_28819,N_28827);
xor U29016 (N_29016,N_28863,N_28959);
nand U29017 (N_29017,N_28829,N_28802);
xnor U29018 (N_29018,N_28855,N_28924);
or U29019 (N_29019,N_28900,N_28991);
xnor U29020 (N_29020,N_28930,N_28834);
nand U29021 (N_29021,N_28977,N_28871);
and U29022 (N_29022,N_28969,N_28962);
nand U29023 (N_29023,N_28953,N_28859);
nor U29024 (N_29024,N_28822,N_28916);
or U29025 (N_29025,N_28961,N_28823);
xnor U29026 (N_29026,N_28801,N_28808);
nor U29027 (N_29027,N_28811,N_28932);
nand U29028 (N_29028,N_28821,N_28975);
xor U29029 (N_29029,N_28848,N_28826);
nor U29030 (N_29030,N_28913,N_28902);
and U29031 (N_29031,N_28899,N_28918);
and U29032 (N_29032,N_28945,N_28814);
nor U29033 (N_29033,N_28816,N_28883);
nor U29034 (N_29034,N_28920,N_28877);
nand U29035 (N_29035,N_28890,N_28867);
and U29036 (N_29036,N_28937,N_28844);
nor U29037 (N_29037,N_28886,N_28864);
or U29038 (N_29038,N_28818,N_28947);
or U29039 (N_29039,N_28838,N_28809);
nor U29040 (N_29040,N_28988,N_28813);
xnor U29041 (N_29041,N_28926,N_28965);
or U29042 (N_29042,N_28831,N_28800);
xnor U29043 (N_29043,N_28939,N_28955);
xnor U29044 (N_29044,N_28887,N_28964);
and U29045 (N_29045,N_28944,N_28990);
xnor U29046 (N_29046,N_28911,N_28989);
and U29047 (N_29047,N_28972,N_28881);
and U29048 (N_29048,N_28815,N_28860);
or U29049 (N_29049,N_28935,N_28922);
nor U29050 (N_29050,N_28936,N_28997);
xor U29051 (N_29051,N_28901,N_28847);
nand U29052 (N_29052,N_28865,N_28830);
nor U29053 (N_29053,N_28869,N_28940);
or U29054 (N_29054,N_28974,N_28912);
nand U29055 (N_29055,N_28839,N_28828);
and U29056 (N_29056,N_28981,N_28966);
nand U29057 (N_29057,N_28982,N_28835);
nand U29058 (N_29058,N_28925,N_28943);
nand U29059 (N_29059,N_28978,N_28885);
or U29060 (N_29060,N_28898,N_28893);
nand U29061 (N_29061,N_28942,N_28986);
or U29062 (N_29062,N_28812,N_28968);
nor U29063 (N_29063,N_28876,N_28904);
or U29064 (N_29064,N_28910,N_28868);
and U29065 (N_29065,N_28907,N_28825);
xnor U29066 (N_29066,N_28908,N_28880);
and U29067 (N_29067,N_28824,N_28843);
xnor U29068 (N_29068,N_28948,N_28906);
or U29069 (N_29069,N_28987,N_28970);
nand U29070 (N_29070,N_28853,N_28983);
and U29071 (N_29071,N_28967,N_28862);
nand U29072 (N_29072,N_28914,N_28857);
nand U29073 (N_29073,N_28804,N_28952);
nand U29074 (N_29074,N_28949,N_28909);
nand U29075 (N_29075,N_28837,N_28973);
xnor U29076 (N_29076,N_28905,N_28810);
and U29077 (N_29077,N_28996,N_28845);
nand U29078 (N_29078,N_28817,N_28861);
nor U29079 (N_29079,N_28971,N_28976);
xnor U29080 (N_29080,N_28846,N_28807);
nand U29081 (N_29081,N_28995,N_28994);
or U29082 (N_29082,N_28985,N_28884);
nand U29083 (N_29083,N_28979,N_28934);
and U29084 (N_29084,N_28938,N_28891);
nor U29085 (N_29085,N_28999,N_28803);
xnor U29086 (N_29086,N_28917,N_28984);
xor U29087 (N_29087,N_28921,N_28919);
or U29088 (N_29088,N_28889,N_28957);
nor U29089 (N_29089,N_28882,N_28851);
or U29090 (N_29090,N_28879,N_28850);
and U29091 (N_29091,N_28927,N_28963);
and U29092 (N_29092,N_28897,N_28928);
nor U29093 (N_29093,N_28960,N_28950);
nand U29094 (N_29094,N_28875,N_28954);
or U29095 (N_29095,N_28929,N_28806);
nand U29096 (N_29096,N_28858,N_28946);
and U29097 (N_29097,N_28842,N_28956);
nor U29098 (N_29098,N_28923,N_28836);
and U29099 (N_29099,N_28993,N_28888);
nand U29100 (N_29100,N_28912,N_28838);
nor U29101 (N_29101,N_28865,N_28812);
xnor U29102 (N_29102,N_28897,N_28980);
nor U29103 (N_29103,N_28944,N_28931);
nand U29104 (N_29104,N_28834,N_28953);
nor U29105 (N_29105,N_28856,N_28813);
nand U29106 (N_29106,N_28856,N_28926);
nand U29107 (N_29107,N_28983,N_28894);
nor U29108 (N_29108,N_28923,N_28855);
and U29109 (N_29109,N_28902,N_28817);
and U29110 (N_29110,N_28803,N_28953);
or U29111 (N_29111,N_28836,N_28963);
and U29112 (N_29112,N_28904,N_28819);
xnor U29113 (N_29113,N_28837,N_28887);
or U29114 (N_29114,N_28965,N_28838);
nand U29115 (N_29115,N_28898,N_28917);
nor U29116 (N_29116,N_28814,N_28976);
xnor U29117 (N_29117,N_28989,N_28982);
xnor U29118 (N_29118,N_28874,N_28855);
and U29119 (N_29119,N_28896,N_28815);
xor U29120 (N_29120,N_28994,N_28859);
and U29121 (N_29121,N_28819,N_28967);
and U29122 (N_29122,N_28885,N_28808);
xor U29123 (N_29123,N_28899,N_28823);
nor U29124 (N_29124,N_28989,N_28844);
or U29125 (N_29125,N_28930,N_28920);
and U29126 (N_29126,N_28907,N_28859);
or U29127 (N_29127,N_28934,N_28846);
nor U29128 (N_29128,N_28801,N_28843);
and U29129 (N_29129,N_28856,N_28950);
and U29130 (N_29130,N_28856,N_28942);
and U29131 (N_29131,N_28906,N_28841);
nand U29132 (N_29132,N_28955,N_28977);
nor U29133 (N_29133,N_28999,N_28953);
or U29134 (N_29134,N_28969,N_28998);
nor U29135 (N_29135,N_28996,N_28906);
and U29136 (N_29136,N_28985,N_28999);
xnor U29137 (N_29137,N_28824,N_28906);
or U29138 (N_29138,N_28985,N_28911);
nand U29139 (N_29139,N_28990,N_28812);
and U29140 (N_29140,N_28929,N_28896);
xnor U29141 (N_29141,N_28895,N_28892);
nand U29142 (N_29142,N_28888,N_28806);
nand U29143 (N_29143,N_28830,N_28952);
and U29144 (N_29144,N_28806,N_28807);
nand U29145 (N_29145,N_28809,N_28944);
xor U29146 (N_29146,N_28930,N_28966);
nand U29147 (N_29147,N_28935,N_28955);
xnor U29148 (N_29148,N_28803,N_28972);
nor U29149 (N_29149,N_28895,N_28883);
nor U29150 (N_29150,N_28884,N_28816);
nand U29151 (N_29151,N_28841,N_28944);
nor U29152 (N_29152,N_28944,N_28995);
nand U29153 (N_29153,N_28926,N_28870);
nor U29154 (N_29154,N_28838,N_28904);
nor U29155 (N_29155,N_28880,N_28832);
or U29156 (N_29156,N_28931,N_28860);
nand U29157 (N_29157,N_28886,N_28945);
xnor U29158 (N_29158,N_28831,N_28809);
and U29159 (N_29159,N_28993,N_28859);
xnor U29160 (N_29160,N_28995,N_28884);
xnor U29161 (N_29161,N_28948,N_28964);
xnor U29162 (N_29162,N_28885,N_28853);
nor U29163 (N_29163,N_28853,N_28865);
and U29164 (N_29164,N_28809,N_28801);
xor U29165 (N_29165,N_28903,N_28998);
nand U29166 (N_29166,N_28964,N_28878);
or U29167 (N_29167,N_28910,N_28821);
nor U29168 (N_29168,N_28819,N_28993);
xor U29169 (N_29169,N_28891,N_28847);
nor U29170 (N_29170,N_28940,N_28814);
nor U29171 (N_29171,N_28830,N_28959);
nand U29172 (N_29172,N_28854,N_28957);
xnor U29173 (N_29173,N_28933,N_28803);
xor U29174 (N_29174,N_28931,N_28929);
nand U29175 (N_29175,N_28864,N_28881);
and U29176 (N_29176,N_28986,N_28813);
or U29177 (N_29177,N_28930,N_28968);
and U29178 (N_29178,N_28935,N_28999);
and U29179 (N_29179,N_28818,N_28994);
xnor U29180 (N_29180,N_28996,N_28877);
or U29181 (N_29181,N_28918,N_28880);
nand U29182 (N_29182,N_28981,N_28967);
xor U29183 (N_29183,N_28977,N_28864);
xor U29184 (N_29184,N_28986,N_28872);
and U29185 (N_29185,N_28925,N_28891);
and U29186 (N_29186,N_28822,N_28891);
nand U29187 (N_29187,N_28963,N_28894);
or U29188 (N_29188,N_28897,N_28997);
nor U29189 (N_29189,N_28800,N_28882);
xor U29190 (N_29190,N_28847,N_28970);
or U29191 (N_29191,N_28840,N_28953);
nand U29192 (N_29192,N_28893,N_28980);
or U29193 (N_29193,N_28959,N_28839);
or U29194 (N_29194,N_28884,N_28903);
and U29195 (N_29195,N_28957,N_28951);
or U29196 (N_29196,N_28884,N_28955);
xor U29197 (N_29197,N_28953,N_28844);
nand U29198 (N_29198,N_28978,N_28956);
and U29199 (N_29199,N_28820,N_28846);
or U29200 (N_29200,N_29057,N_29135);
or U29201 (N_29201,N_29128,N_29015);
nand U29202 (N_29202,N_29031,N_29028);
nor U29203 (N_29203,N_29194,N_29012);
xnor U29204 (N_29204,N_29059,N_29007);
nand U29205 (N_29205,N_29068,N_29101);
or U29206 (N_29206,N_29029,N_29184);
or U29207 (N_29207,N_29083,N_29018);
and U29208 (N_29208,N_29175,N_29017);
and U29209 (N_29209,N_29034,N_29041);
or U29210 (N_29210,N_29095,N_29052);
and U29211 (N_29211,N_29169,N_29192);
xor U29212 (N_29212,N_29180,N_29093);
nor U29213 (N_29213,N_29042,N_29146);
and U29214 (N_29214,N_29092,N_29033);
nor U29215 (N_29215,N_29178,N_29165);
nand U29216 (N_29216,N_29047,N_29051);
xor U29217 (N_29217,N_29069,N_29046);
or U29218 (N_29218,N_29056,N_29049);
and U29219 (N_29219,N_29191,N_29151);
nor U29220 (N_29220,N_29011,N_29127);
or U29221 (N_29221,N_29020,N_29189);
or U29222 (N_29222,N_29013,N_29043);
and U29223 (N_29223,N_29163,N_29140);
and U29224 (N_29224,N_29001,N_29195);
and U29225 (N_29225,N_29008,N_29123);
or U29226 (N_29226,N_29174,N_29155);
xnor U29227 (N_29227,N_29148,N_29177);
nand U29228 (N_29228,N_29153,N_29150);
xnor U29229 (N_29229,N_29118,N_29131);
or U29230 (N_29230,N_29039,N_29027);
and U29231 (N_29231,N_29094,N_29117);
nand U29232 (N_29232,N_29055,N_29136);
nor U29233 (N_29233,N_29138,N_29058);
nand U29234 (N_29234,N_29154,N_29139);
and U29235 (N_29235,N_29010,N_29164);
or U29236 (N_29236,N_29102,N_29084);
nand U29237 (N_29237,N_29103,N_29000);
nand U29238 (N_29238,N_29183,N_29048);
xor U29239 (N_29239,N_29182,N_29014);
or U29240 (N_29240,N_29079,N_29111);
nor U29241 (N_29241,N_29116,N_29040);
nand U29242 (N_29242,N_29145,N_29066);
nand U29243 (N_29243,N_29099,N_29016);
and U29244 (N_29244,N_29075,N_29112);
or U29245 (N_29245,N_29185,N_29002);
nor U29246 (N_29246,N_29085,N_29122);
and U29247 (N_29247,N_29170,N_29035);
and U29248 (N_29248,N_29104,N_29086);
or U29249 (N_29249,N_29050,N_29023);
or U29250 (N_29250,N_29141,N_29114);
nand U29251 (N_29251,N_29108,N_29024);
xnor U29252 (N_29252,N_29067,N_29072);
nor U29253 (N_29253,N_29063,N_29106);
and U29254 (N_29254,N_29162,N_29022);
or U29255 (N_29255,N_29147,N_29082);
nor U29256 (N_29256,N_29149,N_29133);
and U29257 (N_29257,N_29168,N_29097);
and U29258 (N_29258,N_29077,N_29009);
xor U29259 (N_29259,N_29126,N_29152);
and U29260 (N_29260,N_29143,N_29025);
nand U29261 (N_29261,N_29157,N_29030);
nor U29262 (N_29262,N_29088,N_29196);
nor U29263 (N_29263,N_29159,N_29091);
and U29264 (N_29264,N_29044,N_29045);
xnor U29265 (N_29265,N_29193,N_29003);
nor U29266 (N_29266,N_29124,N_29129);
nor U29267 (N_29267,N_29090,N_29032);
nor U29268 (N_29268,N_29021,N_29113);
and U29269 (N_29269,N_29119,N_29125);
nand U29270 (N_29270,N_29074,N_29061);
xor U29271 (N_29271,N_29199,N_29190);
xor U29272 (N_29272,N_29004,N_29076);
nor U29273 (N_29273,N_29062,N_29089);
nor U29274 (N_29274,N_29172,N_29121);
or U29275 (N_29275,N_29037,N_29181);
or U29276 (N_29276,N_29132,N_29142);
and U29277 (N_29277,N_29110,N_29098);
or U29278 (N_29278,N_29171,N_29173);
or U29279 (N_29279,N_29144,N_29060);
xnor U29280 (N_29280,N_29134,N_29158);
nand U29281 (N_29281,N_29078,N_29186);
nand U29282 (N_29282,N_29156,N_29115);
and U29283 (N_29283,N_29107,N_29105);
or U29284 (N_29284,N_29109,N_29176);
nor U29285 (N_29285,N_29019,N_29166);
and U29286 (N_29286,N_29036,N_29054);
xnor U29287 (N_29287,N_29161,N_29187);
nor U29288 (N_29288,N_29197,N_29005);
or U29289 (N_29289,N_29160,N_29080);
and U29290 (N_29290,N_29188,N_29120);
nand U29291 (N_29291,N_29087,N_29053);
or U29292 (N_29292,N_29096,N_29070);
and U29293 (N_29293,N_29130,N_29026);
nor U29294 (N_29294,N_29179,N_29038);
xnor U29295 (N_29295,N_29006,N_29064);
xnor U29296 (N_29296,N_29137,N_29198);
and U29297 (N_29297,N_29071,N_29073);
xnor U29298 (N_29298,N_29065,N_29167);
nor U29299 (N_29299,N_29081,N_29100);
or U29300 (N_29300,N_29058,N_29085);
or U29301 (N_29301,N_29186,N_29144);
and U29302 (N_29302,N_29171,N_29128);
nor U29303 (N_29303,N_29029,N_29088);
and U29304 (N_29304,N_29072,N_29165);
and U29305 (N_29305,N_29186,N_29152);
xor U29306 (N_29306,N_29032,N_29127);
or U29307 (N_29307,N_29184,N_29107);
xor U29308 (N_29308,N_29110,N_29167);
nand U29309 (N_29309,N_29067,N_29038);
and U29310 (N_29310,N_29098,N_29139);
and U29311 (N_29311,N_29131,N_29036);
xor U29312 (N_29312,N_29003,N_29018);
xnor U29313 (N_29313,N_29056,N_29053);
nor U29314 (N_29314,N_29115,N_29077);
xor U29315 (N_29315,N_29149,N_29051);
xor U29316 (N_29316,N_29195,N_29189);
or U29317 (N_29317,N_29184,N_29113);
or U29318 (N_29318,N_29169,N_29159);
nand U29319 (N_29319,N_29018,N_29151);
or U29320 (N_29320,N_29040,N_29140);
nand U29321 (N_29321,N_29144,N_29083);
nor U29322 (N_29322,N_29163,N_29176);
xnor U29323 (N_29323,N_29094,N_29041);
nor U29324 (N_29324,N_29033,N_29099);
nor U29325 (N_29325,N_29147,N_29035);
nor U29326 (N_29326,N_29130,N_29167);
or U29327 (N_29327,N_29189,N_29113);
xor U29328 (N_29328,N_29175,N_29130);
xnor U29329 (N_29329,N_29104,N_29017);
or U29330 (N_29330,N_29154,N_29059);
xnor U29331 (N_29331,N_29022,N_29024);
or U29332 (N_29332,N_29116,N_29167);
nor U29333 (N_29333,N_29169,N_29096);
xor U29334 (N_29334,N_29162,N_29077);
and U29335 (N_29335,N_29125,N_29039);
and U29336 (N_29336,N_29149,N_29143);
xor U29337 (N_29337,N_29176,N_29033);
and U29338 (N_29338,N_29139,N_29066);
nor U29339 (N_29339,N_29106,N_29195);
or U29340 (N_29340,N_29113,N_29050);
xor U29341 (N_29341,N_29179,N_29133);
nor U29342 (N_29342,N_29063,N_29126);
xor U29343 (N_29343,N_29023,N_29102);
xnor U29344 (N_29344,N_29141,N_29069);
xor U29345 (N_29345,N_29007,N_29189);
nor U29346 (N_29346,N_29169,N_29026);
and U29347 (N_29347,N_29015,N_29092);
xnor U29348 (N_29348,N_29180,N_29075);
and U29349 (N_29349,N_29062,N_29171);
nand U29350 (N_29350,N_29005,N_29162);
and U29351 (N_29351,N_29111,N_29124);
nand U29352 (N_29352,N_29083,N_29177);
and U29353 (N_29353,N_29151,N_29100);
nor U29354 (N_29354,N_29110,N_29149);
nor U29355 (N_29355,N_29033,N_29139);
or U29356 (N_29356,N_29109,N_29072);
xnor U29357 (N_29357,N_29097,N_29142);
nand U29358 (N_29358,N_29136,N_29172);
and U29359 (N_29359,N_29083,N_29127);
or U29360 (N_29360,N_29058,N_29073);
or U29361 (N_29361,N_29115,N_29065);
and U29362 (N_29362,N_29034,N_29077);
nand U29363 (N_29363,N_29114,N_29013);
nor U29364 (N_29364,N_29029,N_29081);
and U29365 (N_29365,N_29016,N_29059);
nor U29366 (N_29366,N_29167,N_29111);
or U29367 (N_29367,N_29118,N_29087);
or U29368 (N_29368,N_29095,N_29075);
and U29369 (N_29369,N_29128,N_29180);
nor U29370 (N_29370,N_29170,N_29175);
nor U29371 (N_29371,N_29153,N_29060);
or U29372 (N_29372,N_29177,N_29023);
nand U29373 (N_29373,N_29036,N_29039);
nor U29374 (N_29374,N_29068,N_29166);
and U29375 (N_29375,N_29061,N_29025);
nor U29376 (N_29376,N_29115,N_29124);
and U29377 (N_29377,N_29008,N_29184);
nand U29378 (N_29378,N_29175,N_29148);
nor U29379 (N_29379,N_29150,N_29063);
or U29380 (N_29380,N_29090,N_29078);
nor U29381 (N_29381,N_29175,N_29036);
nor U29382 (N_29382,N_29140,N_29015);
nand U29383 (N_29383,N_29047,N_29135);
xor U29384 (N_29384,N_29062,N_29196);
xor U29385 (N_29385,N_29025,N_29026);
or U29386 (N_29386,N_29108,N_29180);
or U29387 (N_29387,N_29062,N_29099);
nand U29388 (N_29388,N_29053,N_29009);
nand U29389 (N_29389,N_29145,N_29102);
nand U29390 (N_29390,N_29094,N_29070);
and U29391 (N_29391,N_29068,N_29027);
or U29392 (N_29392,N_29117,N_29097);
and U29393 (N_29393,N_29029,N_29181);
and U29394 (N_29394,N_29121,N_29022);
xor U29395 (N_29395,N_29018,N_29088);
and U29396 (N_29396,N_29063,N_29022);
and U29397 (N_29397,N_29102,N_29054);
nor U29398 (N_29398,N_29168,N_29030);
nand U29399 (N_29399,N_29154,N_29067);
and U29400 (N_29400,N_29228,N_29305);
nor U29401 (N_29401,N_29287,N_29306);
and U29402 (N_29402,N_29399,N_29240);
and U29403 (N_29403,N_29344,N_29249);
nor U29404 (N_29404,N_29216,N_29304);
xnor U29405 (N_29405,N_29372,N_29272);
xnor U29406 (N_29406,N_29261,N_29382);
nor U29407 (N_29407,N_29312,N_29346);
or U29408 (N_29408,N_29361,N_29268);
and U29409 (N_29409,N_29381,N_29289);
and U29410 (N_29410,N_29213,N_29284);
and U29411 (N_29411,N_29398,N_29222);
or U29412 (N_29412,N_29277,N_29219);
or U29413 (N_29413,N_29303,N_29229);
and U29414 (N_29414,N_29386,N_29243);
and U29415 (N_29415,N_29297,N_29334);
or U29416 (N_29416,N_29311,N_29373);
nand U29417 (N_29417,N_29244,N_29390);
nand U29418 (N_29418,N_29236,N_29211);
or U29419 (N_29419,N_29365,N_29375);
or U29420 (N_29420,N_29245,N_29354);
or U29421 (N_29421,N_29376,N_29337);
xor U29422 (N_29422,N_29387,N_29391);
nor U29423 (N_29423,N_29350,N_29340);
or U29424 (N_29424,N_29256,N_29274);
nand U29425 (N_29425,N_29320,N_29233);
nor U29426 (N_29426,N_29359,N_29273);
xor U29427 (N_29427,N_29258,N_29336);
nand U29428 (N_29428,N_29267,N_29347);
nor U29429 (N_29429,N_29253,N_29221);
nor U29430 (N_29430,N_29384,N_29369);
and U29431 (N_29431,N_29332,N_29246);
nand U29432 (N_29432,N_29328,N_29353);
or U29433 (N_29433,N_29278,N_29368);
or U29434 (N_29434,N_29371,N_29286);
nor U29435 (N_29435,N_29203,N_29237);
nor U29436 (N_29436,N_29263,N_29314);
and U29437 (N_29437,N_29325,N_29301);
or U29438 (N_29438,N_29271,N_29259);
nand U29439 (N_29439,N_29308,N_29232);
nor U29440 (N_29440,N_29374,N_29338);
and U29441 (N_29441,N_29318,N_29255);
nor U29442 (N_29442,N_29231,N_29342);
nor U29443 (N_29443,N_29279,N_29299);
xor U29444 (N_29444,N_29380,N_29358);
or U29445 (N_29445,N_29357,N_29331);
nand U29446 (N_29446,N_29335,N_29225);
or U29447 (N_29447,N_29351,N_29257);
and U29448 (N_29448,N_29383,N_29247);
xor U29449 (N_29449,N_29241,N_29295);
and U29450 (N_29450,N_29205,N_29223);
nor U29451 (N_29451,N_29300,N_29282);
or U29452 (N_29452,N_29397,N_29339);
and U29453 (N_29453,N_29393,N_29360);
or U29454 (N_29454,N_29234,N_29379);
nand U29455 (N_29455,N_29262,N_29204);
xor U29456 (N_29456,N_29264,N_29209);
nand U29457 (N_29457,N_29227,N_29315);
nor U29458 (N_29458,N_29319,N_29202);
and U29459 (N_29459,N_29329,N_29296);
xnor U29460 (N_29460,N_29355,N_29333);
xnor U29461 (N_29461,N_29276,N_29389);
and U29462 (N_29462,N_29280,N_29298);
and U29463 (N_29463,N_29370,N_29214);
nand U29464 (N_29464,N_29341,N_29201);
or U29465 (N_29465,N_29254,N_29285);
or U29466 (N_29466,N_29349,N_29266);
and U29467 (N_29467,N_29352,N_29293);
or U29468 (N_29468,N_29394,N_29330);
nand U29469 (N_29469,N_29395,N_29200);
or U29470 (N_29470,N_29269,N_29367);
xnor U29471 (N_29471,N_29238,N_29322);
nand U29472 (N_29472,N_29307,N_29388);
and U29473 (N_29473,N_29392,N_29215);
and U29474 (N_29474,N_29378,N_29302);
and U29475 (N_29475,N_29281,N_29324);
and U29476 (N_29476,N_29260,N_29309);
nor U29477 (N_29477,N_29294,N_29317);
and U29478 (N_29478,N_29265,N_29363);
or U29479 (N_29479,N_29345,N_29208);
or U29480 (N_29480,N_29230,N_29226);
and U29481 (N_29481,N_29291,N_29366);
xnor U29482 (N_29482,N_29356,N_29210);
xnor U29483 (N_29483,N_29310,N_29313);
nand U29484 (N_29484,N_29242,N_29239);
or U29485 (N_29485,N_29326,N_29327);
and U29486 (N_29486,N_29364,N_29248);
nor U29487 (N_29487,N_29348,N_29385);
and U29488 (N_29488,N_29220,N_29323);
or U29489 (N_29489,N_29212,N_29343);
nor U29490 (N_29490,N_29362,N_29235);
and U29491 (N_29491,N_29316,N_29251);
or U29492 (N_29492,N_29206,N_29288);
nor U29493 (N_29493,N_29250,N_29218);
nand U29494 (N_29494,N_29207,N_29290);
nor U29495 (N_29495,N_29321,N_29224);
or U29496 (N_29496,N_29283,N_29396);
and U29497 (N_29497,N_29270,N_29275);
nand U29498 (N_29498,N_29292,N_29377);
nand U29499 (N_29499,N_29252,N_29217);
and U29500 (N_29500,N_29305,N_29266);
nor U29501 (N_29501,N_29320,N_29329);
xor U29502 (N_29502,N_29324,N_29250);
nor U29503 (N_29503,N_29345,N_29227);
xor U29504 (N_29504,N_29255,N_29299);
or U29505 (N_29505,N_29222,N_29214);
xor U29506 (N_29506,N_29210,N_29263);
nor U29507 (N_29507,N_29283,N_29297);
or U29508 (N_29508,N_29306,N_29375);
nand U29509 (N_29509,N_29316,N_29242);
nand U29510 (N_29510,N_29242,N_29331);
and U29511 (N_29511,N_29347,N_29317);
xor U29512 (N_29512,N_29286,N_29223);
and U29513 (N_29513,N_29363,N_29294);
nor U29514 (N_29514,N_29240,N_29213);
xor U29515 (N_29515,N_29243,N_29349);
xor U29516 (N_29516,N_29288,N_29332);
or U29517 (N_29517,N_29252,N_29319);
nand U29518 (N_29518,N_29386,N_29359);
nand U29519 (N_29519,N_29228,N_29327);
and U29520 (N_29520,N_29220,N_29264);
xnor U29521 (N_29521,N_29285,N_29222);
or U29522 (N_29522,N_29331,N_29247);
or U29523 (N_29523,N_29395,N_29250);
xnor U29524 (N_29524,N_29368,N_29207);
xor U29525 (N_29525,N_29229,N_29268);
nand U29526 (N_29526,N_29302,N_29355);
nor U29527 (N_29527,N_29318,N_29344);
xor U29528 (N_29528,N_29224,N_29204);
xor U29529 (N_29529,N_29268,N_29262);
or U29530 (N_29530,N_29272,N_29228);
nor U29531 (N_29531,N_29352,N_29358);
nor U29532 (N_29532,N_29244,N_29352);
nor U29533 (N_29533,N_29297,N_29302);
and U29534 (N_29534,N_29237,N_29384);
xor U29535 (N_29535,N_29352,N_29348);
nor U29536 (N_29536,N_29259,N_29269);
or U29537 (N_29537,N_29338,N_29357);
nor U29538 (N_29538,N_29321,N_29206);
xnor U29539 (N_29539,N_29245,N_29220);
and U29540 (N_29540,N_29305,N_29379);
nor U29541 (N_29541,N_29324,N_29265);
nand U29542 (N_29542,N_29342,N_29388);
xnor U29543 (N_29543,N_29375,N_29316);
nand U29544 (N_29544,N_29280,N_29300);
and U29545 (N_29545,N_29355,N_29360);
nor U29546 (N_29546,N_29345,N_29363);
or U29547 (N_29547,N_29320,N_29267);
xnor U29548 (N_29548,N_29308,N_29277);
or U29549 (N_29549,N_29339,N_29247);
and U29550 (N_29550,N_29380,N_29299);
nor U29551 (N_29551,N_29356,N_29307);
nand U29552 (N_29552,N_29264,N_29321);
and U29553 (N_29553,N_29389,N_29249);
and U29554 (N_29554,N_29361,N_29285);
nand U29555 (N_29555,N_29261,N_29361);
nand U29556 (N_29556,N_29376,N_29250);
nand U29557 (N_29557,N_29230,N_29369);
or U29558 (N_29558,N_29339,N_29252);
xnor U29559 (N_29559,N_29204,N_29322);
nand U29560 (N_29560,N_29329,N_29279);
or U29561 (N_29561,N_29298,N_29335);
nor U29562 (N_29562,N_29346,N_29260);
and U29563 (N_29563,N_29380,N_29239);
and U29564 (N_29564,N_29233,N_29361);
or U29565 (N_29565,N_29295,N_29316);
nor U29566 (N_29566,N_29352,N_29368);
nor U29567 (N_29567,N_29204,N_29351);
nor U29568 (N_29568,N_29254,N_29319);
nand U29569 (N_29569,N_29243,N_29373);
nor U29570 (N_29570,N_29301,N_29252);
xnor U29571 (N_29571,N_29365,N_29246);
nor U29572 (N_29572,N_29208,N_29373);
and U29573 (N_29573,N_29369,N_29390);
xor U29574 (N_29574,N_29212,N_29313);
or U29575 (N_29575,N_29334,N_29351);
and U29576 (N_29576,N_29279,N_29264);
xor U29577 (N_29577,N_29312,N_29255);
xor U29578 (N_29578,N_29272,N_29285);
xor U29579 (N_29579,N_29310,N_29275);
nand U29580 (N_29580,N_29320,N_29375);
nor U29581 (N_29581,N_29208,N_29335);
xor U29582 (N_29582,N_29344,N_29365);
and U29583 (N_29583,N_29389,N_29277);
xor U29584 (N_29584,N_29321,N_29389);
nand U29585 (N_29585,N_29327,N_29202);
nand U29586 (N_29586,N_29308,N_29207);
nor U29587 (N_29587,N_29240,N_29357);
xor U29588 (N_29588,N_29265,N_29349);
nor U29589 (N_29589,N_29325,N_29316);
and U29590 (N_29590,N_29294,N_29286);
or U29591 (N_29591,N_29206,N_29265);
xor U29592 (N_29592,N_29255,N_29206);
and U29593 (N_29593,N_29281,N_29285);
and U29594 (N_29594,N_29200,N_29264);
xnor U29595 (N_29595,N_29278,N_29247);
nor U29596 (N_29596,N_29363,N_29341);
nand U29597 (N_29597,N_29387,N_29315);
nand U29598 (N_29598,N_29305,N_29388);
or U29599 (N_29599,N_29322,N_29209);
or U29600 (N_29600,N_29470,N_29488);
nor U29601 (N_29601,N_29409,N_29481);
nor U29602 (N_29602,N_29512,N_29581);
xor U29603 (N_29603,N_29454,N_29477);
nor U29604 (N_29604,N_29460,N_29572);
nand U29605 (N_29605,N_29569,N_29429);
nor U29606 (N_29606,N_29453,N_29549);
xor U29607 (N_29607,N_29515,N_29412);
or U29608 (N_29608,N_29514,N_29579);
and U29609 (N_29609,N_29585,N_29543);
xor U29610 (N_29610,N_29592,N_29523);
or U29611 (N_29611,N_29492,N_29583);
xnor U29612 (N_29612,N_29506,N_29446);
nor U29613 (N_29613,N_29561,N_29433);
nor U29614 (N_29614,N_29465,N_29552);
nor U29615 (N_29615,N_29505,N_29513);
or U29616 (N_29616,N_29559,N_29530);
nor U29617 (N_29617,N_29498,N_29595);
nor U29618 (N_29618,N_29463,N_29575);
nor U29619 (N_29619,N_29430,N_29435);
xnor U29620 (N_29620,N_29422,N_29554);
and U29621 (N_29621,N_29482,N_29527);
or U29622 (N_29622,N_29442,N_29560);
or U29623 (N_29623,N_29594,N_29487);
and U29624 (N_29624,N_29582,N_29591);
and U29625 (N_29625,N_29468,N_29431);
nand U29626 (N_29626,N_29538,N_29516);
nor U29627 (N_29627,N_29474,N_29472);
xnor U29628 (N_29628,N_29455,N_29478);
and U29629 (N_29629,N_29593,N_29459);
or U29630 (N_29630,N_29440,N_29489);
nor U29631 (N_29631,N_29526,N_29562);
nand U29632 (N_29632,N_29504,N_29443);
xnor U29633 (N_29633,N_29404,N_29417);
and U29634 (N_29634,N_29507,N_29425);
or U29635 (N_29635,N_29508,N_29547);
nand U29636 (N_29636,N_29565,N_29419);
or U29637 (N_29637,N_29408,N_29449);
nand U29638 (N_29638,N_29545,N_29503);
or U29639 (N_29639,N_29589,N_29401);
nor U29640 (N_29640,N_29556,N_29416);
nand U29641 (N_29641,N_29520,N_29415);
and U29642 (N_29642,N_29590,N_29518);
nor U29643 (N_29643,N_29580,N_29546);
or U29644 (N_29644,N_29540,N_29548);
or U29645 (N_29645,N_29586,N_29588);
and U29646 (N_29646,N_29536,N_29439);
nor U29647 (N_29647,N_29434,N_29500);
xnor U29648 (N_29648,N_29567,N_29400);
xnor U29649 (N_29649,N_29421,N_29457);
nor U29650 (N_29650,N_29510,N_29406);
nor U29651 (N_29651,N_29564,N_29568);
xor U29652 (N_29652,N_29448,N_29517);
xnor U29653 (N_29653,N_29598,N_29497);
or U29654 (N_29654,N_29420,N_29410);
xnor U29655 (N_29655,N_29553,N_29413);
and U29656 (N_29656,N_29471,N_29432);
nand U29657 (N_29657,N_29466,N_29578);
or U29658 (N_29658,N_29550,N_29555);
nand U29659 (N_29659,N_29524,N_29424);
or U29660 (N_29660,N_29402,N_29494);
nand U29661 (N_29661,N_29576,N_29414);
nor U29662 (N_29662,N_29519,N_29509);
or U29663 (N_29663,N_29462,N_29456);
xor U29664 (N_29664,N_29563,N_29437);
or U29665 (N_29665,N_29473,N_29537);
and U29666 (N_29666,N_29441,N_29438);
nand U29667 (N_29667,N_29491,N_29485);
and U29668 (N_29668,N_29480,N_29447);
nor U29669 (N_29669,N_29428,N_29461);
or U29670 (N_29670,N_29597,N_29534);
nand U29671 (N_29671,N_29493,N_29532);
xor U29672 (N_29672,N_29528,N_29451);
xnor U29673 (N_29673,N_29423,N_29436);
and U29674 (N_29674,N_29502,N_29570);
xnor U29675 (N_29675,N_29476,N_29501);
and U29676 (N_29676,N_29484,N_29587);
nand U29677 (N_29677,N_29574,N_29596);
or U29678 (N_29678,N_29486,N_29426);
nor U29679 (N_29679,N_29557,N_29475);
and U29680 (N_29680,N_29511,N_29467);
xor U29681 (N_29681,N_29411,N_29535);
nor U29682 (N_29682,N_29483,N_29599);
xor U29683 (N_29683,N_29458,N_29539);
xor U29684 (N_29684,N_29496,N_29544);
nand U29685 (N_29685,N_29450,N_29525);
and U29686 (N_29686,N_29495,N_29577);
or U29687 (N_29687,N_29551,N_29418);
or U29688 (N_29688,N_29573,N_29427);
xor U29689 (N_29689,N_29584,N_29479);
xor U29690 (N_29690,N_29490,N_29407);
nor U29691 (N_29691,N_29541,N_29571);
and U29692 (N_29692,N_29531,N_29445);
nand U29693 (N_29693,N_29533,N_29403);
and U29694 (N_29694,N_29469,N_29542);
and U29695 (N_29695,N_29444,N_29558);
and U29696 (N_29696,N_29405,N_29452);
and U29697 (N_29697,N_29499,N_29529);
nor U29698 (N_29698,N_29566,N_29521);
xor U29699 (N_29699,N_29522,N_29464);
xor U29700 (N_29700,N_29468,N_29404);
xor U29701 (N_29701,N_29445,N_29562);
xor U29702 (N_29702,N_29594,N_29426);
nand U29703 (N_29703,N_29500,N_29468);
nand U29704 (N_29704,N_29421,N_29437);
nor U29705 (N_29705,N_29489,N_29402);
xor U29706 (N_29706,N_29556,N_29519);
xnor U29707 (N_29707,N_29578,N_29434);
xor U29708 (N_29708,N_29480,N_29438);
or U29709 (N_29709,N_29458,N_29575);
or U29710 (N_29710,N_29577,N_29440);
or U29711 (N_29711,N_29403,N_29550);
and U29712 (N_29712,N_29480,N_29510);
nor U29713 (N_29713,N_29599,N_29520);
xor U29714 (N_29714,N_29489,N_29508);
and U29715 (N_29715,N_29576,N_29415);
nor U29716 (N_29716,N_29429,N_29535);
nand U29717 (N_29717,N_29490,N_29579);
nor U29718 (N_29718,N_29577,N_29425);
or U29719 (N_29719,N_29597,N_29400);
nand U29720 (N_29720,N_29459,N_29472);
nand U29721 (N_29721,N_29436,N_29468);
nor U29722 (N_29722,N_29414,N_29588);
or U29723 (N_29723,N_29454,N_29404);
and U29724 (N_29724,N_29579,N_29483);
and U29725 (N_29725,N_29409,N_29442);
nor U29726 (N_29726,N_29499,N_29427);
xnor U29727 (N_29727,N_29517,N_29418);
nand U29728 (N_29728,N_29556,N_29483);
and U29729 (N_29729,N_29440,N_29521);
and U29730 (N_29730,N_29501,N_29511);
or U29731 (N_29731,N_29435,N_29417);
and U29732 (N_29732,N_29458,N_29457);
or U29733 (N_29733,N_29507,N_29518);
and U29734 (N_29734,N_29462,N_29415);
xor U29735 (N_29735,N_29411,N_29414);
and U29736 (N_29736,N_29437,N_29574);
xor U29737 (N_29737,N_29425,N_29508);
and U29738 (N_29738,N_29543,N_29470);
or U29739 (N_29739,N_29512,N_29457);
xnor U29740 (N_29740,N_29534,N_29416);
or U29741 (N_29741,N_29530,N_29497);
nor U29742 (N_29742,N_29431,N_29540);
or U29743 (N_29743,N_29563,N_29551);
and U29744 (N_29744,N_29513,N_29580);
nor U29745 (N_29745,N_29432,N_29405);
nand U29746 (N_29746,N_29452,N_29535);
and U29747 (N_29747,N_29465,N_29447);
xnor U29748 (N_29748,N_29590,N_29407);
nand U29749 (N_29749,N_29505,N_29473);
or U29750 (N_29750,N_29405,N_29556);
nor U29751 (N_29751,N_29480,N_29551);
or U29752 (N_29752,N_29435,N_29458);
and U29753 (N_29753,N_29595,N_29471);
or U29754 (N_29754,N_29542,N_29483);
xor U29755 (N_29755,N_29411,N_29483);
nand U29756 (N_29756,N_29499,N_29465);
or U29757 (N_29757,N_29478,N_29583);
nand U29758 (N_29758,N_29441,N_29550);
nor U29759 (N_29759,N_29424,N_29589);
xor U29760 (N_29760,N_29524,N_29467);
or U29761 (N_29761,N_29522,N_29513);
or U29762 (N_29762,N_29415,N_29581);
nor U29763 (N_29763,N_29563,N_29558);
xor U29764 (N_29764,N_29468,N_29506);
and U29765 (N_29765,N_29508,N_29483);
and U29766 (N_29766,N_29564,N_29487);
nand U29767 (N_29767,N_29517,N_29472);
or U29768 (N_29768,N_29409,N_29598);
or U29769 (N_29769,N_29433,N_29589);
nor U29770 (N_29770,N_29438,N_29561);
and U29771 (N_29771,N_29438,N_29464);
nand U29772 (N_29772,N_29502,N_29574);
nor U29773 (N_29773,N_29411,N_29511);
xor U29774 (N_29774,N_29489,N_29507);
and U29775 (N_29775,N_29521,N_29423);
xnor U29776 (N_29776,N_29450,N_29425);
nand U29777 (N_29777,N_29527,N_29578);
and U29778 (N_29778,N_29506,N_29408);
xnor U29779 (N_29779,N_29455,N_29467);
or U29780 (N_29780,N_29419,N_29582);
xnor U29781 (N_29781,N_29532,N_29474);
xor U29782 (N_29782,N_29436,N_29471);
nor U29783 (N_29783,N_29574,N_29576);
nand U29784 (N_29784,N_29594,N_29412);
or U29785 (N_29785,N_29469,N_29504);
nand U29786 (N_29786,N_29569,N_29547);
nand U29787 (N_29787,N_29492,N_29567);
or U29788 (N_29788,N_29513,N_29573);
nand U29789 (N_29789,N_29420,N_29487);
or U29790 (N_29790,N_29485,N_29542);
or U29791 (N_29791,N_29485,N_29504);
xnor U29792 (N_29792,N_29586,N_29559);
xnor U29793 (N_29793,N_29592,N_29418);
or U29794 (N_29794,N_29534,N_29525);
nand U29795 (N_29795,N_29524,N_29565);
nand U29796 (N_29796,N_29404,N_29556);
nand U29797 (N_29797,N_29408,N_29509);
nor U29798 (N_29798,N_29542,N_29418);
and U29799 (N_29799,N_29571,N_29445);
and U29800 (N_29800,N_29763,N_29708);
nand U29801 (N_29801,N_29718,N_29620);
and U29802 (N_29802,N_29787,N_29627);
nand U29803 (N_29803,N_29633,N_29688);
nor U29804 (N_29804,N_29675,N_29640);
nor U29805 (N_29805,N_29734,N_29723);
xnor U29806 (N_29806,N_29741,N_29609);
or U29807 (N_29807,N_29619,N_29656);
or U29808 (N_29808,N_29654,N_29716);
nand U29809 (N_29809,N_29754,N_29702);
or U29810 (N_29810,N_29695,N_29750);
nor U29811 (N_29811,N_29694,N_29696);
nand U29812 (N_29812,N_29612,N_29673);
and U29813 (N_29813,N_29624,N_29739);
or U29814 (N_29814,N_29605,N_29717);
or U29815 (N_29815,N_29626,N_29663);
nand U29816 (N_29816,N_29653,N_29730);
nor U29817 (N_29817,N_29672,N_29700);
xnor U29818 (N_29818,N_29744,N_29639);
and U29819 (N_29819,N_29759,N_29601);
nor U29820 (N_29820,N_29731,N_29666);
nand U29821 (N_29821,N_29707,N_29768);
nor U29822 (N_29822,N_29749,N_29692);
nor U29823 (N_29823,N_29751,N_29722);
nand U29824 (N_29824,N_29714,N_29776);
nand U29825 (N_29825,N_29642,N_29685);
and U29826 (N_29826,N_29784,N_29799);
xor U29827 (N_29827,N_29625,N_29761);
and U29828 (N_29828,N_29764,N_29711);
nor U29829 (N_29829,N_29747,N_29630);
and U29830 (N_29830,N_29636,N_29681);
and U29831 (N_29831,N_29703,N_29745);
and U29832 (N_29832,N_29713,N_29766);
nand U29833 (N_29833,N_29606,N_29682);
or U29834 (N_29834,N_29705,N_29769);
or U29835 (N_29835,N_29641,N_29698);
or U29836 (N_29836,N_29638,N_29680);
or U29837 (N_29837,N_29758,N_29760);
nor U29838 (N_29838,N_29645,N_29632);
nor U29839 (N_29839,N_29660,N_29634);
nor U29840 (N_29840,N_29782,N_29646);
nand U29841 (N_29841,N_29773,N_29793);
xnor U29842 (N_29842,N_29797,N_29756);
nand U29843 (N_29843,N_29603,N_29622);
nand U29844 (N_29844,N_29662,N_29777);
nand U29845 (N_29845,N_29616,N_29795);
nor U29846 (N_29846,N_29790,N_29778);
nand U29847 (N_29847,N_29712,N_29725);
and U29848 (N_29848,N_29623,N_29610);
or U29849 (N_29849,N_29665,N_29737);
nor U29850 (N_29850,N_29691,N_29774);
nand U29851 (N_29851,N_29657,N_29785);
nand U29852 (N_29852,N_29637,N_29789);
nand U29853 (N_29853,N_29686,N_29792);
nand U29854 (N_29854,N_29614,N_29798);
nand U29855 (N_29855,N_29621,N_29659);
nand U29856 (N_29856,N_29693,N_29742);
nor U29857 (N_29857,N_29752,N_29733);
or U29858 (N_29858,N_29677,N_29724);
xor U29859 (N_29859,N_29600,N_29671);
or U29860 (N_29860,N_29736,N_29613);
nand U29861 (N_29861,N_29780,N_29618);
xnor U29862 (N_29862,N_29649,N_29781);
nand U29863 (N_29863,N_29631,N_29729);
and U29864 (N_29864,N_29788,N_29783);
nand U29865 (N_29865,N_29720,N_29755);
and U29866 (N_29866,N_29650,N_29699);
nor U29867 (N_29867,N_29683,N_29779);
nor U29868 (N_29868,N_29628,N_29772);
nor U29869 (N_29869,N_29629,N_29726);
xnor U29870 (N_29870,N_29710,N_29644);
nor U29871 (N_29871,N_29794,N_29669);
xor U29872 (N_29872,N_29753,N_29706);
and U29873 (N_29873,N_29732,N_29604);
xnor U29874 (N_29874,N_29678,N_29635);
and U29875 (N_29875,N_29684,N_29775);
nor U29876 (N_29876,N_29658,N_29715);
or U29877 (N_29877,N_29602,N_29740);
or U29878 (N_29878,N_29608,N_29687);
nand U29879 (N_29879,N_29719,N_29704);
xnor U29880 (N_29880,N_29651,N_29615);
nand U29881 (N_29881,N_29679,N_29786);
and U29882 (N_29882,N_29690,N_29727);
or U29883 (N_29883,N_29767,N_29617);
xnor U29884 (N_29884,N_29689,N_29748);
nand U29885 (N_29885,N_29721,N_29607);
or U29886 (N_29886,N_29796,N_29738);
and U29887 (N_29887,N_29674,N_29661);
nor U29888 (N_29888,N_29647,N_29743);
and U29889 (N_29889,N_29655,N_29676);
nor U29890 (N_29890,N_29667,N_29668);
nand U29891 (N_29891,N_29643,N_29611);
or U29892 (N_29892,N_29701,N_29771);
or U29893 (N_29893,N_29664,N_29757);
xor U29894 (N_29894,N_29648,N_29670);
xor U29895 (N_29895,N_29652,N_29735);
or U29896 (N_29896,N_29791,N_29697);
and U29897 (N_29897,N_29762,N_29746);
nand U29898 (N_29898,N_29770,N_29709);
or U29899 (N_29899,N_29728,N_29765);
or U29900 (N_29900,N_29670,N_29683);
nand U29901 (N_29901,N_29749,N_29744);
nand U29902 (N_29902,N_29693,N_29703);
or U29903 (N_29903,N_29690,N_29782);
nor U29904 (N_29904,N_29651,N_29697);
xnor U29905 (N_29905,N_29719,N_29624);
nor U29906 (N_29906,N_29752,N_29750);
nand U29907 (N_29907,N_29622,N_29645);
nand U29908 (N_29908,N_29776,N_29640);
and U29909 (N_29909,N_29745,N_29761);
and U29910 (N_29910,N_29789,N_29652);
or U29911 (N_29911,N_29757,N_29609);
nand U29912 (N_29912,N_29782,N_29707);
nand U29913 (N_29913,N_29620,N_29683);
nand U29914 (N_29914,N_29632,N_29658);
nand U29915 (N_29915,N_29645,N_29753);
or U29916 (N_29916,N_29651,N_29731);
nor U29917 (N_29917,N_29785,N_29722);
xnor U29918 (N_29918,N_29736,N_29645);
and U29919 (N_29919,N_29696,N_29659);
and U29920 (N_29920,N_29795,N_29725);
or U29921 (N_29921,N_29754,N_29657);
nand U29922 (N_29922,N_29786,N_29609);
xnor U29923 (N_29923,N_29751,N_29656);
and U29924 (N_29924,N_29794,N_29749);
nor U29925 (N_29925,N_29611,N_29667);
and U29926 (N_29926,N_29615,N_29789);
or U29927 (N_29927,N_29749,N_29782);
and U29928 (N_29928,N_29664,N_29659);
and U29929 (N_29929,N_29610,N_29775);
nor U29930 (N_29930,N_29720,N_29798);
nand U29931 (N_29931,N_29702,N_29764);
xor U29932 (N_29932,N_29783,N_29700);
nor U29933 (N_29933,N_29735,N_29708);
or U29934 (N_29934,N_29766,N_29681);
or U29935 (N_29935,N_29692,N_29748);
nand U29936 (N_29936,N_29787,N_29722);
nor U29937 (N_29937,N_29697,N_29603);
and U29938 (N_29938,N_29785,N_29617);
xnor U29939 (N_29939,N_29793,N_29769);
and U29940 (N_29940,N_29667,N_29722);
nand U29941 (N_29941,N_29684,N_29699);
xnor U29942 (N_29942,N_29650,N_29658);
nand U29943 (N_29943,N_29787,N_29657);
or U29944 (N_29944,N_29601,N_29604);
or U29945 (N_29945,N_29771,N_29652);
or U29946 (N_29946,N_29640,N_29752);
and U29947 (N_29947,N_29691,N_29712);
nor U29948 (N_29948,N_29696,N_29627);
xor U29949 (N_29949,N_29716,N_29793);
and U29950 (N_29950,N_29607,N_29711);
xor U29951 (N_29951,N_29777,N_29621);
nand U29952 (N_29952,N_29792,N_29769);
and U29953 (N_29953,N_29647,N_29681);
nand U29954 (N_29954,N_29681,N_29646);
or U29955 (N_29955,N_29611,N_29712);
nand U29956 (N_29956,N_29734,N_29780);
or U29957 (N_29957,N_29652,N_29698);
nor U29958 (N_29958,N_29697,N_29633);
or U29959 (N_29959,N_29628,N_29768);
nand U29960 (N_29960,N_29651,N_29616);
nor U29961 (N_29961,N_29692,N_29741);
and U29962 (N_29962,N_29642,N_29606);
nor U29963 (N_29963,N_29691,N_29696);
or U29964 (N_29964,N_29716,N_29754);
and U29965 (N_29965,N_29775,N_29757);
xor U29966 (N_29966,N_29717,N_29693);
nand U29967 (N_29967,N_29792,N_29607);
nand U29968 (N_29968,N_29714,N_29724);
xor U29969 (N_29969,N_29771,N_29618);
and U29970 (N_29970,N_29766,N_29721);
xor U29971 (N_29971,N_29635,N_29619);
nor U29972 (N_29972,N_29600,N_29771);
nor U29973 (N_29973,N_29789,N_29766);
xor U29974 (N_29974,N_29601,N_29681);
or U29975 (N_29975,N_29704,N_29670);
or U29976 (N_29976,N_29762,N_29678);
nor U29977 (N_29977,N_29645,N_29764);
nor U29978 (N_29978,N_29742,N_29634);
or U29979 (N_29979,N_29631,N_29673);
and U29980 (N_29980,N_29792,N_29673);
or U29981 (N_29981,N_29771,N_29703);
xnor U29982 (N_29982,N_29752,N_29742);
and U29983 (N_29983,N_29674,N_29780);
nand U29984 (N_29984,N_29676,N_29732);
and U29985 (N_29985,N_29618,N_29663);
xnor U29986 (N_29986,N_29685,N_29660);
xnor U29987 (N_29987,N_29616,N_29645);
xnor U29988 (N_29988,N_29706,N_29689);
and U29989 (N_29989,N_29623,N_29727);
or U29990 (N_29990,N_29668,N_29719);
nor U29991 (N_29991,N_29781,N_29691);
or U29992 (N_29992,N_29671,N_29690);
nor U29993 (N_29993,N_29678,N_29766);
nand U29994 (N_29994,N_29630,N_29737);
or U29995 (N_29995,N_29792,N_29705);
nand U29996 (N_29996,N_29651,N_29745);
xor U29997 (N_29997,N_29615,N_29755);
and U29998 (N_29998,N_29742,N_29662);
and U29999 (N_29999,N_29635,N_29782);
or UO_0 (O_0,N_29851,N_29801);
xnor UO_1 (O_1,N_29973,N_29982);
xnor UO_2 (O_2,N_29929,N_29959);
nor UO_3 (O_3,N_29892,N_29930);
and UO_4 (O_4,N_29800,N_29918);
nand UO_5 (O_5,N_29886,N_29839);
or UO_6 (O_6,N_29809,N_29946);
or UO_7 (O_7,N_29951,N_29907);
nand UO_8 (O_8,N_29945,N_29895);
or UO_9 (O_9,N_29854,N_29825);
nand UO_10 (O_10,N_29874,N_29891);
nand UO_11 (O_11,N_29916,N_29957);
or UO_12 (O_12,N_29862,N_29820);
or UO_13 (O_13,N_29981,N_29901);
or UO_14 (O_14,N_29865,N_29936);
and UO_15 (O_15,N_29988,N_29952);
nor UO_16 (O_16,N_29881,N_29822);
xnor UO_17 (O_17,N_29914,N_29921);
and UO_18 (O_18,N_29961,N_29828);
or UO_19 (O_19,N_29938,N_29884);
nor UO_20 (O_20,N_29850,N_29919);
nand UO_21 (O_21,N_29909,N_29831);
nand UO_22 (O_22,N_29812,N_29897);
or UO_23 (O_23,N_29856,N_29913);
xor UO_24 (O_24,N_29910,N_29880);
xnor UO_25 (O_25,N_29821,N_29966);
or UO_26 (O_26,N_29934,N_29948);
nor UO_27 (O_27,N_29836,N_29958);
and UO_28 (O_28,N_29908,N_29894);
nor UO_29 (O_29,N_29816,N_29882);
or UO_30 (O_30,N_29827,N_29920);
and UO_31 (O_31,N_29872,N_29964);
or UO_32 (O_32,N_29833,N_29943);
or UO_33 (O_33,N_29853,N_29876);
or UO_34 (O_34,N_29819,N_29927);
or UO_35 (O_35,N_29896,N_29912);
nor UO_36 (O_36,N_29858,N_29842);
or UO_37 (O_37,N_29994,N_29879);
nand UO_38 (O_38,N_29904,N_29885);
nor UO_39 (O_39,N_29954,N_29911);
nor UO_40 (O_40,N_29840,N_29848);
nor UO_41 (O_41,N_29995,N_29989);
nand UO_42 (O_42,N_29944,N_29997);
nand UO_43 (O_43,N_29939,N_29941);
nor UO_44 (O_44,N_29998,N_29846);
and UO_45 (O_45,N_29926,N_29838);
xor UO_46 (O_46,N_29814,N_29875);
xnor UO_47 (O_47,N_29937,N_29861);
nor UO_48 (O_48,N_29977,N_29815);
nand UO_49 (O_49,N_29843,N_29857);
or UO_50 (O_50,N_29869,N_29983);
or UO_51 (O_51,N_29986,N_29902);
nor UO_52 (O_52,N_29949,N_29855);
nand UO_53 (O_53,N_29878,N_29834);
nand UO_54 (O_54,N_29950,N_29808);
nor UO_55 (O_55,N_29893,N_29978);
xor UO_56 (O_56,N_29942,N_29844);
nand UO_57 (O_57,N_29837,N_29987);
xor UO_58 (O_58,N_29922,N_29849);
nand UO_59 (O_59,N_29889,N_29805);
nand UO_60 (O_60,N_29818,N_29847);
xor UO_61 (O_61,N_29873,N_29992);
and UO_62 (O_62,N_29993,N_29947);
nor UO_63 (O_63,N_29917,N_29860);
xnor UO_64 (O_64,N_29980,N_29804);
nor UO_65 (O_65,N_29979,N_29866);
nand UO_66 (O_66,N_29877,N_29969);
xnor UO_67 (O_67,N_29975,N_29962);
nand UO_68 (O_68,N_29830,N_29803);
xor UO_69 (O_69,N_29806,N_29990);
or UO_70 (O_70,N_29841,N_29924);
xnor UO_71 (O_71,N_29953,N_29906);
nand UO_72 (O_72,N_29972,N_29940);
xnor UO_73 (O_73,N_29932,N_29824);
nand UO_74 (O_74,N_29999,N_29845);
or UO_75 (O_75,N_29963,N_29915);
and UO_76 (O_76,N_29991,N_29903);
and UO_77 (O_77,N_29933,N_29817);
or UO_78 (O_78,N_29900,N_29890);
or UO_79 (O_79,N_29887,N_29955);
nand UO_80 (O_80,N_29870,N_29965);
or UO_81 (O_81,N_29883,N_29863);
or UO_82 (O_82,N_29826,N_29832);
and UO_83 (O_83,N_29871,N_29835);
xor UO_84 (O_84,N_29984,N_29935);
nor UO_85 (O_85,N_29807,N_29899);
xor UO_86 (O_86,N_29970,N_29923);
nor UO_87 (O_87,N_29985,N_29898);
and UO_88 (O_88,N_29956,N_29925);
xnor UO_89 (O_89,N_29867,N_29996);
nand UO_90 (O_90,N_29968,N_29811);
nor UO_91 (O_91,N_29813,N_29859);
nand UO_92 (O_92,N_29928,N_29905);
xnor UO_93 (O_93,N_29810,N_29864);
and UO_94 (O_94,N_29976,N_29974);
nand UO_95 (O_95,N_29802,N_29931);
nand UO_96 (O_96,N_29829,N_29868);
nand UO_97 (O_97,N_29888,N_29823);
nor UO_98 (O_98,N_29960,N_29967);
or UO_99 (O_99,N_29852,N_29971);
or UO_100 (O_100,N_29991,N_29956);
nand UO_101 (O_101,N_29992,N_29946);
and UO_102 (O_102,N_29946,N_29997);
or UO_103 (O_103,N_29862,N_29945);
nor UO_104 (O_104,N_29928,N_29898);
or UO_105 (O_105,N_29936,N_29820);
or UO_106 (O_106,N_29822,N_29889);
xor UO_107 (O_107,N_29874,N_29820);
and UO_108 (O_108,N_29830,N_29997);
xor UO_109 (O_109,N_29868,N_29849);
or UO_110 (O_110,N_29993,N_29819);
xnor UO_111 (O_111,N_29908,N_29941);
or UO_112 (O_112,N_29973,N_29950);
nand UO_113 (O_113,N_29899,N_29816);
nor UO_114 (O_114,N_29935,N_29931);
and UO_115 (O_115,N_29956,N_29947);
or UO_116 (O_116,N_29949,N_29915);
or UO_117 (O_117,N_29822,N_29859);
xnor UO_118 (O_118,N_29893,N_29874);
nand UO_119 (O_119,N_29863,N_29890);
nor UO_120 (O_120,N_29801,N_29875);
or UO_121 (O_121,N_29814,N_29988);
or UO_122 (O_122,N_29961,N_29908);
nand UO_123 (O_123,N_29833,N_29906);
nor UO_124 (O_124,N_29845,N_29945);
xnor UO_125 (O_125,N_29838,N_29887);
and UO_126 (O_126,N_29847,N_29993);
and UO_127 (O_127,N_29970,N_29983);
nor UO_128 (O_128,N_29871,N_29843);
nor UO_129 (O_129,N_29972,N_29923);
nor UO_130 (O_130,N_29874,N_29866);
nand UO_131 (O_131,N_29908,N_29821);
xor UO_132 (O_132,N_29923,N_29945);
nand UO_133 (O_133,N_29830,N_29929);
or UO_134 (O_134,N_29822,N_29812);
xnor UO_135 (O_135,N_29848,N_29946);
nand UO_136 (O_136,N_29800,N_29917);
and UO_137 (O_137,N_29857,N_29824);
or UO_138 (O_138,N_29838,N_29863);
xor UO_139 (O_139,N_29813,N_29896);
or UO_140 (O_140,N_29964,N_29842);
or UO_141 (O_141,N_29829,N_29802);
and UO_142 (O_142,N_29820,N_29954);
nand UO_143 (O_143,N_29802,N_29918);
and UO_144 (O_144,N_29926,N_29841);
and UO_145 (O_145,N_29867,N_29872);
nor UO_146 (O_146,N_29956,N_29821);
or UO_147 (O_147,N_29894,N_29856);
nor UO_148 (O_148,N_29942,N_29824);
or UO_149 (O_149,N_29872,N_29819);
or UO_150 (O_150,N_29902,N_29802);
or UO_151 (O_151,N_29953,N_29872);
xor UO_152 (O_152,N_29958,N_29882);
nor UO_153 (O_153,N_29861,N_29849);
and UO_154 (O_154,N_29950,N_29859);
nand UO_155 (O_155,N_29931,N_29934);
or UO_156 (O_156,N_29944,N_29801);
and UO_157 (O_157,N_29924,N_29894);
nor UO_158 (O_158,N_29955,N_29906);
nor UO_159 (O_159,N_29989,N_29942);
or UO_160 (O_160,N_29845,N_29988);
and UO_161 (O_161,N_29870,N_29979);
or UO_162 (O_162,N_29898,N_29999);
xnor UO_163 (O_163,N_29880,N_29819);
or UO_164 (O_164,N_29807,N_29983);
or UO_165 (O_165,N_29824,N_29902);
and UO_166 (O_166,N_29973,N_29874);
or UO_167 (O_167,N_29850,N_29929);
nand UO_168 (O_168,N_29841,N_29858);
or UO_169 (O_169,N_29911,N_29984);
nor UO_170 (O_170,N_29807,N_29942);
and UO_171 (O_171,N_29844,N_29992);
xor UO_172 (O_172,N_29911,N_29908);
xor UO_173 (O_173,N_29856,N_29815);
or UO_174 (O_174,N_29856,N_29857);
nor UO_175 (O_175,N_29922,N_29831);
nand UO_176 (O_176,N_29925,N_29954);
or UO_177 (O_177,N_29876,N_29806);
or UO_178 (O_178,N_29957,N_29835);
and UO_179 (O_179,N_29996,N_29998);
xnor UO_180 (O_180,N_29925,N_29962);
nand UO_181 (O_181,N_29918,N_29889);
and UO_182 (O_182,N_29903,N_29895);
and UO_183 (O_183,N_29979,N_29933);
nor UO_184 (O_184,N_29825,N_29811);
xor UO_185 (O_185,N_29853,N_29965);
nand UO_186 (O_186,N_29838,N_29982);
xor UO_187 (O_187,N_29859,N_29880);
nor UO_188 (O_188,N_29991,N_29869);
or UO_189 (O_189,N_29836,N_29834);
nor UO_190 (O_190,N_29811,N_29953);
xor UO_191 (O_191,N_29846,N_29865);
nand UO_192 (O_192,N_29986,N_29936);
xnor UO_193 (O_193,N_29934,N_29831);
xor UO_194 (O_194,N_29999,N_29889);
or UO_195 (O_195,N_29973,N_29867);
nand UO_196 (O_196,N_29811,N_29845);
or UO_197 (O_197,N_29950,N_29830);
nor UO_198 (O_198,N_29940,N_29994);
nand UO_199 (O_199,N_29889,N_29865);
or UO_200 (O_200,N_29840,N_29960);
xor UO_201 (O_201,N_29829,N_29964);
and UO_202 (O_202,N_29888,N_29941);
and UO_203 (O_203,N_29822,N_29807);
nor UO_204 (O_204,N_29999,N_29915);
and UO_205 (O_205,N_29915,N_29971);
nor UO_206 (O_206,N_29947,N_29936);
nor UO_207 (O_207,N_29890,N_29901);
xor UO_208 (O_208,N_29989,N_29956);
nor UO_209 (O_209,N_29835,N_29868);
nor UO_210 (O_210,N_29876,N_29807);
xnor UO_211 (O_211,N_29871,N_29967);
nand UO_212 (O_212,N_29948,N_29827);
nand UO_213 (O_213,N_29820,N_29907);
xnor UO_214 (O_214,N_29955,N_29968);
and UO_215 (O_215,N_29852,N_29894);
and UO_216 (O_216,N_29989,N_29950);
xor UO_217 (O_217,N_29903,N_29818);
xnor UO_218 (O_218,N_29968,N_29996);
xor UO_219 (O_219,N_29878,N_29987);
nor UO_220 (O_220,N_29803,N_29832);
xor UO_221 (O_221,N_29991,N_29862);
and UO_222 (O_222,N_29843,N_29878);
xor UO_223 (O_223,N_29832,N_29847);
nand UO_224 (O_224,N_29900,N_29924);
nand UO_225 (O_225,N_29847,N_29831);
nor UO_226 (O_226,N_29838,N_29832);
nor UO_227 (O_227,N_29963,N_29869);
nor UO_228 (O_228,N_29810,N_29935);
xor UO_229 (O_229,N_29956,N_29998);
and UO_230 (O_230,N_29923,N_29958);
and UO_231 (O_231,N_29991,N_29802);
or UO_232 (O_232,N_29805,N_29838);
nor UO_233 (O_233,N_29978,N_29829);
and UO_234 (O_234,N_29874,N_29997);
or UO_235 (O_235,N_29800,N_29836);
or UO_236 (O_236,N_29897,N_29823);
xnor UO_237 (O_237,N_29896,N_29848);
or UO_238 (O_238,N_29892,N_29807);
nor UO_239 (O_239,N_29885,N_29829);
and UO_240 (O_240,N_29944,N_29951);
nor UO_241 (O_241,N_29853,N_29914);
and UO_242 (O_242,N_29838,N_29849);
and UO_243 (O_243,N_29902,N_29875);
xor UO_244 (O_244,N_29961,N_29886);
or UO_245 (O_245,N_29885,N_29811);
and UO_246 (O_246,N_29867,N_29917);
nand UO_247 (O_247,N_29835,N_29839);
or UO_248 (O_248,N_29984,N_29954);
nand UO_249 (O_249,N_29870,N_29859);
xor UO_250 (O_250,N_29989,N_29969);
nor UO_251 (O_251,N_29853,N_29828);
or UO_252 (O_252,N_29832,N_29980);
or UO_253 (O_253,N_29982,N_29942);
nand UO_254 (O_254,N_29830,N_29853);
nand UO_255 (O_255,N_29963,N_29964);
nor UO_256 (O_256,N_29826,N_29829);
and UO_257 (O_257,N_29923,N_29899);
xor UO_258 (O_258,N_29940,N_29906);
nand UO_259 (O_259,N_29876,N_29847);
and UO_260 (O_260,N_29824,N_29922);
nor UO_261 (O_261,N_29963,N_29941);
xnor UO_262 (O_262,N_29932,N_29986);
nand UO_263 (O_263,N_29862,N_29842);
and UO_264 (O_264,N_29974,N_29942);
nor UO_265 (O_265,N_29935,N_29920);
xnor UO_266 (O_266,N_29871,N_29852);
and UO_267 (O_267,N_29838,N_29963);
nand UO_268 (O_268,N_29992,N_29866);
nor UO_269 (O_269,N_29913,N_29843);
nor UO_270 (O_270,N_29861,N_29987);
xor UO_271 (O_271,N_29953,N_29994);
and UO_272 (O_272,N_29862,N_29931);
nor UO_273 (O_273,N_29825,N_29947);
or UO_274 (O_274,N_29919,N_29897);
xor UO_275 (O_275,N_29912,N_29955);
nand UO_276 (O_276,N_29994,N_29820);
nand UO_277 (O_277,N_29944,N_29924);
nor UO_278 (O_278,N_29904,N_29801);
or UO_279 (O_279,N_29945,N_29819);
and UO_280 (O_280,N_29873,N_29823);
nor UO_281 (O_281,N_29815,N_29826);
and UO_282 (O_282,N_29880,N_29929);
nand UO_283 (O_283,N_29872,N_29892);
nand UO_284 (O_284,N_29834,N_29907);
nor UO_285 (O_285,N_29818,N_29848);
and UO_286 (O_286,N_29993,N_29843);
xor UO_287 (O_287,N_29976,N_29964);
nand UO_288 (O_288,N_29872,N_29937);
and UO_289 (O_289,N_29929,N_29808);
or UO_290 (O_290,N_29850,N_29958);
xor UO_291 (O_291,N_29908,N_29925);
or UO_292 (O_292,N_29860,N_29826);
nor UO_293 (O_293,N_29920,N_29998);
or UO_294 (O_294,N_29884,N_29945);
nor UO_295 (O_295,N_29963,N_29829);
xor UO_296 (O_296,N_29941,N_29808);
and UO_297 (O_297,N_29844,N_29856);
or UO_298 (O_298,N_29861,N_29845);
nand UO_299 (O_299,N_29891,N_29823);
nor UO_300 (O_300,N_29962,N_29800);
nor UO_301 (O_301,N_29870,N_29836);
xor UO_302 (O_302,N_29803,N_29981);
and UO_303 (O_303,N_29976,N_29991);
nor UO_304 (O_304,N_29948,N_29867);
nand UO_305 (O_305,N_29868,N_29804);
nor UO_306 (O_306,N_29853,N_29865);
nand UO_307 (O_307,N_29953,N_29998);
nand UO_308 (O_308,N_29952,N_29912);
nand UO_309 (O_309,N_29889,N_29904);
nor UO_310 (O_310,N_29982,N_29936);
or UO_311 (O_311,N_29936,N_29845);
xnor UO_312 (O_312,N_29833,N_29811);
nand UO_313 (O_313,N_29842,N_29969);
and UO_314 (O_314,N_29813,N_29895);
nor UO_315 (O_315,N_29818,N_29813);
or UO_316 (O_316,N_29824,N_29821);
nand UO_317 (O_317,N_29967,N_29942);
and UO_318 (O_318,N_29938,N_29864);
or UO_319 (O_319,N_29848,N_29965);
nand UO_320 (O_320,N_29802,N_29977);
and UO_321 (O_321,N_29803,N_29920);
nand UO_322 (O_322,N_29874,N_29941);
nand UO_323 (O_323,N_29879,N_29808);
nor UO_324 (O_324,N_29944,N_29929);
nand UO_325 (O_325,N_29893,N_29869);
xor UO_326 (O_326,N_29802,N_29821);
and UO_327 (O_327,N_29894,N_29833);
xor UO_328 (O_328,N_29912,N_29878);
and UO_329 (O_329,N_29848,N_29939);
nand UO_330 (O_330,N_29922,N_29853);
nor UO_331 (O_331,N_29860,N_29955);
nand UO_332 (O_332,N_29814,N_29821);
and UO_333 (O_333,N_29993,N_29897);
or UO_334 (O_334,N_29915,N_29808);
or UO_335 (O_335,N_29936,N_29877);
xor UO_336 (O_336,N_29823,N_29883);
and UO_337 (O_337,N_29920,N_29929);
nand UO_338 (O_338,N_29832,N_29902);
xnor UO_339 (O_339,N_29844,N_29889);
nor UO_340 (O_340,N_29854,N_29950);
and UO_341 (O_341,N_29955,N_29845);
nor UO_342 (O_342,N_29801,N_29861);
xnor UO_343 (O_343,N_29880,N_29898);
nor UO_344 (O_344,N_29974,N_29993);
nor UO_345 (O_345,N_29804,N_29852);
nand UO_346 (O_346,N_29917,N_29804);
or UO_347 (O_347,N_29833,N_29823);
nor UO_348 (O_348,N_29878,N_29939);
or UO_349 (O_349,N_29946,N_29818);
or UO_350 (O_350,N_29893,N_29850);
or UO_351 (O_351,N_29923,N_29981);
nor UO_352 (O_352,N_29961,N_29939);
nand UO_353 (O_353,N_29859,N_29988);
or UO_354 (O_354,N_29865,N_29839);
xor UO_355 (O_355,N_29894,N_29945);
nor UO_356 (O_356,N_29862,N_29818);
and UO_357 (O_357,N_29811,N_29959);
xor UO_358 (O_358,N_29973,N_29939);
or UO_359 (O_359,N_29902,N_29939);
or UO_360 (O_360,N_29900,N_29861);
nor UO_361 (O_361,N_29837,N_29959);
nor UO_362 (O_362,N_29959,N_29947);
nand UO_363 (O_363,N_29810,N_29957);
nand UO_364 (O_364,N_29872,N_29908);
or UO_365 (O_365,N_29984,N_29888);
and UO_366 (O_366,N_29993,N_29965);
and UO_367 (O_367,N_29971,N_29883);
and UO_368 (O_368,N_29951,N_29920);
xor UO_369 (O_369,N_29911,N_29930);
and UO_370 (O_370,N_29859,N_29820);
or UO_371 (O_371,N_29845,N_29836);
and UO_372 (O_372,N_29969,N_29932);
xnor UO_373 (O_373,N_29883,N_29830);
xor UO_374 (O_374,N_29860,N_29943);
nand UO_375 (O_375,N_29921,N_29853);
nand UO_376 (O_376,N_29912,N_29950);
nor UO_377 (O_377,N_29850,N_29908);
nand UO_378 (O_378,N_29998,N_29857);
nor UO_379 (O_379,N_29837,N_29839);
xor UO_380 (O_380,N_29909,N_29807);
nor UO_381 (O_381,N_29814,N_29969);
xnor UO_382 (O_382,N_29861,N_29896);
or UO_383 (O_383,N_29884,N_29903);
xor UO_384 (O_384,N_29863,N_29938);
and UO_385 (O_385,N_29815,N_29937);
nand UO_386 (O_386,N_29887,N_29967);
and UO_387 (O_387,N_29926,N_29974);
xor UO_388 (O_388,N_29828,N_29889);
nand UO_389 (O_389,N_29855,N_29925);
or UO_390 (O_390,N_29982,N_29834);
xnor UO_391 (O_391,N_29876,N_29870);
and UO_392 (O_392,N_29904,N_29855);
or UO_393 (O_393,N_29915,N_29907);
and UO_394 (O_394,N_29931,N_29840);
and UO_395 (O_395,N_29958,N_29803);
and UO_396 (O_396,N_29863,N_29893);
nand UO_397 (O_397,N_29852,N_29997);
or UO_398 (O_398,N_29889,N_29924);
xnor UO_399 (O_399,N_29995,N_29987);
xnor UO_400 (O_400,N_29943,N_29992);
nor UO_401 (O_401,N_29873,N_29872);
nand UO_402 (O_402,N_29896,N_29962);
nor UO_403 (O_403,N_29898,N_29981);
nand UO_404 (O_404,N_29933,N_29958);
xnor UO_405 (O_405,N_29923,N_29827);
nand UO_406 (O_406,N_29913,N_29827);
and UO_407 (O_407,N_29888,N_29825);
nor UO_408 (O_408,N_29982,N_29810);
and UO_409 (O_409,N_29823,N_29918);
xnor UO_410 (O_410,N_29962,N_29806);
and UO_411 (O_411,N_29919,N_29865);
nor UO_412 (O_412,N_29821,N_29884);
and UO_413 (O_413,N_29944,N_29810);
and UO_414 (O_414,N_29863,N_29911);
nand UO_415 (O_415,N_29978,N_29819);
nand UO_416 (O_416,N_29832,N_29964);
nand UO_417 (O_417,N_29858,N_29812);
nand UO_418 (O_418,N_29953,N_29926);
nor UO_419 (O_419,N_29821,N_29938);
xor UO_420 (O_420,N_29826,N_29969);
xnor UO_421 (O_421,N_29921,N_29828);
xnor UO_422 (O_422,N_29875,N_29884);
xor UO_423 (O_423,N_29931,N_29854);
nand UO_424 (O_424,N_29845,N_29801);
and UO_425 (O_425,N_29884,N_29949);
or UO_426 (O_426,N_29880,N_29938);
xor UO_427 (O_427,N_29841,N_29827);
nand UO_428 (O_428,N_29825,N_29967);
nor UO_429 (O_429,N_29858,N_29959);
or UO_430 (O_430,N_29964,N_29866);
and UO_431 (O_431,N_29884,N_29977);
and UO_432 (O_432,N_29986,N_29955);
and UO_433 (O_433,N_29965,N_29831);
or UO_434 (O_434,N_29980,N_29976);
or UO_435 (O_435,N_29926,N_29866);
or UO_436 (O_436,N_29824,N_29884);
nand UO_437 (O_437,N_29900,N_29839);
and UO_438 (O_438,N_29971,N_29853);
or UO_439 (O_439,N_29807,N_29802);
and UO_440 (O_440,N_29818,N_29868);
and UO_441 (O_441,N_29906,N_29979);
and UO_442 (O_442,N_29940,N_29997);
nand UO_443 (O_443,N_29900,N_29908);
nand UO_444 (O_444,N_29991,N_29927);
or UO_445 (O_445,N_29928,N_29813);
or UO_446 (O_446,N_29814,N_29974);
nand UO_447 (O_447,N_29923,N_29857);
or UO_448 (O_448,N_29988,N_29862);
nor UO_449 (O_449,N_29816,N_29806);
nand UO_450 (O_450,N_29803,N_29891);
nor UO_451 (O_451,N_29978,N_29952);
nand UO_452 (O_452,N_29857,N_29895);
nand UO_453 (O_453,N_29881,N_29873);
and UO_454 (O_454,N_29931,N_29899);
xor UO_455 (O_455,N_29836,N_29943);
and UO_456 (O_456,N_29802,N_29948);
xor UO_457 (O_457,N_29972,N_29833);
nand UO_458 (O_458,N_29971,N_29986);
nand UO_459 (O_459,N_29997,N_29911);
nand UO_460 (O_460,N_29938,N_29886);
nand UO_461 (O_461,N_29830,N_29843);
nand UO_462 (O_462,N_29971,N_29919);
nand UO_463 (O_463,N_29907,N_29964);
nor UO_464 (O_464,N_29975,N_29808);
nand UO_465 (O_465,N_29811,N_29881);
nand UO_466 (O_466,N_29808,N_29947);
xor UO_467 (O_467,N_29912,N_29939);
or UO_468 (O_468,N_29807,N_29948);
nor UO_469 (O_469,N_29986,N_29975);
nor UO_470 (O_470,N_29906,N_29857);
xnor UO_471 (O_471,N_29896,N_29876);
and UO_472 (O_472,N_29873,N_29847);
or UO_473 (O_473,N_29980,N_29989);
xor UO_474 (O_474,N_29814,N_29861);
or UO_475 (O_475,N_29847,N_29866);
nor UO_476 (O_476,N_29896,N_29999);
nor UO_477 (O_477,N_29833,N_29867);
nor UO_478 (O_478,N_29963,N_29867);
nand UO_479 (O_479,N_29949,N_29984);
xnor UO_480 (O_480,N_29938,N_29802);
nor UO_481 (O_481,N_29988,N_29871);
xor UO_482 (O_482,N_29900,N_29855);
or UO_483 (O_483,N_29852,N_29991);
nor UO_484 (O_484,N_29823,N_29847);
nor UO_485 (O_485,N_29904,N_29860);
nor UO_486 (O_486,N_29904,N_29980);
nor UO_487 (O_487,N_29872,N_29916);
and UO_488 (O_488,N_29981,N_29829);
and UO_489 (O_489,N_29959,N_29984);
nand UO_490 (O_490,N_29849,N_29973);
and UO_491 (O_491,N_29817,N_29956);
and UO_492 (O_492,N_29804,N_29814);
and UO_493 (O_493,N_29946,N_29864);
nand UO_494 (O_494,N_29911,N_29815);
nor UO_495 (O_495,N_29949,N_29905);
xnor UO_496 (O_496,N_29803,N_29860);
or UO_497 (O_497,N_29800,N_29988);
or UO_498 (O_498,N_29839,N_29849);
xor UO_499 (O_499,N_29919,N_29853);
and UO_500 (O_500,N_29954,N_29993);
and UO_501 (O_501,N_29862,N_29887);
or UO_502 (O_502,N_29808,N_29979);
nand UO_503 (O_503,N_29901,N_29953);
xor UO_504 (O_504,N_29873,N_29976);
nand UO_505 (O_505,N_29952,N_29971);
or UO_506 (O_506,N_29937,N_29927);
nand UO_507 (O_507,N_29939,N_29860);
and UO_508 (O_508,N_29965,N_29866);
or UO_509 (O_509,N_29887,N_29931);
and UO_510 (O_510,N_29976,N_29963);
xnor UO_511 (O_511,N_29959,N_29831);
nand UO_512 (O_512,N_29938,N_29997);
nand UO_513 (O_513,N_29868,N_29874);
nor UO_514 (O_514,N_29939,N_29971);
or UO_515 (O_515,N_29897,N_29858);
xor UO_516 (O_516,N_29865,N_29911);
and UO_517 (O_517,N_29825,N_29829);
xor UO_518 (O_518,N_29964,N_29886);
nand UO_519 (O_519,N_29944,N_29910);
or UO_520 (O_520,N_29968,N_29944);
nand UO_521 (O_521,N_29901,N_29941);
xor UO_522 (O_522,N_29984,N_29963);
or UO_523 (O_523,N_29837,N_29971);
nor UO_524 (O_524,N_29978,N_29809);
nand UO_525 (O_525,N_29983,N_29928);
or UO_526 (O_526,N_29980,N_29815);
nand UO_527 (O_527,N_29955,N_29951);
and UO_528 (O_528,N_29934,N_29845);
nor UO_529 (O_529,N_29889,N_29814);
nor UO_530 (O_530,N_29995,N_29941);
and UO_531 (O_531,N_29893,N_29809);
xor UO_532 (O_532,N_29854,N_29922);
nor UO_533 (O_533,N_29827,N_29964);
nor UO_534 (O_534,N_29998,N_29960);
nor UO_535 (O_535,N_29932,N_29945);
nor UO_536 (O_536,N_29822,N_29802);
nand UO_537 (O_537,N_29882,N_29870);
nor UO_538 (O_538,N_29871,N_29965);
or UO_539 (O_539,N_29981,N_29903);
or UO_540 (O_540,N_29888,N_29853);
xor UO_541 (O_541,N_29984,N_29843);
or UO_542 (O_542,N_29938,N_29842);
or UO_543 (O_543,N_29972,N_29939);
and UO_544 (O_544,N_29961,N_29853);
or UO_545 (O_545,N_29960,N_29879);
or UO_546 (O_546,N_29852,N_29818);
nor UO_547 (O_547,N_29923,N_29825);
nand UO_548 (O_548,N_29846,N_29818);
or UO_549 (O_549,N_29872,N_29863);
nor UO_550 (O_550,N_29822,N_29969);
or UO_551 (O_551,N_29922,N_29809);
xor UO_552 (O_552,N_29904,N_29812);
or UO_553 (O_553,N_29983,N_29981);
nand UO_554 (O_554,N_29990,N_29892);
nand UO_555 (O_555,N_29893,N_29993);
nor UO_556 (O_556,N_29963,N_29846);
or UO_557 (O_557,N_29866,N_29943);
nor UO_558 (O_558,N_29842,N_29830);
or UO_559 (O_559,N_29982,N_29947);
or UO_560 (O_560,N_29956,N_29858);
or UO_561 (O_561,N_29884,N_29916);
nor UO_562 (O_562,N_29868,N_29989);
and UO_563 (O_563,N_29937,N_29858);
or UO_564 (O_564,N_29993,N_29809);
nor UO_565 (O_565,N_29943,N_29998);
xnor UO_566 (O_566,N_29979,N_29987);
nand UO_567 (O_567,N_29931,N_29995);
nor UO_568 (O_568,N_29893,N_29912);
or UO_569 (O_569,N_29890,N_29822);
xnor UO_570 (O_570,N_29814,N_29911);
nand UO_571 (O_571,N_29831,N_29936);
and UO_572 (O_572,N_29805,N_29947);
nor UO_573 (O_573,N_29945,N_29806);
xor UO_574 (O_574,N_29800,N_29878);
xor UO_575 (O_575,N_29976,N_29817);
nand UO_576 (O_576,N_29953,N_29960);
xor UO_577 (O_577,N_29914,N_29998);
xnor UO_578 (O_578,N_29861,N_29917);
nand UO_579 (O_579,N_29914,N_29992);
or UO_580 (O_580,N_29948,N_29813);
nand UO_581 (O_581,N_29984,N_29997);
or UO_582 (O_582,N_29820,N_29811);
and UO_583 (O_583,N_29854,N_29878);
nor UO_584 (O_584,N_29979,N_29994);
xor UO_585 (O_585,N_29963,N_29933);
xnor UO_586 (O_586,N_29958,N_29844);
and UO_587 (O_587,N_29945,N_29803);
and UO_588 (O_588,N_29987,N_29989);
nand UO_589 (O_589,N_29845,N_29917);
or UO_590 (O_590,N_29863,N_29820);
nand UO_591 (O_591,N_29839,N_29908);
nand UO_592 (O_592,N_29954,N_29936);
and UO_593 (O_593,N_29965,N_29898);
and UO_594 (O_594,N_29827,N_29981);
nand UO_595 (O_595,N_29861,N_29951);
and UO_596 (O_596,N_29993,N_29992);
or UO_597 (O_597,N_29810,N_29827);
or UO_598 (O_598,N_29954,N_29919);
and UO_599 (O_599,N_29923,N_29878);
xor UO_600 (O_600,N_29942,N_29901);
xnor UO_601 (O_601,N_29970,N_29997);
or UO_602 (O_602,N_29922,N_29841);
nor UO_603 (O_603,N_29879,N_29956);
nand UO_604 (O_604,N_29880,N_29807);
nor UO_605 (O_605,N_29837,N_29880);
or UO_606 (O_606,N_29907,N_29828);
and UO_607 (O_607,N_29931,N_29889);
nand UO_608 (O_608,N_29814,N_29836);
or UO_609 (O_609,N_29955,N_29857);
xnor UO_610 (O_610,N_29937,N_29941);
and UO_611 (O_611,N_29866,N_29870);
nand UO_612 (O_612,N_29948,N_29952);
or UO_613 (O_613,N_29844,N_29981);
xor UO_614 (O_614,N_29905,N_29824);
and UO_615 (O_615,N_29994,N_29886);
or UO_616 (O_616,N_29833,N_29950);
nand UO_617 (O_617,N_29803,N_29997);
xor UO_618 (O_618,N_29999,N_29969);
and UO_619 (O_619,N_29866,N_29805);
or UO_620 (O_620,N_29988,N_29935);
xnor UO_621 (O_621,N_29896,N_29901);
nor UO_622 (O_622,N_29970,N_29823);
nor UO_623 (O_623,N_29837,N_29904);
and UO_624 (O_624,N_29946,N_29957);
nand UO_625 (O_625,N_29898,N_29835);
xor UO_626 (O_626,N_29852,N_29877);
xnor UO_627 (O_627,N_29875,N_29918);
and UO_628 (O_628,N_29861,N_29816);
and UO_629 (O_629,N_29866,N_29917);
xnor UO_630 (O_630,N_29863,N_29909);
and UO_631 (O_631,N_29934,N_29940);
xor UO_632 (O_632,N_29977,N_29890);
xnor UO_633 (O_633,N_29835,N_29934);
and UO_634 (O_634,N_29827,N_29939);
xor UO_635 (O_635,N_29948,N_29907);
nand UO_636 (O_636,N_29824,N_29827);
nand UO_637 (O_637,N_29878,N_29907);
xor UO_638 (O_638,N_29922,N_29820);
or UO_639 (O_639,N_29823,N_29832);
and UO_640 (O_640,N_29880,N_29845);
xnor UO_641 (O_641,N_29982,N_29872);
xnor UO_642 (O_642,N_29823,N_29932);
xor UO_643 (O_643,N_29969,N_29900);
xor UO_644 (O_644,N_29829,N_29822);
nor UO_645 (O_645,N_29873,N_29849);
nor UO_646 (O_646,N_29861,N_29869);
or UO_647 (O_647,N_29982,N_29931);
or UO_648 (O_648,N_29985,N_29810);
xnor UO_649 (O_649,N_29898,N_29946);
nor UO_650 (O_650,N_29922,N_29961);
and UO_651 (O_651,N_29815,N_29835);
and UO_652 (O_652,N_29892,N_29997);
and UO_653 (O_653,N_29848,N_29926);
nor UO_654 (O_654,N_29986,N_29952);
nor UO_655 (O_655,N_29817,N_29913);
and UO_656 (O_656,N_29814,N_29850);
nor UO_657 (O_657,N_29906,N_29824);
xnor UO_658 (O_658,N_29924,N_29987);
or UO_659 (O_659,N_29811,N_29934);
or UO_660 (O_660,N_29868,N_29999);
and UO_661 (O_661,N_29947,N_29995);
nand UO_662 (O_662,N_29809,N_29931);
xor UO_663 (O_663,N_29898,N_29897);
nor UO_664 (O_664,N_29897,N_29819);
xnor UO_665 (O_665,N_29904,N_29911);
or UO_666 (O_666,N_29935,N_29925);
nand UO_667 (O_667,N_29959,N_29890);
nand UO_668 (O_668,N_29887,N_29982);
nand UO_669 (O_669,N_29883,N_29842);
nor UO_670 (O_670,N_29894,N_29961);
nor UO_671 (O_671,N_29969,N_29972);
and UO_672 (O_672,N_29825,N_29844);
and UO_673 (O_673,N_29905,N_29982);
nor UO_674 (O_674,N_29916,N_29923);
nand UO_675 (O_675,N_29943,N_29953);
or UO_676 (O_676,N_29880,N_29983);
or UO_677 (O_677,N_29894,N_29996);
or UO_678 (O_678,N_29807,N_29820);
or UO_679 (O_679,N_29847,N_29943);
and UO_680 (O_680,N_29815,N_29837);
nand UO_681 (O_681,N_29807,N_29843);
nand UO_682 (O_682,N_29995,N_29849);
xnor UO_683 (O_683,N_29929,N_29895);
nor UO_684 (O_684,N_29835,N_29914);
nor UO_685 (O_685,N_29984,N_29821);
nand UO_686 (O_686,N_29927,N_29903);
xor UO_687 (O_687,N_29975,N_29974);
nand UO_688 (O_688,N_29811,N_29985);
nor UO_689 (O_689,N_29999,N_29904);
nor UO_690 (O_690,N_29804,N_29853);
nor UO_691 (O_691,N_29923,N_29886);
nand UO_692 (O_692,N_29941,N_29978);
xor UO_693 (O_693,N_29954,N_29927);
and UO_694 (O_694,N_29881,N_29990);
xnor UO_695 (O_695,N_29868,N_29810);
nor UO_696 (O_696,N_29855,N_29847);
or UO_697 (O_697,N_29955,N_29858);
or UO_698 (O_698,N_29917,N_29846);
or UO_699 (O_699,N_29931,N_29888);
nor UO_700 (O_700,N_29933,N_29907);
xnor UO_701 (O_701,N_29921,N_29881);
and UO_702 (O_702,N_29977,N_29960);
nor UO_703 (O_703,N_29880,N_29868);
nand UO_704 (O_704,N_29912,N_29902);
or UO_705 (O_705,N_29920,N_29925);
nand UO_706 (O_706,N_29843,N_29863);
xnor UO_707 (O_707,N_29966,N_29903);
and UO_708 (O_708,N_29921,N_29808);
or UO_709 (O_709,N_29838,N_29824);
nor UO_710 (O_710,N_29807,N_29980);
nor UO_711 (O_711,N_29876,N_29892);
or UO_712 (O_712,N_29806,N_29980);
and UO_713 (O_713,N_29863,N_29850);
and UO_714 (O_714,N_29803,N_29862);
nor UO_715 (O_715,N_29901,N_29849);
nand UO_716 (O_716,N_29957,N_29988);
xnor UO_717 (O_717,N_29951,N_29889);
and UO_718 (O_718,N_29816,N_29870);
and UO_719 (O_719,N_29895,N_29836);
nor UO_720 (O_720,N_29991,N_29865);
and UO_721 (O_721,N_29852,N_29926);
and UO_722 (O_722,N_29872,N_29947);
nand UO_723 (O_723,N_29893,N_29916);
and UO_724 (O_724,N_29842,N_29913);
xor UO_725 (O_725,N_29879,N_29904);
nand UO_726 (O_726,N_29961,N_29827);
and UO_727 (O_727,N_29913,N_29929);
nand UO_728 (O_728,N_29831,N_29928);
xnor UO_729 (O_729,N_29988,N_29947);
xnor UO_730 (O_730,N_29819,N_29969);
and UO_731 (O_731,N_29970,N_29857);
and UO_732 (O_732,N_29837,N_29884);
or UO_733 (O_733,N_29924,N_29971);
and UO_734 (O_734,N_29862,N_29932);
xor UO_735 (O_735,N_29963,N_29983);
xor UO_736 (O_736,N_29971,N_29866);
nand UO_737 (O_737,N_29869,N_29920);
nor UO_738 (O_738,N_29910,N_29866);
nand UO_739 (O_739,N_29982,N_29945);
nand UO_740 (O_740,N_29906,N_29880);
nand UO_741 (O_741,N_29985,N_29945);
nor UO_742 (O_742,N_29836,N_29929);
and UO_743 (O_743,N_29922,N_29928);
and UO_744 (O_744,N_29845,N_29869);
nand UO_745 (O_745,N_29821,N_29980);
xnor UO_746 (O_746,N_29965,N_29857);
xnor UO_747 (O_747,N_29966,N_29828);
or UO_748 (O_748,N_29976,N_29864);
or UO_749 (O_749,N_29930,N_29940);
xor UO_750 (O_750,N_29993,N_29865);
xor UO_751 (O_751,N_29894,N_29974);
nand UO_752 (O_752,N_29820,N_29999);
or UO_753 (O_753,N_29933,N_29906);
or UO_754 (O_754,N_29885,N_29826);
or UO_755 (O_755,N_29855,N_29878);
xor UO_756 (O_756,N_29896,N_29837);
nand UO_757 (O_757,N_29967,N_29915);
or UO_758 (O_758,N_29965,N_29861);
or UO_759 (O_759,N_29854,N_29892);
nor UO_760 (O_760,N_29872,N_29981);
nand UO_761 (O_761,N_29858,N_29909);
nand UO_762 (O_762,N_29839,N_29948);
or UO_763 (O_763,N_29863,N_29884);
nor UO_764 (O_764,N_29959,N_29901);
xnor UO_765 (O_765,N_29878,N_29883);
nand UO_766 (O_766,N_29892,N_29923);
or UO_767 (O_767,N_29825,N_29963);
or UO_768 (O_768,N_29988,N_29981);
and UO_769 (O_769,N_29937,N_29958);
or UO_770 (O_770,N_29844,N_29937);
nand UO_771 (O_771,N_29844,N_29971);
and UO_772 (O_772,N_29907,N_29902);
nor UO_773 (O_773,N_29936,N_29899);
xor UO_774 (O_774,N_29853,N_29868);
nand UO_775 (O_775,N_29976,N_29843);
or UO_776 (O_776,N_29915,N_29960);
xor UO_777 (O_777,N_29978,N_29975);
and UO_778 (O_778,N_29898,N_29921);
nand UO_779 (O_779,N_29850,N_29874);
and UO_780 (O_780,N_29933,N_29989);
or UO_781 (O_781,N_29899,N_29858);
and UO_782 (O_782,N_29834,N_29867);
or UO_783 (O_783,N_29895,N_29807);
nor UO_784 (O_784,N_29946,N_29959);
nor UO_785 (O_785,N_29954,N_29841);
nor UO_786 (O_786,N_29856,N_29946);
nand UO_787 (O_787,N_29918,N_29820);
nor UO_788 (O_788,N_29896,N_29845);
xor UO_789 (O_789,N_29886,N_29813);
and UO_790 (O_790,N_29833,N_29961);
xnor UO_791 (O_791,N_29888,N_29815);
nor UO_792 (O_792,N_29955,N_29874);
nand UO_793 (O_793,N_29951,N_29999);
nor UO_794 (O_794,N_29852,N_29844);
or UO_795 (O_795,N_29957,N_29950);
or UO_796 (O_796,N_29857,N_29997);
nor UO_797 (O_797,N_29952,N_29944);
nor UO_798 (O_798,N_29979,N_29935);
xnor UO_799 (O_799,N_29987,N_29839);
and UO_800 (O_800,N_29822,N_29942);
and UO_801 (O_801,N_29859,N_29971);
and UO_802 (O_802,N_29995,N_29901);
or UO_803 (O_803,N_29831,N_29806);
xnor UO_804 (O_804,N_29932,N_29933);
nor UO_805 (O_805,N_29995,N_29970);
nand UO_806 (O_806,N_29892,N_29943);
nand UO_807 (O_807,N_29833,N_29904);
or UO_808 (O_808,N_29989,N_29833);
nand UO_809 (O_809,N_29875,N_29979);
nand UO_810 (O_810,N_29930,N_29942);
nor UO_811 (O_811,N_29803,N_29936);
nand UO_812 (O_812,N_29847,N_29875);
or UO_813 (O_813,N_29885,N_29859);
nor UO_814 (O_814,N_29881,N_29844);
and UO_815 (O_815,N_29987,N_29944);
and UO_816 (O_816,N_29897,N_29957);
nor UO_817 (O_817,N_29877,N_29875);
xnor UO_818 (O_818,N_29834,N_29894);
and UO_819 (O_819,N_29929,N_29879);
xnor UO_820 (O_820,N_29993,N_29975);
nand UO_821 (O_821,N_29988,N_29970);
nand UO_822 (O_822,N_29849,N_29840);
xor UO_823 (O_823,N_29924,N_29913);
xnor UO_824 (O_824,N_29988,N_29902);
and UO_825 (O_825,N_29968,N_29904);
and UO_826 (O_826,N_29840,N_29850);
nand UO_827 (O_827,N_29921,N_29884);
nor UO_828 (O_828,N_29908,N_29984);
and UO_829 (O_829,N_29894,N_29966);
nand UO_830 (O_830,N_29837,N_29955);
nand UO_831 (O_831,N_29920,N_29941);
xor UO_832 (O_832,N_29885,N_29819);
nor UO_833 (O_833,N_29867,N_29952);
or UO_834 (O_834,N_29920,N_29833);
nor UO_835 (O_835,N_29968,N_29847);
nor UO_836 (O_836,N_29950,N_29922);
nor UO_837 (O_837,N_29994,N_29856);
and UO_838 (O_838,N_29973,N_29869);
or UO_839 (O_839,N_29927,N_29982);
or UO_840 (O_840,N_29943,N_29935);
nor UO_841 (O_841,N_29867,N_29967);
and UO_842 (O_842,N_29909,N_29827);
or UO_843 (O_843,N_29926,N_29931);
nor UO_844 (O_844,N_29924,N_29931);
and UO_845 (O_845,N_29984,N_29842);
nor UO_846 (O_846,N_29893,N_29806);
xor UO_847 (O_847,N_29855,N_29965);
nor UO_848 (O_848,N_29987,N_29930);
or UO_849 (O_849,N_29886,N_29902);
nor UO_850 (O_850,N_29895,N_29901);
or UO_851 (O_851,N_29847,N_29836);
xnor UO_852 (O_852,N_29966,N_29803);
or UO_853 (O_853,N_29804,N_29839);
nor UO_854 (O_854,N_29964,N_29956);
nand UO_855 (O_855,N_29840,N_29802);
and UO_856 (O_856,N_29944,N_29990);
nand UO_857 (O_857,N_29889,N_29992);
nand UO_858 (O_858,N_29989,N_29901);
or UO_859 (O_859,N_29835,N_29837);
nor UO_860 (O_860,N_29851,N_29836);
xor UO_861 (O_861,N_29822,N_29805);
or UO_862 (O_862,N_29997,N_29972);
or UO_863 (O_863,N_29981,N_29866);
nand UO_864 (O_864,N_29936,N_29956);
nor UO_865 (O_865,N_29815,N_29905);
or UO_866 (O_866,N_29883,N_29906);
xor UO_867 (O_867,N_29963,N_29974);
and UO_868 (O_868,N_29861,N_29904);
or UO_869 (O_869,N_29976,N_29993);
nor UO_870 (O_870,N_29906,N_29865);
or UO_871 (O_871,N_29821,N_29817);
nand UO_872 (O_872,N_29889,N_29911);
xor UO_873 (O_873,N_29897,N_29947);
nor UO_874 (O_874,N_29876,N_29933);
nor UO_875 (O_875,N_29891,N_29904);
or UO_876 (O_876,N_29887,N_29894);
nand UO_877 (O_877,N_29804,N_29854);
nand UO_878 (O_878,N_29941,N_29944);
and UO_879 (O_879,N_29949,N_29979);
nand UO_880 (O_880,N_29883,N_29845);
nor UO_881 (O_881,N_29890,N_29819);
xnor UO_882 (O_882,N_29819,N_29954);
nor UO_883 (O_883,N_29829,N_29976);
or UO_884 (O_884,N_29998,N_29973);
nand UO_885 (O_885,N_29957,N_29846);
nor UO_886 (O_886,N_29984,N_29971);
xnor UO_887 (O_887,N_29817,N_29859);
nand UO_888 (O_888,N_29810,N_29834);
nor UO_889 (O_889,N_29975,N_29818);
xnor UO_890 (O_890,N_29852,N_29830);
and UO_891 (O_891,N_29920,N_29845);
nand UO_892 (O_892,N_29996,N_29954);
or UO_893 (O_893,N_29883,N_29945);
nand UO_894 (O_894,N_29802,N_29962);
nand UO_895 (O_895,N_29956,N_29802);
or UO_896 (O_896,N_29942,N_29886);
nand UO_897 (O_897,N_29869,N_29946);
xnor UO_898 (O_898,N_29834,N_29908);
nor UO_899 (O_899,N_29837,N_29813);
nand UO_900 (O_900,N_29979,N_29806);
nor UO_901 (O_901,N_29930,N_29881);
nand UO_902 (O_902,N_29971,N_29814);
and UO_903 (O_903,N_29944,N_29892);
nand UO_904 (O_904,N_29816,N_29883);
xnor UO_905 (O_905,N_29805,N_29905);
nor UO_906 (O_906,N_29858,N_29869);
nand UO_907 (O_907,N_29965,N_29889);
nand UO_908 (O_908,N_29806,N_29826);
and UO_909 (O_909,N_29802,N_29953);
and UO_910 (O_910,N_29901,N_29923);
or UO_911 (O_911,N_29912,N_29894);
and UO_912 (O_912,N_29800,N_29834);
or UO_913 (O_913,N_29858,N_29878);
xor UO_914 (O_914,N_29899,N_29919);
nand UO_915 (O_915,N_29915,N_29877);
nor UO_916 (O_916,N_29957,N_29832);
or UO_917 (O_917,N_29918,N_29946);
nand UO_918 (O_918,N_29925,N_29921);
and UO_919 (O_919,N_29965,N_29955);
nor UO_920 (O_920,N_29999,N_29902);
and UO_921 (O_921,N_29867,N_29812);
xor UO_922 (O_922,N_29922,N_29974);
and UO_923 (O_923,N_29854,N_29910);
nor UO_924 (O_924,N_29937,N_29830);
nand UO_925 (O_925,N_29862,N_29889);
and UO_926 (O_926,N_29988,N_29898);
nand UO_927 (O_927,N_29877,N_29890);
nor UO_928 (O_928,N_29954,N_29966);
nand UO_929 (O_929,N_29925,N_29941);
and UO_930 (O_930,N_29920,N_29821);
xor UO_931 (O_931,N_29974,N_29883);
xor UO_932 (O_932,N_29841,N_29860);
xnor UO_933 (O_933,N_29877,N_29888);
nand UO_934 (O_934,N_29813,N_29916);
nand UO_935 (O_935,N_29844,N_29945);
nand UO_936 (O_936,N_29918,N_29988);
nor UO_937 (O_937,N_29900,N_29886);
nor UO_938 (O_938,N_29964,N_29857);
nor UO_939 (O_939,N_29925,N_29916);
nor UO_940 (O_940,N_29966,N_29936);
or UO_941 (O_941,N_29973,N_29953);
nand UO_942 (O_942,N_29837,N_29938);
or UO_943 (O_943,N_29964,N_29905);
or UO_944 (O_944,N_29977,N_29951);
nand UO_945 (O_945,N_29805,N_29806);
and UO_946 (O_946,N_29839,N_29869);
nor UO_947 (O_947,N_29823,N_29993);
or UO_948 (O_948,N_29891,N_29860);
and UO_949 (O_949,N_29855,N_29956);
nand UO_950 (O_950,N_29891,N_29813);
xnor UO_951 (O_951,N_29970,N_29846);
and UO_952 (O_952,N_29961,N_29931);
nand UO_953 (O_953,N_29819,N_29866);
and UO_954 (O_954,N_29804,N_29877);
nand UO_955 (O_955,N_29935,N_29855);
nand UO_956 (O_956,N_29817,N_29874);
and UO_957 (O_957,N_29859,N_29964);
nand UO_958 (O_958,N_29969,N_29887);
nand UO_959 (O_959,N_29810,N_29889);
xnor UO_960 (O_960,N_29850,N_29898);
nand UO_961 (O_961,N_29994,N_29840);
nor UO_962 (O_962,N_29882,N_29898);
or UO_963 (O_963,N_29860,N_29856);
xor UO_964 (O_964,N_29937,N_29862);
and UO_965 (O_965,N_29869,N_29928);
nor UO_966 (O_966,N_29963,N_29879);
or UO_967 (O_967,N_29930,N_29995);
xor UO_968 (O_968,N_29920,N_29883);
and UO_969 (O_969,N_29851,N_29804);
nand UO_970 (O_970,N_29835,N_29948);
nand UO_971 (O_971,N_29852,N_29897);
or UO_972 (O_972,N_29995,N_29818);
xnor UO_973 (O_973,N_29899,N_29958);
nand UO_974 (O_974,N_29991,N_29945);
or UO_975 (O_975,N_29904,N_29933);
nand UO_976 (O_976,N_29978,N_29849);
xor UO_977 (O_977,N_29917,N_29820);
nor UO_978 (O_978,N_29915,N_29802);
nand UO_979 (O_979,N_29882,N_29940);
and UO_980 (O_980,N_29989,N_29852);
nand UO_981 (O_981,N_29980,N_29961);
xor UO_982 (O_982,N_29805,N_29921);
and UO_983 (O_983,N_29931,N_29869);
xnor UO_984 (O_984,N_29812,N_29863);
nor UO_985 (O_985,N_29882,N_29838);
nor UO_986 (O_986,N_29950,N_29880);
nand UO_987 (O_987,N_29980,N_29913);
and UO_988 (O_988,N_29831,N_29835);
nor UO_989 (O_989,N_29943,N_29988);
nand UO_990 (O_990,N_29934,N_29902);
nand UO_991 (O_991,N_29995,N_29800);
nand UO_992 (O_992,N_29970,N_29802);
or UO_993 (O_993,N_29834,N_29919);
xor UO_994 (O_994,N_29970,N_29836);
or UO_995 (O_995,N_29861,N_29910);
nor UO_996 (O_996,N_29949,N_29914);
nand UO_997 (O_997,N_29884,N_29827);
or UO_998 (O_998,N_29825,N_29933);
and UO_999 (O_999,N_29884,N_29959);
nand UO_1000 (O_1000,N_29871,N_29954);
and UO_1001 (O_1001,N_29824,N_29939);
or UO_1002 (O_1002,N_29928,N_29899);
nor UO_1003 (O_1003,N_29950,N_29998);
or UO_1004 (O_1004,N_29884,N_29883);
and UO_1005 (O_1005,N_29832,N_29815);
xnor UO_1006 (O_1006,N_29822,N_29837);
and UO_1007 (O_1007,N_29815,N_29833);
or UO_1008 (O_1008,N_29963,N_29968);
nand UO_1009 (O_1009,N_29959,N_29853);
xnor UO_1010 (O_1010,N_29933,N_29914);
xor UO_1011 (O_1011,N_29896,N_29926);
or UO_1012 (O_1012,N_29994,N_29896);
and UO_1013 (O_1013,N_29996,N_29916);
and UO_1014 (O_1014,N_29953,N_29806);
or UO_1015 (O_1015,N_29961,N_29904);
nand UO_1016 (O_1016,N_29868,N_29936);
nand UO_1017 (O_1017,N_29969,N_29864);
xnor UO_1018 (O_1018,N_29872,N_29980);
xor UO_1019 (O_1019,N_29862,N_29881);
or UO_1020 (O_1020,N_29939,N_29897);
nor UO_1021 (O_1021,N_29943,N_29851);
nand UO_1022 (O_1022,N_29870,N_29902);
or UO_1023 (O_1023,N_29854,N_29935);
and UO_1024 (O_1024,N_29921,N_29865);
nor UO_1025 (O_1025,N_29807,N_29861);
or UO_1026 (O_1026,N_29898,N_29802);
xnor UO_1027 (O_1027,N_29866,N_29885);
nor UO_1028 (O_1028,N_29886,N_29823);
nand UO_1029 (O_1029,N_29974,N_29908);
nand UO_1030 (O_1030,N_29843,N_29910);
or UO_1031 (O_1031,N_29823,N_29949);
nand UO_1032 (O_1032,N_29959,N_29843);
nor UO_1033 (O_1033,N_29939,N_29872);
and UO_1034 (O_1034,N_29981,N_29946);
and UO_1035 (O_1035,N_29863,N_29828);
nand UO_1036 (O_1036,N_29921,N_29947);
xor UO_1037 (O_1037,N_29830,N_29806);
xnor UO_1038 (O_1038,N_29891,N_29954);
or UO_1039 (O_1039,N_29827,N_29972);
xnor UO_1040 (O_1040,N_29859,N_29969);
xnor UO_1041 (O_1041,N_29973,N_29856);
and UO_1042 (O_1042,N_29940,N_29804);
or UO_1043 (O_1043,N_29945,N_29843);
nand UO_1044 (O_1044,N_29807,N_29864);
nand UO_1045 (O_1045,N_29986,N_29853);
or UO_1046 (O_1046,N_29927,N_29960);
and UO_1047 (O_1047,N_29968,N_29917);
nand UO_1048 (O_1048,N_29805,N_29893);
nand UO_1049 (O_1049,N_29875,N_29932);
xnor UO_1050 (O_1050,N_29995,N_29888);
and UO_1051 (O_1051,N_29838,N_29831);
nor UO_1052 (O_1052,N_29819,N_29975);
nand UO_1053 (O_1053,N_29914,N_29840);
and UO_1054 (O_1054,N_29860,N_29967);
nand UO_1055 (O_1055,N_29804,N_29924);
xnor UO_1056 (O_1056,N_29911,N_29821);
xnor UO_1057 (O_1057,N_29887,N_29902);
or UO_1058 (O_1058,N_29845,N_29838);
nor UO_1059 (O_1059,N_29977,N_29981);
and UO_1060 (O_1060,N_29951,N_29848);
and UO_1061 (O_1061,N_29988,N_29900);
nand UO_1062 (O_1062,N_29918,N_29972);
or UO_1063 (O_1063,N_29941,N_29841);
and UO_1064 (O_1064,N_29881,N_29843);
nand UO_1065 (O_1065,N_29885,N_29963);
nor UO_1066 (O_1066,N_29880,N_29993);
and UO_1067 (O_1067,N_29834,N_29998);
xnor UO_1068 (O_1068,N_29850,N_29956);
nor UO_1069 (O_1069,N_29849,N_29943);
xnor UO_1070 (O_1070,N_29842,N_29907);
nor UO_1071 (O_1071,N_29879,N_29805);
nor UO_1072 (O_1072,N_29988,N_29973);
and UO_1073 (O_1073,N_29808,N_29886);
nor UO_1074 (O_1074,N_29966,N_29995);
and UO_1075 (O_1075,N_29885,N_29869);
xnor UO_1076 (O_1076,N_29927,N_29969);
or UO_1077 (O_1077,N_29879,N_29866);
xor UO_1078 (O_1078,N_29874,N_29993);
nand UO_1079 (O_1079,N_29828,N_29858);
and UO_1080 (O_1080,N_29988,N_29888);
nand UO_1081 (O_1081,N_29872,N_29866);
nor UO_1082 (O_1082,N_29979,N_29988);
and UO_1083 (O_1083,N_29818,N_29857);
xnor UO_1084 (O_1084,N_29955,N_29846);
xor UO_1085 (O_1085,N_29888,N_29886);
xnor UO_1086 (O_1086,N_29909,N_29882);
and UO_1087 (O_1087,N_29917,N_29953);
nor UO_1088 (O_1088,N_29985,N_29961);
xor UO_1089 (O_1089,N_29916,N_29815);
nand UO_1090 (O_1090,N_29847,N_29879);
nand UO_1091 (O_1091,N_29968,N_29923);
or UO_1092 (O_1092,N_29961,N_29845);
and UO_1093 (O_1093,N_29919,N_29810);
nand UO_1094 (O_1094,N_29874,N_29948);
xnor UO_1095 (O_1095,N_29987,N_29927);
and UO_1096 (O_1096,N_29975,N_29837);
nand UO_1097 (O_1097,N_29858,N_29991);
nand UO_1098 (O_1098,N_29965,N_29872);
or UO_1099 (O_1099,N_29952,N_29810);
or UO_1100 (O_1100,N_29964,N_29911);
and UO_1101 (O_1101,N_29952,N_29914);
or UO_1102 (O_1102,N_29902,N_29983);
and UO_1103 (O_1103,N_29935,N_29970);
xor UO_1104 (O_1104,N_29944,N_29881);
or UO_1105 (O_1105,N_29803,N_29824);
nand UO_1106 (O_1106,N_29907,N_29823);
nand UO_1107 (O_1107,N_29855,N_29953);
xor UO_1108 (O_1108,N_29968,N_29907);
xor UO_1109 (O_1109,N_29977,N_29839);
nand UO_1110 (O_1110,N_29948,N_29882);
xor UO_1111 (O_1111,N_29859,N_29862);
nand UO_1112 (O_1112,N_29803,N_29809);
or UO_1113 (O_1113,N_29939,N_29928);
nand UO_1114 (O_1114,N_29993,N_29883);
and UO_1115 (O_1115,N_29978,N_29912);
xnor UO_1116 (O_1116,N_29986,N_29944);
and UO_1117 (O_1117,N_29951,N_29933);
xor UO_1118 (O_1118,N_29850,N_29967);
or UO_1119 (O_1119,N_29856,N_29832);
and UO_1120 (O_1120,N_29853,N_29973);
nand UO_1121 (O_1121,N_29800,N_29992);
xor UO_1122 (O_1122,N_29955,N_29936);
nand UO_1123 (O_1123,N_29986,N_29874);
or UO_1124 (O_1124,N_29815,N_29930);
nand UO_1125 (O_1125,N_29971,N_29997);
nor UO_1126 (O_1126,N_29991,N_29806);
xor UO_1127 (O_1127,N_29990,N_29816);
nand UO_1128 (O_1128,N_29906,N_29982);
or UO_1129 (O_1129,N_29899,N_29860);
or UO_1130 (O_1130,N_29950,N_29949);
and UO_1131 (O_1131,N_29804,N_29941);
nor UO_1132 (O_1132,N_29965,N_29880);
nor UO_1133 (O_1133,N_29933,N_29871);
nand UO_1134 (O_1134,N_29955,N_29816);
and UO_1135 (O_1135,N_29959,N_29821);
and UO_1136 (O_1136,N_29902,N_29818);
nor UO_1137 (O_1137,N_29990,N_29924);
and UO_1138 (O_1138,N_29911,N_29932);
or UO_1139 (O_1139,N_29981,N_29957);
xnor UO_1140 (O_1140,N_29852,N_29803);
xnor UO_1141 (O_1141,N_29889,N_29957);
nand UO_1142 (O_1142,N_29956,N_29876);
nand UO_1143 (O_1143,N_29807,N_29998);
and UO_1144 (O_1144,N_29990,N_29936);
nand UO_1145 (O_1145,N_29895,N_29907);
nand UO_1146 (O_1146,N_29993,N_29888);
and UO_1147 (O_1147,N_29959,N_29985);
nor UO_1148 (O_1148,N_29876,N_29836);
and UO_1149 (O_1149,N_29869,N_29948);
and UO_1150 (O_1150,N_29984,N_29986);
or UO_1151 (O_1151,N_29920,N_29928);
or UO_1152 (O_1152,N_29825,N_29943);
nor UO_1153 (O_1153,N_29954,N_29968);
or UO_1154 (O_1154,N_29902,N_29942);
or UO_1155 (O_1155,N_29926,N_29911);
xnor UO_1156 (O_1156,N_29871,N_29878);
xnor UO_1157 (O_1157,N_29852,N_29995);
xnor UO_1158 (O_1158,N_29847,N_29841);
xnor UO_1159 (O_1159,N_29957,N_29867);
nand UO_1160 (O_1160,N_29973,N_29804);
nor UO_1161 (O_1161,N_29893,N_29910);
xnor UO_1162 (O_1162,N_29859,N_29900);
nor UO_1163 (O_1163,N_29852,N_29982);
or UO_1164 (O_1164,N_29895,N_29960);
nor UO_1165 (O_1165,N_29904,N_29847);
nor UO_1166 (O_1166,N_29922,N_29842);
xor UO_1167 (O_1167,N_29826,N_29937);
nand UO_1168 (O_1168,N_29913,N_29835);
and UO_1169 (O_1169,N_29821,N_29846);
nor UO_1170 (O_1170,N_29852,N_29854);
xor UO_1171 (O_1171,N_29979,N_29844);
nand UO_1172 (O_1172,N_29834,N_29928);
xor UO_1173 (O_1173,N_29889,N_29842);
nand UO_1174 (O_1174,N_29851,N_29984);
nor UO_1175 (O_1175,N_29813,N_29925);
nor UO_1176 (O_1176,N_29857,N_29959);
xnor UO_1177 (O_1177,N_29863,N_29962);
nor UO_1178 (O_1178,N_29835,N_29900);
nand UO_1179 (O_1179,N_29971,N_29981);
xnor UO_1180 (O_1180,N_29971,N_29807);
and UO_1181 (O_1181,N_29816,N_29862);
or UO_1182 (O_1182,N_29991,N_29957);
nand UO_1183 (O_1183,N_29924,N_29831);
nand UO_1184 (O_1184,N_29808,N_29862);
or UO_1185 (O_1185,N_29976,N_29810);
xor UO_1186 (O_1186,N_29910,N_29943);
nor UO_1187 (O_1187,N_29893,N_29931);
nand UO_1188 (O_1188,N_29804,N_29886);
nand UO_1189 (O_1189,N_29900,N_29977);
nor UO_1190 (O_1190,N_29829,N_29993);
xor UO_1191 (O_1191,N_29864,N_29893);
nand UO_1192 (O_1192,N_29877,N_29813);
nand UO_1193 (O_1193,N_29975,N_29908);
or UO_1194 (O_1194,N_29943,N_29805);
nor UO_1195 (O_1195,N_29938,N_29925);
and UO_1196 (O_1196,N_29884,N_29830);
or UO_1197 (O_1197,N_29905,N_29870);
xnor UO_1198 (O_1198,N_29890,N_29870);
nor UO_1199 (O_1199,N_29904,N_29895);
nand UO_1200 (O_1200,N_29950,N_29817);
or UO_1201 (O_1201,N_29828,N_29833);
xnor UO_1202 (O_1202,N_29831,N_29970);
xor UO_1203 (O_1203,N_29815,N_29870);
nor UO_1204 (O_1204,N_29897,N_29952);
and UO_1205 (O_1205,N_29832,N_29928);
and UO_1206 (O_1206,N_29986,N_29920);
xnor UO_1207 (O_1207,N_29954,N_29836);
nor UO_1208 (O_1208,N_29912,N_29948);
nor UO_1209 (O_1209,N_29823,N_29816);
nor UO_1210 (O_1210,N_29868,N_29915);
nand UO_1211 (O_1211,N_29852,N_29889);
or UO_1212 (O_1212,N_29807,N_29865);
or UO_1213 (O_1213,N_29873,N_29806);
nand UO_1214 (O_1214,N_29948,N_29804);
xnor UO_1215 (O_1215,N_29955,N_29999);
and UO_1216 (O_1216,N_29943,N_29843);
xnor UO_1217 (O_1217,N_29847,N_29961);
and UO_1218 (O_1218,N_29914,N_29837);
or UO_1219 (O_1219,N_29927,N_29891);
or UO_1220 (O_1220,N_29936,N_29931);
or UO_1221 (O_1221,N_29989,N_29850);
nor UO_1222 (O_1222,N_29817,N_29929);
nand UO_1223 (O_1223,N_29818,N_29951);
nand UO_1224 (O_1224,N_29964,N_29939);
xor UO_1225 (O_1225,N_29871,N_29842);
and UO_1226 (O_1226,N_29890,N_29814);
nor UO_1227 (O_1227,N_29841,N_29942);
or UO_1228 (O_1228,N_29903,N_29971);
and UO_1229 (O_1229,N_29907,N_29865);
nor UO_1230 (O_1230,N_29985,N_29910);
nand UO_1231 (O_1231,N_29861,N_29871);
or UO_1232 (O_1232,N_29872,N_29926);
and UO_1233 (O_1233,N_29839,N_29999);
or UO_1234 (O_1234,N_29975,N_29859);
nand UO_1235 (O_1235,N_29865,N_29975);
and UO_1236 (O_1236,N_29891,N_29897);
and UO_1237 (O_1237,N_29807,N_29863);
xor UO_1238 (O_1238,N_29923,N_29882);
or UO_1239 (O_1239,N_29865,N_29827);
nand UO_1240 (O_1240,N_29885,N_29951);
xor UO_1241 (O_1241,N_29864,N_29885);
nand UO_1242 (O_1242,N_29938,N_29989);
and UO_1243 (O_1243,N_29973,N_29833);
and UO_1244 (O_1244,N_29926,N_29809);
xnor UO_1245 (O_1245,N_29808,N_29849);
xor UO_1246 (O_1246,N_29903,N_29866);
and UO_1247 (O_1247,N_29826,N_29903);
and UO_1248 (O_1248,N_29965,N_29998);
or UO_1249 (O_1249,N_29831,N_29956);
nor UO_1250 (O_1250,N_29974,N_29910);
nand UO_1251 (O_1251,N_29870,N_29878);
and UO_1252 (O_1252,N_29881,N_29945);
xnor UO_1253 (O_1253,N_29881,N_29982);
xor UO_1254 (O_1254,N_29864,N_29861);
nor UO_1255 (O_1255,N_29934,N_29973);
xor UO_1256 (O_1256,N_29979,N_29973);
nor UO_1257 (O_1257,N_29814,N_29949);
nand UO_1258 (O_1258,N_29836,N_29955);
xnor UO_1259 (O_1259,N_29994,N_29863);
or UO_1260 (O_1260,N_29812,N_29802);
nor UO_1261 (O_1261,N_29913,N_29939);
nor UO_1262 (O_1262,N_29982,N_29897);
nor UO_1263 (O_1263,N_29895,N_29827);
and UO_1264 (O_1264,N_29895,N_29835);
xor UO_1265 (O_1265,N_29859,N_29994);
or UO_1266 (O_1266,N_29808,N_29908);
and UO_1267 (O_1267,N_29812,N_29993);
nand UO_1268 (O_1268,N_29933,N_29946);
or UO_1269 (O_1269,N_29915,N_29829);
xor UO_1270 (O_1270,N_29905,N_29985);
nor UO_1271 (O_1271,N_29869,N_29832);
nand UO_1272 (O_1272,N_29995,N_29922);
and UO_1273 (O_1273,N_29936,N_29806);
xnor UO_1274 (O_1274,N_29953,N_29857);
or UO_1275 (O_1275,N_29926,N_29923);
or UO_1276 (O_1276,N_29986,N_29998);
and UO_1277 (O_1277,N_29800,N_29844);
or UO_1278 (O_1278,N_29825,N_29840);
xor UO_1279 (O_1279,N_29948,N_29967);
and UO_1280 (O_1280,N_29859,N_29802);
xnor UO_1281 (O_1281,N_29989,N_29959);
xnor UO_1282 (O_1282,N_29831,N_29998);
nor UO_1283 (O_1283,N_29880,N_29941);
nor UO_1284 (O_1284,N_29830,N_29953);
or UO_1285 (O_1285,N_29836,N_29841);
and UO_1286 (O_1286,N_29948,N_29906);
xor UO_1287 (O_1287,N_29995,N_29869);
nand UO_1288 (O_1288,N_29998,N_29903);
nor UO_1289 (O_1289,N_29915,N_29952);
or UO_1290 (O_1290,N_29875,N_29869);
and UO_1291 (O_1291,N_29868,N_29925);
xor UO_1292 (O_1292,N_29901,N_29884);
and UO_1293 (O_1293,N_29983,N_29978);
nor UO_1294 (O_1294,N_29954,N_29950);
and UO_1295 (O_1295,N_29914,N_29954);
nand UO_1296 (O_1296,N_29802,N_29997);
nor UO_1297 (O_1297,N_29887,N_29867);
nand UO_1298 (O_1298,N_29935,N_29954);
nand UO_1299 (O_1299,N_29911,N_29952);
nor UO_1300 (O_1300,N_29855,N_29879);
nand UO_1301 (O_1301,N_29863,N_29974);
xnor UO_1302 (O_1302,N_29830,N_29948);
nand UO_1303 (O_1303,N_29992,N_29885);
xnor UO_1304 (O_1304,N_29926,N_29907);
and UO_1305 (O_1305,N_29895,N_29972);
or UO_1306 (O_1306,N_29971,N_29926);
xor UO_1307 (O_1307,N_29802,N_29818);
and UO_1308 (O_1308,N_29886,N_29957);
xor UO_1309 (O_1309,N_29815,N_29822);
xor UO_1310 (O_1310,N_29892,N_29897);
nand UO_1311 (O_1311,N_29989,N_29883);
and UO_1312 (O_1312,N_29903,N_29926);
nand UO_1313 (O_1313,N_29940,N_29857);
and UO_1314 (O_1314,N_29834,N_29974);
and UO_1315 (O_1315,N_29973,N_29883);
and UO_1316 (O_1316,N_29844,N_29840);
nor UO_1317 (O_1317,N_29951,N_29985);
xnor UO_1318 (O_1318,N_29955,N_29920);
xnor UO_1319 (O_1319,N_29927,N_29957);
or UO_1320 (O_1320,N_29890,N_29889);
or UO_1321 (O_1321,N_29839,N_29818);
or UO_1322 (O_1322,N_29812,N_29917);
and UO_1323 (O_1323,N_29825,N_29924);
nor UO_1324 (O_1324,N_29958,N_29961);
nor UO_1325 (O_1325,N_29848,N_29849);
or UO_1326 (O_1326,N_29835,N_29930);
nor UO_1327 (O_1327,N_29820,N_29966);
nand UO_1328 (O_1328,N_29979,N_29842);
and UO_1329 (O_1329,N_29976,N_29960);
and UO_1330 (O_1330,N_29990,N_29846);
or UO_1331 (O_1331,N_29833,N_29966);
or UO_1332 (O_1332,N_29892,N_29932);
nor UO_1333 (O_1333,N_29888,N_29953);
and UO_1334 (O_1334,N_29921,N_29970);
nor UO_1335 (O_1335,N_29903,N_29871);
nand UO_1336 (O_1336,N_29917,N_29847);
or UO_1337 (O_1337,N_29830,N_29879);
xnor UO_1338 (O_1338,N_29838,N_29877);
xnor UO_1339 (O_1339,N_29927,N_29992);
nand UO_1340 (O_1340,N_29918,N_29877);
or UO_1341 (O_1341,N_29863,N_29830);
xor UO_1342 (O_1342,N_29911,N_29992);
xnor UO_1343 (O_1343,N_29914,N_29843);
nor UO_1344 (O_1344,N_29997,N_29979);
and UO_1345 (O_1345,N_29892,N_29884);
or UO_1346 (O_1346,N_29825,N_29999);
or UO_1347 (O_1347,N_29806,N_29977);
and UO_1348 (O_1348,N_29868,N_29988);
xnor UO_1349 (O_1349,N_29813,N_29878);
or UO_1350 (O_1350,N_29906,N_29834);
and UO_1351 (O_1351,N_29823,N_29913);
and UO_1352 (O_1352,N_29913,N_29829);
nand UO_1353 (O_1353,N_29951,N_29863);
xor UO_1354 (O_1354,N_29893,N_29846);
and UO_1355 (O_1355,N_29829,N_29871);
and UO_1356 (O_1356,N_29970,N_29877);
nor UO_1357 (O_1357,N_29833,N_29856);
xor UO_1358 (O_1358,N_29930,N_29912);
and UO_1359 (O_1359,N_29989,N_29881);
nor UO_1360 (O_1360,N_29932,N_29876);
or UO_1361 (O_1361,N_29997,N_29839);
or UO_1362 (O_1362,N_29945,N_29886);
and UO_1363 (O_1363,N_29939,N_29916);
nor UO_1364 (O_1364,N_29916,N_29904);
nor UO_1365 (O_1365,N_29935,N_29847);
nor UO_1366 (O_1366,N_29839,N_29947);
nand UO_1367 (O_1367,N_29812,N_29896);
xnor UO_1368 (O_1368,N_29976,N_29879);
or UO_1369 (O_1369,N_29974,N_29948);
or UO_1370 (O_1370,N_29994,N_29905);
or UO_1371 (O_1371,N_29887,N_29879);
nand UO_1372 (O_1372,N_29955,N_29871);
nand UO_1373 (O_1373,N_29841,N_29951);
nor UO_1374 (O_1374,N_29882,N_29910);
or UO_1375 (O_1375,N_29886,N_29951);
nor UO_1376 (O_1376,N_29920,N_29816);
nor UO_1377 (O_1377,N_29809,N_29821);
nand UO_1378 (O_1378,N_29911,N_29832);
and UO_1379 (O_1379,N_29822,N_29851);
and UO_1380 (O_1380,N_29808,N_29903);
nand UO_1381 (O_1381,N_29925,N_29919);
xnor UO_1382 (O_1382,N_29935,N_29898);
and UO_1383 (O_1383,N_29883,N_29814);
or UO_1384 (O_1384,N_29909,N_29946);
and UO_1385 (O_1385,N_29981,N_29936);
nand UO_1386 (O_1386,N_29865,N_29961);
or UO_1387 (O_1387,N_29889,N_29806);
xor UO_1388 (O_1388,N_29922,N_29847);
xnor UO_1389 (O_1389,N_29918,N_29807);
nand UO_1390 (O_1390,N_29887,N_29950);
nor UO_1391 (O_1391,N_29805,N_29935);
or UO_1392 (O_1392,N_29806,N_29860);
xnor UO_1393 (O_1393,N_29960,N_29888);
xnor UO_1394 (O_1394,N_29953,N_29865);
or UO_1395 (O_1395,N_29880,N_29961);
xnor UO_1396 (O_1396,N_29879,N_29874);
or UO_1397 (O_1397,N_29820,N_29927);
xor UO_1398 (O_1398,N_29866,N_29969);
nand UO_1399 (O_1399,N_29822,N_29852);
nand UO_1400 (O_1400,N_29846,N_29908);
or UO_1401 (O_1401,N_29813,N_29936);
nand UO_1402 (O_1402,N_29936,N_29833);
xnor UO_1403 (O_1403,N_29813,N_29914);
and UO_1404 (O_1404,N_29868,N_29952);
nand UO_1405 (O_1405,N_29986,N_29884);
nand UO_1406 (O_1406,N_29842,N_29973);
nand UO_1407 (O_1407,N_29973,N_29808);
xor UO_1408 (O_1408,N_29949,N_29986);
nand UO_1409 (O_1409,N_29987,N_29863);
or UO_1410 (O_1410,N_29974,N_29928);
xnor UO_1411 (O_1411,N_29816,N_29805);
nor UO_1412 (O_1412,N_29948,N_29932);
nor UO_1413 (O_1413,N_29869,N_29968);
and UO_1414 (O_1414,N_29989,N_29992);
nand UO_1415 (O_1415,N_29954,N_29892);
nor UO_1416 (O_1416,N_29982,N_29988);
nand UO_1417 (O_1417,N_29912,N_29839);
and UO_1418 (O_1418,N_29988,N_29976);
nor UO_1419 (O_1419,N_29923,N_29854);
xnor UO_1420 (O_1420,N_29864,N_29803);
nand UO_1421 (O_1421,N_29948,N_29977);
and UO_1422 (O_1422,N_29843,N_29992);
nor UO_1423 (O_1423,N_29996,N_29973);
nand UO_1424 (O_1424,N_29859,N_29853);
nor UO_1425 (O_1425,N_29973,N_29944);
nor UO_1426 (O_1426,N_29832,N_29971);
nor UO_1427 (O_1427,N_29802,N_29874);
nor UO_1428 (O_1428,N_29854,N_29821);
xnor UO_1429 (O_1429,N_29847,N_29845);
nor UO_1430 (O_1430,N_29900,N_29854);
or UO_1431 (O_1431,N_29969,N_29891);
nor UO_1432 (O_1432,N_29917,N_29900);
xor UO_1433 (O_1433,N_29879,N_29831);
xnor UO_1434 (O_1434,N_29957,N_29958);
nand UO_1435 (O_1435,N_29847,N_29871);
nand UO_1436 (O_1436,N_29868,N_29864);
or UO_1437 (O_1437,N_29853,N_29955);
nand UO_1438 (O_1438,N_29801,N_29828);
xnor UO_1439 (O_1439,N_29953,N_29803);
nand UO_1440 (O_1440,N_29805,N_29845);
or UO_1441 (O_1441,N_29831,N_29992);
xnor UO_1442 (O_1442,N_29977,N_29994);
xor UO_1443 (O_1443,N_29954,N_29874);
xor UO_1444 (O_1444,N_29845,N_29888);
xnor UO_1445 (O_1445,N_29915,N_29984);
or UO_1446 (O_1446,N_29829,N_29952);
and UO_1447 (O_1447,N_29997,N_29826);
nor UO_1448 (O_1448,N_29823,N_29908);
or UO_1449 (O_1449,N_29870,N_29800);
nor UO_1450 (O_1450,N_29875,N_29961);
nand UO_1451 (O_1451,N_29884,N_29882);
and UO_1452 (O_1452,N_29861,N_29906);
nand UO_1453 (O_1453,N_29968,N_29938);
nand UO_1454 (O_1454,N_29831,N_29864);
or UO_1455 (O_1455,N_29952,N_29973);
and UO_1456 (O_1456,N_29953,N_29908);
nor UO_1457 (O_1457,N_29872,N_29962);
nor UO_1458 (O_1458,N_29930,N_29962);
nor UO_1459 (O_1459,N_29956,N_29957);
nor UO_1460 (O_1460,N_29827,N_29933);
nand UO_1461 (O_1461,N_29848,N_29843);
and UO_1462 (O_1462,N_29871,N_29993);
and UO_1463 (O_1463,N_29910,N_29995);
xor UO_1464 (O_1464,N_29895,N_29871);
and UO_1465 (O_1465,N_29959,N_29976);
xor UO_1466 (O_1466,N_29810,N_29904);
and UO_1467 (O_1467,N_29966,N_29861);
nor UO_1468 (O_1468,N_29905,N_29817);
nand UO_1469 (O_1469,N_29996,N_29899);
xnor UO_1470 (O_1470,N_29863,N_29842);
and UO_1471 (O_1471,N_29921,N_29887);
or UO_1472 (O_1472,N_29885,N_29804);
nand UO_1473 (O_1473,N_29890,N_29884);
and UO_1474 (O_1474,N_29870,N_29808);
or UO_1475 (O_1475,N_29992,N_29985);
and UO_1476 (O_1476,N_29835,N_29963);
and UO_1477 (O_1477,N_29885,N_29853);
xor UO_1478 (O_1478,N_29983,N_29884);
nor UO_1479 (O_1479,N_29919,N_29829);
or UO_1480 (O_1480,N_29943,N_29868);
nor UO_1481 (O_1481,N_29943,N_29944);
and UO_1482 (O_1482,N_29999,N_29985);
or UO_1483 (O_1483,N_29807,N_29842);
or UO_1484 (O_1484,N_29850,N_29935);
xnor UO_1485 (O_1485,N_29850,N_29922);
xnor UO_1486 (O_1486,N_29901,N_29922);
nand UO_1487 (O_1487,N_29869,N_29941);
nor UO_1488 (O_1488,N_29932,N_29890);
and UO_1489 (O_1489,N_29844,N_29953);
nand UO_1490 (O_1490,N_29808,N_29946);
nand UO_1491 (O_1491,N_29907,N_29821);
and UO_1492 (O_1492,N_29999,N_29891);
nand UO_1493 (O_1493,N_29944,N_29843);
nand UO_1494 (O_1494,N_29890,N_29878);
and UO_1495 (O_1495,N_29899,N_29846);
or UO_1496 (O_1496,N_29934,N_29807);
xnor UO_1497 (O_1497,N_29803,N_29880);
nor UO_1498 (O_1498,N_29994,N_29877);
xor UO_1499 (O_1499,N_29853,N_29866);
and UO_1500 (O_1500,N_29992,N_29865);
nor UO_1501 (O_1501,N_29984,N_29977);
nor UO_1502 (O_1502,N_29895,N_29998);
and UO_1503 (O_1503,N_29995,N_29935);
nor UO_1504 (O_1504,N_29998,N_29848);
and UO_1505 (O_1505,N_29941,N_29938);
and UO_1506 (O_1506,N_29974,N_29941);
xor UO_1507 (O_1507,N_29837,N_29819);
and UO_1508 (O_1508,N_29965,N_29868);
xnor UO_1509 (O_1509,N_29917,N_29989);
and UO_1510 (O_1510,N_29993,N_29921);
nor UO_1511 (O_1511,N_29846,N_29815);
nand UO_1512 (O_1512,N_29941,N_29825);
nor UO_1513 (O_1513,N_29812,N_29995);
nand UO_1514 (O_1514,N_29850,N_29947);
nor UO_1515 (O_1515,N_29878,N_29924);
xor UO_1516 (O_1516,N_29875,N_29924);
nand UO_1517 (O_1517,N_29831,N_29984);
nor UO_1518 (O_1518,N_29980,N_29836);
nor UO_1519 (O_1519,N_29844,N_29961);
xor UO_1520 (O_1520,N_29917,N_29894);
or UO_1521 (O_1521,N_29911,N_29907);
nand UO_1522 (O_1522,N_29937,N_29911);
nand UO_1523 (O_1523,N_29912,N_29808);
nand UO_1524 (O_1524,N_29937,N_29984);
and UO_1525 (O_1525,N_29985,N_29930);
and UO_1526 (O_1526,N_29908,N_29903);
nand UO_1527 (O_1527,N_29837,N_29973);
and UO_1528 (O_1528,N_29857,N_29976);
nor UO_1529 (O_1529,N_29863,N_29970);
and UO_1530 (O_1530,N_29832,N_29941);
and UO_1531 (O_1531,N_29939,N_29963);
xor UO_1532 (O_1532,N_29992,N_29884);
and UO_1533 (O_1533,N_29880,N_29930);
or UO_1534 (O_1534,N_29974,N_29879);
and UO_1535 (O_1535,N_29802,N_29866);
nor UO_1536 (O_1536,N_29984,N_29881);
nor UO_1537 (O_1537,N_29975,N_29968);
nor UO_1538 (O_1538,N_29840,N_29930);
nand UO_1539 (O_1539,N_29940,N_29889);
xnor UO_1540 (O_1540,N_29900,N_29901);
nand UO_1541 (O_1541,N_29882,N_29857);
nor UO_1542 (O_1542,N_29812,N_29939);
or UO_1543 (O_1543,N_29893,N_29804);
or UO_1544 (O_1544,N_29902,N_29853);
xnor UO_1545 (O_1545,N_29966,N_29999);
nand UO_1546 (O_1546,N_29926,N_29913);
or UO_1547 (O_1547,N_29947,N_29929);
xnor UO_1548 (O_1548,N_29929,N_29885);
xor UO_1549 (O_1549,N_29961,N_29994);
xor UO_1550 (O_1550,N_29940,N_29969);
or UO_1551 (O_1551,N_29884,N_29964);
and UO_1552 (O_1552,N_29946,N_29916);
xnor UO_1553 (O_1553,N_29971,N_29824);
nor UO_1554 (O_1554,N_29928,N_29978);
nor UO_1555 (O_1555,N_29890,N_29887);
nand UO_1556 (O_1556,N_29807,N_29950);
nand UO_1557 (O_1557,N_29827,N_29975);
nand UO_1558 (O_1558,N_29818,N_29934);
or UO_1559 (O_1559,N_29876,N_29845);
or UO_1560 (O_1560,N_29851,N_29830);
nor UO_1561 (O_1561,N_29987,N_29919);
xnor UO_1562 (O_1562,N_29947,N_29827);
or UO_1563 (O_1563,N_29810,N_29869);
or UO_1564 (O_1564,N_29949,N_29846);
xor UO_1565 (O_1565,N_29886,N_29862);
nand UO_1566 (O_1566,N_29924,N_29930);
or UO_1567 (O_1567,N_29958,N_29984);
and UO_1568 (O_1568,N_29808,N_29806);
nand UO_1569 (O_1569,N_29865,N_29825);
nand UO_1570 (O_1570,N_29881,N_29961);
xor UO_1571 (O_1571,N_29973,N_29862);
xnor UO_1572 (O_1572,N_29803,N_29911);
or UO_1573 (O_1573,N_29949,N_29931);
and UO_1574 (O_1574,N_29955,N_29806);
xor UO_1575 (O_1575,N_29913,N_29891);
and UO_1576 (O_1576,N_29871,N_29882);
xnor UO_1577 (O_1577,N_29979,N_29847);
nand UO_1578 (O_1578,N_29928,N_29860);
or UO_1579 (O_1579,N_29891,N_29854);
or UO_1580 (O_1580,N_29813,N_29880);
and UO_1581 (O_1581,N_29852,N_29977);
nand UO_1582 (O_1582,N_29957,N_29813);
or UO_1583 (O_1583,N_29856,N_29958);
xnor UO_1584 (O_1584,N_29881,N_29957);
and UO_1585 (O_1585,N_29904,N_29988);
and UO_1586 (O_1586,N_29902,N_29810);
nor UO_1587 (O_1587,N_29815,N_29971);
and UO_1588 (O_1588,N_29988,N_29912);
nor UO_1589 (O_1589,N_29899,N_29893);
nor UO_1590 (O_1590,N_29817,N_29934);
nor UO_1591 (O_1591,N_29974,N_29880);
or UO_1592 (O_1592,N_29971,N_29849);
xnor UO_1593 (O_1593,N_29804,N_29922);
or UO_1594 (O_1594,N_29894,N_29936);
and UO_1595 (O_1595,N_29861,N_29934);
or UO_1596 (O_1596,N_29829,N_29882);
nor UO_1597 (O_1597,N_29913,N_29869);
nor UO_1598 (O_1598,N_29890,N_29921);
or UO_1599 (O_1599,N_29867,N_29938);
nand UO_1600 (O_1600,N_29888,N_29865);
nand UO_1601 (O_1601,N_29907,N_29811);
nand UO_1602 (O_1602,N_29803,N_29912);
or UO_1603 (O_1603,N_29978,N_29909);
nand UO_1604 (O_1604,N_29924,N_29885);
xor UO_1605 (O_1605,N_29812,N_29988);
nand UO_1606 (O_1606,N_29910,N_29892);
nand UO_1607 (O_1607,N_29999,N_29874);
and UO_1608 (O_1608,N_29838,N_29923);
nand UO_1609 (O_1609,N_29821,N_29868);
xor UO_1610 (O_1610,N_29945,N_29956);
nor UO_1611 (O_1611,N_29994,N_29923);
nor UO_1612 (O_1612,N_29901,N_29861);
xor UO_1613 (O_1613,N_29921,N_29979);
nand UO_1614 (O_1614,N_29999,N_29826);
xnor UO_1615 (O_1615,N_29897,N_29817);
xnor UO_1616 (O_1616,N_29977,N_29933);
nor UO_1617 (O_1617,N_29820,N_29814);
xor UO_1618 (O_1618,N_29865,N_29819);
nand UO_1619 (O_1619,N_29968,N_29802);
nor UO_1620 (O_1620,N_29893,N_29939);
and UO_1621 (O_1621,N_29853,N_29849);
or UO_1622 (O_1622,N_29851,N_29869);
nand UO_1623 (O_1623,N_29872,N_29912);
xnor UO_1624 (O_1624,N_29976,N_29828);
xor UO_1625 (O_1625,N_29831,N_29882);
nor UO_1626 (O_1626,N_29958,N_29995);
nor UO_1627 (O_1627,N_29841,N_29894);
xnor UO_1628 (O_1628,N_29924,N_29997);
or UO_1629 (O_1629,N_29882,N_29968);
and UO_1630 (O_1630,N_29887,N_29861);
nor UO_1631 (O_1631,N_29823,N_29922);
or UO_1632 (O_1632,N_29923,N_29842);
and UO_1633 (O_1633,N_29907,N_29972);
nor UO_1634 (O_1634,N_29873,N_29800);
and UO_1635 (O_1635,N_29894,N_29957);
nand UO_1636 (O_1636,N_29943,N_29982);
and UO_1637 (O_1637,N_29938,N_29874);
nand UO_1638 (O_1638,N_29881,N_29979);
nand UO_1639 (O_1639,N_29859,N_29904);
nor UO_1640 (O_1640,N_29936,N_29848);
and UO_1641 (O_1641,N_29845,N_29976);
nor UO_1642 (O_1642,N_29939,N_29802);
and UO_1643 (O_1643,N_29844,N_29883);
xor UO_1644 (O_1644,N_29990,N_29810);
nor UO_1645 (O_1645,N_29999,N_29989);
and UO_1646 (O_1646,N_29918,N_29925);
nor UO_1647 (O_1647,N_29938,N_29935);
xnor UO_1648 (O_1648,N_29849,N_29989);
or UO_1649 (O_1649,N_29841,N_29903);
xor UO_1650 (O_1650,N_29867,N_29899);
nor UO_1651 (O_1651,N_29958,N_29897);
and UO_1652 (O_1652,N_29842,N_29915);
or UO_1653 (O_1653,N_29944,N_29976);
nand UO_1654 (O_1654,N_29941,N_29929);
nor UO_1655 (O_1655,N_29903,N_29909);
nand UO_1656 (O_1656,N_29921,N_29817);
and UO_1657 (O_1657,N_29928,N_29998);
nor UO_1658 (O_1658,N_29824,N_29823);
nand UO_1659 (O_1659,N_29919,N_29910);
xnor UO_1660 (O_1660,N_29800,N_29948);
nand UO_1661 (O_1661,N_29824,N_29873);
xor UO_1662 (O_1662,N_29951,N_29964);
nor UO_1663 (O_1663,N_29982,N_29832);
and UO_1664 (O_1664,N_29871,N_29877);
xor UO_1665 (O_1665,N_29964,N_29922);
and UO_1666 (O_1666,N_29865,N_29840);
or UO_1667 (O_1667,N_29952,N_29804);
nand UO_1668 (O_1668,N_29933,N_29947);
and UO_1669 (O_1669,N_29865,N_29973);
xor UO_1670 (O_1670,N_29949,N_29880);
nor UO_1671 (O_1671,N_29888,N_29833);
or UO_1672 (O_1672,N_29859,N_29875);
xnor UO_1673 (O_1673,N_29886,N_29869);
nand UO_1674 (O_1674,N_29922,N_29993);
nor UO_1675 (O_1675,N_29808,N_29944);
or UO_1676 (O_1676,N_29800,N_29996);
or UO_1677 (O_1677,N_29836,N_29981);
or UO_1678 (O_1678,N_29917,N_29859);
nor UO_1679 (O_1679,N_29816,N_29863);
nand UO_1680 (O_1680,N_29985,N_29978);
nand UO_1681 (O_1681,N_29928,N_29923);
or UO_1682 (O_1682,N_29933,N_29937);
nor UO_1683 (O_1683,N_29977,N_29967);
nand UO_1684 (O_1684,N_29991,N_29871);
nor UO_1685 (O_1685,N_29961,N_29914);
xor UO_1686 (O_1686,N_29956,N_29954);
nor UO_1687 (O_1687,N_29817,N_29935);
nand UO_1688 (O_1688,N_29951,N_29825);
and UO_1689 (O_1689,N_29952,N_29954);
or UO_1690 (O_1690,N_29896,N_29924);
xnor UO_1691 (O_1691,N_29895,N_29978);
nand UO_1692 (O_1692,N_29990,N_29970);
nor UO_1693 (O_1693,N_29822,N_29981);
xor UO_1694 (O_1694,N_29916,N_29956);
or UO_1695 (O_1695,N_29960,N_29851);
xor UO_1696 (O_1696,N_29920,N_29902);
or UO_1697 (O_1697,N_29911,N_29950);
xnor UO_1698 (O_1698,N_29952,N_29881);
or UO_1699 (O_1699,N_29954,N_29959);
and UO_1700 (O_1700,N_29934,N_29965);
nor UO_1701 (O_1701,N_29833,N_29804);
and UO_1702 (O_1702,N_29939,N_29801);
or UO_1703 (O_1703,N_29888,N_29885);
or UO_1704 (O_1704,N_29939,N_29965);
and UO_1705 (O_1705,N_29902,N_29958);
and UO_1706 (O_1706,N_29880,N_29872);
and UO_1707 (O_1707,N_29801,N_29818);
xor UO_1708 (O_1708,N_29831,N_29953);
nor UO_1709 (O_1709,N_29975,N_29917);
nand UO_1710 (O_1710,N_29981,N_29823);
xnor UO_1711 (O_1711,N_29849,N_29887);
nor UO_1712 (O_1712,N_29902,N_29974);
nor UO_1713 (O_1713,N_29857,N_29816);
or UO_1714 (O_1714,N_29810,N_29949);
nand UO_1715 (O_1715,N_29885,N_29936);
nor UO_1716 (O_1716,N_29876,N_29975);
xnor UO_1717 (O_1717,N_29820,N_29945);
nand UO_1718 (O_1718,N_29853,N_29953);
nor UO_1719 (O_1719,N_29827,N_29941);
and UO_1720 (O_1720,N_29906,N_29966);
and UO_1721 (O_1721,N_29919,N_29911);
nor UO_1722 (O_1722,N_29811,N_29922);
nor UO_1723 (O_1723,N_29946,N_29812);
nor UO_1724 (O_1724,N_29945,N_29818);
nand UO_1725 (O_1725,N_29872,N_29928);
xnor UO_1726 (O_1726,N_29817,N_29894);
xor UO_1727 (O_1727,N_29872,N_29956);
or UO_1728 (O_1728,N_29968,N_29839);
nor UO_1729 (O_1729,N_29933,N_29967);
and UO_1730 (O_1730,N_29869,N_29843);
nor UO_1731 (O_1731,N_29906,N_29976);
or UO_1732 (O_1732,N_29875,N_29867);
xor UO_1733 (O_1733,N_29990,N_29917);
and UO_1734 (O_1734,N_29860,N_29979);
nor UO_1735 (O_1735,N_29931,N_29919);
or UO_1736 (O_1736,N_29962,N_29873);
xor UO_1737 (O_1737,N_29803,N_29910);
xor UO_1738 (O_1738,N_29885,N_29822);
xnor UO_1739 (O_1739,N_29870,N_29907);
nand UO_1740 (O_1740,N_29941,N_29815);
nor UO_1741 (O_1741,N_29918,N_29966);
and UO_1742 (O_1742,N_29881,N_29951);
nor UO_1743 (O_1743,N_29937,N_29914);
and UO_1744 (O_1744,N_29973,N_29937);
nor UO_1745 (O_1745,N_29888,N_29913);
nand UO_1746 (O_1746,N_29812,N_29869);
and UO_1747 (O_1747,N_29843,N_29809);
nor UO_1748 (O_1748,N_29933,N_29886);
and UO_1749 (O_1749,N_29809,N_29823);
nand UO_1750 (O_1750,N_29920,N_29933);
or UO_1751 (O_1751,N_29872,N_29805);
or UO_1752 (O_1752,N_29982,N_29804);
nand UO_1753 (O_1753,N_29870,N_29804);
xor UO_1754 (O_1754,N_29945,N_29965);
nand UO_1755 (O_1755,N_29843,N_29990);
nor UO_1756 (O_1756,N_29825,N_29935);
and UO_1757 (O_1757,N_29823,N_29954);
xnor UO_1758 (O_1758,N_29937,N_29909);
or UO_1759 (O_1759,N_29937,N_29974);
xor UO_1760 (O_1760,N_29963,N_29858);
and UO_1761 (O_1761,N_29946,N_29852);
nor UO_1762 (O_1762,N_29920,N_29879);
nor UO_1763 (O_1763,N_29901,N_29910);
xor UO_1764 (O_1764,N_29888,N_29827);
nor UO_1765 (O_1765,N_29863,N_29857);
or UO_1766 (O_1766,N_29888,N_29936);
xor UO_1767 (O_1767,N_29907,N_29910);
xnor UO_1768 (O_1768,N_29862,N_29978);
nand UO_1769 (O_1769,N_29874,N_29965);
and UO_1770 (O_1770,N_29826,N_29902);
and UO_1771 (O_1771,N_29862,N_29972);
and UO_1772 (O_1772,N_29947,N_29912);
xor UO_1773 (O_1773,N_29946,N_29888);
and UO_1774 (O_1774,N_29946,N_29883);
nand UO_1775 (O_1775,N_29952,N_29892);
and UO_1776 (O_1776,N_29932,N_29872);
or UO_1777 (O_1777,N_29927,N_29900);
nor UO_1778 (O_1778,N_29868,N_29882);
or UO_1779 (O_1779,N_29892,N_29907);
nand UO_1780 (O_1780,N_29817,N_29918);
and UO_1781 (O_1781,N_29899,N_29891);
and UO_1782 (O_1782,N_29962,N_29807);
or UO_1783 (O_1783,N_29827,N_29963);
nand UO_1784 (O_1784,N_29824,N_29937);
nor UO_1785 (O_1785,N_29821,N_29850);
or UO_1786 (O_1786,N_29841,N_29832);
nand UO_1787 (O_1787,N_29961,N_29969);
nand UO_1788 (O_1788,N_29958,N_29874);
or UO_1789 (O_1789,N_29926,N_29855);
xor UO_1790 (O_1790,N_29893,N_29995);
or UO_1791 (O_1791,N_29942,N_29896);
xor UO_1792 (O_1792,N_29890,N_29974);
nor UO_1793 (O_1793,N_29936,N_29804);
and UO_1794 (O_1794,N_29987,N_29833);
and UO_1795 (O_1795,N_29965,N_29800);
and UO_1796 (O_1796,N_29928,N_29956);
xor UO_1797 (O_1797,N_29802,N_29916);
xnor UO_1798 (O_1798,N_29831,N_29888);
xnor UO_1799 (O_1799,N_29804,N_29921);
nand UO_1800 (O_1800,N_29857,N_29835);
nor UO_1801 (O_1801,N_29810,N_29913);
xor UO_1802 (O_1802,N_29932,N_29976);
nand UO_1803 (O_1803,N_29992,N_29837);
or UO_1804 (O_1804,N_29915,N_29909);
nand UO_1805 (O_1805,N_29869,N_29904);
or UO_1806 (O_1806,N_29832,N_29881);
and UO_1807 (O_1807,N_29944,N_29902);
nor UO_1808 (O_1808,N_29965,N_29969);
nand UO_1809 (O_1809,N_29901,N_29936);
or UO_1810 (O_1810,N_29962,N_29965);
or UO_1811 (O_1811,N_29896,N_29992);
or UO_1812 (O_1812,N_29839,N_29844);
xnor UO_1813 (O_1813,N_29878,N_29891);
nor UO_1814 (O_1814,N_29994,N_29883);
nor UO_1815 (O_1815,N_29855,N_29934);
nor UO_1816 (O_1816,N_29969,N_29841);
and UO_1817 (O_1817,N_29838,N_29864);
xor UO_1818 (O_1818,N_29966,N_29825);
and UO_1819 (O_1819,N_29871,N_29828);
nor UO_1820 (O_1820,N_29895,N_29870);
or UO_1821 (O_1821,N_29955,N_29855);
nand UO_1822 (O_1822,N_29976,N_29863);
nor UO_1823 (O_1823,N_29926,N_29849);
nand UO_1824 (O_1824,N_29880,N_29857);
or UO_1825 (O_1825,N_29965,N_29966);
nand UO_1826 (O_1826,N_29923,N_29841);
nor UO_1827 (O_1827,N_29905,N_29846);
xor UO_1828 (O_1828,N_29940,N_29891);
and UO_1829 (O_1829,N_29997,N_29977);
xnor UO_1830 (O_1830,N_29926,N_29856);
nor UO_1831 (O_1831,N_29864,N_29843);
nor UO_1832 (O_1832,N_29941,N_29811);
or UO_1833 (O_1833,N_29919,N_29848);
nor UO_1834 (O_1834,N_29852,N_29812);
nand UO_1835 (O_1835,N_29980,N_29886);
or UO_1836 (O_1836,N_29987,N_29969);
nand UO_1837 (O_1837,N_29850,N_29931);
nor UO_1838 (O_1838,N_29961,N_29874);
and UO_1839 (O_1839,N_29863,N_29960);
xor UO_1840 (O_1840,N_29891,N_29848);
nand UO_1841 (O_1841,N_29842,N_29853);
and UO_1842 (O_1842,N_29898,N_29895);
or UO_1843 (O_1843,N_29844,N_29851);
nor UO_1844 (O_1844,N_29873,N_29819);
nand UO_1845 (O_1845,N_29898,N_29836);
and UO_1846 (O_1846,N_29882,N_29895);
or UO_1847 (O_1847,N_29948,N_29972);
nor UO_1848 (O_1848,N_29823,N_29865);
or UO_1849 (O_1849,N_29855,N_29819);
or UO_1850 (O_1850,N_29806,N_29987);
and UO_1851 (O_1851,N_29882,N_29927);
xor UO_1852 (O_1852,N_29805,N_29912);
or UO_1853 (O_1853,N_29974,N_29862);
and UO_1854 (O_1854,N_29867,N_29988);
xnor UO_1855 (O_1855,N_29906,N_29952);
xor UO_1856 (O_1856,N_29949,N_29853);
nand UO_1857 (O_1857,N_29943,N_29826);
nand UO_1858 (O_1858,N_29862,N_29935);
and UO_1859 (O_1859,N_29947,N_29898);
xnor UO_1860 (O_1860,N_29969,N_29832);
nor UO_1861 (O_1861,N_29858,N_29814);
and UO_1862 (O_1862,N_29909,N_29861);
or UO_1863 (O_1863,N_29959,N_29973);
nor UO_1864 (O_1864,N_29976,N_29849);
and UO_1865 (O_1865,N_29974,N_29866);
nor UO_1866 (O_1866,N_29908,N_29907);
nor UO_1867 (O_1867,N_29891,N_29828);
xor UO_1868 (O_1868,N_29985,N_29933);
and UO_1869 (O_1869,N_29899,N_29972);
nor UO_1870 (O_1870,N_29952,N_29967);
xnor UO_1871 (O_1871,N_29857,N_29986);
xnor UO_1872 (O_1872,N_29935,N_29916);
nand UO_1873 (O_1873,N_29849,N_29867);
or UO_1874 (O_1874,N_29927,N_29863);
nand UO_1875 (O_1875,N_29989,N_29848);
or UO_1876 (O_1876,N_29846,N_29876);
or UO_1877 (O_1877,N_29833,N_29805);
nand UO_1878 (O_1878,N_29800,N_29820);
nor UO_1879 (O_1879,N_29862,N_29870);
xor UO_1880 (O_1880,N_29934,N_29999);
nor UO_1881 (O_1881,N_29882,N_29955);
or UO_1882 (O_1882,N_29857,N_29967);
or UO_1883 (O_1883,N_29941,N_29943);
nand UO_1884 (O_1884,N_29811,N_29993);
xor UO_1885 (O_1885,N_29921,N_29905);
and UO_1886 (O_1886,N_29843,N_29900);
xor UO_1887 (O_1887,N_29867,N_29925);
nand UO_1888 (O_1888,N_29893,N_29922);
nand UO_1889 (O_1889,N_29919,N_29856);
nor UO_1890 (O_1890,N_29888,N_29814);
and UO_1891 (O_1891,N_29952,N_29880);
and UO_1892 (O_1892,N_29991,N_29851);
nor UO_1893 (O_1893,N_29854,N_29932);
or UO_1894 (O_1894,N_29973,N_29851);
nand UO_1895 (O_1895,N_29972,N_29802);
xnor UO_1896 (O_1896,N_29952,N_29872);
and UO_1897 (O_1897,N_29924,N_29892);
and UO_1898 (O_1898,N_29906,N_29942);
nand UO_1899 (O_1899,N_29874,N_29988);
nor UO_1900 (O_1900,N_29831,N_29899);
nand UO_1901 (O_1901,N_29897,N_29824);
and UO_1902 (O_1902,N_29809,N_29881);
xor UO_1903 (O_1903,N_29889,N_29863);
nand UO_1904 (O_1904,N_29931,N_29822);
nor UO_1905 (O_1905,N_29882,N_29920);
xor UO_1906 (O_1906,N_29955,N_29950);
xnor UO_1907 (O_1907,N_29961,N_29941);
nand UO_1908 (O_1908,N_29957,N_29978);
or UO_1909 (O_1909,N_29905,N_29910);
xor UO_1910 (O_1910,N_29926,N_29836);
xor UO_1911 (O_1911,N_29939,N_29975);
xnor UO_1912 (O_1912,N_29906,N_29849);
xor UO_1913 (O_1913,N_29881,N_29839);
xor UO_1914 (O_1914,N_29981,N_29991);
or UO_1915 (O_1915,N_29874,N_29824);
or UO_1916 (O_1916,N_29805,N_29881);
or UO_1917 (O_1917,N_29931,N_29861);
nand UO_1918 (O_1918,N_29989,N_29940);
nand UO_1919 (O_1919,N_29922,N_29894);
nand UO_1920 (O_1920,N_29803,N_29975);
or UO_1921 (O_1921,N_29892,N_29837);
and UO_1922 (O_1922,N_29824,N_29956);
nor UO_1923 (O_1923,N_29966,N_29996);
and UO_1924 (O_1924,N_29950,N_29831);
xnor UO_1925 (O_1925,N_29946,N_29810);
nor UO_1926 (O_1926,N_29860,N_29832);
xnor UO_1927 (O_1927,N_29870,N_29916);
and UO_1928 (O_1928,N_29842,N_29968);
or UO_1929 (O_1929,N_29813,N_29879);
nor UO_1930 (O_1930,N_29815,N_29933);
nand UO_1931 (O_1931,N_29845,N_29942);
or UO_1932 (O_1932,N_29873,N_29910);
or UO_1933 (O_1933,N_29932,N_29991);
and UO_1934 (O_1934,N_29971,N_29941);
and UO_1935 (O_1935,N_29983,N_29888);
nor UO_1936 (O_1936,N_29890,N_29882);
xnor UO_1937 (O_1937,N_29989,N_29870);
or UO_1938 (O_1938,N_29965,N_29920);
nor UO_1939 (O_1939,N_29939,N_29901);
nand UO_1940 (O_1940,N_29926,N_29898);
or UO_1941 (O_1941,N_29890,N_29912);
nor UO_1942 (O_1942,N_29928,N_29950);
xor UO_1943 (O_1943,N_29887,N_29814);
xnor UO_1944 (O_1944,N_29840,N_29833);
or UO_1945 (O_1945,N_29893,N_29838);
nand UO_1946 (O_1946,N_29899,N_29962);
xor UO_1947 (O_1947,N_29928,N_29937);
or UO_1948 (O_1948,N_29908,N_29882);
nand UO_1949 (O_1949,N_29986,N_29870);
or UO_1950 (O_1950,N_29976,N_29833);
and UO_1951 (O_1951,N_29959,N_29855);
and UO_1952 (O_1952,N_29839,N_29934);
or UO_1953 (O_1953,N_29844,N_29838);
nor UO_1954 (O_1954,N_29836,N_29960);
and UO_1955 (O_1955,N_29946,N_29926);
xnor UO_1956 (O_1956,N_29868,N_29854);
xor UO_1957 (O_1957,N_29959,N_29978);
or UO_1958 (O_1958,N_29893,N_29820);
xor UO_1959 (O_1959,N_29844,N_29863);
or UO_1960 (O_1960,N_29852,N_29970);
xor UO_1961 (O_1961,N_29960,N_29988);
xor UO_1962 (O_1962,N_29960,N_29910);
and UO_1963 (O_1963,N_29969,N_29992);
and UO_1964 (O_1964,N_29962,N_29902);
and UO_1965 (O_1965,N_29834,N_29910);
xor UO_1966 (O_1966,N_29881,N_29918);
nand UO_1967 (O_1967,N_29991,N_29837);
or UO_1968 (O_1968,N_29861,N_29960);
or UO_1969 (O_1969,N_29951,N_29937);
xor UO_1970 (O_1970,N_29977,N_29803);
and UO_1971 (O_1971,N_29848,N_29869);
xnor UO_1972 (O_1972,N_29868,N_29809);
nor UO_1973 (O_1973,N_29878,N_29866);
or UO_1974 (O_1974,N_29923,N_29814);
nand UO_1975 (O_1975,N_29811,N_29906);
nand UO_1976 (O_1976,N_29992,N_29988);
or UO_1977 (O_1977,N_29987,N_29840);
nand UO_1978 (O_1978,N_29954,N_29883);
xnor UO_1979 (O_1979,N_29882,N_29800);
or UO_1980 (O_1980,N_29875,N_29883);
nor UO_1981 (O_1981,N_29880,N_29945);
or UO_1982 (O_1982,N_29982,N_29817);
and UO_1983 (O_1983,N_29908,N_29844);
nor UO_1984 (O_1984,N_29944,N_29958);
xnor UO_1985 (O_1985,N_29804,N_29985);
or UO_1986 (O_1986,N_29958,N_29905);
and UO_1987 (O_1987,N_29859,N_29920);
nor UO_1988 (O_1988,N_29976,N_29867);
nor UO_1989 (O_1989,N_29891,N_29847);
nor UO_1990 (O_1990,N_29851,N_29823);
nand UO_1991 (O_1991,N_29808,N_29855);
nor UO_1992 (O_1992,N_29883,N_29999);
nor UO_1993 (O_1993,N_29873,N_29885);
xnor UO_1994 (O_1994,N_29888,N_29889);
nor UO_1995 (O_1995,N_29813,N_29990);
or UO_1996 (O_1996,N_29952,N_29853);
xnor UO_1997 (O_1997,N_29949,N_29983);
and UO_1998 (O_1998,N_29974,N_29844);
or UO_1999 (O_1999,N_29869,N_29979);
and UO_2000 (O_2000,N_29992,N_29997);
or UO_2001 (O_2001,N_29935,N_29972);
or UO_2002 (O_2002,N_29970,N_29981);
and UO_2003 (O_2003,N_29932,N_29973);
or UO_2004 (O_2004,N_29850,N_29879);
or UO_2005 (O_2005,N_29952,N_29893);
nand UO_2006 (O_2006,N_29933,N_29887);
or UO_2007 (O_2007,N_29880,N_29839);
nand UO_2008 (O_2008,N_29968,N_29997);
xor UO_2009 (O_2009,N_29840,N_29842);
and UO_2010 (O_2010,N_29969,N_29984);
xor UO_2011 (O_2011,N_29991,N_29973);
and UO_2012 (O_2012,N_29975,N_29851);
nor UO_2013 (O_2013,N_29947,N_29927);
nand UO_2014 (O_2014,N_29936,N_29984);
nor UO_2015 (O_2015,N_29932,N_29924);
nor UO_2016 (O_2016,N_29908,N_29861);
nor UO_2017 (O_2017,N_29983,N_29873);
nand UO_2018 (O_2018,N_29988,N_29886);
or UO_2019 (O_2019,N_29822,N_29838);
or UO_2020 (O_2020,N_29952,N_29966);
and UO_2021 (O_2021,N_29932,N_29881);
nor UO_2022 (O_2022,N_29802,N_29899);
nand UO_2023 (O_2023,N_29813,N_29861);
or UO_2024 (O_2024,N_29950,N_29947);
or UO_2025 (O_2025,N_29806,N_29901);
nor UO_2026 (O_2026,N_29930,N_29931);
or UO_2027 (O_2027,N_29819,N_29949);
or UO_2028 (O_2028,N_29911,N_29955);
xor UO_2029 (O_2029,N_29962,N_29878);
nand UO_2030 (O_2030,N_29990,N_29893);
xnor UO_2031 (O_2031,N_29910,N_29820);
nand UO_2032 (O_2032,N_29885,N_29891);
and UO_2033 (O_2033,N_29867,N_29878);
and UO_2034 (O_2034,N_29821,N_29946);
and UO_2035 (O_2035,N_29872,N_29949);
xor UO_2036 (O_2036,N_29808,N_29803);
nor UO_2037 (O_2037,N_29852,N_29891);
nand UO_2038 (O_2038,N_29889,N_29804);
or UO_2039 (O_2039,N_29922,N_29873);
nor UO_2040 (O_2040,N_29997,N_29869);
and UO_2041 (O_2041,N_29811,N_29896);
xor UO_2042 (O_2042,N_29826,N_29891);
nor UO_2043 (O_2043,N_29974,N_29994);
nand UO_2044 (O_2044,N_29937,N_29803);
or UO_2045 (O_2045,N_29885,N_29993);
nand UO_2046 (O_2046,N_29941,N_29835);
nand UO_2047 (O_2047,N_29969,N_29882);
and UO_2048 (O_2048,N_29952,N_29982);
nand UO_2049 (O_2049,N_29958,N_29885);
xor UO_2050 (O_2050,N_29913,N_29886);
or UO_2051 (O_2051,N_29811,N_29964);
and UO_2052 (O_2052,N_29852,N_29921);
xor UO_2053 (O_2053,N_29911,N_29877);
and UO_2054 (O_2054,N_29891,N_29827);
nand UO_2055 (O_2055,N_29812,N_29859);
and UO_2056 (O_2056,N_29993,N_29857);
and UO_2057 (O_2057,N_29900,N_29826);
or UO_2058 (O_2058,N_29885,N_29983);
nor UO_2059 (O_2059,N_29888,N_29854);
xor UO_2060 (O_2060,N_29925,N_29823);
and UO_2061 (O_2061,N_29996,N_29958);
xor UO_2062 (O_2062,N_29998,N_29882);
and UO_2063 (O_2063,N_29938,N_29877);
and UO_2064 (O_2064,N_29856,N_29881);
and UO_2065 (O_2065,N_29970,N_29979);
and UO_2066 (O_2066,N_29922,N_29877);
xor UO_2067 (O_2067,N_29987,N_29977);
and UO_2068 (O_2068,N_29993,N_29926);
nand UO_2069 (O_2069,N_29984,N_29993);
and UO_2070 (O_2070,N_29858,N_29873);
and UO_2071 (O_2071,N_29966,N_29905);
xor UO_2072 (O_2072,N_29993,N_29837);
and UO_2073 (O_2073,N_29983,N_29875);
and UO_2074 (O_2074,N_29904,N_29989);
nand UO_2075 (O_2075,N_29971,N_29931);
and UO_2076 (O_2076,N_29868,N_29867);
xor UO_2077 (O_2077,N_29939,N_29988);
or UO_2078 (O_2078,N_29982,N_29967);
nand UO_2079 (O_2079,N_29986,N_29862);
nand UO_2080 (O_2080,N_29887,N_29995);
and UO_2081 (O_2081,N_29928,N_29969);
nor UO_2082 (O_2082,N_29882,N_29991);
nor UO_2083 (O_2083,N_29942,N_29819);
nand UO_2084 (O_2084,N_29998,N_29840);
nor UO_2085 (O_2085,N_29980,N_29853);
and UO_2086 (O_2086,N_29879,N_29902);
xnor UO_2087 (O_2087,N_29969,N_29995);
or UO_2088 (O_2088,N_29843,N_29870);
or UO_2089 (O_2089,N_29835,N_29855);
or UO_2090 (O_2090,N_29858,N_29914);
nand UO_2091 (O_2091,N_29878,N_29928);
xor UO_2092 (O_2092,N_29930,N_29875);
xnor UO_2093 (O_2093,N_29949,N_29932);
or UO_2094 (O_2094,N_29868,N_29865);
nand UO_2095 (O_2095,N_29856,N_29842);
or UO_2096 (O_2096,N_29991,N_29922);
nand UO_2097 (O_2097,N_29979,N_29951);
and UO_2098 (O_2098,N_29916,N_29910);
xor UO_2099 (O_2099,N_29860,N_29910);
and UO_2100 (O_2100,N_29888,N_29982);
or UO_2101 (O_2101,N_29966,N_29979);
and UO_2102 (O_2102,N_29912,N_29870);
nand UO_2103 (O_2103,N_29943,N_29846);
nand UO_2104 (O_2104,N_29902,N_29975);
nand UO_2105 (O_2105,N_29857,N_29941);
nor UO_2106 (O_2106,N_29813,N_29890);
and UO_2107 (O_2107,N_29934,N_29935);
and UO_2108 (O_2108,N_29843,N_29948);
nand UO_2109 (O_2109,N_29833,N_29965);
xor UO_2110 (O_2110,N_29904,N_29850);
xor UO_2111 (O_2111,N_29902,N_29913);
xor UO_2112 (O_2112,N_29815,N_29825);
or UO_2113 (O_2113,N_29993,N_29939);
nor UO_2114 (O_2114,N_29809,N_29962);
nand UO_2115 (O_2115,N_29961,N_29890);
or UO_2116 (O_2116,N_29873,N_29950);
and UO_2117 (O_2117,N_29912,N_29919);
xnor UO_2118 (O_2118,N_29984,N_29979);
or UO_2119 (O_2119,N_29976,N_29807);
nand UO_2120 (O_2120,N_29899,N_29938);
xor UO_2121 (O_2121,N_29919,N_29831);
xnor UO_2122 (O_2122,N_29947,N_29896);
and UO_2123 (O_2123,N_29808,N_29884);
nand UO_2124 (O_2124,N_29986,N_29888);
xnor UO_2125 (O_2125,N_29843,N_29901);
or UO_2126 (O_2126,N_29848,N_29883);
or UO_2127 (O_2127,N_29918,N_29810);
xnor UO_2128 (O_2128,N_29877,N_29937);
or UO_2129 (O_2129,N_29933,N_29900);
or UO_2130 (O_2130,N_29965,N_29839);
nor UO_2131 (O_2131,N_29888,N_29997);
and UO_2132 (O_2132,N_29810,N_29960);
nor UO_2133 (O_2133,N_29868,N_29986);
or UO_2134 (O_2134,N_29897,N_29907);
nor UO_2135 (O_2135,N_29893,N_29851);
xor UO_2136 (O_2136,N_29936,N_29985);
nand UO_2137 (O_2137,N_29977,N_29941);
and UO_2138 (O_2138,N_29914,N_29987);
nor UO_2139 (O_2139,N_29820,N_29892);
and UO_2140 (O_2140,N_29820,N_29958);
nor UO_2141 (O_2141,N_29909,N_29982);
and UO_2142 (O_2142,N_29830,N_29913);
nor UO_2143 (O_2143,N_29989,N_29826);
nand UO_2144 (O_2144,N_29922,N_29829);
or UO_2145 (O_2145,N_29969,N_29848);
or UO_2146 (O_2146,N_29939,N_29884);
and UO_2147 (O_2147,N_29923,N_29977);
or UO_2148 (O_2148,N_29975,N_29989);
nand UO_2149 (O_2149,N_29983,N_29917);
or UO_2150 (O_2150,N_29978,N_29859);
or UO_2151 (O_2151,N_29816,N_29934);
xor UO_2152 (O_2152,N_29930,N_29813);
and UO_2153 (O_2153,N_29919,N_29845);
or UO_2154 (O_2154,N_29966,N_29846);
nand UO_2155 (O_2155,N_29963,N_29960);
xor UO_2156 (O_2156,N_29837,N_29851);
and UO_2157 (O_2157,N_29929,N_29810);
nor UO_2158 (O_2158,N_29869,N_29880);
nor UO_2159 (O_2159,N_29944,N_29893);
nand UO_2160 (O_2160,N_29868,N_29815);
or UO_2161 (O_2161,N_29914,N_29990);
and UO_2162 (O_2162,N_29942,N_29984);
nand UO_2163 (O_2163,N_29950,N_29983);
nand UO_2164 (O_2164,N_29851,N_29877);
xnor UO_2165 (O_2165,N_29863,N_29869);
and UO_2166 (O_2166,N_29865,N_29965);
nor UO_2167 (O_2167,N_29823,N_29843);
and UO_2168 (O_2168,N_29804,N_29963);
nand UO_2169 (O_2169,N_29846,N_29956);
and UO_2170 (O_2170,N_29927,N_29975);
nand UO_2171 (O_2171,N_29971,N_29816);
and UO_2172 (O_2172,N_29919,N_29815);
or UO_2173 (O_2173,N_29928,N_29979);
nand UO_2174 (O_2174,N_29823,N_29884);
and UO_2175 (O_2175,N_29808,N_29982);
or UO_2176 (O_2176,N_29864,N_29912);
nor UO_2177 (O_2177,N_29958,N_29881);
or UO_2178 (O_2178,N_29853,N_29819);
nand UO_2179 (O_2179,N_29998,N_29819);
nand UO_2180 (O_2180,N_29959,N_29817);
nand UO_2181 (O_2181,N_29864,N_29847);
nand UO_2182 (O_2182,N_29861,N_29862);
xor UO_2183 (O_2183,N_29930,N_29878);
xnor UO_2184 (O_2184,N_29990,N_29820);
or UO_2185 (O_2185,N_29999,N_29924);
nor UO_2186 (O_2186,N_29846,N_29866);
and UO_2187 (O_2187,N_29874,N_29813);
and UO_2188 (O_2188,N_29980,N_29996);
nor UO_2189 (O_2189,N_29801,N_29858);
and UO_2190 (O_2190,N_29987,N_29871);
nor UO_2191 (O_2191,N_29887,N_29830);
xnor UO_2192 (O_2192,N_29911,N_29846);
xor UO_2193 (O_2193,N_29981,N_29890);
xnor UO_2194 (O_2194,N_29996,N_29895);
and UO_2195 (O_2195,N_29800,N_29830);
nor UO_2196 (O_2196,N_29853,N_29844);
nand UO_2197 (O_2197,N_29935,N_29857);
or UO_2198 (O_2198,N_29970,N_29910);
and UO_2199 (O_2199,N_29854,N_29838);
or UO_2200 (O_2200,N_29880,N_29856);
and UO_2201 (O_2201,N_29802,N_29943);
nor UO_2202 (O_2202,N_29999,N_29843);
xnor UO_2203 (O_2203,N_29852,N_29929);
and UO_2204 (O_2204,N_29920,N_29909);
xnor UO_2205 (O_2205,N_29996,N_29967);
nor UO_2206 (O_2206,N_29982,N_29959);
and UO_2207 (O_2207,N_29940,N_29862);
nand UO_2208 (O_2208,N_29818,N_29924);
or UO_2209 (O_2209,N_29829,N_29887);
nor UO_2210 (O_2210,N_29933,N_29879);
xor UO_2211 (O_2211,N_29824,N_29883);
or UO_2212 (O_2212,N_29977,N_29831);
nor UO_2213 (O_2213,N_29825,N_29833);
nand UO_2214 (O_2214,N_29862,N_29882);
or UO_2215 (O_2215,N_29985,N_29982);
nand UO_2216 (O_2216,N_29948,N_29944);
nand UO_2217 (O_2217,N_29946,N_29840);
nor UO_2218 (O_2218,N_29851,N_29805);
xnor UO_2219 (O_2219,N_29920,N_29903);
or UO_2220 (O_2220,N_29911,N_29828);
and UO_2221 (O_2221,N_29901,N_29902);
nor UO_2222 (O_2222,N_29857,N_29995);
nand UO_2223 (O_2223,N_29926,N_29977);
and UO_2224 (O_2224,N_29912,N_29818);
and UO_2225 (O_2225,N_29984,N_29801);
nor UO_2226 (O_2226,N_29883,N_29905);
or UO_2227 (O_2227,N_29828,N_29899);
xnor UO_2228 (O_2228,N_29915,N_29809);
xnor UO_2229 (O_2229,N_29933,N_29840);
nor UO_2230 (O_2230,N_29832,N_29877);
xnor UO_2231 (O_2231,N_29818,N_29855);
nor UO_2232 (O_2232,N_29925,N_29934);
nand UO_2233 (O_2233,N_29998,N_29812);
xnor UO_2234 (O_2234,N_29805,N_29987);
nor UO_2235 (O_2235,N_29970,N_29908);
nand UO_2236 (O_2236,N_29898,N_29828);
or UO_2237 (O_2237,N_29831,N_29871);
or UO_2238 (O_2238,N_29823,N_29818);
nor UO_2239 (O_2239,N_29822,N_29961);
xor UO_2240 (O_2240,N_29889,N_29974);
and UO_2241 (O_2241,N_29918,N_29863);
or UO_2242 (O_2242,N_29856,N_29956);
or UO_2243 (O_2243,N_29800,N_29915);
and UO_2244 (O_2244,N_29958,N_29990);
nor UO_2245 (O_2245,N_29985,N_29824);
or UO_2246 (O_2246,N_29897,N_29888);
or UO_2247 (O_2247,N_29968,N_29862);
and UO_2248 (O_2248,N_29914,N_29967);
nor UO_2249 (O_2249,N_29882,N_29907);
or UO_2250 (O_2250,N_29913,N_29909);
nor UO_2251 (O_2251,N_29915,N_29910);
nor UO_2252 (O_2252,N_29889,N_29845);
xor UO_2253 (O_2253,N_29899,N_29875);
nor UO_2254 (O_2254,N_29931,N_29912);
xor UO_2255 (O_2255,N_29959,N_29807);
nand UO_2256 (O_2256,N_29842,N_29886);
nor UO_2257 (O_2257,N_29843,N_29884);
nand UO_2258 (O_2258,N_29849,N_29948);
xor UO_2259 (O_2259,N_29813,N_29940);
xor UO_2260 (O_2260,N_29936,N_29920);
nand UO_2261 (O_2261,N_29987,N_29966);
xnor UO_2262 (O_2262,N_29904,N_29913);
and UO_2263 (O_2263,N_29930,N_29913);
and UO_2264 (O_2264,N_29974,N_29842);
nand UO_2265 (O_2265,N_29928,N_29894);
nand UO_2266 (O_2266,N_29821,N_29867);
xnor UO_2267 (O_2267,N_29822,N_29839);
xor UO_2268 (O_2268,N_29804,N_29974);
and UO_2269 (O_2269,N_29894,N_29913);
nor UO_2270 (O_2270,N_29842,N_29812);
or UO_2271 (O_2271,N_29867,N_29935);
nor UO_2272 (O_2272,N_29953,N_29814);
nor UO_2273 (O_2273,N_29972,N_29876);
xor UO_2274 (O_2274,N_29903,N_29937);
nor UO_2275 (O_2275,N_29821,N_29967);
nor UO_2276 (O_2276,N_29884,N_29907);
or UO_2277 (O_2277,N_29822,N_29954);
xor UO_2278 (O_2278,N_29824,N_29930);
xor UO_2279 (O_2279,N_29978,N_29892);
and UO_2280 (O_2280,N_29952,N_29960);
nand UO_2281 (O_2281,N_29857,N_29900);
nand UO_2282 (O_2282,N_29988,N_29965);
and UO_2283 (O_2283,N_29853,N_29827);
nor UO_2284 (O_2284,N_29854,N_29911);
nor UO_2285 (O_2285,N_29818,N_29887);
nand UO_2286 (O_2286,N_29899,N_29900);
nor UO_2287 (O_2287,N_29961,N_29855);
xor UO_2288 (O_2288,N_29813,N_29804);
and UO_2289 (O_2289,N_29999,N_29895);
nor UO_2290 (O_2290,N_29955,N_29994);
and UO_2291 (O_2291,N_29899,N_29935);
nand UO_2292 (O_2292,N_29912,N_29884);
nand UO_2293 (O_2293,N_29939,N_29931);
or UO_2294 (O_2294,N_29835,N_29844);
and UO_2295 (O_2295,N_29975,N_29894);
nor UO_2296 (O_2296,N_29858,N_29908);
nand UO_2297 (O_2297,N_29840,N_29877);
xnor UO_2298 (O_2298,N_29802,N_29914);
nor UO_2299 (O_2299,N_29945,N_29859);
nand UO_2300 (O_2300,N_29810,N_29993);
nor UO_2301 (O_2301,N_29885,N_29965);
nor UO_2302 (O_2302,N_29840,N_29975);
xor UO_2303 (O_2303,N_29890,N_29818);
nor UO_2304 (O_2304,N_29977,N_29939);
xnor UO_2305 (O_2305,N_29820,N_29813);
and UO_2306 (O_2306,N_29812,N_29847);
xnor UO_2307 (O_2307,N_29964,N_29921);
xnor UO_2308 (O_2308,N_29845,N_29837);
or UO_2309 (O_2309,N_29817,N_29850);
nand UO_2310 (O_2310,N_29959,N_29906);
nor UO_2311 (O_2311,N_29855,N_29824);
or UO_2312 (O_2312,N_29839,N_29820);
and UO_2313 (O_2313,N_29999,N_29897);
or UO_2314 (O_2314,N_29964,N_29845);
or UO_2315 (O_2315,N_29807,N_29989);
nor UO_2316 (O_2316,N_29977,N_29867);
nor UO_2317 (O_2317,N_29975,N_29944);
or UO_2318 (O_2318,N_29800,N_29933);
nand UO_2319 (O_2319,N_29824,N_29943);
xor UO_2320 (O_2320,N_29949,N_29994);
nand UO_2321 (O_2321,N_29817,N_29969);
or UO_2322 (O_2322,N_29929,N_29847);
and UO_2323 (O_2323,N_29935,N_29894);
nor UO_2324 (O_2324,N_29834,N_29891);
and UO_2325 (O_2325,N_29827,N_29890);
and UO_2326 (O_2326,N_29884,N_29819);
nand UO_2327 (O_2327,N_29873,N_29975);
nand UO_2328 (O_2328,N_29850,N_29884);
nand UO_2329 (O_2329,N_29962,N_29928);
nor UO_2330 (O_2330,N_29811,N_29967);
xor UO_2331 (O_2331,N_29805,N_29985);
and UO_2332 (O_2332,N_29904,N_29903);
and UO_2333 (O_2333,N_29852,N_29805);
and UO_2334 (O_2334,N_29881,N_29964);
and UO_2335 (O_2335,N_29917,N_29830);
xor UO_2336 (O_2336,N_29804,N_29856);
and UO_2337 (O_2337,N_29861,N_29956);
or UO_2338 (O_2338,N_29915,N_29841);
and UO_2339 (O_2339,N_29829,N_29878);
or UO_2340 (O_2340,N_29848,N_29899);
nor UO_2341 (O_2341,N_29960,N_29908);
nand UO_2342 (O_2342,N_29941,N_29992);
nand UO_2343 (O_2343,N_29903,N_29951);
xor UO_2344 (O_2344,N_29923,N_29821);
nor UO_2345 (O_2345,N_29865,N_29987);
or UO_2346 (O_2346,N_29833,N_29846);
xor UO_2347 (O_2347,N_29855,N_29936);
nand UO_2348 (O_2348,N_29849,N_29982);
nor UO_2349 (O_2349,N_29981,N_29861);
or UO_2350 (O_2350,N_29995,N_29885);
and UO_2351 (O_2351,N_29856,N_29855);
and UO_2352 (O_2352,N_29993,N_29923);
xnor UO_2353 (O_2353,N_29905,N_29884);
xnor UO_2354 (O_2354,N_29842,N_29982);
and UO_2355 (O_2355,N_29822,N_29907);
or UO_2356 (O_2356,N_29956,N_29803);
xor UO_2357 (O_2357,N_29998,N_29810);
nor UO_2358 (O_2358,N_29853,N_29945);
xor UO_2359 (O_2359,N_29842,N_29989);
nor UO_2360 (O_2360,N_29996,N_29817);
and UO_2361 (O_2361,N_29846,N_29934);
nand UO_2362 (O_2362,N_29866,N_29907);
or UO_2363 (O_2363,N_29966,N_29842);
nand UO_2364 (O_2364,N_29886,N_29844);
or UO_2365 (O_2365,N_29806,N_29957);
nand UO_2366 (O_2366,N_29915,N_29821);
nor UO_2367 (O_2367,N_29998,N_29967);
or UO_2368 (O_2368,N_29966,N_29928);
xnor UO_2369 (O_2369,N_29980,N_29930);
xnor UO_2370 (O_2370,N_29999,N_29988);
or UO_2371 (O_2371,N_29935,N_29952);
xor UO_2372 (O_2372,N_29964,N_29983);
nor UO_2373 (O_2373,N_29926,N_29902);
or UO_2374 (O_2374,N_29937,N_29940);
nand UO_2375 (O_2375,N_29820,N_29840);
nor UO_2376 (O_2376,N_29963,N_29970);
nor UO_2377 (O_2377,N_29940,N_29883);
nor UO_2378 (O_2378,N_29946,N_29902);
nor UO_2379 (O_2379,N_29892,N_29898);
xnor UO_2380 (O_2380,N_29914,N_29801);
and UO_2381 (O_2381,N_29802,N_29868);
or UO_2382 (O_2382,N_29953,N_29849);
nor UO_2383 (O_2383,N_29890,N_29838);
xor UO_2384 (O_2384,N_29895,N_29954);
nand UO_2385 (O_2385,N_29910,N_29853);
nor UO_2386 (O_2386,N_29832,N_29846);
and UO_2387 (O_2387,N_29986,N_29866);
nor UO_2388 (O_2388,N_29906,N_29943);
or UO_2389 (O_2389,N_29953,N_29897);
xor UO_2390 (O_2390,N_29926,N_29912);
or UO_2391 (O_2391,N_29883,N_29819);
nor UO_2392 (O_2392,N_29990,N_29957);
or UO_2393 (O_2393,N_29887,N_29824);
and UO_2394 (O_2394,N_29938,N_29908);
and UO_2395 (O_2395,N_29970,N_29919);
nor UO_2396 (O_2396,N_29863,N_29846);
or UO_2397 (O_2397,N_29855,N_29836);
nand UO_2398 (O_2398,N_29805,N_29904);
nand UO_2399 (O_2399,N_29844,N_29946);
nand UO_2400 (O_2400,N_29825,N_29886);
and UO_2401 (O_2401,N_29838,N_29961);
nand UO_2402 (O_2402,N_29994,N_29899);
xor UO_2403 (O_2403,N_29866,N_29835);
nor UO_2404 (O_2404,N_29905,N_29837);
and UO_2405 (O_2405,N_29996,N_29962);
nand UO_2406 (O_2406,N_29993,N_29977);
and UO_2407 (O_2407,N_29926,N_29988);
xnor UO_2408 (O_2408,N_29997,N_29987);
nor UO_2409 (O_2409,N_29944,N_29878);
xnor UO_2410 (O_2410,N_29926,N_29880);
nor UO_2411 (O_2411,N_29982,N_29926);
nor UO_2412 (O_2412,N_29835,N_29877);
nor UO_2413 (O_2413,N_29974,N_29977);
or UO_2414 (O_2414,N_29963,N_29805);
or UO_2415 (O_2415,N_29970,N_29954);
nor UO_2416 (O_2416,N_29839,N_29856);
nor UO_2417 (O_2417,N_29816,N_29803);
xnor UO_2418 (O_2418,N_29846,N_29946);
or UO_2419 (O_2419,N_29865,N_29963);
or UO_2420 (O_2420,N_29811,N_29863);
xor UO_2421 (O_2421,N_29910,N_29979);
or UO_2422 (O_2422,N_29846,N_29827);
nand UO_2423 (O_2423,N_29916,N_29983);
and UO_2424 (O_2424,N_29927,N_29862);
and UO_2425 (O_2425,N_29828,N_29842);
xor UO_2426 (O_2426,N_29825,N_29858);
or UO_2427 (O_2427,N_29882,N_29823);
nand UO_2428 (O_2428,N_29975,N_29805);
nor UO_2429 (O_2429,N_29811,N_29812);
xnor UO_2430 (O_2430,N_29973,N_29901);
and UO_2431 (O_2431,N_29915,N_29998);
and UO_2432 (O_2432,N_29982,N_29814);
and UO_2433 (O_2433,N_29855,N_29919);
nand UO_2434 (O_2434,N_29927,N_29948);
nand UO_2435 (O_2435,N_29852,N_29893);
nor UO_2436 (O_2436,N_29907,N_29934);
and UO_2437 (O_2437,N_29885,N_29812);
nand UO_2438 (O_2438,N_29872,N_29954);
and UO_2439 (O_2439,N_29840,N_29891);
or UO_2440 (O_2440,N_29958,N_29949);
xnor UO_2441 (O_2441,N_29946,N_29977);
or UO_2442 (O_2442,N_29919,N_29893);
nand UO_2443 (O_2443,N_29935,N_29826);
xor UO_2444 (O_2444,N_29864,N_29820);
nor UO_2445 (O_2445,N_29874,N_29951);
or UO_2446 (O_2446,N_29819,N_29858);
xnor UO_2447 (O_2447,N_29822,N_29834);
or UO_2448 (O_2448,N_29806,N_29908);
and UO_2449 (O_2449,N_29810,N_29891);
nand UO_2450 (O_2450,N_29916,N_29886);
xor UO_2451 (O_2451,N_29804,N_29808);
nand UO_2452 (O_2452,N_29914,N_29810);
nor UO_2453 (O_2453,N_29968,N_29858);
nand UO_2454 (O_2454,N_29855,N_29837);
xnor UO_2455 (O_2455,N_29812,N_29918);
xnor UO_2456 (O_2456,N_29816,N_29919);
or UO_2457 (O_2457,N_29840,N_29990);
or UO_2458 (O_2458,N_29871,N_29990);
xnor UO_2459 (O_2459,N_29977,N_29979);
and UO_2460 (O_2460,N_29874,N_29903);
nand UO_2461 (O_2461,N_29966,N_29886);
xor UO_2462 (O_2462,N_29845,N_29946);
or UO_2463 (O_2463,N_29869,N_29874);
and UO_2464 (O_2464,N_29922,N_29863);
and UO_2465 (O_2465,N_29835,N_29806);
and UO_2466 (O_2466,N_29979,N_29919);
xnor UO_2467 (O_2467,N_29918,N_29879);
nand UO_2468 (O_2468,N_29841,N_29901);
or UO_2469 (O_2469,N_29948,N_29946);
nand UO_2470 (O_2470,N_29999,N_29823);
or UO_2471 (O_2471,N_29829,N_29941);
or UO_2472 (O_2472,N_29880,N_29881);
nand UO_2473 (O_2473,N_29994,N_29847);
and UO_2474 (O_2474,N_29825,N_29891);
xnor UO_2475 (O_2475,N_29963,N_29953);
nand UO_2476 (O_2476,N_29946,N_29944);
nand UO_2477 (O_2477,N_29860,N_29871);
nor UO_2478 (O_2478,N_29822,N_29841);
nor UO_2479 (O_2479,N_29897,N_29992);
and UO_2480 (O_2480,N_29899,N_29943);
nand UO_2481 (O_2481,N_29813,N_29934);
or UO_2482 (O_2482,N_29873,N_29937);
nor UO_2483 (O_2483,N_29951,N_29899);
and UO_2484 (O_2484,N_29967,N_29920);
nor UO_2485 (O_2485,N_29834,N_29849);
nor UO_2486 (O_2486,N_29992,N_29878);
and UO_2487 (O_2487,N_29909,N_29999);
nor UO_2488 (O_2488,N_29870,N_29856);
nand UO_2489 (O_2489,N_29843,N_29814);
nand UO_2490 (O_2490,N_29977,N_29902);
and UO_2491 (O_2491,N_29939,N_29842);
xor UO_2492 (O_2492,N_29997,N_29807);
and UO_2493 (O_2493,N_29910,N_29989);
and UO_2494 (O_2494,N_29903,N_29892);
or UO_2495 (O_2495,N_29902,N_29996);
and UO_2496 (O_2496,N_29932,N_29963);
nor UO_2497 (O_2497,N_29884,N_29906);
nand UO_2498 (O_2498,N_29958,N_29978);
nor UO_2499 (O_2499,N_29839,N_29828);
nand UO_2500 (O_2500,N_29972,N_29975);
and UO_2501 (O_2501,N_29850,N_29962);
or UO_2502 (O_2502,N_29884,N_29832);
nand UO_2503 (O_2503,N_29804,N_29842);
nand UO_2504 (O_2504,N_29999,N_29903);
and UO_2505 (O_2505,N_29979,N_29915);
xnor UO_2506 (O_2506,N_29838,N_29995);
and UO_2507 (O_2507,N_29888,N_29912);
nand UO_2508 (O_2508,N_29960,N_29820);
or UO_2509 (O_2509,N_29976,N_29956);
xor UO_2510 (O_2510,N_29998,N_29863);
or UO_2511 (O_2511,N_29993,N_29911);
nand UO_2512 (O_2512,N_29999,N_29899);
or UO_2513 (O_2513,N_29837,N_29979);
or UO_2514 (O_2514,N_29948,N_29959);
nand UO_2515 (O_2515,N_29843,N_29800);
or UO_2516 (O_2516,N_29846,N_29869);
and UO_2517 (O_2517,N_29951,N_29834);
nand UO_2518 (O_2518,N_29854,N_29991);
xnor UO_2519 (O_2519,N_29820,N_29915);
nand UO_2520 (O_2520,N_29910,N_29992);
xnor UO_2521 (O_2521,N_29917,N_29802);
nor UO_2522 (O_2522,N_29894,N_29831);
nor UO_2523 (O_2523,N_29820,N_29971);
and UO_2524 (O_2524,N_29898,N_29911);
nand UO_2525 (O_2525,N_29966,N_29913);
xnor UO_2526 (O_2526,N_29977,N_29843);
xor UO_2527 (O_2527,N_29933,N_29973);
and UO_2528 (O_2528,N_29923,N_29861);
nor UO_2529 (O_2529,N_29866,N_29901);
nor UO_2530 (O_2530,N_29893,N_29969);
nor UO_2531 (O_2531,N_29956,N_29966);
nand UO_2532 (O_2532,N_29943,N_29852);
and UO_2533 (O_2533,N_29819,N_29989);
xor UO_2534 (O_2534,N_29910,N_29934);
nor UO_2535 (O_2535,N_29955,N_29883);
nand UO_2536 (O_2536,N_29932,N_29880);
xor UO_2537 (O_2537,N_29896,N_29858);
nand UO_2538 (O_2538,N_29943,N_29994);
or UO_2539 (O_2539,N_29991,N_29917);
nor UO_2540 (O_2540,N_29916,N_29995);
or UO_2541 (O_2541,N_29904,N_29920);
or UO_2542 (O_2542,N_29863,N_29917);
or UO_2543 (O_2543,N_29994,N_29839);
nor UO_2544 (O_2544,N_29868,N_29845);
nor UO_2545 (O_2545,N_29979,N_29880);
nor UO_2546 (O_2546,N_29978,N_29800);
nand UO_2547 (O_2547,N_29984,N_29961);
nand UO_2548 (O_2548,N_29819,N_29800);
xor UO_2549 (O_2549,N_29963,N_29921);
xor UO_2550 (O_2550,N_29914,N_29966);
nand UO_2551 (O_2551,N_29974,N_29991);
nor UO_2552 (O_2552,N_29970,N_29880);
nor UO_2553 (O_2553,N_29951,N_29969);
or UO_2554 (O_2554,N_29810,N_29987);
nor UO_2555 (O_2555,N_29854,N_29969);
nand UO_2556 (O_2556,N_29929,N_29826);
and UO_2557 (O_2557,N_29951,N_29909);
nand UO_2558 (O_2558,N_29941,N_29959);
nand UO_2559 (O_2559,N_29911,N_29924);
xor UO_2560 (O_2560,N_29984,N_29875);
xor UO_2561 (O_2561,N_29937,N_29814);
xnor UO_2562 (O_2562,N_29915,N_29932);
or UO_2563 (O_2563,N_29926,N_29981);
nor UO_2564 (O_2564,N_29917,N_29919);
or UO_2565 (O_2565,N_29978,N_29891);
nor UO_2566 (O_2566,N_29935,N_29923);
and UO_2567 (O_2567,N_29963,N_29999);
and UO_2568 (O_2568,N_29968,N_29962);
xor UO_2569 (O_2569,N_29842,N_29848);
xnor UO_2570 (O_2570,N_29946,N_29939);
nand UO_2571 (O_2571,N_29905,N_29984);
xor UO_2572 (O_2572,N_29834,N_29929);
xnor UO_2573 (O_2573,N_29914,N_29922);
xor UO_2574 (O_2574,N_29832,N_29829);
xor UO_2575 (O_2575,N_29994,N_29934);
or UO_2576 (O_2576,N_29911,N_29986);
nor UO_2577 (O_2577,N_29908,N_29950);
and UO_2578 (O_2578,N_29857,N_29918);
nor UO_2579 (O_2579,N_29873,N_29989);
and UO_2580 (O_2580,N_29906,N_29969);
nand UO_2581 (O_2581,N_29973,N_29843);
or UO_2582 (O_2582,N_29878,N_29823);
nor UO_2583 (O_2583,N_29949,N_29917);
nor UO_2584 (O_2584,N_29834,N_29926);
and UO_2585 (O_2585,N_29807,N_29894);
and UO_2586 (O_2586,N_29994,N_29874);
and UO_2587 (O_2587,N_29815,N_29913);
xor UO_2588 (O_2588,N_29906,N_29891);
and UO_2589 (O_2589,N_29919,N_29827);
or UO_2590 (O_2590,N_29970,N_29951);
or UO_2591 (O_2591,N_29828,N_29993);
and UO_2592 (O_2592,N_29822,N_29904);
and UO_2593 (O_2593,N_29929,N_29818);
or UO_2594 (O_2594,N_29998,N_29880);
xor UO_2595 (O_2595,N_29822,N_29803);
or UO_2596 (O_2596,N_29875,N_29825);
nor UO_2597 (O_2597,N_29986,N_29885);
nand UO_2598 (O_2598,N_29864,N_29812);
or UO_2599 (O_2599,N_29825,N_29979);
nand UO_2600 (O_2600,N_29919,N_29874);
and UO_2601 (O_2601,N_29820,N_29890);
and UO_2602 (O_2602,N_29816,N_29901);
nor UO_2603 (O_2603,N_29872,N_29853);
and UO_2604 (O_2604,N_29965,N_29937);
or UO_2605 (O_2605,N_29914,N_29999);
xor UO_2606 (O_2606,N_29836,N_29982);
nand UO_2607 (O_2607,N_29955,N_29907);
or UO_2608 (O_2608,N_29889,N_29977);
nor UO_2609 (O_2609,N_29906,N_29998);
nor UO_2610 (O_2610,N_29831,N_29867);
nor UO_2611 (O_2611,N_29897,N_29938);
and UO_2612 (O_2612,N_29944,N_29887);
xor UO_2613 (O_2613,N_29912,N_29895);
and UO_2614 (O_2614,N_29810,N_29848);
and UO_2615 (O_2615,N_29959,N_29945);
nand UO_2616 (O_2616,N_29905,N_29991);
nor UO_2617 (O_2617,N_29906,N_29862);
nor UO_2618 (O_2618,N_29937,N_29825);
and UO_2619 (O_2619,N_29980,N_29993);
or UO_2620 (O_2620,N_29919,N_29864);
nand UO_2621 (O_2621,N_29901,N_29960);
xnor UO_2622 (O_2622,N_29895,N_29840);
nand UO_2623 (O_2623,N_29898,N_29970);
and UO_2624 (O_2624,N_29813,N_29909);
nand UO_2625 (O_2625,N_29849,N_29934);
xor UO_2626 (O_2626,N_29889,N_29873);
or UO_2627 (O_2627,N_29968,N_29916);
and UO_2628 (O_2628,N_29802,N_29805);
and UO_2629 (O_2629,N_29867,N_29892);
xnor UO_2630 (O_2630,N_29927,N_29976);
xor UO_2631 (O_2631,N_29828,N_29994);
xnor UO_2632 (O_2632,N_29872,N_29864);
or UO_2633 (O_2633,N_29848,N_29902);
xnor UO_2634 (O_2634,N_29980,N_29931);
or UO_2635 (O_2635,N_29870,N_29855);
or UO_2636 (O_2636,N_29823,N_29976);
xnor UO_2637 (O_2637,N_29842,N_29880);
xor UO_2638 (O_2638,N_29850,N_29851);
nand UO_2639 (O_2639,N_29912,N_29951);
nand UO_2640 (O_2640,N_29898,N_29830);
or UO_2641 (O_2641,N_29976,N_29968);
nor UO_2642 (O_2642,N_29916,N_29838);
nor UO_2643 (O_2643,N_29907,N_29806);
and UO_2644 (O_2644,N_29982,N_29806);
xor UO_2645 (O_2645,N_29866,N_29803);
nand UO_2646 (O_2646,N_29938,N_29840);
or UO_2647 (O_2647,N_29824,N_29822);
nand UO_2648 (O_2648,N_29873,N_29977);
and UO_2649 (O_2649,N_29849,N_29990);
xnor UO_2650 (O_2650,N_29966,N_29917);
xor UO_2651 (O_2651,N_29832,N_29822);
or UO_2652 (O_2652,N_29844,N_29810);
nor UO_2653 (O_2653,N_29870,N_29956);
or UO_2654 (O_2654,N_29924,N_29882);
or UO_2655 (O_2655,N_29972,N_29932);
nand UO_2656 (O_2656,N_29848,N_29915);
xnor UO_2657 (O_2657,N_29843,N_29805);
or UO_2658 (O_2658,N_29971,N_29871);
nor UO_2659 (O_2659,N_29859,N_29907);
and UO_2660 (O_2660,N_29815,N_29921);
xor UO_2661 (O_2661,N_29873,N_29883);
or UO_2662 (O_2662,N_29875,N_29820);
xnor UO_2663 (O_2663,N_29961,N_29892);
nor UO_2664 (O_2664,N_29901,N_29878);
nor UO_2665 (O_2665,N_29807,N_29977);
nand UO_2666 (O_2666,N_29856,N_29909);
xor UO_2667 (O_2667,N_29923,N_29828);
xnor UO_2668 (O_2668,N_29957,N_29975);
nor UO_2669 (O_2669,N_29953,N_29909);
nor UO_2670 (O_2670,N_29951,N_29943);
xor UO_2671 (O_2671,N_29816,N_29834);
or UO_2672 (O_2672,N_29945,N_29841);
nand UO_2673 (O_2673,N_29821,N_29851);
nand UO_2674 (O_2674,N_29932,N_29928);
or UO_2675 (O_2675,N_29917,N_29865);
nand UO_2676 (O_2676,N_29817,N_29928);
and UO_2677 (O_2677,N_29970,N_29885);
xnor UO_2678 (O_2678,N_29990,N_29900);
and UO_2679 (O_2679,N_29857,N_29892);
or UO_2680 (O_2680,N_29892,N_29909);
xnor UO_2681 (O_2681,N_29990,N_29941);
or UO_2682 (O_2682,N_29967,N_29957);
nor UO_2683 (O_2683,N_29898,N_29993);
xor UO_2684 (O_2684,N_29800,N_29916);
xor UO_2685 (O_2685,N_29904,N_29932);
and UO_2686 (O_2686,N_29818,N_29906);
nor UO_2687 (O_2687,N_29984,N_29990);
nand UO_2688 (O_2688,N_29859,N_29974);
or UO_2689 (O_2689,N_29851,N_29966);
nand UO_2690 (O_2690,N_29907,N_29896);
nand UO_2691 (O_2691,N_29985,N_29817);
or UO_2692 (O_2692,N_29856,N_29906);
xnor UO_2693 (O_2693,N_29926,N_29991);
nand UO_2694 (O_2694,N_29975,N_29817);
and UO_2695 (O_2695,N_29951,N_29831);
and UO_2696 (O_2696,N_29891,N_29856);
nor UO_2697 (O_2697,N_29807,N_29906);
nor UO_2698 (O_2698,N_29961,N_29932);
nor UO_2699 (O_2699,N_29823,N_29940);
or UO_2700 (O_2700,N_29922,N_29858);
and UO_2701 (O_2701,N_29998,N_29827);
nand UO_2702 (O_2702,N_29954,N_29921);
xor UO_2703 (O_2703,N_29996,N_29911);
and UO_2704 (O_2704,N_29944,N_29898);
nor UO_2705 (O_2705,N_29889,N_29896);
xnor UO_2706 (O_2706,N_29949,N_29904);
or UO_2707 (O_2707,N_29898,N_29994);
xor UO_2708 (O_2708,N_29892,N_29982);
xnor UO_2709 (O_2709,N_29849,N_29994);
nor UO_2710 (O_2710,N_29864,N_29873);
or UO_2711 (O_2711,N_29876,N_29830);
and UO_2712 (O_2712,N_29872,N_29909);
or UO_2713 (O_2713,N_29952,N_29859);
or UO_2714 (O_2714,N_29967,N_29941);
nor UO_2715 (O_2715,N_29919,N_29959);
xor UO_2716 (O_2716,N_29999,N_29836);
and UO_2717 (O_2717,N_29991,N_29896);
and UO_2718 (O_2718,N_29850,N_29885);
nand UO_2719 (O_2719,N_29850,N_29965);
nand UO_2720 (O_2720,N_29933,N_29851);
and UO_2721 (O_2721,N_29958,N_29938);
nor UO_2722 (O_2722,N_29889,N_29991);
or UO_2723 (O_2723,N_29820,N_29962);
and UO_2724 (O_2724,N_29876,N_29865);
nor UO_2725 (O_2725,N_29811,N_29923);
and UO_2726 (O_2726,N_29967,N_29904);
and UO_2727 (O_2727,N_29871,N_29814);
nand UO_2728 (O_2728,N_29802,N_29838);
and UO_2729 (O_2729,N_29821,N_29943);
nand UO_2730 (O_2730,N_29867,N_29835);
nand UO_2731 (O_2731,N_29984,N_29879);
and UO_2732 (O_2732,N_29912,N_29940);
and UO_2733 (O_2733,N_29834,N_29840);
xor UO_2734 (O_2734,N_29956,N_29931);
nor UO_2735 (O_2735,N_29894,N_29868);
or UO_2736 (O_2736,N_29912,N_29971);
nor UO_2737 (O_2737,N_29872,N_29941);
and UO_2738 (O_2738,N_29830,N_29802);
or UO_2739 (O_2739,N_29897,N_29976);
nor UO_2740 (O_2740,N_29986,N_29822);
nand UO_2741 (O_2741,N_29983,N_29848);
xnor UO_2742 (O_2742,N_29987,N_29820);
nor UO_2743 (O_2743,N_29805,N_29825);
nand UO_2744 (O_2744,N_29901,N_29885);
nor UO_2745 (O_2745,N_29925,N_29943);
nand UO_2746 (O_2746,N_29917,N_29841);
nor UO_2747 (O_2747,N_29880,N_29946);
and UO_2748 (O_2748,N_29890,N_29934);
or UO_2749 (O_2749,N_29903,N_29990);
xnor UO_2750 (O_2750,N_29921,N_29915);
or UO_2751 (O_2751,N_29826,N_29916);
nor UO_2752 (O_2752,N_29858,N_29989);
nor UO_2753 (O_2753,N_29802,N_29848);
nand UO_2754 (O_2754,N_29902,N_29837);
and UO_2755 (O_2755,N_29906,N_29964);
nand UO_2756 (O_2756,N_29863,N_29867);
nor UO_2757 (O_2757,N_29823,N_29945);
nor UO_2758 (O_2758,N_29998,N_29814);
and UO_2759 (O_2759,N_29886,N_29978);
and UO_2760 (O_2760,N_29998,N_29988);
nor UO_2761 (O_2761,N_29944,N_29821);
or UO_2762 (O_2762,N_29872,N_29904);
xor UO_2763 (O_2763,N_29957,N_29980);
xnor UO_2764 (O_2764,N_29804,N_29806);
xnor UO_2765 (O_2765,N_29985,N_29825);
and UO_2766 (O_2766,N_29937,N_29987);
xor UO_2767 (O_2767,N_29860,N_29912);
and UO_2768 (O_2768,N_29850,N_29900);
nand UO_2769 (O_2769,N_29972,N_29884);
and UO_2770 (O_2770,N_29841,N_29928);
and UO_2771 (O_2771,N_29909,N_29895);
nand UO_2772 (O_2772,N_29906,N_29971);
xor UO_2773 (O_2773,N_29984,N_29975);
nand UO_2774 (O_2774,N_29965,N_29820);
nand UO_2775 (O_2775,N_29989,N_29889);
xor UO_2776 (O_2776,N_29949,N_29836);
xnor UO_2777 (O_2777,N_29819,N_29891);
or UO_2778 (O_2778,N_29808,N_29889);
and UO_2779 (O_2779,N_29977,N_29989);
and UO_2780 (O_2780,N_29870,N_29861);
or UO_2781 (O_2781,N_29991,N_29978);
xor UO_2782 (O_2782,N_29925,N_29899);
nor UO_2783 (O_2783,N_29875,N_29923);
and UO_2784 (O_2784,N_29995,N_29972);
nor UO_2785 (O_2785,N_29979,N_29848);
and UO_2786 (O_2786,N_29875,N_29893);
or UO_2787 (O_2787,N_29859,N_29877);
nand UO_2788 (O_2788,N_29870,N_29929);
or UO_2789 (O_2789,N_29977,N_29874);
nand UO_2790 (O_2790,N_29889,N_29910);
xnor UO_2791 (O_2791,N_29821,N_29961);
or UO_2792 (O_2792,N_29928,N_29964);
or UO_2793 (O_2793,N_29960,N_29936);
xnor UO_2794 (O_2794,N_29907,N_29850);
nand UO_2795 (O_2795,N_29856,N_29961);
and UO_2796 (O_2796,N_29857,N_29860);
nand UO_2797 (O_2797,N_29885,N_29803);
nand UO_2798 (O_2798,N_29969,N_29909);
xor UO_2799 (O_2799,N_29902,N_29861);
nor UO_2800 (O_2800,N_29805,N_29844);
xnor UO_2801 (O_2801,N_29940,N_29957);
or UO_2802 (O_2802,N_29810,N_29856);
and UO_2803 (O_2803,N_29839,N_29885);
nor UO_2804 (O_2804,N_29828,N_29913);
and UO_2805 (O_2805,N_29906,N_29815);
nand UO_2806 (O_2806,N_29925,N_29831);
xnor UO_2807 (O_2807,N_29937,N_29811);
nand UO_2808 (O_2808,N_29804,N_29995);
and UO_2809 (O_2809,N_29908,N_29946);
and UO_2810 (O_2810,N_29971,N_29937);
and UO_2811 (O_2811,N_29888,N_29934);
nor UO_2812 (O_2812,N_29911,N_29808);
or UO_2813 (O_2813,N_29912,N_29968);
nor UO_2814 (O_2814,N_29837,N_29801);
nor UO_2815 (O_2815,N_29893,N_29881);
and UO_2816 (O_2816,N_29871,N_29926);
nand UO_2817 (O_2817,N_29961,N_29919);
nand UO_2818 (O_2818,N_29894,N_29947);
xnor UO_2819 (O_2819,N_29816,N_29979);
nand UO_2820 (O_2820,N_29910,N_29940);
nor UO_2821 (O_2821,N_29856,N_29859);
or UO_2822 (O_2822,N_29902,N_29914);
xnor UO_2823 (O_2823,N_29985,N_29986);
nor UO_2824 (O_2824,N_29972,N_29998);
xor UO_2825 (O_2825,N_29851,N_29847);
nor UO_2826 (O_2826,N_29881,N_29943);
nand UO_2827 (O_2827,N_29863,N_29882);
xor UO_2828 (O_2828,N_29903,N_29915);
or UO_2829 (O_2829,N_29802,N_29993);
or UO_2830 (O_2830,N_29906,N_29947);
nand UO_2831 (O_2831,N_29835,N_29841);
and UO_2832 (O_2832,N_29897,N_29905);
xor UO_2833 (O_2833,N_29838,N_29848);
nor UO_2834 (O_2834,N_29985,N_29834);
xnor UO_2835 (O_2835,N_29814,N_29892);
and UO_2836 (O_2836,N_29879,N_29935);
and UO_2837 (O_2837,N_29884,N_29985);
and UO_2838 (O_2838,N_29818,N_29928);
and UO_2839 (O_2839,N_29891,N_29926);
nand UO_2840 (O_2840,N_29900,N_29980);
xor UO_2841 (O_2841,N_29968,N_29969);
xor UO_2842 (O_2842,N_29967,N_29985);
xnor UO_2843 (O_2843,N_29990,N_29858);
nand UO_2844 (O_2844,N_29991,N_29825);
xnor UO_2845 (O_2845,N_29921,N_29842);
or UO_2846 (O_2846,N_29967,N_29987);
nor UO_2847 (O_2847,N_29845,N_29866);
nor UO_2848 (O_2848,N_29898,N_29956);
or UO_2849 (O_2849,N_29992,N_29938);
and UO_2850 (O_2850,N_29875,N_29977);
and UO_2851 (O_2851,N_29929,N_29940);
nor UO_2852 (O_2852,N_29980,N_29831);
nand UO_2853 (O_2853,N_29830,N_29927);
and UO_2854 (O_2854,N_29910,N_29942);
and UO_2855 (O_2855,N_29868,N_29962);
or UO_2856 (O_2856,N_29835,N_29986);
or UO_2857 (O_2857,N_29976,N_29865);
xor UO_2858 (O_2858,N_29934,N_29943);
and UO_2859 (O_2859,N_29988,N_29993);
or UO_2860 (O_2860,N_29975,N_29853);
nor UO_2861 (O_2861,N_29970,N_29850);
nor UO_2862 (O_2862,N_29914,N_29923);
nor UO_2863 (O_2863,N_29887,N_29802);
nand UO_2864 (O_2864,N_29903,N_29899);
and UO_2865 (O_2865,N_29955,N_29949);
nor UO_2866 (O_2866,N_29899,N_29895);
nand UO_2867 (O_2867,N_29997,N_29811);
and UO_2868 (O_2868,N_29909,N_29889);
and UO_2869 (O_2869,N_29917,N_29840);
and UO_2870 (O_2870,N_29988,N_29811);
xor UO_2871 (O_2871,N_29978,N_29922);
xnor UO_2872 (O_2872,N_29841,N_29843);
xnor UO_2873 (O_2873,N_29871,N_29918);
and UO_2874 (O_2874,N_29887,N_29993);
or UO_2875 (O_2875,N_29889,N_29823);
and UO_2876 (O_2876,N_29803,N_29952);
and UO_2877 (O_2877,N_29967,N_29859);
and UO_2878 (O_2878,N_29807,N_29986);
nor UO_2879 (O_2879,N_29915,N_29853);
or UO_2880 (O_2880,N_29995,N_29805);
nor UO_2881 (O_2881,N_29867,N_29881);
and UO_2882 (O_2882,N_29994,N_29922);
nand UO_2883 (O_2883,N_29935,N_29821);
or UO_2884 (O_2884,N_29995,N_29878);
xor UO_2885 (O_2885,N_29813,N_29843);
and UO_2886 (O_2886,N_29888,N_29817);
nor UO_2887 (O_2887,N_29815,N_29831);
or UO_2888 (O_2888,N_29809,N_29825);
and UO_2889 (O_2889,N_29988,N_29936);
nor UO_2890 (O_2890,N_29955,N_29941);
nor UO_2891 (O_2891,N_29894,N_29875);
nor UO_2892 (O_2892,N_29895,N_29893);
and UO_2893 (O_2893,N_29959,N_29997);
and UO_2894 (O_2894,N_29996,N_29923);
and UO_2895 (O_2895,N_29819,N_29813);
and UO_2896 (O_2896,N_29868,N_29888);
and UO_2897 (O_2897,N_29873,N_29941);
nor UO_2898 (O_2898,N_29900,N_29973);
nand UO_2899 (O_2899,N_29986,N_29895);
nand UO_2900 (O_2900,N_29862,N_29829);
nor UO_2901 (O_2901,N_29828,N_29910);
nand UO_2902 (O_2902,N_29957,N_29874);
nor UO_2903 (O_2903,N_29806,N_29884);
or UO_2904 (O_2904,N_29807,N_29933);
xor UO_2905 (O_2905,N_29972,N_29974);
nand UO_2906 (O_2906,N_29895,N_29884);
and UO_2907 (O_2907,N_29905,N_29965);
and UO_2908 (O_2908,N_29957,N_29891);
and UO_2909 (O_2909,N_29912,N_29821);
and UO_2910 (O_2910,N_29960,N_29984);
nor UO_2911 (O_2911,N_29936,N_29971);
or UO_2912 (O_2912,N_29828,N_29973);
or UO_2913 (O_2913,N_29978,N_29850);
nand UO_2914 (O_2914,N_29875,N_29998);
nor UO_2915 (O_2915,N_29832,N_29962);
and UO_2916 (O_2916,N_29858,N_29997);
and UO_2917 (O_2917,N_29982,N_29983);
and UO_2918 (O_2918,N_29938,N_29819);
xnor UO_2919 (O_2919,N_29898,N_29915);
xor UO_2920 (O_2920,N_29927,N_29870);
or UO_2921 (O_2921,N_29897,N_29876);
xor UO_2922 (O_2922,N_29835,N_29951);
and UO_2923 (O_2923,N_29853,N_29920);
nand UO_2924 (O_2924,N_29840,N_29890);
and UO_2925 (O_2925,N_29922,N_29954);
and UO_2926 (O_2926,N_29941,N_29838);
nor UO_2927 (O_2927,N_29877,N_29802);
or UO_2928 (O_2928,N_29917,N_29937);
or UO_2929 (O_2929,N_29952,N_29821);
or UO_2930 (O_2930,N_29909,N_29875);
xor UO_2931 (O_2931,N_29932,N_29956);
or UO_2932 (O_2932,N_29833,N_29940);
nand UO_2933 (O_2933,N_29881,N_29994);
and UO_2934 (O_2934,N_29858,N_29851);
xnor UO_2935 (O_2935,N_29918,N_29992);
xor UO_2936 (O_2936,N_29868,N_29984);
or UO_2937 (O_2937,N_29940,N_29931);
or UO_2938 (O_2938,N_29940,N_29915);
or UO_2939 (O_2939,N_29854,N_29940);
nand UO_2940 (O_2940,N_29870,N_29806);
xor UO_2941 (O_2941,N_29862,N_29817);
xnor UO_2942 (O_2942,N_29809,N_29806);
or UO_2943 (O_2943,N_29806,N_29988);
or UO_2944 (O_2944,N_29898,N_29950);
nand UO_2945 (O_2945,N_29948,N_29938);
xnor UO_2946 (O_2946,N_29909,N_29942);
or UO_2947 (O_2947,N_29903,N_29975);
xor UO_2948 (O_2948,N_29871,N_29923);
or UO_2949 (O_2949,N_29878,N_29973);
nor UO_2950 (O_2950,N_29862,N_29971);
xnor UO_2951 (O_2951,N_29878,N_29804);
nand UO_2952 (O_2952,N_29979,N_29863);
and UO_2953 (O_2953,N_29837,N_29841);
nor UO_2954 (O_2954,N_29922,N_29909);
nor UO_2955 (O_2955,N_29951,N_29942);
and UO_2956 (O_2956,N_29801,N_29948);
nand UO_2957 (O_2957,N_29803,N_29998);
or UO_2958 (O_2958,N_29933,N_29960);
nand UO_2959 (O_2959,N_29905,N_29919);
and UO_2960 (O_2960,N_29973,N_29871);
and UO_2961 (O_2961,N_29819,N_29893);
or UO_2962 (O_2962,N_29909,N_29916);
xor UO_2963 (O_2963,N_29952,N_29949);
or UO_2964 (O_2964,N_29839,N_29813);
nor UO_2965 (O_2965,N_29826,N_29958);
or UO_2966 (O_2966,N_29848,N_29887);
xnor UO_2967 (O_2967,N_29853,N_29871);
nor UO_2968 (O_2968,N_29942,N_29859);
and UO_2969 (O_2969,N_29879,N_29844);
xnor UO_2970 (O_2970,N_29997,N_29951);
nand UO_2971 (O_2971,N_29813,N_29884);
nand UO_2972 (O_2972,N_29838,N_29801);
nand UO_2973 (O_2973,N_29942,N_29868);
or UO_2974 (O_2974,N_29992,N_29835);
and UO_2975 (O_2975,N_29995,N_29923);
or UO_2976 (O_2976,N_29960,N_29857);
xnor UO_2977 (O_2977,N_29999,N_29936);
nand UO_2978 (O_2978,N_29967,N_29921);
nor UO_2979 (O_2979,N_29986,N_29970);
and UO_2980 (O_2980,N_29825,N_29994);
nand UO_2981 (O_2981,N_29958,N_29976);
nor UO_2982 (O_2982,N_29937,N_29860);
or UO_2983 (O_2983,N_29906,N_29852);
nor UO_2984 (O_2984,N_29952,N_29910);
or UO_2985 (O_2985,N_29970,N_29842);
and UO_2986 (O_2986,N_29839,N_29966);
or UO_2987 (O_2987,N_29888,N_29860);
nand UO_2988 (O_2988,N_29929,N_29887);
and UO_2989 (O_2989,N_29850,N_29997);
and UO_2990 (O_2990,N_29838,N_29964);
and UO_2991 (O_2991,N_29908,N_29854);
nor UO_2992 (O_2992,N_29816,N_29839);
xnor UO_2993 (O_2993,N_29821,N_29840);
or UO_2994 (O_2994,N_29909,N_29952);
nand UO_2995 (O_2995,N_29805,N_29969);
or UO_2996 (O_2996,N_29879,N_29908);
nand UO_2997 (O_2997,N_29854,N_29887);
nand UO_2998 (O_2998,N_29816,N_29877);
nand UO_2999 (O_2999,N_29930,N_29957);
nand UO_3000 (O_3000,N_29940,N_29951);
nand UO_3001 (O_3001,N_29969,N_29916);
and UO_3002 (O_3002,N_29870,N_29988);
or UO_3003 (O_3003,N_29841,N_29825);
and UO_3004 (O_3004,N_29897,N_29960);
nor UO_3005 (O_3005,N_29805,N_29828);
and UO_3006 (O_3006,N_29943,N_29949);
or UO_3007 (O_3007,N_29934,N_29937);
and UO_3008 (O_3008,N_29986,N_29811);
and UO_3009 (O_3009,N_29851,N_29995);
nor UO_3010 (O_3010,N_29889,N_29903);
xor UO_3011 (O_3011,N_29848,N_29811);
nor UO_3012 (O_3012,N_29951,N_29862);
xor UO_3013 (O_3013,N_29894,N_29821);
and UO_3014 (O_3014,N_29838,N_29886);
or UO_3015 (O_3015,N_29854,N_29860);
or UO_3016 (O_3016,N_29974,N_29958);
xor UO_3017 (O_3017,N_29961,N_29834);
xor UO_3018 (O_3018,N_29952,N_29857);
nand UO_3019 (O_3019,N_29835,N_29813);
xnor UO_3020 (O_3020,N_29996,N_29822);
xnor UO_3021 (O_3021,N_29856,N_29852);
and UO_3022 (O_3022,N_29884,N_29885);
and UO_3023 (O_3023,N_29979,N_29894);
and UO_3024 (O_3024,N_29910,N_29811);
nor UO_3025 (O_3025,N_29809,N_29835);
nand UO_3026 (O_3026,N_29874,N_29846);
nand UO_3027 (O_3027,N_29939,N_29935);
nor UO_3028 (O_3028,N_29863,N_29810);
nand UO_3029 (O_3029,N_29967,N_29932);
xnor UO_3030 (O_3030,N_29829,N_29970);
xnor UO_3031 (O_3031,N_29918,N_29995);
nand UO_3032 (O_3032,N_29808,N_29945);
xor UO_3033 (O_3033,N_29942,N_29953);
nor UO_3034 (O_3034,N_29957,N_29979);
or UO_3035 (O_3035,N_29886,N_29998);
nand UO_3036 (O_3036,N_29899,N_29849);
nand UO_3037 (O_3037,N_29959,N_29882);
nand UO_3038 (O_3038,N_29803,N_29916);
nor UO_3039 (O_3039,N_29801,N_29991);
nand UO_3040 (O_3040,N_29843,N_29893);
xor UO_3041 (O_3041,N_29850,N_29901);
nand UO_3042 (O_3042,N_29832,N_29998);
nor UO_3043 (O_3043,N_29949,N_29883);
nand UO_3044 (O_3044,N_29948,N_29899);
nor UO_3045 (O_3045,N_29883,N_29899);
nor UO_3046 (O_3046,N_29960,N_29941);
and UO_3047 (O_3047,N_29860,N_29853);
and UO_3048 (O_3048,N_29886,N_29807);
xor UO_3049 (O_3049,N_29805,N_29972);
nor UO_3050 (O_3050,N_29844,N_29842);
or UO_3051 (O_3051,N_29956,N_29910);
or UO_3052 (O_3052,N_29841,N_29936);
and UO_3053 (O_3053,N_29857,N_29874);
nor UO_3054 (O_3054,N_29941,N_29949);
nand UO_3055 (O_3055,N_29855,N_29851);
xnor UO_3056 (O_3056,N_29812,N_29921);
xnor UO_3057 (O_3057,N_29991,N_29809);
nor UO_3058 (O_3058,N_29869,N_29929);
and UO_3059 (O_3059,N_29933,N_29824);
xor UO_3060 (O_3060,N_29838,N_29998);
or UO_3061 (O_3061,N_29990,N_29965);
or UO_3062 (O_3062,N_29959,N_29921);
nor UO_3063 (O_3063,N_29824,N_29833);
or UO_3064 (O_3064,N_29802,N_29803);
or UO_3065 (O_3065,N_29839,N_29864);
nand UO_3066 (O_3066,N_29836,N_29893);
xor UO_3067 (O_3067,N_29972,N_29890);
nor UO_3068 (O_3068,N_29894,N_29952);
xor UO_3069 (O_3069,N_29894,N_29830);
nand UO_3070 (O_3070,N_29892,N_29873);
or UO_3071 (O_3071,N_29802,N_29982);
and UO_3072 (O_3072,N_29957,N_29934);
nand UO_3073 (O_3073,N_29801,N_29899);
or UO_3074 (O_3074,N_29988,N_29984);
or UO_3075 (O_3075,N_29903,N_29986);
nor UO_3076 (O_3076,N_29869,N_29981);
nand UO_3077 (O_3077,N_29925,N_29877);
or UO_3078 (O_3078,N_29952,N_29806);
nor UO_3079 (O_3079,N_29987,N_29900);
or UO_3080 (O_3080,N_29900,N_29853);
xor UO_3081 (O_3081,N_29995,N_29998);
xor UO_3082 (O_3082,N_29998,N_29921);
or UO_3083 (O_3083,N_29925,N_29857);
nor UO_3084 (O_3084,N_29891,N_29879);
nand UO_3085 (O_3085,N_29825,N_29826);
and UO_3086 (O_3086,N_29931,N_29902);
nand UO_3087 (O_3087,N_29817,N_29805);
nor UO_3088 (O_3088,N_29904,N_29877);
nand UO_3089 (O_3089,N_29903,N_29935);
and UO_3090 (O_3090,N_29995,N_29872);
and UO_3091 (O_3091,N_29966,N_29834);
xor UO_3092 (O_3092,N_29816,N_29843);
xnor UO_3093 (O_3093,N_29991,N_29908);
and UO_3094 (O_3094,N_29897,N_29899);
or UO_3095 (O_3095,N_29896,N_29838);
nor UO_3096 (O_3096,N_29999,N_29997);
nor UO_3097 (O_3097,N_29965,N_29807);
nor UO_3098 (O_3098,N_29827,N_29995);
and UO_3099 (O_3099,N_29836,N_29994);
or UO_3100 (O_3100,N_29810,N_29989);
xnor UO_3101 (O_3101,N_29947,N_29810);
and UO_3102 (O_3102,N_29821,N_29960);
nor UO_3103 (O_3103,N_29971,N_29830);
xor UO_3104 (O_3104,N_29858,N_29925);
nor UO_3105 (O_3105,N_29818,N_29840);
xnor UO_3106 (O_3106,N_29868,N_29808);
and UO_3107 (O_3107,N_29970,N_29894);
nand UO_3108 (O_3108,N_29886,N_29822);
nor UO_3109 (O_3109,N_29962,N_29861);
nand UO_3110 (O_3110,N_29979,N_29947);
and UO_3111 (O_3111,N_29833,N_29919);
or UO_3112 (O_3112,N_29868,N_29995);
or UO_3113 (O_3113,N_29949,N_29857);
xor UO_3114 (O_3114,N_29849,N_29932);
or UO_3115 (O_3115,N_29869,N_29912);
nor UO_3116 (O_3116,N_29972,N_29801);
xnor UO_3117 (O_3117,N_29837,N_29950);
and UO_3118 (O_3118,N_29980,N_29852);
nand UO_3119 (O_3119,N_29837,N_29937);
and UO_3120 (O_3120,N_29991,N_29915);
xor UO_3121 (O_3121,N_29800,N_29814);
or UO_3122 (O_3122,N_29904,N_29972);
and UO_3123 (O_3123,N_29957,N_29843);
and UO_3124 (O_3124,N_29814,N_29815);
and UO_3125 (O_3125,N_29918,N_29859);
and UO_3126 (O_3126,N_29823,N_29875);
nand UO_3127 (O_3127,N_29958,N_29810);
nor UO_3128 (O_3128,N_29830,N_29947);
xnor UO_3129 (O_3129,N_29810,N_29912);
or UO_3130 (O_3130,N_29892,N_29908);
nor UO_3131 (O_3131,N_29836,N_29840);
nand UO_3132 (O_3132,N_29874,N_29921);
nand UO_3133 (O_3133,N_29910,N_29928);
or UO_3134 (O_3134,N_29990,N_29925);
or UO_3135 (O_3135,N_29987,N_29887);
xor UO_3136 (O_3136,N_29809,N_29804);
nor UO_3137 (O_3137,N_29830,N_29893);
nor UO_3138 (O_3138,N_29809,N_29810);
xnor UO_3139 (O_3139,N_29808,N_29858);
or UO_3140 (O_3140,N_29861,N_29824);
xnor UO_3141 (O_3141,N_29849,N_29959);
xor UO_3142 (O_3142,N_29897,N_29857);
or UO_3143 (O_3143,N_29853,N_29938);
nand UO_3144 (O_3144,N_29938,N_29845);
nand UO_3145 (O_3145,N_29934,N_29990);
nand UO_3146 (O_3146,N_29945,N_29941);
or UO_3147 (O_3147,N_29940,N_29800);
xor UO_3148 (O_3148,N_29810,N_29858);
xor UO_3149 (O_3149,N_29807,N_29816);
and UO_3150 (O_3150,N_29864,N_29925);
nor UO_3151 (O_3151,N_29822,N_29920);
and UO_3152 (O_3152,N_29999,N_29804);
nand UO_3153 (O_3153,N_29937,N_29966);
xnor UO_3154 (O_3154,N_29966,N_29896);
nand UO_3155 (O_3155,N_29913,N_29987);
or UO_3156 (O_3156,N_29893,N_29937);
and UO_3157 (O_3157,N_29858,N_29816);
nor UO_3158 (O_3158,N_29874,N_29978);
xor UO_3159 (O_3159,N_29946,N_29985);
and UO_3160 (O_3160,N_29971,N_29805);
xor UO_3161 (O_3161,N_29891,N_29964);
or UO_3162 (O_3162,N_29955,N_29821);
xnor UO_3163 (O_3163,N_29983,N_29972);
and UO_3164 (O_3164,N_29946,N_29817);
or UO_3165 (O_3165,N_29813,N_29966);
nand UO_3166 (O_3166,N_29812,N_29930);
or UO_3167 (O_3167,N_29976,N_29804);
nand UO_3168 (O_3168,N_29899,N_29904);
and UO_3169 (O_3169,N_29882,N_29822);
or UO_3170 (O_3170,N_29855,N_29983);
or UO_3171 (O_3171,N_29823,N_29982);
xnor UO_3172 (O_3172,N_29902,N_29847);
or UO_3173 (O_3173,N_29909,N_29947);
or UO_3174 (O_3174,N_29844,N_29923);
xor UO_3175 (O_3175,N_29967,N_29992);
or UO_3176 (O_3176,N_29859,N_29940);
and UO_3177 (O_3177,N_29933,N_29846);
xor UO_3178 (O_3178,N_29953,N_29848);
or UO_3179 (O_3179,N_29986,N_29871);
nor UO_3180 (O_3180,N_29805,N_29897);
or UO_3181 (O_3181,N_29951,N_29989);
nor UO_3182 (O_3182,N_29984,N_29999);
nand UO_3183 (O_3183,N_29917,N_29970);
nand UO_3184 (O_3184,N_29827,N_29931);
and UO_3185 (O_3185,N_29966,N_29893);
nand UO_3186 (O_3186,N_29802,N_29817);
and UO_3187 (O_3187,N_29894,N_29904);
or UO_3188 (O_3188,N_29913,N_29841);
nand UO_3189 (O_3189,N_29977,N_29881);
and UO_3190 (O_3190,N_29824,N_29801);
nor UO_3191 (O_3191,N_29993,N_29989);
nand UO_3192 (O_3192,N_29971,N_29822);
xnor UO_3193 (O_3193,N_29985,N_29921);
or UO_3194 (O_3194,N_29960,N_29983);
xor UO_3195 (O_3195,N_29951,N_29876);
nand UO_3196 (O_3196,N_29898,N_29899);
and UO_3197 (O_3197,N_29957,N_29822);
or UO_3198 (O_3198,N_29823,N_29910);
nand UO_3199 (O_3199,N_29952,N_29907);
xnor UO_3200 (O_3200,N_29820,N_29846);
nor UO_3201 (O_3201,N_29903,N_29834);
or UO_3202 (O_3202,N_29895,N_29891);
nor UO_3203 (O_3203,N_29805,N_29876);
nor UO_3204 (O_3204,N_29964,N_29961);
xnor UO_3205 (O_3205,N_29881,N_29991);
and UO_3206 (O_3206,N_29873,N_29822);
and UO_3207 (O_3207,N_29990,N_29979);
or UO_3208 (O_3208,N_29885,N_29985);
and UO_3209 (O_3209,N_29918,N_29929);
nor UO_3210 (O_3210,N_29939,N_29891);
xnor UO_3211 (O_3211,N_29890,N_29988);
nand UO_3212 (O_3212,N_29910,N_29902);
nand UO_3213 (O_3213,N_29942,N_29959);
xnor UO_3214 (O_3214,N_29844,N_29829);
nor UO_3215 (O_3215,N_29964,N_29870);
or UO_3216 (O_3216,N_29837,N_29966);
and UO_3217 (O_3217,N_29860,N_29830);
or UO_3218 (O_3218,N_29905,N_29868);
nand UO_3219 (O_3219,N_29844,N_29951);
or UO_3220 (O_3220,N_29833,N_29970);
or UO_3221 (O_3221,N_29938,N_29901);
and UO_3222 (O_3222,N_29849,N_29927);
xnor UO_3223 (O_3223,N_29847,N_29899);
nand UO_3224 (O_3224,N_29843,N_29874);
nand UO_3225 (O_3225,N_29883,N_29805);
nor UO_3226 (O_3226,N_29890,N_29910);
and UO_3227 (O_3227,N_29867,N_29837);
nor UO_3228 (O_3228,N_29801,N_29896);
xnor UO_3229 (O_3229,N_29841,N_29880);
xnor UO_3230 (O_3230,N_29951,N_29929);
nor UO_3231 (O_3231,N_29896,N_29804);
or UO_3232 (O_3232,N_29982,N_29914);
xnor UO_3233 (O_3233,N_29877,N_29854);
nand UO_3234 (O_3234,N_29872,N_29992);
nor UO_3235 (O_3235,N_29934,N_29962);
nand UO_3236 (O_3236,N_29806,N_29900);
xnor UO_3237 (O_3237,N_29896,N_29978);
or UO_3238 (O_3238,N_29996,N_29934);
xor UO_3239 (O_3239,N_29992,N_29822);
nand UO_3240 (O_3240,N_29932,N_29958);
xnor UO_3241 (O_3241,N_29851,N_29813);
xor UO_3242 (O_3242,N_29877,N_29846);
nand UO_3243 (O_3243,N_29877,N_29916);
or UO_3244 (O_3244,N_29814,N_29876);
xor UO_3245 (O_3245,N_29875,N_29850);
nand UO_3246 (O_3246,N_29823,N_29938);
and UO_3247 (O_3247,N_29874,N_29930);
xnor UO_3248 (O_3248,N_29832,N_29899);
and UO_3249 (O_3249,N_29989,N_29841);
nand UO_3250 (O_3250,N_29946,N_29889);
or UO_3251 (O_3251,N_29829,N_29814);
or UO_3252 (O_3252,N_29815,N_29869);
nor UO_3253 (O_3253,N_29923,N_29884);
and UO_3254 (O_3254,N_29893,N_29808);
and UO_3255 (O_3255,N_29820,N_29899);
nor UO_3256 (O_3256,N_29918,N_29811);
nand UO_3257 (O_3257,N_29881,N_29865);
nor UO_3258 (O_3258,N_29852,N_29968);
nor UO_3259 (O_3259,N_29847,N_29803);
and UO_3260 (O_3260,N_29842,N_29866);
and UO_3261 (O_3261,N_29840,N_29875);
nand UO_3262 (O_3262,N_29914,N_29928);
nand UO_3263 (O_3263,N_29897,N_29844);
and UO_3264 (O_3264,N_29848,N_29922);
nor UO_3265 (O_3265,N_29912,N_29901);
nor UO_3266 (O_3266,N_29967,N_29802);
nand UO_3267 (O_3267,N_29858,N_29952);
nor UO_3268 (O_3268,N_29824,N_29963);
nand UO_3269 (O_3269,N_29885,N_29990);
nor UO_3270 (O_3270,N_29879,N_29811);
nand UO_3271 (O_3271,N_29810,N_29967);
or UO_3272 (O_3272,N_29821,N_29989);
and UO_3273 (O_3273,N_29993,N_29956);
and UO_3274 (O_3274,N_29948,N_29956);
nand UO_3275 (O_3275,N_29842,N_29895);
or UO_3276 (O_3276,N_29853,N_29996);
nor UO_3277 (O_3277,N_29866,N_29960);
xnor UO_3278 (O_3278,N_29863,N_29989);
nor UO_3279 (O_3279,N_29837,N_29968);
xor UO_3280 (O_3280,N_29917,N_29813);
nand UO_3281 (O_3281,N_29942,N_29881);
nor UO_3282 (O_3282,N_29915,N_29879);
xor UO_3283 (O_3283,N_29892,N_29859);
and UO_3284 (O_3284,N_29851,N_29997);
xnor UO_3285 (O_3285,N_29980,N_29896);
or UO_3286 (O_3286,N_29991,N_29803);
or UO_3287 (O_3287,N_29986,N_29840);
xor UO_3288 (O_3288,N_29926,N_29800);
and UO_3289 (O_3289,N_29894,N_29892);
and UO_3290 (O_3290,N_29849,N_29961);
or UO_3291 (O_3291,N_29833,N_29907);
nand UO_3292 (O_3292,N_29896,N_29948);
nand UO_3293 (O_3293,N_29815,N_29823);
nand UO_3294 (O_3294,N_29913,N_29903);
or UO_3295 (O_3295,N_29898,N_29941);
nand UO_3296 (O_3296,N_29857,N_29849);
or UO_3297 (O_3297,N_29923,N_29895);
nor UO_3298 (O_3298,N_29958,N_29801);
nand UO_3299 (O_3299,N_29872,N_29911);
nand UO_3300 (O_3300,N_29997,N_29936);
and UO_3301 (O_3301,N_29905,N_29939);
nor UO_3302 (O_3302,N_29830,N_29920);
and UO_3303 (O_3303,N_29806,N_29823);
nand UO_3304 (O_3304,N_29973,N_29923);
or UO_3305 (O_3305,N_29890,N_29874);
and UO_3306 (O_3306,N_29984,N_29980);
and UO_3307 (O_3307,N_29919,N_29840);
nor UO_3308 (O_3308,N_29954,N_29818);
and UO_3309 (O_3309,N_29868,N_29885);
nand UO_3310 (O_3310,N_29890,N_29943);
nor UO_3311 (O_3311,N_29911,N_29862);
and UO_3312 (O_3312,N_29991,N_29942);
or UO_3313 (O_3313,N_29883,N_29925);
nor UO_3314 (O_3314,N_29828,N_29992);
nor UO_3315 (O_3315,N_29803,N_29907);
or UO_3316 (O_3316,N_29896,N_29956);
or UO_3317 (O_3317,N_29940,N_29974);
nand UO_3318 (O_3318,N_29977,N_29866);
or UO_3319 (O_3319,N_29975,N_29823);
or UO_3320 (O_3320,N_29950,N_29844);
nand UO_3321 (O_3321,N_29909,N_29852);
xnor UO_3322 (O_3322,N_29996,N_29889);
or UO_3323 (O_3323,N_29932,N_29975);
nand UO_3324 (O_3324,N_29865,N_29856);
nor UO_3325 (O_3325,N_29975,N_29831);
nor UO_3326 (O_3326,N_29939,N_29937);
nor UO_3327 (O_3327,N_29979,N_29849);
or UO_3328 (O_3328,N_29874,N_29911);
nand UO_3329 (O_3329,N_29894,N_29948);
xnor UO_3330 (O_3330,N_29832,N_29892);
xnor UO_3331 (O_3331,N_29825,N_29956);
and UO_3332 (O_3332,N_29846,N_29915);
nor UO_3333 (O_3333,N_29896,N_29883);
and UO_3334 (O_3334,N_29921,N_29816);
nand UO_3335 (O_3335,N_29875,N_29934);
nand UO_3336 (O_3336,N_29924,N_29991);
and UO_3337 (O_3337,N_29896,N_29960);
or UO_3338 (O_3338,N_29888,N_29881);
and UO_3339 (O_3339,N_29823,N_29842);
or UO_3340 (O_3340,N_29991,N_29921);
nand UO_3341 (O_3341,N_29926,N_29862);
xnor UO_3342 (O_3342,N_29843,N_29868);
and UO_3343 (O_3343,N_29903,N_29988);
xnor UO_3344 (O_3344,N_29986,N_29968);
xnor UO_3345 (O_3345,N_29949,N_29974);
xnor UO_3346 (O_3346,N_29894,N_29850);
xor UO_3347 (O_3347,N_29911,N_29981);
or UO_3348 (O_3348,N_29808,N_29888);
and UO_3349 (O_3349,N_29925,N_29800);
or UO_3350 (O_3350,N_29939,N_29921);
xnor UO_3351 (O_3351,N_29984,N_29867);
nor UO_3352 (O_3352,N_29982,N_29895);
nor UO_3353 (O_3353,N_29819,N_29915);
or UO_3354 (O_3354,N_29879,N_29897);
and UO_3355 (O_3355,N_29996,N_29928);
xnor UO_3356 (O_3356,N_29878,N_29845);
nand UO_3357 (O_3357,N_29852,N_29825);
xnor UO_3358 (O_3358,N_29899,N_29896);
xor UO_3359 (O_3359,N_29831,N_29868);
nor UO_3360 (O_3360,N_29832,N_29978);
xnor UO_3361 (O_3361,N_29990,N_29938);
nand UO_3362 (O_3362,N_29817,N_29936);
and UO_3363 (O_3363,N_29994,N_29971);
or UO_3364 (O_3364,N_29959,N_29934);
nand UO_3365 (O_3365,N_29998,N_29899);
nor UO_3366 (O_3366,N_29933,N_29842);
xor UO_3367 (O_3367,N_29816,N_29972);
xor UO_3368 (O_3368,N_29926,N_29934);
xnor UO_3369 (O_3369,N_29854,N_29926);
and UO_3370 (O_3370,N_29939,N_29903);
xnor UO_3371 (O_3371,N_29955,N_29822);
xor UO_3372 (O_3372,N_29827,N_29880);
nor UO_3373 (O_3373,N_29809,N_29951);
nand UO_3374 (O_3374,N_29965,N_29851);
nand UO_3375 (O_3375,N_29811,N_29974);
or UO_3376 (O_3376,N_29864,N_29980);
xor UO_3377 (O_3377,N_29818,N_29851);
nand UO_3378 (O_3378,N_29954,N_29964);
or UO_3379 (O_3379,N_29952,N_29968);
or UO_3380 (O_3380,N_29944,N_29961);
nor UO_3381 (O_3381,N_29934,N_29980);
and UO_3382 (O_3382,N_29916,N_29806);
and UO_3383 (O_3383,N_29935,N_29816);
and UO_3384 (O_3384,N_29889,N_29902);
xor UO_3385 (O_3385,N_29808,N_29928);
nand UO_3386 (O_3386,N_29875,N_29844);
and UO_3387 (O_3387,N_29923,N_29837);
nor UO_3388 (O_3388,N_29938,N_29969);
xor UO_3389 (O_3389,N_29918,N_29904);
and UO_3390 (O_3390,N_29957,N_29827);
nor UO_3391 (O_3391,N_29838,N_29858);
and UO_3392 (O_3392,N_29835,N_29977);
and UO_3393 (O_3393,N_29878,N_29811);
nor UO_3394 (O_3394,N_29823,N_29803);
xor UO_3395 (O_3395,N_29921,N_29969);
and UO_3396 (O_3396,N_29887,N_29895);
nand UO_3397 (O_3397,N_29894,N_29876);
xor UO_3398 (O_3398,N_29876,N_29874);
nor UO_3399 (O_3399,N_29895,N_29826);
and UO_3400 (O_3400,N_29970,N_29874);
nor UO_3401 (O_3401,N_29961,N_29911);
and UO_3402 (O_3402,N_29989,N_29834);
and UO_3403 (O_3403,N_29893,N_29996);
and UO_3404 (O_3404,N_29816,N_29945);
xor UO_3405 (O_3405,N_29825,N_29808);
xor UO_3406 (O_3406,N_29845,N_29853);
nand UO_3407 (O_3407,N_29944,N_29931);
nand UO_3408 (O_3408,N_29823,N_29902);
nand UO_3409 (O_3409,N_29895,N_29844);
and UO_3410 (O_3410,N_29897,N_29946);
or UO_3411 (O_3411,N_29978,N_29843);
and UO_3412 (O_3412,N_29992,N_29939);
nor UO_3413 (O_3413,N_29865,N_29971);
nor UO_3414 (O_3414,N_29849,N_29854);
and UO_3415 (O_3415,N_29970,N_29886);
nand UO_3416 (O_3416,N_29812,N_29961);
xor UO_3417 (O_3417,N_29931,N_29918);
or UO_3418 (O_3418,N_29814,N_29967);
nor UO_3419 (O_3419,N_29812,N_29980);
and UO_3420 (O_3420,N_29992,N_29935);
nand UO_3421 (O_3421,N_29975,N_29862);
xor UO_3422 (O_3422,N_29981,N_29876);
nand UO_3423 (O_3423,N_29870,N_29880);
xor UO_3424 (O_3424,N_29955,N_29838);
xor UO_3425 (O_3425,N_29963,N_29839);
or UO_3426 (O_3426,N_29997,N_29954);
nor UO_3427 (O_3427,N_29885,N_29876);
xor UO_3428 (O_3428,N_29860,N_29873);
and UO_3429 (O_3429,N_29860,N_29935);
xnor UO_3430 (O_3430,N_29831,N_29940);
xor UO_3431 (O_3431,N_29832,N_29864);
xor UO_3432 (O_3432,N_29879,N_29996);
and UO_3433 (O_3433,N_29895,N_29981);
nand UO_3434 (O_3434,N_29958,N_29924);
and UO_3435 (O_3435,N_29831,N_29839);
nor UO_3436 (O_3436,N_29920,N_29852);
and UO_3437 (O_3437,N_29974,N_29829);
or UO_3438 (O_3438,N_29957,N_29907);
and UO_3439 (O_3439,N_29838,N_29900);
xnor UO_3440 (O_3440,N_29883,N_29832);
nor UO_3441 (O_3441,N_29927,N_29964);
nand UO_3442 (O_3442,N_29983,N_29921);
xor UO_3443 (O_3443,N_29836,N_29809);
or UO_3444 (O_3444,N_29900,N_29831);
and UO_3445 (O_3445,N_29967,N_29837);
and UO_3446 (O_3446,N_29885,N_29897);
and UO_3447 (O_3447,N_29824,N_29895);
xor UO_3448 (O_3448,N_29965,N_29869);
xor UO_3449 (O_3449,N_29889,N_29807);
nor UO_3450 (O_3450,N_29819,N_29947);
or UO_3451 (O_3451,N_29836,N_29911);
xnor UO_3452 (O_3452,N_29812,N_29970);
and UO_3453 (O_3453,N_29916,N_29865);
and UO_3454 (O_3454,N_29862,N_29828);
xnor UO_3455 (O_3455,N_29938,N_29862);
or UO_3456 (O_3456,N_29868,N_29985);
and UO_3457 (O_3457,N_29803,N_29933);
nand UO_3458 (O_3458,N_29852,N_29951);
nand UO_3459 (O_3459,N_29839,N_29866);
and UO_3460 (O_3460,N_29829,N_29881);
xor UO_3461 (O_3461,N_29826,N_29886);
nor UO_3462 (O_3462,N_29888,N_29925);
nor UO_3463 (O_3463,N_29891,N_29986);
nor UO_3464 (O_3464,N_29856,N_29868);
nand UO_3465 (O_3465,N_29854,N_29975);
nor UO_3466 (O_3466,N_29935,N_29808);
nor UO_3467 (O_3467,N_29921,N_29928);
or UO_3468 (O_3468,N_29981,N_29927);
and UO_3469 (O_3469,N_29898,N_29865);
or UO_3470 (O_3470,N_29815,N_29883);
nor UO_3471 (O_3471,N_29926,N_29865);
xnor UO_3472 (O_3472,N_29987,N_29875);
xor UO_3473 (O_3473,N_29861,N_29846);
nor UO_3474 (O_3474,N_29832,N_29922);
nand UO_3475 (O_3475,N_29961,N_29962);
and UO_3476 (O_3476,N_29960,N_29868);
or UO_3477 (O_3477,N_29921,N_29838);
and UO_3478 (O_3478,N_29839,N_29938);
nor UO_3479 (O_3479,N_29981,N_29825);
or UO_3480 (O_3480,N_29951,N_29858);
nand UO_3481 (O_3481,N_29996,N_29858);
nand UO_3482 (O_3482,N_29919,N_29851);
and UO_3483 (O_3483,N_29989,N_29944);
nor UO_3484 (O_3484,N_29934,N_29960);
xor UO_3485 (O_3485,N_29888,N_29965);
or UO_3486 (O_3486,N_29870,N_29992);
xor UO_3487 (O_3487,N_29809,N_29829);
nor UO_3488 (O_3488,N_29906,N_29851);
nand UO_3489 (O_3489,N_29840,N_29805);
or UO_3490 (O_3490,N_29912,N_29925);
nor UO_3491 (O_3491,N_29834,N_29869);
or UO_3492 (O_3492,N_29860,N_29852);
nor UO_3493 (O_3493,N_29833,N_29814);
and UO_3494 (O_3494,N_29811,N_29875);
xnor UO_3495 (O_3495,N_29802,N_29926);
xnor UO_3496 (O_3496,N_29989,N_29984);
nand UO_3497 (O_3497,N_29863,N_29892);
nand UO_3498 (O_3498,N_29992,N_29806);
nor UO_3499 (O_3499,N_29874,N_29968);
endmodule