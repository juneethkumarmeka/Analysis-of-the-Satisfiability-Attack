module basic_2500_25000_3000_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_2301,In_1912);
or U1 (N_1,In_455,In_290);
and U2 (N_2,In_1340,In_1937);
nand U3 (N_3,In_2462,In_389);
nand U4 (N_4,In_1395,In_2325);
nor U5 (N_5,In_2167,In_502);
and U6 (N_6,In_774,In_754);
nand U7 (N_7,In_858,In_1301);
xor U8 (N_8,In_1190,In_970);
nand U9 (N_9,In_558,In_1413);
nor U10 (N_10,In_904,In_815);
nor U11 (N_11,In_2045,In_788);
and U12 (N_12,In_478,In_1795);
and U13 (N_13,In_2148,In_972);
and U14 (N_14,In_1172,In_2409);
or U15 (N_15,In_308,In_1794);
nor U16 (N_16,In_2171,In_1982);
or U17 (N_17,In_1809,In_941);
or U18 (N_18,In_2401,In_2473);
and U19 (N_19,In_805,In_2156);
and U20 (N_20,In_613,In_2264);
nor U21 (N_21,In_861,In_2039);
nor U22 (N_22,In_32,In_2211);
nor U23 (N_23,In_566,In_72);
nor U24 (N_24,In_895,In_2097);
and U25 (N_25,In_2221,In_2475);
and U26 (N_26,In_2217,In_2165);
nor U27 (N_27,In_827,In_2437);
or U28 (N_28,In_2499,In_706);
nor U29 (N_29,In_1827,In_954);
nand U30 (N_30,In_2418,In_1957);
nor U31 (N_31,In_581,In_95);
nand U32 (N_32,In_1730,In_907);
xnor U33 (N_33,In_764,In_1160);
nand U34 (N_34,In_2210,In_987);
nor U35 (N_35,In_1662,In_283);
nand U36 (N_36,In_1023,In_409);
nand U37 (N_37,In_2372,In_610);
nor U38 (N_38,In_977,In_1867);
or U39 (N_39,In_2207,In_894);
xor U40 (N_40,In_2255,In_380);
or U41 (N_41,In_2061,In_1818);
nor U42 (N_42,In_946,In_1669);
nor U43 (N_43,In_371,In_119);
or U44 (N_44,In_29,In_1067);
or U45 (N_45,In_778,In_199);
nand U46 (N_46,In_410,In_235);
xnor U47 (N_47,In_2104,In_1799);
nand U48 (N_48,In_1053,In_1749);
and U49 (N_49,In_746,In_278);
nor U50 (N_50,In_39,In_497);
nor U51 (N_51,In_1876,In_953);
nand U52 (N_52,In_2294,In_137);
nor U53 (N_53,In_2016,In_265);
or U54 (N_54,In_2223,In_848);
or U55 (N_55,In_1112,In_1570);
xnor U56 (N_56,In_401,In_2429);
or U57 (N_57,In_865,In_479);
or U58 (N_58,In_997,In_1543);
nand U59 (N_59,In_1556,In_1544);
or U60 (N_60,In_1477,In_1904);
nor U61 (N_61,In_2295,In_1065);
nor U62 (N_62,In_792,In_664);
or U63 (N_63,In_794,In_1316);
nand U64 (N_64,In_1616,In_2007);
xnor U65 (N_65,In_1962,In_2428);
nand U66 (N_66,In_2214,In_940);
or U67 (N_67,In_1906,In_147);
nor U68 (N_68,In_768,In_884);
xnor U69 (N_69,In_806,In_173);
xor U70 (N_70,In_1357,In_1322);
or U71 (N_71,In_1502,In_2395);
nor U72 (N_72,In_1341,In_446);
xnor U73 (N_73,In_780,In_918);
nor U74 (N_74,In_703,In_966);
nor U75 (N_75,In_334,In_1949);
nor U76 (N_76,In_1823,In_512);
nor U77 (N_77,In_1927,In_916);
nor U78 (N_78,In_973,In_546);
xor U79 (N_79,In_1014,In_1678);
nand U80 (N_80,In_59,In_728);
nor U81 (N_81,In_1924,In_3);
and U82 (N_82,In_1946,In_1455);
nor U83 (N_83,In_212,In_1295);
or U84 (N_84,In_2312,In_177);
or U85 (N_85,In_574,In_1038);
or U86 (N_86,In_2309,In_2164);
nand U87 (N_87,In_1396,In_926);
nand U88 (N_88,In_258,In_1448);
nor U89 (N_89,In_1165,In_2087);
or U90 (N_90,In_14,In_342);
nand U91 (N_91,In_312,In_1049);
xor U92 (N_92,In_2206,In_1120);
and U93 (N_93,In_451,In_922);
xnor U94 (N_94,In_1028,In_2052);
or U95 (N_95,In_723,In_362);
nand U96 (N_96,In_40,In_866);
nand U97 (N_97,In_1926,In_1353);
xor U98 (N_98,In_1964,In_1457);
xnor U99 (N_99,In_2240,In_180);
nor U100 (N_100,In_201,In_629);
and U101 (N_101,In_717,In_1251);
or U102 (N_102,In_2055,In_1785);
nand U103 (N_103,In_2178,In_1360);
and U104 (N_104,In_1131,In_208);
nor U105 (N_105,In_697,In_1725);
and U106 (N_106,In_698,In_1822);
and U107 (N_107,In_1540,In_416);
nand U108 (N_108,In_915,In_87);
and U109 (N_109,In_30,In_252);
or U110 (N_110,In_183,In_2476);
or U111 (N_111,In_1772,In_795);
nand U112 (N_112,In_1441,In_507);
nand U113 (N_113,In_1105,In_1266);
and U114 (N_114,In_1337,In_114);
or U115 (N_115,In_2226,In_2440);
and U116 (N_116,In_1447,In_2062);
xor U117 (N_117,In_831,In_442);
and U118 (N_118,In_669,In_317);
nor U119 (N_119,In_653,In_309);
nand U120 (N_120,In_1327,In_149);
nand U121 (N_121,In_696,In_1109);
xnor U122 (N_122,In_1950,In_2023);
or U123 (N_123,In_472,In_1967);
nor U124 (N_124,In_73,In_2352);
and U125 (N_125,In_1330,In_631);
nor U126 (N_126,In_1536,In_1599);
xor U127 (N_127,In_286,In_1205);
nor U128 (N_128,In_2291,In_2026);
nand U129 (N_129,In_677,In_656);
nor U130 (N_130,In_514,In_1042);
and U131 (N_131,In_2387,In_590);
nand U132 (N_132,In_383,In_247);
or U133 (N_133,In_2031,In_2154);
xnor U134 (N_134,In_2050,In_693);
nor U135 (N_135,In_1731,In_1796);
or U136 (N_136,In_898,In_1667);
xnor U137 (N_137,In_1636,In_187);
or U138 (N_138,In_575,In_1035);
and U139 (N_139,In_1377,In_474);
nand U140 (N_140,In_1405,In_428);
nand U141 (N_141,In_2285,In_1635);
and U142 (N_142,In_1138,In_412);
and U143 (N_143,In_877,In_226);
and U144 (N_144,In_280,In_2200);
or U145 (N_145,In_2172,In_2105);
and U146 (N_146,In_1249,In_1496);
nand U147 (N_147,In_1420,In_1722);
and U148 (N_148,In_1717,In_569);
or U149 (N_149,In_1270,In_2474);
and U150 (N_150,In_246,In_985);
xor U151 (N_151,In_468,In_1090);
or U152 (N_152,In_108,In_243);
nor U153 (N_153,In_1917,In_896);
and U154 (N_154,In_1506,In_1861);
and U155 (N_155,In_1673,In_709);
nor U156 (N_156,In_879,In_1750);
or U157 (N_157,In_2009,In_829);
nand U158 (N_158,In_1782,In_1524);
and U159 (N_159,In_1974,In_90);
and U160 (N_160,In_1039,In_85);
and U161 (N_161,In_1527,In_415);
xor U162 (N_162,In_2002,In_1983);
nor U163 (N_163,In_583,In_1256);
and U164 (N_164,In_78,In_390);
or U165 (N_165,In_94,In_1808);
and U166 (N_166,In_2355,In_2419);
nor U167 (N_167,In_1993,In_36);
or U168 (N_168,In_294,In_191);
xor U169 (N_169,In_370,In_135);
and U170 (N_170,In_1651,In_1179);
nor U171 (N_171,In_110,In_288);
nand U172 (N_172,In_500,In_2072);
nor U173 (N_173,In_1215,In_27);
nor U174 (N_174,In_1031,In_777);
nor U175 (N_175,In_1850,In_820);
nand U176 (N_176,In_1415,In_2361);
or U177 (N_177,In_144,In_1142);
or U178 (N_178,In_152,In_1541);
nor U179 (N_179,In_1201,In_1253);
and U180 (N_180,In_911,In_945);
and U181 (N_181,In_251,In_2160);
and U182 (N_182,In_2458,In_2296);
nand U183 (N_183,In_1155,In_647);
nand U184 (N_184,In_1248,In_2140);
and U185 (N_185,In_485,In_151);
and U186 (N_186,In_1365,In_337);
and U187 (N_187,In_526,In_622);
or U188 (N_188,In_281,In_2324);
xor U189 (N_189,In_1989,In_2477);
nand U190 (N_190,In_611,In_2470);
and U191 (N_191,In_75,In_1431);
nand U192 (N_192,In_1021,In_1735);
nand U193 (N_193,In_399,In_2189);
and U194 (N_194,In_1319,In_716);
nand U195 (N_195,In_249,In_1774);
and U196 (N_196,In_2251,In_1836);
and U197 (N_197,In_2006,In_419);
or U198 (N_198,In_1871,In_239);
nand U199 (N_199,In_938,In_2193);
xor U200 (N_200,In_453,In_1378);
nor U201 (N_201,In_845,In_1857);
xor U202 (N_202,In_2430,In_1777);
or U203 (N_203,In_878,In_737);
nand U204 (N_204,In_1840,In_2205);
and U205 (N_205,In_1211,In_804);
and U206 (N_206,In_1282,In_530);
or U207 (N_207,In_1855,In_2224);
and U208 (N_208,In_1884,In_2414);
xor U209 (N_209,In_1469,In_157);
nor U210 (N_210,In_494,In_2333);
or U211 (N_211,In_505,In_434);
nor U212 (N_212,In_1079,In_908);
xnor U213 (N_213,In_687,In_1640);
xor U214 (N_214,In_1243,In_106);
nor U215 (N_215,In_341,In_639);
or U216 (N_216,In_1553,In_1700);
nor U217 (N_217,In_2485,In_699);
nand U218 (N_218,In_2405,In_955);
nor U219 (N_219,In_1334,In_1689);
nor U220 (N_220,In_19,In_1901);
nor U221 (N_221,In_1846,In_655);
nand U222 (N_222,In_1606,In_385);
nor U223 (N_223,In_327,In_1728);
nand U224 (N_224,In_1970,In_1308);
and U225 (N_225,In_695,In_1117);
xor U226 (N_226,In_1602,In_842);
or U227 (N_227,In_2273,In_328);
nand U228 (N_228,In_515,In_2199);
and U229 (N_229,In_734,In_21);
and U230 (N_230,In_521,In_807);
nand U231 (N_231,In_1767,In_2111);
nor U232 (N_232,In_793,In_189);
xnor U233 (N_233,In_440,In_1289);
and U234 (N_234,In_1603,In_2010);
nand U235 (N_235,In_1699,In_1189);
xor U236 (N_236,In_1978,In_1586);
nand U237 (N_237,In_2252,In_2481);
and U238 (N_238,In_2351,In_57);
nand U239 (N_239,In_1947,In_772);
nor U240 (N_240,In_22,In_274);
and U241 (N_241,In_2371,In_939);
and U242 (N_242,In_220,In_359);
and U243 (N_243,In_1193,In_2220);
xor U244 (N_244,In_2368,In_437);
nor U245 (N_245,In_1481,In_123);
nor U246 (N_246,In_1775,In_2202);
or U247 (N_247,In_2276,In_762);
nor U248 (N_248,In_2425,In_1787);
xnor U249 (N_249,In_1886,In_1006);
or U250 (N_250,In_196,In_2259);
or U251 (N_251,In_720,In_1139);
or U252 (N_252,In_1575,In_1597);
or U253 (N_253,In_1012,In_1870);
or U254 (N_254,In_2439,In_1727);
nor U255 (N_255,In_64,In_1943);
nand U256 (N_256,In_1625,In_1746);
and U257 (N_257,In_2162,In_96);
or U258 (N_258,In_1621,In_168);
or U259 (N_259,In_1979,In_2054);
and U260 (N_260,In_1492,In_1806);
or U261 (N_261,In_227,In_1310);
nor U262 (N_262,In_1881,In_2246);
nor U263 (N_263,In_2118,In_457);
and U264 (N_264,In_0,In_958);
and U265 (N_265,In_751,In_1280);
nand U266 (N_266,In_1019,In_1116);
nand U267 (N_267,In_2161,In_1841);
or U268 (N_268,In_931,In_1241);
nand U269 (N_269,In_992,In_1362);
and U270 (N_270,In_593,In_158);
or U271 (N_271,In_2121,In_2478);
and U272 (N_272,In_60,In_1615);
nor U273 (N_273,In_2179,In_1686);
nor U274 (N_274,In_1712,In_1545);
and U275 (N_275,In_1748,In_279);
nor U276 (N_276,In_663,In_287);
or U277 (N_277,In_481,In_612);
or U278 (N_278,In_2168,In_1095);
and U279 (N_279,In_830,In_1834);
nand U280 (N_280,In_1733,In_2422);
or U281 (N_281,In_678,In_1565);
and U282 (N_282,In_2091,In_1093);
nor U283 (N_283,In_1157,In_998);
or U284 (N_284,In_1317,In_2131);
and U285 (N_285,In_850,In_426);
nor U286 (N_286,In_1896,In_1017);
xor U287 (N_287,In_1567,In_1088);
nand U288 (N_288,In_1790,In_591);
nor U289 (N_289,In_2185,In_844);
nor U290 (N_290,In_2175,In_1315);
nor U291 (N_291,In_914,In_1258);
nor U292 (N_292,In_2053,In_943);
or U293 (N_293,In_232,In_439);
xnor U294 (N_294,In_11,In_93);
or U295 (N_295,In_1569,In_368);
nand U296 (N_296,In_156,In_2346);
nand U297 (N_297,In_122,In_1410);
nand U298 (N_298,In_285,In_1302);
and U299 (N_299,In_933,In_1493);
and U300 (N_300,In_336,In_1532);
xnor U301 (N_301,In_219,In_418);
and U302 (N_302,In_2347,In_1652);
nand U303 (N_303,In_2298,In_937);
and U304 (N_304,In_26,In_1343);
xor U305 (N_305,In_739,In_2399);
nand U306 (N_306,In_2353,In_892);
nand U307 (N_307,In_2424,In_2377);
xnor U308 (N_308,In_1885,In_833);
and U309 (N_309,In_198,In_1339);
nor U310 (N_310,In_2433,In_15);
nand U311 (N_311,In_260,In_97);
or U312 (N_312,In_1745,In_1223);
nor U313 (N_313,In_745,In_310);
nand U314 (N_314,In_1872,In_1366);
xor U315 (N_315,In_1512,In_2426);
nor U316 (N_316,In_1170,In_1966);
and U317 (N_317,In_2283,In_563);
and U318 (N_318,In_2113,In_1096);
and U319 (N_319,In_1761,In_1259);
nand U320 (N_320,In_2059,In_2230);
or U321 (N_321,In_47,In_2404);
nand U322 (N_322,In_159,In_2281);
and U323 (N_323,In_1626,In_1008);
nor U324 (N_324,In_1007,In_1134);
nand U325 (N_325,In_1274,In_74);
or U326 (N_326,In_1037,In_802);
nor U327 (N_327,In_143,In_1734);
or U328 (N_328,In_1789,In_1875);
and U329 (N_329,In_1480,In_519);
xor U330 (N_330,In_1336,In_1212);
or U331 (N_331,In_1941,In_771);
or U332 (N_332,In_595,In_615);
or U333 (N_333,In_1601,In_917);
or U334 (N_334,In_1425,In_1788);
nor U335 (N_335,In_400,In_588);
or U336 (N_336,In_2015,In_467);
nor U337 (N_337,In_568,In_1406);
xor U338 (N_338,In_2146,In_1491);
nand U339 (N_339,In_9,In_1972);
xor U340 (N_340,In_424,In_1558);
nor U341 (N_341,In_1408,In_466);
and U342 (N_342,In_1400,In_1698);
and U343 (N_343,In_387,In_1679);
and U344 (N_344,In_2106,In_2108);
and U345 (N_345,In_819,In_1342);
xnor U346 (N_346,In_107,In_1309);
and U347 (N_347,In_1844,In_1898);
and U348 (N_348,In_1034,In_184);
nor U349 (N_349,In_2034,In_1);
nor U350 (N_350,In_195,In_432);
nor U351 (N_351,In_978,In_1272);
nor U352 (N_352,In_465,In_1487);
nor U353 (N_353,In_705,In_2212);
nand U354 (N_354,In_1838,In_1675);
and U355 (N_355,In_203,In_111);
xor U356 (N_356,In_1650,In_1287);
and U357 (N_357,In_1304,In_1268);
or U358 (N_358,In_2332,In_1600);
xnor U359 (N_359,In_68,In_525);
nor U360 (N_360,In_1835,In_379);
nand U361 (N_361,In_1375,In_2367);
or U362 (N_362,In_361,In_891);
or U363 (N_363,In_200,In_641);
nand U364 (N_364,In_407,In_298);
nor U365 (N_365,In_901,In_2345);
nor U366 (N_366,In_2443,In_810);
nor U367 (N_367,In_1998,In_1364);
or U368 (N_368,In_2065,In_1637);
and U369 (N_369,In_2003,In_2147);
nand U370 (N_370,In_1323,In_523);
nand U371 (N_371,In_315,In_1299);
and U372 (N_372,In_1475,In_2288);
nand U373 (N_373,In_33,In_1345);
and U374 (N_374,In_1032,In_1837);
and U375 (N_375,In_599,In_1991);
and U376 (N_376,In_165,In_1184);
or U377 (N_377,In_2423,In_2466);
nor U378 (N_378,In_2303,In_1664);
or U379 (N_379,In_1624,In_1780);
nand U380 (N_380,In_822,In_394);
nand U381 (N_381,In_2051,In_2103);
nor U382 (N_382,In_1942,In_2384);
and U383 (N_383,In_726,In_2075);
xnor U384 (N_384,In_2231,In_809);
and U385 (N_385,In_1704,In_702);
nor U386 (N_386,In_503,In_1737);
nand U387 (N_387,In_162,In_871);
and U388 (N_388,In_1374,In_2304);
xnor U389 (N_389,In_690,In_221);
nand U390 (N_390,In_1203,In_1436);
or U391 (N_391,In_1376,In_344);
nand U392 (N_392,In_1511,In_1427);
and U393 (N_393,In_531,In_2127);
and U394 (N_394,In_242,In_1706);
nor U395 (N_395,In_1312,In_1368);
and U396 (N_396,In_1951,In_2037);
nor U397 (N_397,In_2300,In_417);
nor U398 (N_398,In_707,In_1275);
and U399 (N_399,In_1645,In_190);
or U400 (N_400,In_2013,In_1468);
or U401 (N_401,In_1716,In_1338);
or U402 (N_402,In_1288,In_1617);
or U403 (N_403,In_1784,In_598);
or U404 (N_404,In_2469,In_2014);
nor U405 (N_405,In_1546,In_269);
xor U406 (N_406,In_2479,In_617);
nand U407 (N_407,In_2115,In_1000);
and U408 (N_408,In_99,In_729);
nor U409 (N_409,In_828,In_1005);
nand U410 (N_410,In_2484,In_2307);
nor U411 (N_411,In_1084,In_749);
and U412 (N_412,In_1634,In_2095);
xnor U413 (N_413,In_1646,In_1352);
nand U414 (N_414,In_2394,In_1981);
or U415 (N_415,In_495,In_392);
nand U416 (N_416,In_930,In_24);
and U417 (N_417,In_1654,In_1026);
and U418 (N_418,In_2397,In_2084);
nor U419 (N_419,In_1618,In_1015);
xnor U420 (N_420,In_2227,In_1622);
nor U421 (N_421,In_1925,In_1828);
nor U422 (N_422,In_1639,In_37);
and U423 (N_423,In_471,In_2079);
xnor U424 (N_424,In_112,In_218);
nor U425 (N_425,In_1713,In_231);
and U426 (N_426,In_719,In_711);
nor U427 (N_427,In_2086,In_1574);
xnor U428 (N_428,In_303,In_547);
or U429 (N_429,In_967,In_1633);
xor U430 (N_430,In_211,In_2044);
xnor U431 (N_431,In_347,In_2310);
nor U432 (N_432,In_1144,In_999);
nand U433 (N_433,In_1895,In_983);
or U434 (N_434,In_420,In_592);
xor U435 (N_435,In_1490,In_1619);
xnor U436 (N_436,In_1968,In_1303);
nor U437 (N_437,In_2092,In_1409);
xnor U438 (N_438,In_305,In_1999);
and U439 (N_439,In_769,In_619);
or U440 (N_440,In_799,In_1324);
and U441 (N_441,In_533,In_2378);
and U442 (N_442,In_2237,In_1451);
and U443 (N_443,In_854,In_1389);
and U444 (N_444,In_1507,In_1629);
or U445 (N_445,In_863,In_2391);
nor U446 (N_446,In_2434,In_880);
and U447 (N_447,In_534,In_1632);
xor U448 (N_448,In_607,In_1161);
and U449 (N_449,In_52,In_637);
and U450 (N_450,In_1052,In_1379);
nand U451 (N_451,In_1099,In_657);
nor U452 (N_452,In_976,In_1430);
nand U453 (N_453,In_2001,In_1938);
and U454 (N_454,In_1214,In_1198);
nand U455 (N_455,In_2432,In_779);
nand U456 (N_456,In_1786,In_1504);
nor U457 (N_457,In_2363,In_975);
or U458 (N_458,In_1125,In_1584);
nor U459 (N_459,In_2228,In_766);
and U460 (N_460,In_755,In_1519);
nor U461 (N_461,In_1221,In_89);
nand U462 (N_462,In_694,In_1935);
nand U463 (N_463,In_1228,In_1412);
nand U464 (N_464,In_783,In_2017);
and U465 (N_465,In_121,In_1182);
or U466 (N_466,In_2201,In_2317);
nand U467 (N_467,In_2491,In_510);
nor U468 (N_468,In_244,In_1663);
nor U469 (N_469,In_2155,In_704);
nor U470 (N_470,In_2472,In_463);
nor U471 (N_471,In_1798,In_2305);
nand U472 (N_472,In_1394,In_322);
nor U473 (N_473,In_1894,In_1812);
nor U474 (N_474,In_2166,In_7);
or U475 (N_475,In_913,In_760);
and U476 (N_476,In_798,In_2225);
and U477 (N_477,In_561,In_2339);
nor U478 (N_478,In_1577,In_348);
and U479 (N_479,In_1236,In_1768);
nand U480 (N_480,In_98,In_1252);
nor U481 (N_481,In_2257,In_364);
nand U482 (N_482,In_773,In_23);
or U483 (N_483,In_857,In_1525);
nand U484 (N_484,In_2270,In_2327);
nand U485 (N_485,In_1561,In_665);
and U486 (N_486,In_1354,In_787);
and U487 (N_487,In_834,In_950);
xnor U488 (N_488,In_1089,In_1571);
nand U489 (N_489,In_1220,In_2457);
or U490 (N_490,In_585,In_589);
nand U491 (N_491,In_268,In_2020);
nand U492 (N_492,In_1370,In_736);
nor U493 (N_493,In_2186,In_375);
or U494 (N_494,In_2452,In_947);
or U495 (N_495,In_2323,In_722);
and U496 (N_496,In_763,In_326);
nand U497 (N_497,In_1444,In_2046);
nand U498 (N_498,In_353,In_5);
or U499 (N_499,In_1534,In_867);
nor U500 (N_500,In_1802,In_1631);
nand U501 (N_501,In_2322,In_381);
nand U502 (N_502,In_2018,In_1063);
nor U503 (N_503,In_271,In_735);
nor U504 (N_504,In_2187,In_1910);
nor U505 (N_505,In_539,In_56);
xor U506 (N_506,In_1489,In_2450);
or U507 (N_507,In_1911,In_586);
nand U508 (N_508,In_1889,In_1714);
or U509 (N_509,In_2278,In_1174);
and U510 (N_510,In_2321,In_1756);
or U511 (N_511,In_346,In_2336);
and U512 (N_512,In_1801,In_142);
or U513 (N_513,In_504,In_1992);
nor U514 (N_514,In_275,In_1783);
and U515 (N_515,In_1583,In_357);
nand U516 (N_516,In_2157,In_1743);
and U517 (N_517,In_781,In_360);
and U518 (N_518,In_1773,In_1554);
nor U519 (N_519,In_113,In_1080);
and U520 (N_520,In_1564,In_2128);
nand U521 (N_521,In_484,In_1133);
nand U522 (N_522,In_597,In_276);
or U523 (N_523,In_2453,In_1391);
nor U524 (N_524,In_529,In_2181);
nor U525 (N_525,In_2239,In_1175);
xnor U526 (N_526,In_571,In_927);
nand U527 (N_527,In_942,In_1437);
nor U528 (N_528,In_461,In_145);
and U529 (N_529,In_1533,In_1563);
and U530 (N_530,In_1030,In_2151);
nand U531 (N_531,In_800,In_1180);
or U532 (N_532,In_1851,In_4);
and U533 (N_533,In_1074,In_58);
nand U534 (N_534,In_1903,In_2070);
and U535 (N_535,In_1588,In_1043);
or U536 (N_536,In_1859,In_160);
nand U537 (N_537,In_363,In_2431);
xor U538 (N_538,In_1426,In_1335);
xor U539 (N_539,In_1776,In_166);
and U540 (N_540,In_2004,In_373);
and U541 (N_541,In_1411,In_1542);
and U542 (N_542,In_2033,In_2057);
nand U543 (N_543,In_2027,In_2169);
or U544 (N_544,In_84,In_2269);
or U545 (N_545,In_120,In_1548);
xor U546 (N_546,In_1445,In_559);
nor U547 (N_547,In_1505,In_626);
and U548 (N_548,In_2150,In_701);
and U549 (N_549,In_1458,In_910);
xor U550 (N_550,In_759,In_1705);
or U551 (N_551,In_1207,In_1510);
nor U552 (N_552,In_1181,In_614);
nand U553 (N_553,In_724,In_1351);
nor U554 (N_554,In_1143,In_445);
and U555 (N_555,In_1158,In_1146);
nand U556 (N_556,In_1693,In_254);
nor U557 (N_557,In_1291,In_1658);
and U558 (N_558,In_1056,In_1865);
nor U559 (N_559,In_470,In_382);
and U560 (N_560,In_2083,In_1909);
and U561 (N_561,In_225,In_1129);
or U562 (N_562,In_54,In_1726);
nand U563 (N_563,In_1036,In_215);
nor U564 (N_564,In_623,In_450);
xor U565 (N_565,In_2293,In_662);
nand U566 (N_566,In_1149,In_2144);
nand U567 (N_567,In_1422,In_126);
or U568 (N_568,In_272,In_1108);
or U569 (N_569,In_2445,In_493);
and U570 (N_570,In_2344,In_1551);
or U571 (N_571,In_1804,In_1959);
nor U572 (N_572,In_1847,In_730);
nand U573 (N_573,In_2385,In_104);
and U574 (N_574,In_2012,In_163);
xnor U575 (N_575,In_2388,In_2334);
and U576 (N_576,In_282,In_971);
xnor U577 (N_577,In_1209,In_369);
nor U578 (N_578,In_1246,In_1676);
or U579 (N_579,In_1046,In_140);
and U580 (N_580,In_2341,In_1568);
nand U581 (N_581,In_2261,In_1845);
and U582 (N_582,In_2328,In_443);
nor U583 (N_583,In_1332,In_2005);
or U584 (N_584,In_1098,In_2060);
nand U585 (N_585,In_262,In_169);
and U586 (N_586,In_366,In_584);
nor U587 (N_587,In_1986,In_1763);
nor U588 (N_588,In_2125,In_13);
or U589 (N_589,In_1944,In_899);
and U590 (N_590,In_1643,In_1418);
or U591 (N_591,In_1119,In_430);
nand U592 (N_592,In_1358,In_2149);
and U593 (N_593,In_1744,In_2386);
nor U594 (N_594,In_2064,In_2250);
nand U595 (N_595,In_621,In_193);
nor U596 (N_596,In_367,In_1916);
or U597 (N_597,In_352,In_349);
and U598 (N_598,In_840,In_127);
or U599 (N_599,In_109,In_1987);
nor U600 (N_600,In_2258,In_1024);
nor U601 (N_601,In_2292,In_1753);
nand U602 (N_602,In_1459,In_80);
xor U603 (N_603,In_2209,In_31);
or U604 (N_604,In_2408,In_1852);
and U605 (N_605,In_1649,In_2098);
or U606 (N_606,In_1709,In_1385);
and U607 (N_607,In_2043,In_961);
nor U608 (N_608,In_436,In_1856);
or U609 (N_609,In_1883,In_44);
nand U610 (N_610,In_2253,In_2000);
and U611 (N_611,In_2197,In_1694);
xnor U612 (N_612,In_1874,In_1176);
or U613 (N_613,In_393,In_1419);
xnor U614 (N_614,In_2286,In_1869);
xnor U615 (N_615,In_757,In_1933);
nor U616 (N_616,In_1839,In_949);
nor U617 (N_617,In_138,In_25);
nor U618 (N_618,In_2152,In_1196);
xnor U619 (N_619,In_2195,In_981);
and U620 (N_620,In_649,In_887);
and U621 (N_621,In_172,In_230);
nand U622 (N_622,In_2329,In_883);
nor U623 (N_623,In_638,In_2343);
xnor U624 (N_624,In_1123,In_1825);
xnor U625 (N_625,In_422,In_83);
or U626 (N_626,In_1297,In_345);
and U627 (N_627,In_164,In_2159);
or U628 (N_628,In_413,In_1860);
nand U629 (N_629,In_1393,In_1905);
xor U630 (N_630,In_1216,In_1347);
nand U631 (N_631,In_2102,In_1596);
or U632 (N_632,In_1075,In_161);
or U633 (N_633,In_1724,In_1306);
or U634 (N_634,In_1446,In_1107);
nor U635 (N_635,In_508,In_873);
nor U636 (N_636,In_1665,In_823);
nor U637 (N_637,In_1826,In_2486);
nor U638 (N_638,In_1238,In_2208);
or U639 (N_639,In_291,In_270);
and U640 (N_640,In_544,In_1882);
and U641 (N_641,In_600,In_452);
and U642 (N_642,In_1578,In_102);
nand U643 (N_643,In_969,In_1399);
nor U644 (N_644,In_1269,In_2435);
nand U645 (N_645,In_2085,In_684);
and U646 (N_646,In_1740,In_1115);
nand U647 (N_647,In_1589,In_1738);
nand U648 (N_648,In_50,In_1050);
nand U649 (N_649,In_1580,In_1244);
or U650 (N_650,In_1305,In_1791);
or U651 (N_651,In_1614,In_761);
xnor U652 (N_652,In_1279,In_1325);
nand U653 (N_653,In_889,In_1055);
or U654 (N_654,In_2058,In_194);
and U655 (N_655,In_1057,In_1975);
or U656 (N_656,In_1832,In_594);
nor U657 (N_657,In_209,In_909);
nor U658 (N_658,In_1990,In_1781);
xnor U659 (N_659,In_2066,In_738);
or U660 (N_660,In_213,In_1539);
nand U661 (N_661,In_1326,In_289);
and U662 (N_662,In_306,In_537);
and U663 (N_663,In_689,In_527);
nand U664 (N_664,In_1058,In_2247);
xnor U665 (N_665,In_2137,In_1918);
or U666 (N_666,In_606,In_372);
nand U667 (N_667,In_1083,In_296);
nand U668 (N_668,In_1206,In_188);
nor U669 (N_669,In_2390,In_1113);
or U670 (N_670,In_1450,In_2460);
nor U671 (N_671,In_1939,In_1778);
and U672 (N_672,In_1276,In_1091);
and U673 (N_673,In_1923,In_2268);
or U674 (N_674,In_1222,In_1456);
nand U675 (N_675,In_1429,In_1521);
nand U676 (N_676,In_2348,In_646);
or U677 (N_677,In_580,In_1495);
or U678 (N_678,In_2331,In_1403);
nor U679 (N_679,In_2267,In_797);
or U680 (N_680,In_782,In_2126);
and U681 (N_681,In_1819,In_8);
and U682 (N_682,In_1473,In_1638);
nor U683 (N_683,In_1815,In_2373);
xnor U684 (N_684,In_1518,In_2272);
nor U685 (N_685,In_2074,In_1764);
nor U686 (N_686,In_1854,In_1520);
nor U687 (N_687,In_2360,In_905);
or U688 (N_688,In_1922,In_217);
nor U689 (N_689,In_2441,In_1264);
or U690 (N_690,In_1278,In_1723);
and U691 (N_691,In_1141,In_1585);
xor U692 (N_692,In_1668,In_386);
nand U693 (N_693,In_2133,In_1217);
nor U694 (N_694,In_1497,In_1611);
nand U695 (N_695,In_101,In_1284);
xnor U696 (N_696,In_2280,In_2238);
nand U697 (N_697,In_1842,In_2145);
xor U698 (N_698,In_549,In_192);
and U699 (N_699,In_35,In_1156);
and U700 (N_700,In_124,In_1087);
nand U701 (N_701,In_1690,In_438);
and U702 (N_702,In_2383,In_676);
nor U703 (N_703,In_811,In_538);
and U704 (N_704,In_1111,In_1077);
nand U705 (N_705,In_605,In_1188);
and U706 (N_706,In_1702,In_919);
nand U707 (N_707,In_785,In_1535);
nand U708 (N_708,In_1522,In_2071);
and U709 (N_709,In_1286,In_499);
and U710 (N_710,In_2342,In_2364);
or U711 (N_711,In_2335,In_301);
nor U712 (N_712,In_1824,In_181);
nand U713 (N_713,In_2421,In_167);
or U714 (N_714,In_1516,In_365);
or U715 (N_715,In_2311,In_849);
nor U716 (N_716,In_959,In_1609);
nand U717 (N_717,In_1879,In_1566);
or U718 (N_718,In_2184,In_963);
nand U719 (N_719,In_673,In_1594);
and U720 (N_720,In_10,In_2029);
nand U721 (N_721,In_1598,In_572);
or U722 (N_722,In_1194,In_1402);
nand U723 (N_723,In_216,In_2381);
or U724 (N_724,In_1682,In_557);
and U725 (N_725,In_1915,In_578);
or U726 (N_726,In_1661,In_2244);
nand U727 (N_727,In_1177,In_6);
nor U728 (N_728,In_1136,In_292);
xor U729 (N_729,In_2493,In_2011);
nand U730 (N_730,In_444,In_2492);
nor U731 (N_731,In_1963,In_1386);
nand U732 (N_732,In_1159,In_1262);
nand U733 (N_733,In_423,In_903);
nand U734 (N_734,In_321,In_1033);
nor U735 (N_735,In_1687,In_994);
nand U736 (N_736,In_408,In_1692);
and U737 (N_737,In_1311,In_1423);
or U738 (N_738,In_1210,In_1320);
or U739 (N_739,In_1380,In_2213);
nor U740 (N_740,In_1440,In_801);
nand U741 (N_741,In_1392,In_1200);
xor U742 (N_742,In_1404,In_1439);
xnor U743 (N_743,In_2056,In_618);
and U744 (N_744,In_1674,In_2448);
nand U745 (N_745,In_2359,In_1054);
nor U746 (N_746,In_1929,In_255);
or U747 (N_747,In_2287,In_1514);
or U748 (N_748,In_920,In_948);
and U749 (N_749,In_924,In_934);
or U750 (N_750,In_46,In_2024);
xor U751 (N_751,In_555,In_814);
nand U752 (N_752,In_1833,In_1830);
and U753 (N_753,In_1659,In_1656);
and U754 (N_754,In_2289,In_2315);
nor U755 (N_755,In_263,In_1752);
xor U756 (N_756,In_1250,In_765);
nand U757 (N_757,In_2094,In_1529);
nor U758 (N_758,In_1573,In_1478);
nor U759 (N_759,In_770,In_1234);
or U760 (N_760,In_552,In_1498);
or U761 (N_761,In_1528,In_2035);
xnor U762 (N_762,In_2194,In_17);
xnor U763 (N_763,In_1025,In_1292);
xor U764 (N_764,In_1434,In_154);
nand U765 (N_765,In_1041,In_253);
nor U766 (N_766,In_1137,In_1729);
nand U767 (N_767,In_18,In_2494);
or U768 (N_768,In_775,In_388);
nand U769 (N_769,In_2249,In_460);
nor U770 (N_770,In_1736,In_391);
nor U771 (N_771,In_1562,In_2402);
nor U772 (N_772,In_2297,In_233);
nand U773 (N_773,In_2090,In_900);
nand U774 (N_774,In_812,In_1988);
or U775 (N_775,In_1930,In_307);
and U776 (N_776,In_492,In_1281);
or U777 (N_777,In_425,In_67);
and U778 (N_778,In_2136,In_870);
nand U779 (N_779,In_2109,In_324);
nand U780 (N_780,In_1483,In_1464);
xor U781 (N_781,In_1371,In_2314);
and U782 (N_782,In_293,In_632);
and U783 (N_783,In_1460,In_2482);
and U784 (N_784,In_2480,In_1612);
and U785 (N_785,In_875,In_634);
nor U786 (N_786,In_2379,In_1681);
nand U787 (N_787,In_2416,In_1265);
nor U788 (N_788,In_2077,In_1466);
and U789 (N_789,In_2410,In_1164);
or U790 (N_790,In_2417,In_1106);
or U791 (N_791,In_16,In_936);
nand U792 (N_792,In_441,In_986);
and U793 (N_793,In_990,In_486);
nor U794 (N_794,In_1173,In_316);
nor U795 (N_795,In_989,In_535);
nor U796 (N_796,In_1711,In_397);
nand U797 (N_797,In_582,In_2313);
or U798 (N_798,In_1240,In_1047);
nor U799 (N_799,In_602,In_2319);
nor U800 (N_800,In_1858,In_2497);
and U801 (N_801,In_186,In_1103);
and U802 (N_802,In_1018,In_1344);
nand U803 (N_803,In_1620,In_1071);
nor U804 (N_804,In_259,In_2369);
and U805 (N_805,In_650,In_1688);
or U806 (N_806,In_536,In_691);
nand U807 (N_807,In_951,In_1064);
nor U808 (N_808,In_708,In_1428);
and U809 (N_809,In_1670,In_1537);
and U810 (N_810,In_1742,In_1307);
and U811 (N_811,In_674,In_63);
nor U812 (N_812,In_1421,In_509);
xnor U813 (N_813,In_1011,In_1022);
and U814 (N_814,In_2021,In_1013);
nor U815 (N_815,In_141,In_1934);
or U816 (N_816,In_1226,In_1820);
nor U817 (N_817,In_2290,In_1432);
or U818 (N_818,In_128,In_1442);
nor U819 (N_819,In_1230,In_224);
and U820 (N_820,In_1931,In_921);
nand U821 (N_821,In_517,In_1239);
xnor U822 (N_822,In_1576,In_516);
nand U823 (N_823,In_996,In_1233);
and U824 (N_824,In_2455,In_1081);
and U825 (N_825,In_587,In_2177);
and U826 (N_826,In_1192,In_758);
xnor U827 (N_827,In_1593,In_2114);
nor U828 (N_828,In_2248,In_2204);
nor U829 (N_829,In_1500,In_340);
or U830 (N_830,In_843,In_1849);
or U831 (N_831,In_1443,In_2495);
nand U832 (N_832,In_1610,In_1218);
and U833 (N_833,In_1069,In_570);
or U834 (N_834,In_573,In_2170);
nor U835 (N_835,In_2076,In_257);
or U836 (N_836,In_1607,In_1293);
or U837 (N_837,In_489,In_876);
or U838 (N_838,In_988,In_1314);
nor U839 (N_839,In_1199,In_601);
or U840 (N_840,In_1001,In_1465);
nor U841 (N_841,In_635,In_553);
nor U842 (N_842,In_1720,In_744);
or U843 (N_843,In_1004,In_100);
nor U844 (N_844,In_2374,In_1277);
or U845 (N_845,In_1759,In_1973);
or U846 (N_846,In_1094,In_912);
nor U847 (N_847,In_1648,In_952);
nor U848 (N_848,In_2407,In_1061);
xor U849 (N_849,In_682,In_1739);
nor U850 (N_850,In_1769,In_2132);
nor U851 (N_851,In_932,In_2349);
or U852 (N_852,In_414,In_240);
nand U853 (N_853,In_825,In_2337);
nand U854 (N_854,In_171,In_1467);
and U855 (N_855,In_1066,In_784);
nor U856 (N_856,In_1685,In_1044);
nor U857 (N_857,In_49,In_2442);
or U858 (N_858,In_1592,In_577);
and U859 (N_859,In_2260,In_1140);
and U860 (N_860,In_714,In_609);
nand U861 (N_861,In_1641,In_477);
nor U862 (N_862,In_1333,In_2153);
nor U863 (N_863,In_897,In_1710);
or U864 (N_864,In_715,In_1398);
and U865 (N_865,In_202,In_2229);
and U866 (N_866,In_45,In_2365);
or U867 (N_867,In_902,In_1997);
nor U868 (N_868,In_395,In_311);
nand U869 (N_869,In_402,In_335);
nor U870 (N_870,In_1765,In_1866);
nor U871 (N_871,In_2110,In_562);
xor U872 (N_872,In_543,In_1073);
nor U873 (N_873,In_648,In_2420);
and U874 (N_874,In_1471,In_241);
nand U875 (N_875,In_1484,In_753);
nor U876 (N_876,In_882,In_925);
or U877 (N_877,In_65,In_747);
nand U878 (N_878,In_354,In_2129);
or U879 (N_879,In_2263,In_838);
and U880 (N_880,In_604,In_150);
and U881 (N_881,In_1132,In_1102);
or U882 (N_882,In_132,In_266);
nor U883 (N_883,In_750,In_2182);
nand U884 (N_884,In_207,In_906);
and U885 (N_885,In_480,In_672);
nor U886 (N_886,In_980,In_153);
or U887 (N_887,In_733,In_1232);
nor U888 (N_888,In_2218,In_851);
nand U889 (N_889,In_1985,In_2256);
and U890 (N_890,In_1242,In_2107);
nor U891 (N_891,In_603,In_129);
and U892 (N_892,In_1914,In_628);
nand U893 (N_893,In_1868,In_796);
and U894 (N_894,In_2490,In_458);
xor U895 (N_895,In_378,In_743);
and U896 (N_896,In_853,In_1863);
nor U897 (N_897,In_645,In_1070);
or U898 (N_898,In_2173,In_1653);
nor U899 (N_899,In_28,In_1355);
xnor U900 (N_900,In_1604,In_860);
nand U901 (N_901,In_1118,In_1817);
and U902 (N_902,In_2116,In_974);
nor U903 (N_903,In_1581,In_1696);
nor U904 (N_904,In_376,In_1273);
or U905 (N_905,In_1697,In_476);
or U906 (N_906,In_264,In_1891);
or U907 (N_907,In_616,In_483);
nor U908 (N_908,In_1862,In_178);
nand U909 (N_909,In_313,In_1453);
and U910 (N_910,In_522,In_1816);
nor U911 (N_911,In_2,In_204);
nand U912 (N_912,In_1779,In_816);
nor U913 (N_913,In_1848,In_1187);
and U914 (N_914,In_1363,In_2362);
nor U915 (N_915,In_1407,In_2068);
or U916 (N_916,In_2463,In_214);
or U917 (N_917,In_1147,In_1488);
or U918 (N_918,In_1958,In_1900);
xor U919 (N_919,In_42,In_2139);
xor U920 (N_920,In_404,In_2356);
nand U921 (N_921,In_69,In_1104);
nand U922 (N_922,In_767,In_2019);
nand U923 (N_923,In_2236,In_222);
nor U924 (N_924,In_1557,In_82);
nand U925 (N_925,In_473,In_2483);
nor U926 (N_926,In_732,In_1913);
or U927 (N_927,In_314,In_1538);
xnor U928 (N_928,In_2142,In_41);
and U929 (N_929,In_491,In_1227);
nand U930 (N_930,In_1741,In_2245);
nand U931 (N_931,In_1237,In_2444);
and U932 (N_932,In_1971,In_1328);
and U933 (N_933,In_545,In_2464);
and U934 (N_934,In_1029,In_1100);
nor U935 (N_935,In_12,In_134);
and U936 (N_936,In_429,In_1953);
and U937 (N_937,In_1919,In_670);
and U938 (N_938,In_528,In_1461);
and U939 (N_939,In_1153,In_482);
nor U940 (N_940,In_1695,In_1762);
and U941 (N_941,In_1245,In_1559);
nand U942 (N_942,In_2036,In_1549);
nor U943 (N_943,In_1254,In_1045);
and U944 (N_944,In_1474,In_62);
nand U945 (N_945,In_2163,In_2096);
or U946 (N_946,In_1068,In_700);
and U947 (N_947,In_331,In_333);
nand U948 (N_948,In_1126,In_92);
and U949 (N_949,In_139,In_2080);
nor U950 (N_950,In_2047,In_791);
and U951 (N_951,In_1873,In_1127);
nand U952 (N_952,In_105,In_643);
nand U953 (N_953,In_740,In_1644);
nor U954 (N_954,In_1555,In_2396);
and U955 (N_955,In_1145,In_725);
and U956 (N_956,In_20,In_2176);
nor U957 (N_957,In_1294,In_2082);
nor U958 (N_958,In_520,In_459);
nand U959 (N_959,In_1263,In_350);
nand U960 (N_960,In_651,In_2338);
or U961 (N_961,In_1082,In_496);
and U962 (N_962,In_1792,In_742);
nand U963 (N_963,In_2048,In_76);
nand U964 (N_964,In_1130,In_1010);
xnor U965 (N_965,In_1965,In_2040);
nand U966 (N_966,In_2318,In_1367);
and U967 (N_967,In_1318,In_2498);
or U968 (N_968,In_273,In_1899);
nor U969 (N_969,In_320,In_727);
nor U970 (N_970,In_1721,In_1387);
nor U971 (N_971,In_862,In_338);
xor U972 (N_972,In_789,In_1897);
and U973 (N_973,In_1452,In_872);
and U974 (N_974,In_2271,In_435);
and U975 (N_975,In_596,In_1290);
nor U976 (N_976,In_403,In_620);
nor U977 (N_977,In_2412,In_1811);
nor U978 (N_978,In_1952,In_2254);
nand U979 (N_979,In_2191,In_1300);
nor U980 (N_980,In_118,In_1121);
and U981 (N_981,In_2465,In_642);
nand U982 (N_982,In_852,In_1349);
nor U983 (N_983,In_685,In_1002);
nand U984 (N_984,In_1800,In_1920);
nand U985 (N_985,In_965,In_1503);
and U986 (N_986,In_1313,In_835);
xnor U987 (N_987,In_433,In_1195);
nor U988 (N_988,In_2487,In_238);
or U989 (N_989,In_2188,In_2030);
and U990 (N_990,In_2427,In_1627);
xor U991 (N_991,In_1152,In_1948);
and U992 (N_992,In_1283,In_556);
or U993 (N_993,In_1151,In_431);
and U994 (N_994,In_302,In_130);
nor U995 (N_995,In_2122,In_692);
nand U996 (N_996,In_170,In_1508);
xnor U997 (N_997,In_1976,In_1671);
nand U998 (N_998,In_355,In_1329);
or U999 (N_999,In_2117,In_929);
and U1000 (N_1000,In_1085,In_1062);
xnor U1001 (N_1001,In_935,In_2265);
or U1002 (N_1002,In_608,In_229);
nand U1003 (N_1003,In_1719,In_2219);
and U1004 (N_1004,In_2192,In_1754);
or U1005 (N_1005,In_667,In_1016);
xor U1006 (N_1006,In_1417,In_748);
nor U1007 (N_1007,In_1051,In_2436);
nand U1008 (N_1008,In_984,In_551);
nor U1009 (N_1009,In_1169,In_1433);
nor U1010 (N_1010,In_133,In_1167);
or U1011 (N_1011,In_824,In_817);
and U1012 (N_1012,In_487,In_2042);
nor U1013 (N_1013,In_2063,In_464);
nor U1014 (N_1014,In_688,In_2235);
nand U1015 (N_1015,In_2398,In_2446);
nand U1016 (N_1016,In_2354,In_131);
xnor U1017 (N_1017,In_837,In_1660);
nor U1018 (N_1018,In_228,In_1135);
or U1019 (N_1019,In_1902,In_982);
and U1020 (N_1020,In_2262,In_1797);
and U1021 (N_1021,In_1261,In_893);
nand U1022 (N_1022,In_721,In_396);
nor U1023 (N_1023,In_2067,In_297);
nand U1024 (N_1024,In_675,In_923);
and U1025 (N_1025,In_1229,In_1285);
or U1026 (N_1026,In_2134,In_1666);
nand U1027 (N_1027,In_1486,In_1482);
xnor U1028 (N_1028,In_1476,In_1163);
and U1029 (N_1029,In_48,In_2456);
nand U1030 (N_1030,In_2049,In_627);
or U1031 (N_1031,In_511,In_1590);
nor U1032 (N_1032,In_1231,In_1128);
or U1033 (N_1033,In_1515,In_1877);
and U1034 (N_1034,In_1110,In_1388);
and U1035 (N_1035,In_234,In_2299);
nor U1036 (N_1036,In_2382,In_462);
or U1037 (N_1037,In_1150,In_960);
and U1038 (N_1038,In_1384,In_1766);
or U1039 (N_1039,In_2022,In_839);
nor U1040 (N_1040,In_1438,In_2454);
nand U1041 (N_1041,In_1219,In_668);
nor U1042 (N_1042,In_1435,In_356);
xor U1043 (N_1043,In_1701,In_2196);
and U1044 (N_1044,In_2101,In_125);
nand U1045 (N_1045,In_1691,In_1928);
or U1046 (N_1046,In_1331,In_1853);
nand U1047 (N_1047,In_1628,In_405);
nand U1048 (N_1048,In_1463,In_325);
nor U1049 (N_1049,In_411,In_579);
and U1050 (N_1050,In_1961,In_300);
nor U1051 (N_1051,In_1994,In_1122);
or U1052 (N_1052,In_1523,In_2008);
xor U1053 (N_1053,In_1582,In_1009);
nor U1054 (N_1054,In_886,In_2069);
or U1055 (N_1055,In_1888,In_1864);
xnor U1056 (N_1056,In_223,In_66);
nor U1057 (N_1057,In_1703,In_2411);
and U1058 (N_1058,In_91,In_469);
nand U1059 (N_1059,In_560,In_1591);
nand U1060 (N_1060,In_2158,In_2028);
or U1061 (N_1061,In_957,In_928);
nand U1062 (N_1062,In_1124,In_2216);
or U1063 (N_1063,In_756,In_2459);
or U1064 (N_1064,In_661,In_1623);
nor U1065 (N_1065,In_1003,In_786);
xor U1066 (N_1066,In_377,In_88);
nand U1067 (N_1067,In_1908,In_448);
or U1068 (N_1068,In_654,In_1552);
and U1069 (N_1069,In_1513,In_1579);
and U1070 (N_1070,In_1346,In_550);
xnor U1071 (N_1071,In_524,In_995);
xor U1072 (N_1072,In_1984,In_1166);
nor U1073 (N_1073,In_1185,In_1397);
nor U1074 (N_1074,In_2389,In_874);
and U1075 (N_1075,In_2233,In_1076);
xor U1076 (N_1076,In_1955,In_1509);
or U1077 (N_1077,In_176,In_71);
xnor U1078 (N_1078,In_864,In_1247);
or U1079 (N_1079,In_206,In_248);
or U1080 (N_1080,In_61,In_449);
xnor U1081 (N_1081,In_1878,In_1996);
nand U1082 (N_1082,In_329,In_1097);
xor U1083 (N_1083,In_427,In_2330);
or U1084 (N_1084,In_1027,In_1747);
nor U1085 (N_1085,In_1213,In_1708);
and U1086 (N_1086,In_518,In_1642);
nand U1087 (N_1087,In_859,In_1980);
or U1088 (N_1088,In_2471,In_813);
or U1089 (N_1089,In_1372,In_821);
or U1090 (N_1090,In_2447,In_565);
and U1091 (N_1091,In_1390,In_658);
nor U1092 (N_1092,In_680,In_2266);
and U1093 (N_1093,In_1560,In_1807);
xor U1094 (N_1094,In_1954,In_1755);
and U1095 (N_1095,In_1977,In_1880);
nand U1096 (N_1096,In_2088,In_261);
or U1097 (N_1097,In_2138,In_501);
nand U1098 (N_1098,In_846,In_2141);
xor U1099 (N_1099,In_1225,In_34);
nand U1100 (N_1100,In_1183,In_542);
nor U1101 (N_1101,In_1760,In_2112);
or U1102 (N_1102,In_1298,In_2392);
or U1103 (N_1103,In_2124,In_1718);
nand U1104 (N_1104,In_2340,In_2215);
nor U1105 (N_1105,In_1940,In_541);
nand U1106 (N_1106,In_2174,In_1831);
xnor U1107 (N_1107,In_2284,In_236);
nand U1108 (N_1108,In_1887,In_2496);
nand U1109 (N_1109,In_2073,In_332);
and U1110 (N_1110,In_1547,In_1995);
xnor U1111 (N_1111,In_1517,In_343);
nor U1112 (N_1112,In_1414,In_1605);
or U1113 (N_1113,In_636,In_1657);
or U1114 (N_1114,In_1771,In_2403);
nand U1115 (N_1115,In_1680,In_710);
nor U1116 (N_1116,In_1630,In_197);
and U1117 (N_1117,In_1197,In_1060);
nor U1118 (N_1118,In_38,In_1020);
nor U1119 (N_1119,In_1383,In_1178);
xor U1120 (N_1120,In_856,In_2282);
and U1121 (N_1121,In_1683,In_1587);
nor U1122 (N_1122,In_681,In_731);
and U1123 (N_1123,In_2081,In_1810);
nand U1124 (N_1124,In_1171,In_868);
or U1125 (N_1125,In_2393,In_2038);
nor U1126 (N_1126,In_2099,In_148);
or U1127 (N_1127,In_712,In_1078);
or U1128 (N_1128,In_358,In_1829);
or U1129 (N_1129,In_1893,In_1373);
nand U1130 (N_1130,In_1356,In_174);
xor U1131 (N_1131,In_2180,In_456);
nor U1132 (N_1132,In_2234,In_1969);
or U1133 (N_1133,In_1793,In_1296);
or U1134 (N_1134,In_1191,In_1485);
nor U1135 (N_1135,In_1803,In_284);
nand U1136 (N_1136,In_2415,In_2041);
and U1137 (N_1137,In_115,In_2277);
or U1138 (N_1138,In_776,In_1224);
or U1139 (N_1139,In_1813,In_1499);
and U1140 (N_1140,In_679,In_299);
or U1141 (N_1141,In_1454,In_1424);
nor U1142 (N_1142,In_1501,In_1072);
and U1143 (N_1143,In_2376,In_2190);
nand U1144 (N_1144,In_836,In_1821);
and U1145 (N_1145,In_2130,In_1462);
nand U1146 (N_1146,In_847,In_2203);
nor U1147 (N_1147,In_1805,In_790);
or U1148 (N_1148,In_103,In_245);
nor U1149 (N_1149,In_421,In_2358);
and U1150 (N_1150,In_179,In_318);
nor U1151 (N_1151,In_885,In_1843);
nand U1152 (N_1152,In_81,In_117);
and U1153 (N_1153,In_1162,In_1204);
nor U1154 (N_1154,In_2461,In_624);
nor U1155 (N_1155,In_175,In_633);
nand U1156 (N_1156,In_532,In_406);
and U1157 (N_1157,In_79,In_2320);
and U1158 (N_1158,In_1613,In_1208);
nor U1159 (N_1159,In_2366,In_116);
nor U1160 (N_1160,In_43,In_686);
or U1161 (N_1161,In_277,In_818);
or U1162 (N_1162,In_1101,In_2279);
nand U1163 (N_1163,In_826,In_323);
and U1164 (N_1164,In_295,In_1757);
and U1165 (N_1165,In_1040,In_671);
or U1166 (N_1166,In_2119,In_713);
nor U1167 (N_1167,In_1770,In_2400);
or U1168 (N_1168,In_2243,In_498);
or U1169 (N_1169,In_962,In_2093);
or U1170 (N_1170,In_1595,In_1271);
xor U1171 (N_1171,In_256,In_454);
nand U1172 (N_1172,In_660,In_2489);
nand U1173 (N_1173,In_1647,In_855);
nand U1174 (N_1174,In_2308,In_1260);
nand U1175 (N_1175,In_513,In_1531);
nand U1176 (N_1176,In_1186,In_2274);
nor U1177 (N_1177,In_384,In_490);
nor U1178 (N_1178,In_304,In_1572);
nor U1179 (N_1179,In_1059,In_86);
nand U1180 (N_1180,In_540,In_1907);
or U1181 (N_1181,In_554,In_644);
or U1182 (N_1182,In_2135,In_1369);
or U1183 (N_1183,In_1890,In_77);
nand U1184 (N_1184,In_2451,In_51);
or U1185 (N_1185,In_1751,In_956);
nand U1186 (N_1186,In_1168,In_2326);
or U1187 (N_1187,In_1655,In_625);
nor U1188 (N_1188,In_2370,In_1956);
and U1189 (N_1189,In_136,In_2183);
xor U1190 (N_1190,In_339,In_683);
nor U1191 (N_1191,In_1321,In_2089);
nand U1192 (N_1192,In_1348,In_1715);
and U1193 (N_1193,In_1255,In_808);
and U1194 (N_1194,In_979,In_475);
nor U1195 (N_1195,In_2143,In_2467);
or U1196 (N_1196,In_2375,In_1267);
xor U1197 (N_1197,In_506,In_2413);
or U1198 (N_1198,In_630,In_1814);
xor U1199 (N_1199,In_146,In_1936);
and U1200 (N_1200,In_888,In_993);
nor U1201 (N_1201,In_1092,In_2025);
and U1202 (N_1202,In_2488,In_398);
nor U1203 (N_1203,In_1707,In_1677);
nand U1204 (N_1204,In_881,In_1945);
nand U1205 (N_1205,In_1401,In_1470);
and U1206 (N_1206,In_1960,In_1672);
nand U1207 (N_1207,In_267,In_1114);
or U1208 (N_1208,In_548,In_351);
nand U1209 (N_1209,In_1892,In_964);
nand U1210 (N_1210,In_250,In_2316);
nor U1211 (N_1211,In_2232,In_2032);
or U1212 (N_1212,In_1449,In_718);
or U1213 (N_1213,In_1758,In_2302);
and U1214 (N_1214,In_2275,In_944);
or U1215 (N_1215,In_1526,In_155);
and U1216 (N_1216,In_2078,In_330);
xnor U1217 (N_1217,In_210,In_1550);
nand U1218 (N_1218,In_2468,In_1608);
or U1219 (N_1219,In_832,In_1382);
nand U1220 (N_1220,In_1148,In_576);
or U1221 (N_1221,In_1732,In_2120);
nor U1222 (N_1222,In_1086,In_1530);
or U1223 (N_1223,In_1257,In_2357);
nand U1224 (N_1224,In_1202,In_2350);
nand U1225 (N_1225,In_1684,In_2438);
and U1226 (N_1226,In_803,In_752);
nand U1227 (N_1227,In_2100,In_567);
and U1228 (N_1228,In_237,In_841);
or U1229 (N_1229,In_2222,In_1381);
or U1230 (N_1230,In_2306,In_968);
or U1231 (N_1231,In_1361,In_1932);
nor U1232 (N_1232,In_652,In_447);
nor U1233 (N_1233,In_991,In_1350);
or U1234 (N_1234,In_2406,In_659);
nand U1235 (N_1235,In_182,In_488);
and U1236 (N_1236,In_1479,In_70);
and U1237 (N_1237,In_2242,In_2241);
xor U1238 (N_1238,In_1359,In_55);
and U1239 (N_1239,In_1921,In_2123);
and U1240 (N_1240,In_205,In_374);
or U1241 (N_1241,In_1154,In_869);
nor U1242 (N_1242,In_319,In_1494);
or U1243 (N_1243,In_53,In_1048);
nor U1244 (N_1244,In_185,In_1472);
or U1245 (N_1245,In_564,In_666);
or U1246 (N_1246,In_2380,In_2449);
nand U1247 (N_1247,In_2198,In_1416);
or U1248 (N_1248,In_890,In_741);
nand U1249 (N_1249,In_1235,In_640);
nor U1250 (N_1250,In_1580,In_2128);
nand U1251 (N_1251,In_809,In_639);
xor U1252 (N_1252,In_965,In_1628);
nor U1253 (N_1253,In_251,In_1459);
nor U1254 (N_1254,In_2206,In_925);
or U1255 (N_1255,In_882,In_668);
or U1256 (N_1256,In_533,In_1836);
xor U1257 (N_1257,In_556,In_956);
and U1258 (N_1258,In_1836,In_2187);
and U1259 (N_1259,In_2010,In_586);
or U1260 (N_1260,In_271,In_446);
or U1261 (N_1261,In_1753,In_1729);
or U1262 (N_1262,In_535,In_684);
and U1263 (N_1263,In_2047,In_97);
and U1264 (N_1264,In_974,In_571);
xor U1265 (N_1265,In_2416,In_46);
xnor U1266 (N_1266,In_1048,In_946);
nor U1267 (N_1267,In_1401,In_620);
and U1268 (N_1268,In_1530,In_347);
nand U1269 (N_1269,In_2183,In_1092);
nand U1270 (N_1270,In_891,In_482);
nor U1271 (N_1271,In_485,In_1632);
and U1272 (N_1272,In_2478,In_146);
and U1273 (N_1273,In_2242,In_93);
nand U1274 (N_1274,In_1200,In_1221);
and U1275 (N_1275,In_636,In_1877);
and U1276 (N_1276,In_1726,In_2476);
or U1277 (N_1277,In_324,In_148);
nor U1278 (N_1278,In_1983,In_2460);
nor U1279 (N_1279,In_53,In_687);
nand U1280 (N_1280,In_2222,In_2393);
and U1281 (N_1281,In_570,In_479);
or U1282 (N_1282,In_840,In_2125);
xor U1283 (N_1283,In_1647,In_1869);
or U1284 (N_1284,In_299,In_891);
nor U1285 (N_1285,In_1560,In_829);
nand U1286 (N_1286,In_2128,In_2456);
or U1287 (N_1287,In_39,In_684);
and U1288 (N_1288,In_1355,In_2225);
or U1289 (N_1289,In_939,In_2324);
or U1290 (N_1290,In_2462,In_2206);
nand U1291 (N_1291,In_1993,In_1048);
and U1292 (N_1292,In_2409,In_853);
or U1293 (N_1293,In_2039,In_2331);
and U1294 (N_1294,In_1687,In_702);
xnor U1295 (N_1295,In_586,In_907);
or U1296 (N_1296,In_2155,In_2279);
and U1297 (N_1297,In_1940,In_1402);
xnor U1298 (N_1298,In_1148,In_1910);
and U1299 (N_1299,In_2240,In_1978);
and U1300 (N_1300,In_2460,In_1952);
nand U1301 (N_1301,In_83,In_942);
or U1302 (N_1302,In_2423,In_1879);
nand U1303 (N_1303,In_1300,In_2152);
or U1304 (N_1304,In_800,In_1381);
or U1305 (N_1305,In_938,In_2365);
and U1306 (N_1306,In_675,In_60);
and U1307 (N_1307,In_1199,In_1512);
nand U1308 (N_1308,In_920,In_2324);
nor U1309 (N_1309,In_2409,In_2255);
nand U1310 (N_1310,In_1591,In_1479);
nor U1311 (N_1311,In_993,In_2073);
and U1312 (N_1312,In_1983,In_588);
or U1313 (N_1313,In_510,In_1618);
xor U1314 (N_1314,In_44,In_1125);
xnor U1315 (N_1315,In_113,In_1096);
nand U1316 (N_1316,In_38,In_2330);
nand U1317 (N_1317,In_767,In_1553);
or U1318 (N_1318,In_1504,In_456);
xnor U1319 (N_1319,In_1664,In_94);
or U1320 (N_1320,In_1548,In_1384);
nor U1321 (N_1321,In_1153,In_1087);
xor U1322 (N_1322,In_176,In_778);
nand U1323 (N_1323,In_1996,In_1004);
and U1324 (N_1324,In_1959,In_1365);
nand U1325 (N_1325,In_1243,In_1327);
nand U1326 (N_1326,In_640,In_664);
nand U1327 (N_1327,In_603,In_529);
and U1328 (N_1328,In_718,In_2473);
or U1329 (N_1329,In_173,In_260);
nand U1330 (N_1330,In_816,In_971);
nor U1331 (N_1331,In_1504,In_70);
nor U1332 (N_1332,In_1518,In_697);
nand U1333 (N_1333,In_399,In_538);
nand U1334 (N_1334,In_1270,In_1487);
or U1335 (N_1335,In_574,In_426);
nor U1336 (N_1336,In_2060,In_400);
nor U1337 (N_1337,In_2330,In_1740);
nand U1338 (N_1338,In_1112,In_1379);
nor U1339 (N_1339,In_898,In_727);
xor U1340 (N_1340,In_1575,In_1814);
or U1341 (N_1341,In_2009,In_1694);
nor U1342 (N_1342,In_535,In_540);
or U1343 (N_1343,In_907,In_2101);
and U1344 (N_1344,In_974,In_90);
nand U1345 (N_1345,In_1497,In_1693);
and U1346 (N_1346,In_1749,In_2021);
nor U1347 (N_1347,In_1335,In_889);
or U1348 (N_1348,In_1396,In_1681);
and U1349 (N_1349,In_589,In_304);
nand U1350 (N_1350,In_1854,In_684);
nand U1351 (N_1351,In_1694,In_1277);
or U1352 (N_1352,In_616,In_2401);
or U1353 (N_1353,In_635,In_1487);
and U1354 (N_1354,In_940,In_709);
nor U1355 (N_1355,In_309,In_1153);
or U1356 (N_1356,In_73,In_1418);
nor U1357 (N_1357,In_82,In_1921);
and U1358 (N_1358,In_1771,In_257);
and U1359 (N_1359,In_565,In_1518);
xor U1360 (N_1360,In_1885,In_735);
nor U1361 (N_1361,In_205,In_2184);
and U1362 (N_1362,In_551,In_92);
and U1363 (N_1363,In_1947,In_1058);
nand U1364 (N_1364,In_188,In_2411);
nand U1365 (N_1365,In_2136,In_214);
nand U1366 (N_1366,In_153,In_1789);
and U1367 (N_1367,In_2224,In_1130);
or U1368 (N_1368,In_1405,In_873);
nand U1369 (N_1369,In_464,In_82);
nor U1370 (N_1370,In_1810,In_2366);
and U1371 (N_1371,In_2366,In_2435);
and U1372 (N_1372,In_2497,In_1643);
xor U1373 (N_1373,In_2061,In_109);
nor U1374 (N_1374,In_1072,In_5);
nor U1375 (N_1375,In_670,In_1288);
or U1376 (N_1376,In_2265,In_1244);
or U1377 (N_1377,In_1687,In_2);
and U1378 (N_1378,In_649,In_1009);
or U1379 (N_1379,In_1038,In_117);
nor U1380 (N_1380,In_1399,In_220);
or U1381 (N_1381,In_2278,In_1789);
nor U1382 (N_1382,In_275,In_2216);
or U1383 (N_1383,In_527,In_428);
and U1384 (N_1384,In_2050,In_627);
or U1385 (N_1385,In_595,In_1411);
xor U1386 (N_1386,In_661,In_2108);
or U1387 (N_1387,In_1287,In_2475);
nor U1388 (N_1388,In_1266,In_1453);
nor U1389 (N_1389,In_153,In_1707);
or U1390 (N_1390,In_752,In_420);
nor U1391 (N_1391,In_1894,In_698);
or U1392 (N_1392,In_1401,In_1879);
nand U1393 (N_1393,In_524,In_1779);
and U1394 (N_1394,In_720,In_2214);
nor U1395 (N_1395,In_1519,In_2382);
nor U1396 (N_1396,In_1841,In_171);
nand U1397 (N_1397,In_312,In_2352);
and U1398 (N_1398,In_1565,In_806);
nand U1399 (N_1399,In_286,In_1013);
or U1400 (N_1400,In_1789,In_886);
and U1401 (N_1401,In_1401,In_1445);
nand U1402 (N_1402,In_2477,In_1647);
nand U1403 (N_1403,In_1124,In_88);
or U1404 (N_1404,In_2088,In_549);
nand U1405 (N_1405,In_744,In_1825);
nand U1406 (N_1406,In_1430,In_1983);
and U1407 (N_1407,In_777,In_1539);
nor U1408 (N_1408,In_538,In_1733);
and U1409 (N_1409,In_578,In_2418);
or U1410 (N_1410,In_2176,In_2279);
nor U1411 (N_1411,In_21,In_1810);
nor U1412 (N_1412,In_1931,In_1603);
nor U1413 (N_1413,In_382,In_2456);
nand U1414 (N_1414,In_503,In_261);
nand U1415 (N_1415,In_269,In_2363);
xor U1416 (N_1416,In_830,In_2458);
nand U1417 (N_1417,In_1024,In_1729);
nand U1418 (N_1418,In_1352,In_427);
and U1419 (N_1419,In_451,In_1159);
and U1420 (N_1420,In_554,In_507);
and U1421 (N_1421,In_896,In_1280);
or U1422 (N_1422,In_581,In_1001);
nand U1423 (N_1423,In_1490,In_1177);
xor U1424 (N_1424,In_1123,In_538);
nand U1425 (N_1425,In_1294,In_727);
nor U1426 (N_1426,In_287,In_77);
nor U1427 (N_1427,In_971,In_2212);
and U1428 (N_1428,In_690,In_1330);
nor U1429 (N_1429,In_1375,In_675);
and U1430 (N_1430,In_2131,In_721);
and U1431 (N_1431,In_1515,In_2098);
nor U1432 (N_1432,In_722,In_975);
nor U1433 (N_1433,In_646,In_1629);
or U1434 (N_1434,In_2014,In_2106);
nand U1435 (N_1435,In_2399,In_2035);
nor U1436 (N_1436,In_825,In_1921);
or U1437 (N_1437,In_1114,In_1615);
and U1438 (N_1438,In_1556,In_276);
xor U1439 (N_1439,In_925,In_1793);
xnor U1440 (N_1440,In_2291,In_319);
nor U1441 (N_1441,In_1016,In_759);
or U1442 (N_1442,In_1,In_2373);
or U1443 (N_1443,In_707,In_525);
nor U1444 (N_1444,In_1996,In_234);
and U1445 (N_1445,In_1096,In_912);
and U1446 (N_1446,In_1523,In_765);
and U1447 (N_1447,In_1456,In_2299);
nand U1448 (N_1448,In_990,In_786);
or U1449 (N_1449,In_1669,In_212);
nand U1450 (N_1450,In_21,In_732);
or U1451 (N_1451,In_1235,In_1265);
and U1452 (N_1452,In_2404,In_913);
or U1453 (N_1453,In_921,In_2395);
nor U1454 (N_1454,In_1018,In_1337);
nor U1455 (N_1455,In_1006,In_1656);
nor U1456 (N_1456,In_605,In_625);
nand U1457 (N_1457,In_802,In_1421);
or U1458 (N_1458,In_492,In_1218);
nand U1459 (N_1459,In_728,In_942);
nand U1460 (N_1460,In_604,In_1367);
or U1461 (N_1461,In_1436,In_1127);
and U1462 (N_1462,In_1516,In_337);
xnor U1463 (N_1463,In_407,In_1961);
or U1464 (N_1464,In_1708,In_991);
nand U1465 (N_1465,In_1092,In_570);
nand U1466 (N_1466,In_388,In_1980);
and U1467 (N_1467,In_2031,In_2223);
nor U1468 (N_1468,In_887,In_1894);
xor U1469 (N_1469,In_2103,In_2340);
or U1470 (N_1470,In_1725,In_1987);
and U1471 (N_1471,In_1015,In_5);
and U1472 (N_1472,In_917,In_1415);
nand U1473 (N_1473,In_1739,In_2267);
and U1474 (N_1474,In_939,In_541);
xor U1475 (N_1475,In_1297,In_2241);
and U1476 (N_1476,In_1575,In_565);
nand U1477 (N_1477,In_1698,In_1014);
nor U1478 (N_1478,In_1656,In_1534);
nor U1479 (N_1479,In_1482,In_322);
xnor U1480 (N_1480,In_1212,In_455);
and U1481 (N_1481,In_639,In_680);
and U1482 (N_1482,In_978,In_2);
and U1483 (N_1483,In_1483,In_771);
or U1484 (N_1484,In_1080,In_1973);
or U1485 (N_1485,In_368,In_1400);
nand U1486 (N_1486,In_1620,In_2230);
and U1487 (N_1487,In_1948,In_1552);
xor U1488 (N_1488,In_429,In_128);
nor U1489 (N_1489,In_138,In_570);
nand U1490 (N_1490,In_2262,In_1420);
xnor U1491 (N_1491,In_326,In_2199);
and U1492 (N_1492,In_1419,In_1319);
or U1493 (N_1493,In_648,In_1907);
or U1494 (N_1494,In_2191,In_536);
nand U1495 (N_1495,In_1936,In_1420);
nand U1496 (N_1496,In_864,In_929);
and U1497 (N_1497,In_194,In_1877);
nand U1498 (N_1498,In_1310,In_1087);
nor U1499 (N_1499,In_398,In_1715);
nor U1500 (N_1500,In_2295,In_1987);
nor U1501 (N_1501,In_569,In_117);
nand U1502 (N_1502,In_303,In_1297);
nand U1503 (N_1503,In_729,In_885);
nand U1504 (N_1504,In_1280,In_1788);
xnor U1505 (N_1505,In_102,In_581);
and U1506 (N_1506,In_652,In_893);
nor U1507 (N_1507,In_812,In_1559);
or U1508 (N_1508,In_758,In_662);
nand U1509 (N_1509,In_887,In_546);
nand U1510 (N_1510,In_1734,In_1514);
xnor U1511 (N_1511,In_460,In_1629);
nand U1512 (N_1512,In_304,In_1702);
nor U1513 (N_1513,In_1382,In_783);
nor U1514 (N_1514,In_847,In_1402);
and U1515 (N_1515,In_1029,In_1980);
or U1516 (N_1516,In_912,In_1348);
and U1517 (N_1517,In_2289,In_328);
nor U1518 (N_1518,In_1674,In_1652);
nor U1519 (N_1519,In_1829,In_1626);
and U1520 (N_1520,In_2420,In_1201);
and U1521 (N_1521,In_2143,In_924);
nand U1522 (N_1522,In_1659,In_628);
or U1523 (N_1523,In_303,In_2320);
nor U1524 (N_1524,In_1632,In_1855);
nand U1525 (N_1525,In_293,In_252);
or U1526 (N_1526,In_226,In_373);
and U1527 (N_1527,In_1645,In_510);
nor U1528 (N_1528,In_294,In_1904);
nor U1529 (N_1529,In_412,In_59);
and U1530 (N_1530,In_2027,In_402);
and U1531 (N_1531,In_1867,In_2080);
nand U1532 (N_1532,In_2045,In_1518);
nand U1533 (N_1533,In_1853,In_1305);
xnor U1534 (N_1534,In_1781,In_229);
nor U1535 (N_1535,In_1943,In_1093);
or U1536 (N_1536,In_2318,In_533);
nor U1537 (N_1537,In_1078,In_52);
nor U1538 (N_1538,In_1874,In_624);
and U1539 (N_1539,In_1564,In_316);
and U1540 (N_1540,In_1758,In_1191);
and U1541 (N_1541,In_544,In_202);
and U1542 (N_1542,In_2324,In_198);
and U1543 (N_1543,In_739,In_2360);
nand U1544 (N_1544,In_723,In_2153);
and U1545 (N_1545,In_1125,In_1652);
xnor U1546 (N_1546,In_326,In_296);
nand U1547 (N_1547,In_439,In_1510);
or U1548 (N_1548,In_2415,In_2056);
and U1549 (N_1549,In_1178,In_2477);
nand U1550 (N_1550,In_915,In_1594);
nor U1551 (N_1551,In_203,In_555);
and U1552 (N_1552,In_551,In_1674);
xnor U1553 (N_1553,In_2248,In_1373);
nand U1554 (N_1554,In_1876,In_1960);
or U1555 (N_1555,In_2060,In_985);
and U1556 (N_1556,In_1230,In_1781);
nand U1557 (N_1557,In_2175,In_2480);
nor U1558 (N_1558,In_2126,In_595);
nand U1559 (N_1559,In_1588,In_465);
nand U1560 (N_1560,In_930,In_1168);
or U1561 (N_1561,In_1749,In_641);
or U1562 (N_1562,In_1225,In_403);
nand U1563 (N_1563,In_1787,In_961);
or U1564 (N_1564,In_1676,In_1019);
xor U1565 (N_1565,In_1071,In_1254);
nor U1566 (N_1566,In_1479,In_2471);
or U1567 (N_1567,In_1451,In_515);
and U1568 (N_1568,In_2018,In_1237);
nor U1569 (N_1569,In_2045,In_1675);
nand U1570 (N_1570,In_2251,In_1667);
and U1571 (N_1571,In_2448,In_2239);
nand U1572 (N_1572,In_6,In_517);
and U1573 (N_1573,In_823,In_480);
nand U1574 (N_1574,In_2090,In_2050);
nand U1575 (N_1575,In_196,In_452);
nor U1576 (N_1576,In_204,In_1456);
nand U1577 (N_1577,In_305,In_1564);
and U1578 (N_1578,In_2347,In_1075);
xnor U1579 (N_1579,In_525,In_259);
xnor U1580 (N_1580,In_2156,In_1447);
xnor U1581 (N_1581,In_97,In_2017);
nor U1582 (N_1582,In_2172,In_1952);
and U1583 (N_1583,In_2067,In_411);
and U1584 (N_1584,In_1669,In_1113);
or U1585 (N_1585,In_317,In_2038);
or U1586 (N_1586,In_677,In_1013);
nor U1587 (N_1587,In_1717,In_2485);
nor U1588 (N_1588,In_389,In_1761);
nor U1589 (N_1589,In_2131,In_2380);
and U1590 (N_1590,In_815,In_1422);
nand U1591 (N_1591,In_744,In_2429);
nor U1592 (N_1592,In_1123,In_2401);
or U1593 (N_1593,In_1894,In_2081);
and U1594 (N_1594,In_2363,In_1041);
nor U1595 (N_1595,In_913,In_1258);
nor U1596 (N_1596,In_276,In_1793);
nor U1597 (N_1597,In_1720,In_1318);
xor U1598 (N_1598,In_634,In_1096);
and U1599 (N_1599,In_507,In_1174);
nor U1600 (N_1600,In_2238,In_2104);
and U1601 (N_1601,In_705,In_1775);
nor U1602 (N_1602,In_2293,In_1884);
and U1603 (N_1603,In_1803,In_2063);
xnor U1604 (N_1604,In_920,In_1109);
nand U1605 (N_1605,In_803,In_2235);
nor U1606 (N_1606,In_1862,In_1432);
xor U1607 (N_1607,In_313,In_487);
or U1608 (N_1608,In_1728,In_1872);
nor U1609 (N_1609,In_721,In_728);
nand U1610 (N_1610,In_26,In_969);
and U1611 (N_1611,In_633,In_2051);
nor U1612 (N_1612,In_1703,In_319);
and U1613 (N_1613,In_402,In_1237);
and U1614 (N_1614,In_2251,In_139);
nand U1615 (N_1615,In_826,In_111);
or U1616 (N_1616,In_1940,In_1757);
nand U1617 (N_1617,In_1921,In_991);
nand U1618 (N_1618,In_1511,In_2447);
and U1619 (N_1619,In_2404,In_2194);
nor U1620 (N_1620,In_1463,In_615);
or U1621 (N_1621,In_1528,In_1857);
nor U1622 (N_1622,In_766,In_733);
and U1623 (N_1623,In_1629,In_2238);
xor U1624 (N_1624,In_949,In_1984);
or U1625 (N_1625,In_90,In_1172);
or U1626 (N_1626,In_714,In_1027);
nor U1627 (N_1627,In_2328,In_1846);
nand U1628 (N_1628,In_2314,In_1919);
or U1629 (N_1629,In_637,In_1620);
and U1630 (N_1630,In_47,In_1547);
nor U1631 (N_1631,In_211,In_16);
or U1632 (N_1632,In_405,In_1146);
nor U1633 (N_1633,In_1138,In_2264);
nor U1634 (N_1634,In_1871,In_1911);
nor U1635 (N_1635,In_655,In_2275);
nor U1636 (N_1636,In_913,In_490);
nand U1637 (N_1637,In_919,In_1447);
nand U1638 (N_1638,In_2013,In_1166);
and U1639 (N_1639,In_464,In_1744);
or U1640 (N_1640,In_787,In_654);
nor U1641 (N_1641,In_2152,In_274);
or U1642 (N_1642,In_1266,In_1579);
or U1643 (N_1643,In_833,In_1376);
nor U1644 (N_1644,In_627,In_1796);
nor U1645 (N_1645,In_72,In_1176);
nor U1646 (N_1646,In_1738,In_1466);
nand U1647 (N_1647,In_212,In_2350);
nor U1648 (N_1648,In_2071,In_2290);
or U1649 (N_1649,In_2026,In_1121);
nand U1650 (N_1650,In_2149,In_1638);
xnor U1651 (N_1651,In_423,In_2264);
xor U1652 (N_1652,In_1809,In_1821);
nor U1653 (N_1653,In_2254,In_2454);
nand U1654 (N_1654,In_548,In_1132);
nand U1655 (N_1655,In_45,In_1334);
xnor U1656 (N_1656,In_265,In_465);
nand U1657 (N_1657,In_1801,In_2201);
nor U1658 (N_1658,In_525,In_1856);
nand U1659 (N_1659,In_1001,In_1271);
or U1660 (N_1660,In_1040,In_500);
or U1661 (N_1661,In_2017,In_682);
or U1662 (N_1662,In_173,In_1699);
nand U1663 (N_1663,In_2234,In_687);
nor U1664 (N_1664,In_731,In_1935);
or U1665 (N_1665,In_2300,In_815);
and U1666 (N_1666,In_1477,In_1804);
xnor U1667 (N_1667,In_1942,In_1883);
nor U1668 (N_1668,In_855,In_2326);
and U1669 (N_1669,In_2488,In_1692);
nand U1670 (N_1670,In_262,In_1322);
and U1671 (N_1671,In_614,In_1472);
and U1672 (N_1672,In_575,In_2010);
and U1673 (N_1673,In_1590,In_1192);
nand U1674 (N_1674,In_1577,In_104);
or U1675 (N_1675,In_85,In_1631);
nor U1676 (N_1676,In_1644,In_560);
or U1677 (N_1677,In_46,In_2151);
and U1678 (N_1678,In_928,In_1792);
and U1679 (N_1679,In_201,In_233);
nand U1680 (N_1680,In_991,In_2137);
and U1681 (N_1681,In_1922,In_2183);
or U1682 (N_1682,In_1469,In_257);
or U1683 (N_1683,In_1550,In_2393);
or U1684 (N_1684,In_1067,In_2401);
nor U1685 (N_1685,In_2288,In_49);
xor U1686 (N_1686,In_1319,In_2212);
xnor U1687 (N_1687,In_117,In_39);
nand U1688 (N_1688,In_475,In_980);
and U1689 (N_1689,In_1450,In_1743);
nor U1690 (N_1690,In_1425,In_2249);
nor U1691 (N_1691,In_955,In_896);
nor U1692 (N_1692,In_1922,In_1410);
or U1693 (N_1693,In_1793,In_511);
nor U1694 (N_1694,In_985,In_1767);
nor U1695 (N_1695,In_327,In_1552);
nand U1696 (N_1696,In_1517,In_425);
nand U1697 (N_1697,In_250,In_1650);
nand U1698 (N_1698,In_1450,In_747);
and U1699 (N_1699,In_711,In_409);
or U1700 (N_1700,In_235,In_1441);
nand U1701 (N_1701,In_1264,In_1022);
and U1702 (N_1702,In_665,In_1696);
nor U1703 (N_1703,In_1309,In_1690);
xnor U1704 (N_1704,In_1478,In_1404);
nor U1705 (N_1705,In_2386,In_325);
and U1706 (N_1706,In_1183,In_612);
xor U1707 (N_1707,In_608,In_688);
nor U1708 (N_1708,In_926,In_1643);
nor U1709 (N_1709,In_320,In_389);
nand U1710 (N_1710,In_1325,In_773);
and U1711 (N_1711,In_1088,In_104);
nor U1712 (N_1712,In_2041,In_1689);
and U1713 (N_1713,In_2473,In_1787);
nand U1714 (N_1714,In_2149,In_1781);
and U1715 (N_1715,In_1055,In_279);
xnor U1716 (N_1716,In_325,In_922);
xor U1717 (N_1717,In_1382,In_2272);
or U1718 (N_1718,In_1333,In_801);
nor U1719 (N_1719,In_2226,In_2397);
xnor U1720 (N_1720,In_1292,In_519);
and U1721 (N_1721,In_1165,In_2057);
nand U1722 (N_1722,In_2168,In_2351);
xor U1723 (N_1723,In_1423,In_2384);
xor U1724 (N_1724,In_2172,In_1521);
xor U1725 (N_1725,In_1975,In_714);
nor U1726 (N_1726,In_188,In_2370);
nor U1727 (N_1727,In_2206,In_787);
and U1728 (N_1728,In_2447,In_2407);
nor U1729 (N_1729,In_1054,In_1318);
or U1730 (N_1730,In_517,In_1562);
and U1731 (N_1731,In_1116,In_475);
and U1732 (N_1732,In_794,In_1695);
nor U1733 (N_1733,In_2094,In_1736);
nor U1734 (N_1734,In_709,In_1489);
nand U1735 (N_1735,In_666,In_623);
nor U1736 (N_1736,In_794,In_1413);
nor U1737 (N_1737,In_1331,In_841);
and U1738 (N_1738,In_2456,In_1081);
and U1739 (N_1739,In_1829,In_1666);
nand U1740 (N_1740,In_349,In_2209);
or U1741 (N_1741,In_1688,In_646);
nor U1742 (N_1742,In_1659,In_1641);
or U1743 (N_1743,In_350,In_245);
nor U1744 (N_1744,In_1763,In_1384);
nand U1745 (N_1745,In_907,In_1331);
and U1746 (N_1746,In_1332,In_1337);
nand U1747 (N_1747,In_1511,In_810);
or U1748 (N_1748,In_1367,In_2209);
or U1749 (N_1749,In_1748,In_1094);
nand U1750 (N_1750,In_1678,In_708);
nor U1751 (N_1751,In_2347,In_1354);
and U1752 (N_1752,In_2315,In_354);
or U1753 (N_1753,In_2180,In_549);
xnor U1754 (N_1754,In_1265,In_1748);
nor U1755 (N_1755,In_2415,In_1447);
nand U1756 (N_1756,In_1000,In_104);
and U1757 (N_1757,In_436,In_1891);
nand U1758 (N_1758,In_1719,In_194);
and U1759 (N_1759,In_287,In_1720);
nand U1760 (N_1760,In_1302,In_2060);
and U1761 (N_1761,In_1309,In_1298);
or U1762 (N_1762,In_1793,In_1858);
and U1763 (N_1763,In_1116,In_1000);
xor U1764 (N_1764,In_566,In_1954);
xnor U1765 (N_1765,In_492,In_1534);
or U1766 (N_1766,In_1489,In_2);
nand U1767 (N_1767,In_662,In_2299);
nor U1768 (N_1768,In_394,In_1936);
nand U1769 (N_1769,In_106,In_1664);
nand U1770 (N_1770,In_2249,In_99);
and U1771 (N_1771,In_2313,In_2409);
xnor U1772 (N_1772,In_1292,In_1740);
nor U1773 (N_1773,In_148,In_83);
nor U1774 (N_1774,In_1518,In_2405);
xnor U1775 (N_1775,In_289,In_1420);
xor U1776 (N_1776,In_527,In_1211);
nand U1777 (N_1777,In_374,In_1655);
or U1778 (N_1778,In_1524,In_1822);
xnor U1779 (N_1779,In_587,In_719);
and U1780 (N_1780,In_1072,In_2084);
or U1781 (N_1781,In_176,In_167);
or U1782 (N_1782,In_237,In_199);
nor U1783 (N_1783,In_82,In_1017);
nor U1784 (N_1784,In_754,In_442);
nand U1785 (N_1785,In_603,In_1009);
nand U1786 (N_1786,In_1946,In_2495);
or U1787 (N_1787,In_679,In_1559);
nand U1788 (N_1788,In_2344,In_272);
or U1789 (N_1789,In_243,In_795);
nor U1790 (N_1790,In_327,In_1650);
and U1791 (N_1791,In_1106,In_394);
nand U1792 (N_1792,In_2240,In_778);
nor U1793 (N_1793,In_460,In_903);
and U1794 (N_1794,In_152,In_898);
nor U1795 (N_1795,In_212,In_198);
and U1796 (N_1796,In_1672,In_1642);
or U1797 (N_1797,In_810,In_1623);
or U1798 (N_1798,In_1447,In_1304);
nor U1799 (N_1799,In_500,In_1532);
nand U1800 (N_1800,In_2075,In_500);
xnor U1801 (N_1801,In_895,In_1153);
or U1802 (N_1802,In_72,In_420);
nand U1803 (N_1803,In_649,In_195);
and U1804 (N_1804,In_2407,In_1183);
nor U1805 (N_1805,In_947,In_2152);
and U1806 (N_1806,In_2467,In_603);
and U1807 (N_1807,In_477,In_49);
nand U1808 (N_1808,In_971,In_2053);
nand U1809 (N_1809,In_117,In_1205);
nor U1810 (N_1810,In_530,In_2496);
or U1811 (N_1811,In_1746,In_1686);
and U1812 (N_1812,In_2158,In_1151);
and U1813 (N_1813,In_2007,In_1948);
or U1814 (N_1814,In_1245,In_866);
nand U1815 (N_1815,In_845,In_350);
nor U1816 (N_1816,In_2047,In_1252);
nor U1817 (N_1817,In_2440,In_1373);
and U1818 (N_1818,In_2156,In_1042);
or U1819 (N_1819,In_1690,In_2067);
or U1820 (N_1820,In_976,In_1687);
nor U1821 (N_1821,In_510,In_1609);
nor U1822 (N_1822,In_1304,In_309);
or U1823 (N_1823,In_1265,In_753);
nor U1824 (N_1824,In_2478,In_1579);
nor U1825 (N_1825,In_1646,In_1831);
and U1826 (N_1826,In_1092,In_2478);
and U1827 (N_1827,In_1419,In_2147);
nor U1828 (N_1828,In_1180,In_2244);
nor U1829 (N_1829,In_2291,In_1615);
or U1830 (N_1830,In_612,In_1844);
nand U1831 (N_1831,In_1095,In_306);
nor U1832 (N_1832,In_1455,In_240);
and U1833 (N_1833,In_220,In_369);
and U1834 (N_1834,In_1355,In_1207);
xnor U1835 (N_1835,In_1959,In_1657);
nand U1836 (N_1836,In_967,In_552);
nand U1837 (N_1837,In_1352,In_1704);
nor U1838 (N_1838,In_540,In_1210);
xor U1839 (N_1839,In_1108,In_2434);
nand U1840 (N_1840,In_33,In_1592);
nand U1841 (N_1841,In_2415,In_407);
or U1842 (N_1842,In_13,In_2338);
and U1843 (N_1843,In_281,In_879);
xnor U1844 (N_1844,In_1732,In_1543);
nand U1845 (N_1845,In_339,In_1814);
nand U1846 (N_1846,In_1539,In_2180);
nand U1847 (N_1847,In_1568,In_1793);
xnor U1848 (N_1848,In_587,In_2289);
or U1849 (N_1849,In_1195,In_1754);
nor U1850 (N_1850,In_1835,In_1688);
or U1851 (N_1851,In_641,In_997);
nor U1852 (N_1852,In_2403,In_1405);
xnor U1853 (N_1853,In_2316,In_2025);
or U1854 (N_1854,In_905,In_644);
and U1855 (N_1855,In_1382,In_2304);
nor U1856 (N_1856,In_1436,In_308);
nor U1857 (N_1857,In_577,In_1724);
or U1858 (N_1858,In_275,In_604);
nand U1859 (N_1859,In_312,In_684);
or U1860 (N_1860,In_2073,In_351);
xnor U1861 (N_1861,In_1428,In_1774);
and U1862 (N_1862,In_1040,In_1772);
nand U1863 (N_1863,In_1432,In_2012);
nand U1864 (N_1864,In_530,In_330);
and U1865 (N_1865,In_143,In_812);
xor U1866 (N_1866,In_2311,In_749);
and U1867 (N_1867,In_854,In_2011);
nand U1868 (N_1868,In_513,In_1122);
and U1869 (N_1869,In_632,In_64);
nor U1870 (N_1870,In_2434,In_2344);
xor U1871 (N_1871,In_244,In_192);
or U1872 (N_1872,In_536,In_222);
nand U1873 (N_1873,In_1136,In_1297);
and U1874 (N_1874,In_1672,In_2375);
nand U1875 (N_1875,In_1,In_922);
nand U1876 (N_1876,In_1325,In_572);
and U1877 (N_1877,In_58,In_193);
xnor U1878 (N_1878,In_1462,In_2380);
nor U1879 (N_1879,In_2202,In_634);
or U1880 (N_1880,In_1993,In_1223);
xor U1881 (N_1881,In_802,In_425);
xnor U1882 (N_1882,In_244,In_2222);
nor U1883 (N_1883,In_915,In_58);
and U1884 (N_1884,In_947,In_2382);
and U1885 (N_1885,In_727,In_2112);
nor U1886 (N_1886,In_2213,In_723);
nor U1887 (N_1887,In_113,In_1832);
or U1888 (N_1888,In_1148,In_244);
and U1889 (N_1889,In_598,In_661);
or U1890 (N_1890,In_1487,In_2305);
nand U1891 (N_1891,In_2263,In_489);
nor U1892 (N_1892,In_1085,In_1811);
or U1893 (N_1893,In_498,In_914);
and U1894 (N_1894,In_1382,In_314);
nand U1895 (N_1895,In_525,In_428);
or U1896 (N_1896,In_760,In_408);
xnor U1897 (N_1897,In_296,In_2369);
and U1898 (N_1898,In_541,In_1596);
or U1899 (N_1899,In_983,In_252);
nand U1900 (N_1900,In_2337,In_183);
nand U1901 (N_1901,In_19,In_918);
nor U1902 (N_1902,In_1514,In_1827);
xor U1903 (N_1903,In_1560,In_1995);
or U1904 (N_1904,In_1607,In_72);
or U1905 (N_1905,In_1161,In_2405);
nor U1906 (N_1906,In_631,In_1841);
and U1907 (N_1907,In_453,In_414);
nand U1908 (N_1908,In_2025,In_346);
nor U1909 (N_1909,In_1567,In_2114);
xnor U1910 (N_1910,In_2441,In_922);
and U1911 (N_1911,In_1051,In_2401);
or U1912 (N_1912,In_685,In_495);
nor U1913 (N_1913,In_2167,In_425);
or U1914 (N_1914,In_920,In_622);
nor U1915 (N_1915,In_829,In_2158);
or U1916 (N_1916,In_1222,In_865);
or U1917 (N_1917,In_2214,In_1823);
or U1918 (N_1918,In_243,In_59);
and U1919 (N_1919,In_985,In_2394);
xnor U1920 (N_1920,In_1851,In_2367);
nor U1921 (N_1921,In_1483,In_1264);
or U1922 (N_1922,In_1882,In_824);
and U1923 (N_1923,In_2076,In_1695);
nand U1924 (N_1924,In_2465,In_390);
nand U1925 (N_1925,In_1871,In_2011);
nand U1926 (N_1926,In_2221,In_500);
or U1927 (N_1927,In_773,In_2112);
and U1928 (N_1928,In_2133,In_1959);
and U1929 (N_1929,In_1674,In_462);
and U1930 (N_1930,In_173,In_782);
or U1931 (N_1931,In_842,In_2163);
and U1932 (N_1932,In_708,In_2453);
or U1933 (N_1933,In_2066,In_2009);
nand U1934 (N_1934,In_2144,In_2329);
and U1935 (N_1935,In_2297,In_2036);
or U1936 (N_1936,In_850,In_1821);
and U1937 (N_1937,In_2400,In_2413);
and U1938 (N_1938,In_1632,In_1198);
nand U1939 (N_1939,In_1869,In_470);
and U1940 (N_1940,In_806,In_801);
xor U1941 (N_1941,In_1298,In_2425);
and U1942 (N_1942,In_559,In_49);
nand U1943 (N_1943,In_646,In_458);
and U1944 (N_1944,In_918,In_2132);
xor U1945 (N_1945,In_1382,In_1282);
and U1946 (N_1946,In_1770,In_1746);
and U1947 (N_1947,In_2109,In_1169);
nor U1948 (N_1948,In_2276,In_772);
nand U1949 (N_1949,In_1276,In_2102);
nand U1950 (N_1950,In_1669,In_217);
and U1951 (N_1951,In_1848,In_1025);
or U1952 (N_1952,In_647,In_849);
and U1953 (N_1953,In_944,In_285);
nor U1954 (N_1954,In_1650,In_2324);
nor U1955 (N_1955,In_2382,In_2267);
or U1956 (N_1956,In_2132,In_2407);
and U1957 (N_1957,In_153,In_2387);
nand U1958 (N_1958,In_1156,In_1441);
nand U1959 (N_1959,In_384,In_243);
nand U1960 (N_1960,In_44,In_641);
or U1961 (N_1961,In_406,In_101);
or U1962 (N_1962,In_1971,In_811);
and U1963 (N_1963,In_1380,In_2311);
and U1964 (N_1964,In_771,In_1003);
and U1965 (N_1965,In_376,In_746);
or U1966 (N_1966,In_661,In_1055);
or U1967 (N_1967,In_1320,In_1886);
nand U1968 (N_1968,In_1889,In_1785);
and U1969 (N_1969,In_976,In_2337);
xor U1970 (N_1970,In_1915,In_159);
nor U1971 (N_1971,In_43,In_898);
and U1972 (N_1972,In_325,In_761);
nand U1973 (N_1973,In_517,In_2348);
xor U1974 (N_1974,In_65,In_1125);
nor U1975 (N_1975,In_1312,In_2484);
nand U1976 (N_1976,In_2350,In_1068);
nand U1977 (N_1977,In_2220,In_1642);
nand U1978 (N_1978,In_409,In_1578);
or U1979 (N_1979,In_1315,In_1732);
nand U1980 (N_1980,In_265,In_663);
or U1981 (N_1981,In_1689,In_1745);
xor U1982 (N_1982,In_2072,In_1481);
and U1983 (N_1983,In_1205,In_93);
nand U1984 (N_1984,In_1409,In_1923);
nor U1985 (N_1985,In_163,In_250);
and U1986 (N_1986,In_1886,In_383);
nor U1987 (N_1987,In_771,In_1283);
nand U1988 (N_1988,In_1905,In_1115);
xnor U1989 (N_1989,In_149,In_843);
or U1990 (N_1990,In_1850,In_867);
nand U1991 (N_1991,In_1910,In_1827);
nand U1992 (N_1992,In_1608,In_590);
or U1993 (N_1993,In_2345,In_430);
or U1994 (N_1994,In_1512,In_808);
nand U1995 (N_1995,In_1773,In_891);
nand U1996 (N_1996,In_657,In_1462);
or U1997 (N_1997,In_2060,In_1053);
nor U1998 (N_1998,In_528,In_2326);
nand U1999 (N_1999,In_439,In_966);
and U2000 (N_2000,In_1916,In_1530);
and U2001 (N_2001,In_584,In_99);
and U2002 (N_2002,In_1735,In_149);
xor U2003 (N_2003,In_584,In_338);
nor U2004 (N_2004,In_723,In_1382);
nor U2005 (N_2005,In_1931,In_1066);
nand U2006 (N_2006,In_926,In_325);
or U2007 (N_2007,In_1554,In_813);
nor U2008 (N_2008,In_2088,In_917);
and U2009 (N_2009,In_448,In_1330);
nor U2010 (N_2010,In_2314,In_1071);
and U2011 (N_2011,In_1930,In_576);
nand U2012 (N_2012,In_174,In_81);
nand U2013 (N_2013,In_1981,In_858);
xor U2014 (N_2014,In_2139,In_2307);
or U2015 (N_2015,In_426,In_1623);
nor U2016 (N_2016,In_1765,In_1444);
nor U2017 (N_2017,In_26,In_1586);
nor U2018 (N_2018,In_1549,In_345);
and U2019 (N_2019,In_2036,In_767);
and U2020 (N_2020,In_927,In_1958);
nor U2021 (N_2021,In_1418,In_863);
and U2022 (N_2022,In_1114,In_1904);
and U2023 (N_2023,In_2428,In_2287);
nor U2024 (N_2024,In_421,In_2277);
or U2025 (N_2025,In_2419,In_253);
xor U2026 (N_2026,In_2436,In_1605);
and U2027 (N_2027,In_1065,In_478);
or U2028 (N_2028,In_1477,In_505);
and U2029 (N_2029,In_2450,In_1550);
nor U2030 (N_2030,In_1703,In_818);
xnor U2031 (N_2031,In_1266,In_1165);
nand U2032 (N_2032,In_1128,In_527);
or U2033 (N_2033,In_518,In_2222);
or U2034 (N_2034,In_2215,In_2029);
or U2035 (N_2035,In_694,In_2363);
and U2036 (N_2036,In_2271,In_677);
nand U2037 (N_2037,In_1523,In_625);
and U2038 (N_2038,In_466,In_1367);
and U2039 (N_2039,In_1133,In_220);
nor U2040 (N_2040,In_313,In_279);
and U2041 (N_2041,In_245,In_2111);
or U2042 (N_2042,In_1993,In_1363);
or U2043 (N_2043,In_566,In_2259);
nand U2044 (N_2044,In_886,In_906);
or U2045 (N_2045,In_211,In_853);
and U2046 (N_2046,In_399,In_1684);
nor U2047 (N_2047,In_2345,In_944);
nor U2048 (N_2048,In_1546,In_2006);
and U2049 (N_2049,In_302,In_1001);
xor U2050 (N_2050,In_1065,In_1792);
and U2051 (N_2051,In_2034,In_1192);
nor U2052 (N_2052,In_700,In_16);
or U2053 (N_2053,In_22,In_1530);
and U2054 (N_2054,In_389,In_2091);
nand U2055 (N_2055,In_566,In_2439);
nand U2056 (N_2056,In_1059,In_1354);
or U2057 (N_2057,In_284,In_246);
nand U2058 (N_2058,In_2201,In_1352);
nand U2059 (N_2059,In_1909,In_1606);
nand U2060 (N_2060,In_2154,In_1360);
nand U2061 (N_2061,In_1639,In_347);
and U2062 (N_2062,In_1856,In_2015);
or U2063 (N_2063,In_695,In_91);
nor U2064 (N_2064,In_778,In_63);
nand U2065 (N_2065,In_1403,In_1625);
nor U2066 (N_2066,In_2428,In_1668);
or U2067 (N_2067,In_1171,In_1727);
or U2068 (N_2068,In_2177,In_1817);
and U2069 (N_2069,In_85,In_169);
xor U2070 (N_2070,In_269,In_1187);
nor U2071 (N_2071,In_1302,In_562);
and U2072 (N_2072,In_2020,In_588);
or U2073 (N_2073,In_546,In_181);
and U2074 (N_2074,In_2259,In_603);
nand U2075 (N_2075,In_466,In_1441);
nor U2076 (N_2076,In_1002,In_1897);
nand U2077 (N_2077,In_1041,In_1668);
and U2078 (N_2078,In_376,In_1930);
or U2079 (N_2079,In_2465,In_2330);
or U2080 (N_2080,In_85,In_490);
nor U2081 (N_2081,In_868,In_2311);
and U2082 (N_2082,In_2271,In_94);
nand U2083 (N_2083,In_762,In_561);
or U2084 (N_2084,In_1514,In_1794);
or U2085 (N_2085,In_241,In_593);
or U2086 (N_2086,In_2161,In_794);
nand U2087 (N_2087,In_538,In_408);
xnor U2088 (N_2088,In_644,In_407);
nand U2089 (N_2089,In_389,In_1278);
and U2090 (N_2090,In_1117,In_359);
and U2091 (N_2091,In_1055,In_1301);
nand U2092 (N_2092,In_2246,In_698);
nor U2093 (N_2093,In_271,In_40);
nand U2094 (N_2094,In_844,In_1456);
nand U2095 (N_2095,In_1230,In_1086);
xor U2096 (N_2096,In_1842,In_103);
nand U2097 (N_2097,In_2137,In_1351);
or U2098 (N_2098,In_1344,In_516);
nand U2099 (N_2099,In_80,In_2312);
and U2100 (N_2100,In_1089,In_723);
and U2101 (N_2101,In_1110,In_1660);
or U2102 (N_2102,In_1267,In_473);
or U2103 (N_2103,In_504,In_948);
nand U2104 (N_2104,In_1957,In_1471);
nor U2105 (N_2105,In_657,In_1076);
and U2106 (N_2106,In_1678,In_2279);
or U2107 (N_2107,In_1218,In_1461);
or U2108 (N_2108,In_1027,In_2423);
or U2109 (N_2109,In_1800,In_2162);
and U2110 (N_2110,In_457,In_907);
nand U2111 (N_2111,In_2319,In_536);
and U2112 (N_2112,In_939,In_2130);
nor U2113 (N_2113,In_2401,In_1594);
and U2114 (N_2114,In_2112,In_1731);
xnor U2115 (N_2115,In_1135,In_1424);
or U2116 (N_2116,In_947,In_1586);
or U2117 (N_2117,In_1905,In_299);
nand U2118 (N_2118,In_1380,In_809);
and U2119 (N_2119,In_2062,In_369);
xor U2120 (N_2120,In_1647,In_163);
or U2121 (N_2121,In_310,In_1418);
nand U2122 (N_2122,In_482,In_1319);
and U2123 (N_2123,In_745,In_1150);
xor U2124 (N_2124,In_1262,In_473);
nand U2125 (N_2125,In_714,In_864);
nor U2126 (N_2126,In_686,In_948);
nor U2127 (N_2127,In_1237,In_2112);
and U2128 (N_2128,In_2182,In_1903);
or U2129 (N_2129,In_561,In_2360);
nand U2130 (N_2130,In_1455,In_1294);
and U2131 (N_2131,In_1230,In_1025);
nand U2132 (N_2132,In_105,In_2264);
or U2133 (N_2133,In_2177,In_425);
nor U2134 (N_2134,In_612,In_1744);
and U2135 (N_2135,In_115,In_661);
nor U2136 (N_2136,In_437,In_2329);
or U2137 (N_2137,In_2005,In_594);
and U2138 (N_2138,In_545,In_1977);
and U2139 (N_2139,In_1717,In_1252);
xor U2140 (N_2140,In_1344,In_2437);
and U2141 (N_2141,In_31,In_1643);
nand U2142 (N_2142,In_271,In_1421);
or U2143 (N_2143,In_845,In_1742);
and U2144 (N_2144,In_1387,In_1776);
and U2145 (N_2145,In_1380,In_2103);
or U2146 (N_2146,In_355,In_398);
or U2147 (N_2147,In_1429,In_1830);
nand U2148 (N_2148,In_2493,In_1756);
xnor U2149 (N_2149,In_1278,In_717);
nor U2150 (N_2150,In_1984,In_559);
nor U2151 (N_2151,In_699,In_1406);
or U2152 (N_2152,In_961,In_112);
nor U2153 (N_2153,In_1576,In_1986);
or U2154 (N_2154,In_2393,In_170);
nor U2155 (N_2155,In_1981,In_1276);
and U2156 (N_2156,In_1789,In_1396);
nor U2157 (N_2157,In_1255,In_1733);
nor U2158 (N_2158,In_486,In_129);
nand U2159 (N_2159,In_2110,In_237);
xor U2160 (N_2160,In_1443,In_2387);
nand U2161 (N_2161,In_1608,In_1483);
nand U2162 (N_2162,In_990,In_2427);
nor U2163 (N_2163,In_1377,In_314);
nor U2164 (N_2164,In_1963,In_845);
nor U2165 (N_2165,In_1020,In_1206);
nand U2166 (N_2166,In_1739,In_869);
nor U2167 (N_2167,In_536,In_810);
nor U2168 (N_2168,In_551,In_2427);
and U2169 (N_2169,In_1554,In_1071);
nand U2170 (N_2170,In_2492,In_1865);
nand U2171 (N_2171,In_1940,In_1650);
and U2172 (N_2172,In_2416,In_1873);
or U2173 (N_2173,In_2008,In_918);
nor U2174 (N_2174,In_1476,In_1968);
and U2175 (N_2175,In_1056,In_1730);
or U2176 (N_2176,In_697,In_1840);
nand U2177 (N_2177,In_2100,In_1995);
nor U2178 (N_2178,In_2404,In_562);
nand U2179 (N_2179,In_1623,In_605);
xor U2180 (N_2180,In_983,In_2031);
and U2181 (N_2181,In_1099,In_465);
and U2182 (N_2182,In_2450,In_1834);
nand U2183 (N_2183,In_2088,In_1661);
and U2184 (N_2184,In_1101,In_745);
xnor U2185 (N_2185,In_2075,In_1402);
nand U2186 (N_2186,In_1144,In_1550);
or U2187 (N_2187,In_1617,In_781);
or U2188 (N_2188,In_272,In_2299);
or U2189 (N_2189,In_2123,In_901);
or U2190 (N_2190,In_363,In_915);
nor U2191 (N_2191,In_497,In_518);
or U2192 (N_2192,In_652,In_41);
nor U2193 (N_2193,In_1083,In_2203);
and U2194 (N_2194,In_929,In_1671);
nor U2195 (N_2195,In_2194,In_301);
or U2196 (N_2196,In_2081,In_1719);
or U2197 (N_2197,In_1828,In_1621);
nand U2198 (N_2198,In_492,In_1650);
nor U2199 (N_2199,In_1400,In_562);
or U2200 (N_2200,In_320,In_2235);
nor U2201 (N_2201,In_1737,In_441);
or U2202 (N_2202,In_1646,In_2377);
and U2203 (N_2203,In_1805,In_579);
xor U2204 (N_2204,In_1784,In_790);
or U2205 (N_2205,In_399,In_1028);
nor U2206 (N_2206,In_1314,In_274);
or U2207 (N_2207,In_583,In_430);
xor U2208 (N_2208,In_162,In_1457);
and U2209 (N_2209,In_1589,In_1969);
or U2210 (N_2210,In_257,In_2077);
nor U2211 (N_2211,In_623,In_1520);
and U2212 (N_2212,In_1544,In_50);
nor U2213 (N_2213,In_828,In_777);
xnor U2214 (N_2214,In_659,In_2360);
nand U2215 (N_2215,In_1004,In_570);
or U2216 (N_2216,In_2020,In_151);
nor U2217 (N_2217,In_1493,In_86);
or U2218 (N_2218,In_2164,In_419);
nor U2219 (N_2219,In_2276,In_1736);
nand U2220 (N_2220,In_1672,In_2409);
nor U2221 (N_2221,In_2170,In_952);
xor U2222 (N_2222,In_2449,In_2066);
nand U2223 (N_2223,In_1455,In_15);
or U2224 (N_2224,In_1036,In_1234);
nor U2225 (N_2225,In_1166,In_433);
nor U2226 (N_2226,In_2078,In_1026);
nor U2227 (N_2227,In_1917,In_2063);
nor U2228 (N_2228,In_560,In_2131);
xor U2229 (N_2229,In_1,In_2138);
xor U2230 (N_2230,In_450,In_1737);
nand U2231 (N_2231,In_795,In_88);
or U2232 (N_2232,In_909,In_1915);
or U2233 (N_2233,In_1551,In_784);
nand U2234 (N_2234,In_464,In_1606);
xnor U2235 (N_2235,In_723,In_2033);
or U2236 (N_2236,In_1072,In_2474);
nor U2237 (N_2237,In_810,In_585);
nor U2238 (N_2238,In_2238,In_254);
xor U2239 (N_2239,In_2237,In_2214);
nor U2240 (N_2240,In_1306,In_333);
nand U2241 (N_2241,In_1739,In_1149);
nor U2242 (N_2242,In_1498,In_716);
or U2243 (N_2243,In_697,In_245);
or U2244 (N_2244,In_848,In_2024);
and U2245 (N_2245,In_1270,In_2106);
nor U2246 (N_2246,In_365,In_1990);
or U2247 (N_2247,In_534,In_2139);
and U2248 (N_2248,In_1663,In_2144);
nor U2249 (N_2249,In_1148,In_1165);
nor U2250 (N_2250,In_546,In_544);
xor U2251 (N_2251,In_1405,In_2160);
nand U2252 (N_2252,In_174,In_316);
and U2253 (N_2253,In_61,In_2114);
or U2254 (N_2254,In_1947,In_1046);
nor U2255 (N_2255,In_2260,In_1281);
and U2256 (N_2256,In_1220,In_1928);
and U2257 (N_2257,In_1483,In_783);
nor U2258 (N_2258,In_1969,In_1145);
or U2259 (N_2259,In_605,In_1392);
or U2260 (N_2260,In_565,In_628);
nor U2261 (N_2261,In_1191,In_1111);
nand U2262 (N_2262,In_684,In_456);
xor U2263 (N_2263,In_2091,In_194);
nor U2264 (N_2264,In_745,In_2101);
or U2265 (N_2265,In_846,In_658);
nand U2266 (N_2266,In_2457,In_1957);
and U2267 (N_2267,In_212,In_368);
or U2268 (N_2268,In_784,In_1928);
and U2269 (N_2269,In_1328,In_697);
nand U2270 (N_2270,In_529,In_1166);
or U2271 (N_2271,In_1915,In_2355);
xnor U2272 (N_2272,In_2236,In_1729);
nand U2273 (N_2273,In_669,In_472);
or U2274 (N_2274,In_2215,In_136);
or U2275 (N_2275,In_2047,In_1466);
nand U2276 (N_2276,In_1009,In_1811);
and U2277 (N_2277,In_2132,In_45);
or U2278 (N_2278,In_2368,In_721);
or U2279 (N_2279,In_1081,In_1493);
and U2280 (N_2280,In_826,In_2303);
nor U2281 (N_2281,In_95,In_630);
nand U2282 (N_2282,In_2015,In_1392);
and U2283 (N_2283,In_697,In_2492);
and U2284 (N_2284,In_1628,In_2115);
or U2285 (N_2285,In_191,In_575);
xor U2286 (N_2286,In_1744,In_1010);
nor U2287 (N_2287,In_1528,In_2251);
nand U2288 (N_2288,In_646,In_1393);
nor U2289 (N_2289,In_342,In_1795);
nor U2290 (N_2290,In_850,In_699);
xnor U2291 (N_2291,In_1762,In_133);
nor U2292 (N_2292,In_392,In_232);
and U2293 (N_2293,In_972,In_834);
nor U2294 (N_2294,In_612,In_1676);
xor U2295 (N_2295,In_138,In_2272);
and U2296 (N_2296,In_1260,In_35);
or U2297 (N_2297,In_1810,In_541);
nand U2298 (N_2298,In_2476,In_846);
and U2299 (N_2299,In_259,In_538);
or U2300 (N_2300,In_1920,In_603);
xor U2301 (N_2301,In_1303,In_1533);
nand U2302 (N_2302,In_763,In_670);
nand U2303 (N_2303,In_2166,In_2198);
nor U2304 (N_2304,In_1154,In_939);
nand U2305 (N_2305,In_1426,In_1144);
nand U2306 (N_2306,In_2245,In_1348);
nor U2307 (N_2307,In_1538,In_1490);
and U2308 (N_2308,In_2287,In_797);
nor U2309 (N_2309,In_986,In_314);
or U2310 (N_2310,In_2405,In_2136);
nor U2311 (N_2311,In_96,In_1692);
and U2312 (N_2312,In_341,In_2328);
nand U2313 (N_2313,In_284,In_2250);
nor U2314 (N_2314,In_1224,In_1573);
nand U2315 (N_2315,In_1726,In_2055);
nand U2316 (N_2316,In_154,In_484);
and U2317 (N_2317,In_1541,In_785);
nand U2318 (N_2318,In_900,In_1720);
or U2319 (N_2319,In_853,In_708);
nor U2320 (N_2320,In_763,In_1374);
and U2321 (N_2321,In_279,In_884);
nand U2322 (N_2322,In_1875,In_1553);
or U2323 (N_2323,In_2091,In_1919);
nor U2324 (N_2324,In_781,In_854);
nor U2325 (N_2325,In_1228,In_1186);
or U2326 (N_2326,In_2412,In_1184);
and U2327 (N_2327,In_541,In_2350);
xnor U2328 (N_2328,In_1531,In_1906);
nor U2329 (N_2329,In_1553,In_896);
nor U2330 (N_2330,In_1789,In_1305);
xnor U2331 (N_2331,In_1329,In_2443);
nand U2332 (N_2332,In_1193,In_2490);
or U2333 (N_2333,In_2124,In_1874);
nand U2334 (N_2334,In_566,In_361);
or U2335 (N_2335,In_915,In_1836);
nand U2336 (N_2336,In_1244,In_1087);
or U2337 (N_2337,In_75,In_2061);
nor U2338 (N_2338,In_2178,In_966);
and U2339 (N_2339,In_1646,In_434);
nand U2340 (N_2340,In_203,In_2332);
nor U2341 (N_2341,In_1253,In_298);
or U2342 (N_2342,In_1493,In_380);
or U2343 (N_2343,In_2019,In_2055);
nor U2344 (N_2344,In_1238,In_1678);
nand U2345 (N_2345,In_1870,In_1084);
or U2346 (N_2346,In_1922,In_1801);
or U2347 (N_2347,In_824,In_1717);
nor U2348 (N_2348,In_725,In_741);
and U2349 (N_2349,In_1026,In_659);
and U2350 (N_2350,In_1924,In_480);
and U2351 (N_2351,In_1796,In_2168);
nand U2352 (N_2352,In_908,In_647);
xnor U2353 (N_2353,In_1333,In_1765);
and U2354 (N_2354,In_2151,In_854);
and U2355 (N_2355,In_1836,In_902);
or U2356 (N_2356,In_248,In_1415);
xor U2357 (N_2357,In_1115,In_1858);
and U2358 (N_2358,In_1774,In_617);
and U2359 (N_2359,In_1798,In_292);
and U2360 (N_2360,In_163,In_1584);
or U2361 (N_2361,In_973,In_2270);
nand U2362 (N_2362,In_1168,In_308);
or U2363 (N_2363,In_1499,In_103);
xor U2364 (N_2364,In_2148,In_1160);
nand U2365 (N_2365,In_735,In_1557);
or U2366 (N_2366,In_2495,In_1943);
or U2367 (N_2367,In_840,In_572);
nand U2368 (N_2368,In_2156,In_1166);
or U2369 (N_2369,In_706,In_1325);
or U2370 (N_2370,In_450,In_2121);
nand U2371 (N_2371,In_1200,In_807);
and U2372 (N_2372,In_1595,In_439);
xnor U2373 (N_2373,In_921,In_681);
and U2374 (N_2374,In_1598,In_1178);
and U2375 (N_2375,In_1228,In_1923);
nor U2376 (N_2376,In_444,In_1860);
or U2377 (N_2377,In_2272,In_2138);
nand U2378 (N_2378,In_255,In_337);
nand U2379 (N_2379,In_809,In_1053);
or U2380 (N_2380,In_2368,In_2418);
nor U2381 (N_2381,In_531,In_1545);
or U2382 (N_2382,In_1699,In_1628);
nor U2383 (N_2383,In_2292,In_2455);
nand U2384 (N_2384,In_735,In_714);
or U2385 (N_2385,In_2159,In_2132);
nand U2386 (N_2386,In_2003,In_1748);
nand U2387 (N_2387,In_854,In_2253);
nor U2388 (N_2388,In_957,In_1082);
nand U2389 (N_2389,In_1626,In_1333);
xnor U2390 (N_2390,In_1963,In_723);
and U2391 (N_2391,In_320,In_1943);
nor U2392 (N_2392,In_928,In_1757);
and U2393 (N_2393,In_156,In_1986);
nor U2394 (N_2394,In_1402,In_354);
and U2395 (N_2395,In_956,In_1871);
nand U2396 (N_2396,In_1886,In_1447);
and U2397 (N_2397,In_164,In_2123);
nor U2398 (N_2398,In_1082,In_385);
nor U2399 (N_2399,In_65,In_1457);
nand U2400 (N_2400,In_1439,In_2204);
and U2401 (N_2401,In_1207,In_939);
nor U2402 (N_2402,In_1373,In_361);
or U2403 (N_2403,In_1503,In_198);
and U2404 (N_2404,In_1240,In_1316);
and U2405 (N_2405,In_599,In_1145);
nor U2406 (N_2406,In_1085,In_1718);
nand U2407 (N_2407,In_2490,In_1923);
nor U2408 (N_2408,In_897,In_141);
nand U2409 (N_2409,In_153,In_2202);
or U2410 (N_2410,In_1934,In_1362);
nor U2411 (N_2411,In_557,In_1761);
nor U2412 (N_2412,In_1861,In_1779);
and U2413 (N_2413,In_728,In_67);
nand U2414 (N_2414,In_204,In_830);
xnor U2415 (N_2415,In_970,In_1397);
or U2416 (N_2416,In_336,In_1003);
or U2417 (N_2417,In_378,In_147);
and U2418 (N_2418,In_2202,In_44);
or U2419 (N_2419,In_1179,In_1101);
nand U2420 (N_2420,In_2174,In_1082);
xor U2421 (N_2421,In_1906,In_886);
and U2422 (N_2422,In_2183,In_1358);
or U2423 (N_2423,In_1500,In_566);
and U2424 (N_2424,In_2361,In_2485);
nor U2425 (N_2425,In_1542,In_598);
nand U2426 (N_2426,In_1295,In_848);
nor U2427 (N_2427,In_1298,In_9);
nand U2428 (N_2428,In_464,In_2246);
nor U2429 (N_2429,In_1701,In_1672);
and U2430 (N_2430,In_1522,In_1764);
or U2431 (N_2431,In_1703,In_97);
nand U2432 (N_2432,In_1237,In_1175);
nand U2433 (N_2433,In_1753,In_1305);
nor U2434 (N_2434,In_1616,In_2035);
nand U2435 (N_2435,In_675,In_2063);
xnor U2436 (N_2436,In_585,In_2324);
nand U2437 (N_2437,In_109,In_242);
or U2438 (N_2438,In_602,In_282);
nand U2439 (N_2439,In_461,In_2250);
or U2440 (N_2440,In_1375,In_2003);
and U2441 (N_2441,In_1202,In_895);
nor U2442 (N_2442,In_16,In_1538);
and U2443 (N_2443,In_1086,In_992);
or U2444 (N_2444,In_309,In_1127);
xnor U2445 (N_2445,In_2366,In_1997);
nand U2446 (N_2446,In_2234,In_1562);
and U2447 (N_2447,In_749,In_934);
xnor U2448 (N_2448,In_1500,In_2354);
or U2449 (N_2449,In_2253,In_1887);
nor U2450 (N_2450,In_149,In_815);
nor U2451 (N_2451,In_1471,In_69);
nor U2452 (N_2452,In_1090,In_1453);
nor U2453 (N_2453,In_382,In_161);
nor U2454 (N_2454,In_1257,In_2460);
and U2455 (N_2455,In_2296,In_2198);
xnor U2456 (N_2456,In_891,In_124);
nand U2457 (N_2457,In_648,In_2280);
and U2458 (N_2458,In_901,In_628);
nand U2459 (N_2459,In_2190,In_1261);
nor U2460 (N_2460,In_285,In_1208);
or U2461 (N_2461,In_343,In_540);
nor U2462 (N_2462,In_1366,In_1966);
nor U2463 (N_2463,In_2075,In_1808);
nand U2464 (N_2464,In_2170,In_2376);
or U2465 (N_2465,In_202,In_2450);
and U2466 (N_2466,In_1621,In_2341);
and U2467 (N_2467,In_1259,In_512);
nand U2468 (N_2468,In_1273,In_2074);
nand U2469 (N_2469,In_2039,In_2006);
or U2470 (N_2470,In_933,In_952);
nor U2471 (N_2471,In_792,In_1141);
and U2472 (N_2472,In_690,In_241);
and U2473 (N_2473,In_1019,In_1232);
or U2474 (N_2474,In_1864,In_364);
or U2475 (N_2475,In_2014,In_2067);
nand U2476 (N_2476,In_1941,In_1914);
xnor U2477 (N_2477,In_880,In_413);
nand U2478 (N_2478,In_1119,In_2045);
or U2479 (N_2479,In_2122,In_439);
or U2480 (N_2480,In_524,In_2230);
and U2481 (N_2481,In_1911,In_95);
and U2482 (N_2482,In_1344,In_462);
nor U2483 (N_2483,In_499,In_4);
nand U2484 (N_2484,In_1512,In_401);
and U2485 (N_2485,In_2464,In_644);
xnor U2486 (N_2486,In_685,In_1978);
nand U2487 (N_2487,In_219,In_2283);
nand U2488 (N_2488,In_2210,In_495);
and U2489 (N_2489,In_532,In_1996);
or U2490 (N_2490,In_615,In_385);
nor U2491 (N_2491,In_273,In_2040);
or U2492 (N_2492,In_585,In_67);
nand U2493 (N_2493,In_1019,In_1195);
and U2494 (N_2494,In_1414,In_2332);
and U2495 (N_2495,In_2163,In_281);
or U2496 (N_2496,In_1873,In_2242);
or U2497 (N_2497,In_109,In_1919);
and U2498 (N_2498,In_871,In_1774);
nand U2499 (N_2499,In_1871,In_2033);
nand U2500 (N_2500,In_674,In_1591);
nand U2501 (N_2501,In_2340,In_2087);
nand U2502 (N_2502,In_1847,In_1355);
or U2503 (N_2503,In_1988,In_2094);
and U2504 (N_2504,In_1181,In_1446);
or U2505 (N_2505,In_54,In_1468);
nand U2506 (N_2506,In_601,In_948);
xnor U2507 (N_2507,In_1933,In_2126);
nand U2508 (N_2508,In_1509,In_581);
or U2509 (N_2509,In_1496,In_956);
or U2510 (N_2510,In_1379,In_1629);
and U2511 (N_2511,In_1947,In_2359);
nor U2512 (N_2512,In_150,In_1653);
nor U2513 (N_2513,In_350,In_1209);
nand U2514 (N_2514,In_1517,In_1258);
nand U2515 (N_2515,In_507,In_1391);
and U2516 (N_2516,In_1143,In_353);
or U2517 (N_2517,In_307,In_458);
nor U2518 (N_2518,In_893,In_934);
xnor U2519 (N_2519,In_633,In_679);
and U2520 (N_2520,In_1631,In_1923);
nor U2521 (N_2521,In_2033,In_520);
and U2522 (N_2522,In_853,In_1904);
and U2523 (N_2523,In_728,In_1745);
nor U2524 (N_2524,In_1428,In_1476);
or U2525 (N_2525,In_38,In_378);
xnor U2526 (N_2526,In_470,In_1264);
xor U2527 (N_2527,In_2176,In_493);
nand U2528 (N_2528,In_264,In_833);
nor U2529 (N_2529,In_1248,In_2068);
and U2530 (N_2530,In_2380,In_465);
and U2531 (N_2531,In_556,In_239);
nand U2532 (N_2532,In_2325,In_1990);
and U2533 (N_2533,In_359,In_2291);
and U2534 (N_2534,In_1020,In_1659);
nor U2535 (N_2535,In_671,In_804);
nor U2536 (N_2536,In_2172,In_1787);
nor U2537 (N_2537,In_1129,In_1713);
and U2538 (N_2538,In_205,In_1011);
xnor U2539 (N_2539,In_808,In_2169);
or U2540 (N_2540,In_721,In_979);
or U2541 (N_2541,In_1255,In_1468);
nor U2542 (N_2542,In_1001,In_1207);
nand U2543 (N_2543,In_1203,In_2447);
and U2544 (N_2544,In_1007,In_778);
xnor U2545 (N_2545,In_1458,In_279);
nand U2546 (N_2546,In_86,In_561);
nor U2547 (N_2547,In_722,In_1131);
nand U2548 (N_2548,In_869,In_753);
nand U2549 (N_2549,In_1103,In_2121);
or U2550 (N_2550,In_217,In_2391);
nand U2551 (N_2551,In_2342,In_1113);
nor U2552 (N_2552,In_572,In_1043);
nor U2553 (N_2553,In_2286,In_2469);
or U2554 (N_2554,In_1371,In_1961);
nand U2555 (N_2555,In_71,In_573);
nor U2556 (N_2556,In_1904,In_592);
nand U2557 (N_2557,In_366,In_2041);
or U2558 (N_2558,In_1578,In_570);
nor U2559 (N_2559,In_226,In_1382);
xnor U2560 (N_2560,In_2111,In_867);
nand U2561 (N_2561,In_376,In_588);
or U2562 (N_2562,In_127,In_1960);
nor U2563 (N_2563,In_5,In_2369);
nor U2564 (N_2564,In_154,In_2106);
nor U2565 (N_2565,In_2111,In_1372);
nor U2566 (N_2566,In_1254,In_1293);
nor U2567 (N_2567,In_2051,In_613);
and U2568 (N_2568,In_111,In_2498);
nor U2569 (N_2569,In_1733,In_2214);
or U2570 (N_2570,In_796,In_774);
and U2571 (N_2571,In_1673,In_689);
or U2572 (N_2572,In_2082,In_447);
nand U2573 (N_2573,In_2414,In_332);
nand U2574 (N_2574,In_2008,In_1640);
and U2575 (N_2575,In_729,In_2314);
or U2576 (N_2576,In_555,In_2396);
nand U2577 (N_2577,In_1878,In_142);
nand U2578 (N_2578,In_1607,In_1739);
or U2579 (N_2579,In_1157,In_148);
or U2580 (N_2580,In_2128,In_1085);
and U2581 (N_2581,In_848,In_845);
nand U2582 (N_2582,In_1407,In_1431);
and U2583 (N_2583,In_1302,In_1718);
nand U2584 (N_2584,In_1338,In_264);
nor U2585 (N_2585,In_906,In_2139);
nand U2586 (N_2586,In_669,In_1670);
and U2587 (N_2587,In_2386,In_1315);
or U2588 (N_2588,In_390,In_1154);
or U2589 (N_2589,In_1938,In_470);
or U2590 (N_2590,In_732,In_290);
nor U2591 (N_2591,In_2478,In_2090);
or U2592 (N_2592,In_626,In_558);
nor U2593 (N_2593,In_223,In_614);
nand U2594 (N_2594,In_1594,In_592);
xnor U2595 (N_2595,In_7,In_965);
nand U2596 (N_2596,In_319,In_778);
or U2597 (N_2597,In_352,In_998);
nor U2598 (N_2598,In_178,In_2118);
nand U2599 (N_2599,In_1514,In_251);
and U2600 (N_2600,In_1194,In_1199);
nand U2601 (N_2601,In_1225,In_1513);
or U2602 (N_2602,In_1071,In_2319);
nand U2603 (N_2603,In_1666,In_552);
nor U2604 (N_2604,In_150,In_2141);
and U2605 (N_2605,In_1826,In_1497);
and U2606 (N_2606,In_1790,In_1735);
or U2607 (N_2607,In_1305,In_2208);
or U2608 (N_2608,In_2120,In_568);
or U2609 (N_2609,In_1604,In_2431);
nor U2610 (N_2610,In_96,In_1716);
nor U2611 (N_2611,In_373,In_189);
and U2612 (N_2612,In_2331,In_1149);
and U2613 (N_2613,In_1665,In_2414);
nand U2614 (N_2614,In_110,In_2249);
nand U2615 (N_2615,In_1922,In_937);
or U2616 (N_2616,In_1555,In_1473);
nand U2617 (N_2617,In_1479,In_1874);
nand U2618 (N_2618,In_688,In_997);
nor U2619 (N_2619,In_2282,In_1007);
or U2620 (N_2620,In_952,In_1411);
and U2621 (N_2621,In_1395,In_1266);
xor U2622 (N_2622,In_87,In_2081);
and U2623 (N_2623,In_778,In_740);
nand U2624 (N_2624,In_1996,In_2467);
nor U2625 (N_2625,In_442,In_228);
nand U2626 (N_2626,In_1809,In_1046);
and U2627 (N_2627,In_164,In_622);
and U2628 (N_2628,In_1028,In_1931);
nor U2629 (N_2629,In_1792,In_662);
and U2630 (N_2630,In_774,In_1060);
nor U2631 (N_2631,In_446,In_2295);
nor U2632 (N_2632,In_2259,In_1953);
nand U2633 (N_2633,In_1164,In_498);
or U2634 (N_2634,In_385,In_1297);
nor U2635 (N_2635,In_1944,In_625);
nor U2636 (N_2636,In_611,In_2445);
nor U2637 (N_2637,In_410,In_2182);
nand U2638 (N_2638,In_1152,In_293);
or U2639 (N_2639,In_367,In_1597);
nor U2640 (N_2640,In_1917,In_618);
and U2641 (N_2641,In_1226,In_255);
and U2642 (N_2642,In_168,In_2318);
or U2643 (N_2643,In_1733,In_1913);
nor U2644 (N_2644,In_2474,In_1475);
or U2645 (N_2645,In_2107,In_1);
nor U2646 (N_2646,In_597,In_971);
and U2647 (N_2647,In_1314,In_340);
or U2648 (N_2648,In_2148,In_564);
nor U2649 (N_2649,In_472,In_985);
nand U2650 (N_2650,In_912,In_1494);
nand U2651 (N_2651,In_2108,In_608);
or U2652 (N_2652,In_1013,In_1321);
or U2653 (N_2653,In_2362,In_1816);
or U2654 (N_2654,In_427,In_1283);
or U2655 (N_2655,In_1086,In_188);
or U2656 (N_2656,In_1285,In_44);
nand U2657 (N_2657,In_139,In_619);
or U2658 (N_2658,In_950,In_348);
nor U2659 (N_2659,In_1059,In_709);
and U2660 (N_2660,In_969,In_1147);
nor U2661 (N_2661,In_2349,In_2339);
or U2662 (N_2662,In_1829,In_35);
xnor U2663 (N_2663,In_469,In_268);
and U2664 (N_2664,In_2155,In_2462);
nand U2665 (N_2665,In_1717,In_771);
nand U2666 (N_2666,In_1050,In_476);
xor U2667 (N_2667,In_81,In_2485);
nor U2668 (N_2668,In_545,In_1064);
or U2669 (N_2669,In_2325,In_316);
nor U2670 (N_2670,In_2241,In_914);
or U2671 (N_2671,In_1880,In_1164);
nand U2672 (N_2672,In_2076,In_1335);
nor U2673 (N_2673,In_873,In_49);
nor U2674 (N_2674,In_2245,In_1301);
xnor U2675 (N_2675,In_216,In_2418);
xnor U2676 (N_2676,In_2142,In_541);
and U2677 (N_2677,In_1370,In_2099);
or U2678 (N_2678,In_500,In_2038);
nor U2679 (N_2679,In_1088,In_1914);
nor U2680 (N_2680,In_804,In_1166);
or U2681 (N_2681,In_63,In_2405);
or U2682 (N_2682,In_492,In_2411);
xnor U2683 (N_2683,In_1083,In_1688);
and U2684 (N_2684,In_2328,In_238);
or U2685 (N_2685,In_2307,In_623);
and U2686 (N_2686,In_2440,In_1248);
nor U2687 (N_2687,In_2341,In_2085);
and U2688 (N_2688,In_2183,In_473);
or U2689 (N_2689,In_1560,In_2142);
nor U2690 (N_2690,In_2272,In_645);
nand U2691 (N_2691,In_113,In_1905);
nand U2692 (N_2692,In_2275,In_712);
xor U2693 (N_2693,In_541,In_1549);
xnor U2694 (N_2694,In_2315,In_2270);
and U2695 (N_2695,In_72,In_762);
or U2696 (N_2696,In_2207,In_252);
or U2697 (N_2697,In_2356,In_2177);
and U2698 (N_2698,In_362,In_810);
nand U2699 (N_2699,In_2313,In_1400);
nand U2700 (N_2700,In_2304,In_964);
nor U2701 (N_2701,In_1019,In_1021);
xor U2702 (N_2702,In_325,In_1083);
nand U2703 (N_2703,In_1252,In_193);
xnor U2704 (N_2704,In_111,In_178);
and U2705 (N_2705,In_1232,In_875);
or U2706 (N_2706,In_5,In_2489);
nand U2707 (N_2707,In_2216,In_2252);
or U2708 (N_2708,In_1939,In_80);
and U2709 (N_2709,In_1242,In_2013);
and U2710 (N_2710,In_1783,In_660);
xnor U2711 (N_2711,In_1740,In_2265);
nand U2712 (N_2712,In_1347,In_1328);
nand U2713 (N_2713,In_651,In_848);
and U2714 (N_2714,In_589,In_1268);
xnor U2715 (N_2715,In_135,In_71);
nand U2716 (N_2716,In_397,In_1398);
or U2717 (N_2717,In_152,In_470);
or U2718 (N_2718,In_457,In_1817);
and U2719 (N_2719,In_57,In_1944);
nor U2720 (N_2720,In_1359,In_398);
nor U2721 (N_2721,In_1793,In_2258);
xor U2722 (N_2722,In_2155,In_2398);
xor U2723 (N_2723,In_1099,In_939);
xor U2724 (N_2724,In_2038,In_2279);
nand U2725 (N_2725,In_1205,In_2390);
nor U2726 (N_2726,In_2260,In_2403);
xor U2727 (N_2727,In_429,In_2241);
nor U2728 (N_2728,In_79,In_553);
and U2729 (N_2729,In_995,In_205);
or U2730 (N_2730,In_63,In_2364);
xor U2731 (N_2731,In_2120,In_1239);
nor U2732 (N_2732,In_649,In_1770);
or U2733 (N_2733,In_644,In_1657);
xor U2734 (N_2734,In_1274,In_2174);
nand U2735 (N_2735,In_1982,In_878);
nand U2736 (N_2736,In_210,In_1534);
and U2737 (N_2737,In_2131,In_1303);
xor U2738 (N_2738,In_479,In_478);
xnor U2739 (N_2739,In_604,In_1163);
nor U2740 (N_2740,In_1975,In_2491);
nor U2741 (N_2741,In_1909,In_1788);
nand U2742 (N_2742,In_1282,In_2377);
or U2743 (N_2743,In_1015,In_691);
xnor U2744 (N_2744,In_2009,In_1213);
or U2745 (N_2745,In_1595,In_1593);
nor U2746 (N_2746,In_1234,In_213);
nand U2747 (N_2747,In_359,In_1876);
and U2748 (N_2748,In_1976,In_1381);
and U2749 (N_2749,In_1213,In_2236);
and U2750 (N_2750,In_2231,In_2439);
nor U2751 (N_2751,In_2214,In_943);
nand U2752 (N_2752,In_131,In_1414);
nor U2753 (N_2753,In_24,In_443);
nor U2754 (N_2754,In_1705,In_806);
or U2755 (N_2755,In_2109,In_2269);
xnor U2756 (N_2756,In_15,In_1616);
nand U2757 (N_2757,In_527,In_735);
nor U2758 (N_2758,In_513,In_434);
xor U2759 (N_2759,In_1600,In_594);
and U2760 (N_2760,In_2092,In_463);
and U2761 (N_2761,In_1013,In_2169);
and U2762 (N_2762,In_1814,In_1558);
nor U2763 (N_2763,In_553,In_1111);
nor U2764 (N_2764,In_368,In_1956);
nand U2765 (N_2765,In_2431,In_1301);
or U2766 (N_2766,In_2051,In_804);
or U2767 (N_2767,In_1926,In_826);
nor U2768 (N_2768,In_1217,In_2316);
nand U2769 (N_2769,In_1552,In_1055);
nor U2770 (N_2770,In_494,In_1179);
nand U2771 (N_2771,In_654,In_710);
or U2772 (N_2772,In_529,In_1428);
nand U2773 (N_2773,In_2258,In_1891);
or U2774 (N_2774,In_2428,In_1450);
nand U2775 (N_2775,In_1721,In_1748);
nor U2776 (N_2776,In_1849,In_1494);
or U2777 (N_2777,In_1619,In_588);
nor U2778 (N_2778,In_1870,In_124);
nand U2779 (N_2779,In_2432,In_1843);
xnor U2780 (N_2780,In_1940,In_160);
nand U2781 (N_2781,In_1458,In_767);
and U2782 (N_2782,In_1393,In_1975);
nand U2783 (N_2783,In_2068,In_1579);
xnor U2784 (N_2784,In_463,In_2109);
and U2785 (N_2785,In_38,In_2450);
nor U2786 (N_2786,In_960,In_2034);
nor U2787 (N_2787,In_2099,In_1098);
nand U2788 (N_2788,In_1356,In_1256);
nor U2789 (N_2789,In_543,In_1298);
nor U2790 (N_2790,In_276,In_1288);
nand U2791 (N_2791,In_844,In_97);
nor U2792 (N_2792,In_187,In_1703);
nand U2793 (N_2793,In_1638,In_2064);
and U2794 (N_2794,In_644,In_667);
and U2795 (N_2795,In_2436,In_1231);
and U2796 (N_2796,In_1217,In_1113);
nand U2797 (N_2797,In_801,In_550);
nor U2798 (N_2798,In_2427,In_2475);
nor U2799 (N_2799,In_99,In_2037);
xnor U2800 (N_2800,In_775,In_1296);
nand U2801 (N_2801,In_2155,In_234);
and U2802 (N_2802,In_2411,In_2475);
and U2803 (N_2803,In_127,In_2149);
and U2804 (N_2804,In_680,In_656);
and U2805 (N_2805,In_322,In_692);
nor U2806 (N_2806,In_407,In_613);
nand U2807 (N_2807,In_603,In_1345);
nand U2808 (N_2808,In_523,In_1064);
and U2809 (N_2809,In_1408,In_1644);
and U2810 (N_2810,In_532,In_1583);
nand U2811 (N_2811,In_4,In_432);
and U2812 (N_2812,In_1072,In_2319);
nor U2813 (N_2813,In_1629,In_1282);
and U2814 (N_2814,In_1655,In_254);
nor U2815 (N_2815,In_416,In_2214);
nor U2816 (N_2816,In_2470,In_382);
or U2817 (N_2817,In_1012,In_2417);
and U2818 (N_2818,In_2265,In_1453);
xnor U2819 (N_2819,In_2154,In_1143);
and U2820 (N_2820,In_2349,In_1960);
nor U2821 (N_2821,In_2479,In_223);
and U2822 (N_2822,In_400,In_1788);
nor U2823 (N_2823,In_642,In_1620);
nand U2824 (N_2824,In_2411,In_1176);
nor U2825 (N_2825,In_478,In_1687);
and U2826 (N_2826,In_1660,In_373);
or U2827 (N_2827,In_1541,In_801);
nor U2828 (N_2828,In_1873,In_1718);
nor U2829 (N_2829,In_1819,In_1889);
nor U2830 (N_2830,In_1791,In_572);
nand U2831 (N_2831,In_1577,In_2282);
or U2832 (N_2832,In_1510,In_745);
or U2833 (N_2833,In_2306,In_1752);
nor U2834 (N_2834,In_624,In_2276);
or U2835 (N_2835,In_1500,In_1478);
nand U2836 (N_2836,In_1972,In_2237);
nand U2837 (N_2837,In_2137,In_1435);
or U2838 (N_2838,In_1054,In_435);
or U2839 (N_2839,In_397,In_960);
and U2840 (N_2840,In_1247,In_882);
nand U2841 (N_2841,In_34,In_1943);
nand U2842 (N_2842,In_1596,In_381);
nor U2843 (N_2843,In_1566,In_1746);
and U2844 (N_2844,In_1560,In_2124);
nand U2845 (N_2845,In_236,In_453);
nor U2846 (N_2846,In_1047,In_1726);
or U2847 (N_2847,In_2198,In_2117);
or U2848 (N_2848,In_1231,In_120);
and U2849 (N_2849,In_1569,In_2441);
nor U2850 (N_2850,In_1875,In_1726);
nand U2851 (N_2851,In_1376,In_1003);
and U2852 (N_2852,In_803,In_498);
xor U2853 (N_2853,In_161,In_721);
nand U2854 (N_2854,In_326,In_2399);
xor U2855 (N_2855,In_1331,In_842);
and U2856 (N_2856,In_1007,In_1572);
or U2857 (N_2857,In_674,In_998);
and U2858 (N_2858,In_423,In_1165);
or U2859 (N_2859,In_2377,In_1727);
xnor U2860 (N_2860,In_1815,In_801);
and U2861 (N_2861,In_137,In_2429);
and U2862 (N_2862,In_125,In_1439);
nand U2863 (N_2863,In_476,In_715);
or U2864 (N_2864,In_283,In_1040);
or U2865 (N_2865,In_1154,In_647);
or U2866 (N_2866,In_330,In_714);
nor U2867 (N_2867,In_403,In_2488);
or U2868 (N_2868,In_2201,In_1946);
and U2869 (N_2869,In_2074,In_819);
nor U2870 (N_2870,In_1092,In_1763);
nand U2871 (N_2871,In_288,In_1240);
and U2872 (N_2872,In_900,In_2498);
or U2873 (N_2873,In_1449,In_730);
nor U2874 (N_2874,In_390,In_930);
nand U2875 (N_2875,In_1637,In_464);
nand U2876 (N_2876,In_1711,In_1297);
nor U2877 (N_2877,In_815,In_2405);
and U2878 (N_2878,In_2057,In_1781);
nand U2879 (N_2879,In_770,In_2154);
nor U2880 (N_2880,In_926,In_2497);
nor U2881 (N_2881,In_1951,In_474);
nor U2882 (N_2882,In_2110,In_107);
or U2883 (N_2883,In_608,In_2276);
or U2884 (N_2884,In_11,In_1651);
xor U2885 (N_2885,In_344,In_496);
nor U2886 (N_2886,In_1702,In_1278);
nor U2887 (N_2887,In_2323,In_2409);
nand U2888 (N_2888,In_72,In_1545);
nand U2889 (N_2889,In_1001,In_2369);
and U2890 (N_2890,In_493,In_1637);
nor U2891 (N_2891,In_1248,In_690);
and U2892 (N_2892,In_488,In_214);
and U2893 (N_2893,In_2312,In_1553);
or U2894 (N_2894,In_1358,In_1240);
or U2895 (N_2895,In_89,In_1856);
nor U2896 (N_2896,In_1469,In_971);
nor U2897 (N_2897,In_11,In_12);
and U2898 (N_2898,In_1064,In_1681);
or U2899 (N_2899,In_2259,In_1950);
or U2900 (N_2900,In_2101,In_2483);
nand U2901 (N_2901,In_450,In_2379);
nand U2902 (N_2902,In_8,In_2490);
or U2903 (N_2903,In_745,In_1736);
nor U2904 (N_2904,In_1133,In_886);
xor U2905 (N_2905,In_1413,In_105);
and U2906 (N_2906,In_838,In_2453);
nor U2907 (N_2907,In_261,In_612);
and U2908 (N_2908,In_1389,In_2249);
nor U2909 (N_2909,In_351,In_1683);
nor U2910 (N_2910,In_2001,In_2152);
xnor U2911 (N_2911,In_2110,In_139);
nor U2912 (N_2912,In_693,In_1047);
and U2913 (N_2913,In_1392,In_1699);
or U2914 (N_2914,In_1030,In_1539);
nor U2915 (N_2915,In_825,In_1007);
xor U2916 (N_2916,In_792,In_1347);
nor U2917 (N_2917,In_1521,In_991);
nand U2918 (N_2918,In_2101,In_1694);
and U2919 (N_2919,In_1191,In_1317);
or U2920 (N_2920,In_1779,In_1214);
xnor U2921 (N_2921,In_1559,In_2362);
and U2922 (N_2922,In_1581,In_2180);
nand U2923 (N_2923,In_1971,In_683);
nor U2924 (N_2924,In_1257,In_1275);
and U2925 (N_2925,In_971,In_634);
and U2926 (N_2926,In_960,In_1171);
and U2927 (N_2927,In_2392,In_978);
or U2928 (N_2928,In_1703,In_707);
or U2929 (N_2929,In_2435,In_1809);
nand U2930 (N_2930,In_785,In_461);
nor U2931 (N_2931,In_1997,In_435);
and U2932 (N_2932,In_1076,In_2200);
nand U2933 (N_2933,In_1155,In_1241);
or U2934 (N_2934,In_623,In_652);
nand U2935 (N_2935,In_1071,In_657);
or U2936 (N_2936,In_2326,In_1104);
and U2937 (N_2937,In_1157,In_2437);
xor U2938 (N_2938,In_2122,In_12);
nor U2939 (N_2939,In_1407,In_1790);
nor U2940 (N_2940,In_96,In_1269);
and U2941 (N_2941,In_2227,In_2285);
nand U2942 (N_2942,In_336,In_928);
or U2943 (N_2943,In_634,In_1531);
nand U2944 (N_2944,In_1939,In_885);
xor U2945 (N_2945,In_1080,In_22);
or U2946 (N_2946,In_619,In_499);
xnor U2947 (N_2947,In_347,In_1258);
or U2948 (N_2948,In_770,In_1181);
nor U2949 (N_2949,In_1423,In_215);
or U2950 (N_2950,In_10,In_92);
nand U2951 (N_2951,In_1527,In_372);
nor U2952 (N_2952,In_1980,In_22);
nand U2953 (N_2953,In_274,In_2150);
nor U2954 (N_2954,In_2266,In_362);
or U2955 (N_2955,In_1711,In_1213);
nand U2956 (N_2956,In_477,In_1324);
or U2957 (N_2957,In_2155,In_37);
nand U2958 (N_2958,In_2357,In_2297);
nand U2959 (N_2959,In_793,In_366);
or U2960 (N_2960,In_1199,In_354);
xnor U2961 (N_2961,In_1580,In_669);
nand U2962 (N_2962,In_192,In_1650);
and U2963 (N_2963,In_6,In_426);
and U2964 (N_2964,In_417,In_522);
nor U2965 (N_2965,In_2070,In_423);
nand U2966 (N_2966,In_2379,In_47);
nand U2967 (N_2967,In_859,In_626);
nor U2968 (N_2968,In_1565,In_1136);
and U2969 (N_2969,In_2129,In_388);
and U2970 (N_2970,In_495,In_2267);
nor U2971 (N_2971,In_244,In_2495);
nor U2972 (N_2972,In_2246,In_1263);
or U2973 (N_2973,In_1980,In_1366);
and U2974 (N_2974,In_1824,In_1339);
or U2975 (N_2975,In_2436,In_2203);
or U2976 (N_2976,In_1005,In_2305);
nand U2977 (N_2977,In_1176,In_573);
and U2978 (N_2978,In_2119,In_1271);
nor U2979 (N_2979,In_673,In_1416);
nand U2980 (N_2980,In_270,In_1263);
and U2981 (N_2981,In_198,In_1563);
nand U2982 (N_2982,In_1657,In_24);
nand U2983 (N_2983,In_1487,In_559);
or U2984 (N_2984,In_2380,In_2472);
nor U2985 (N_2985,In_1716,In_624);
and U2986 (N_2986,In_1294,In_2338);
and U2987 (N_2987,In_129,In_116);
nor U2988 (N_2988,In_1710,In_2422);
or U2989 (N_2989,In_1754,In_828);
nor U2990 (N_2990,In_24,In_1443);
or U2991 (N_2991,In_1537,In_2121);
and U2992 (N_2992,In_1653,In_1727);
and U2993 (N_2993,In_604,In_224);
nand U2994 (N_2994,In_1117,In_748);
nand U2995 (N_2995,In_2150,In_123);
nor U2996 (N_2996,In_488,In_2104);
nor U2997 (N_2997,In_1311,In_625);
or U2998 (N_2998,In_377,In_1627);
nand U2999 (N_2999,In_1663,In_1584);
xnor U3000 (N_3000,In_192,In_962);
and U3001 (N_3001,In_1956,In_503);
xor U3002 (N_3002,In_797,In_2477);
xnor U3003 (N_3003,In_1765,In_1568);
nand U3004 (N_3004,In_1962,In_37);
or U3005 (N_3005,In_2377,In_494);
and U3006 (N_3006,In_1604,In_929);
xor U3007 (N_3007,In_1490,In_2459);
nand U3008 (N_3008,In_86,In_1737);
nor U3009 (N_3009,In_685,In_702);
nor U3010 (N_3010,In_1008,In_1540);
nor U3011 (N_3011,In_2337,In_1910);
or U3012 (N_3012,In_2005,In_477);
or U3013 (N_3013,In_937,In_894);
nand U3014 (N_3014,In_1155,In_253);
and U3015 (N_3015,In_1368,In_2004);
or U3016 (N_3016,In_1113,In_1033);
or U3017 (N_3017,In_159,In_2246);
nand U3018 (N_3018,In_900,In_792);
nor U3019 (N_3019,In_784,In_1460);
or U3020 (N_3020,In_1003,In_443);
nor U3021 (N_3021,In_1209,In_2349);
or U3022 (N_3022,In_1051,In_1670);
nor U3023 (N_3023,In_1034,In_1171);
or U3024 (N_3024,In_1089,In_180);
xor U3025 (N_3025,In_677,In_1023);
or U3026 (N_3026,In_111,In_1986);
nand U3027 (N_3027,In_1999,In_954);
and U3028 (N_3028,In_681,In_1798);
and U3029 (N_3029,In_368,In_834);
or U3030 (N_3030,In_358,In_2151);
xor U3031 (N_3031,In_2049,In_27);
or U3032 (N_3032,In_301,In_1556);
and U3033 (N_3033,In_244,In_2107);
or U3034 (N_3034,In_1809,In_405);
nand U3035 (N_3035,In_156,In_1300);
nand U3036 (N_3036,In_1157,In_875);
and U3037 (N_3037,In_640,In_757);
nor U3038 (N_3038,In_1931,In_2210);
nor U3039 (N_3039,In_2405,In_212);
nor U3040 (N_3040,In_2298,In_2430);
and U3041 (N_3041,In_687,In_1010);
nor U3042 (N_3042,In_2493,In_1440);
nand U3043 (N_3043,In_1958,In_2122);
or U3044 (N_3044,In_483,In_417);
or U3045 (N_3045,In_639,In_1123);
and U3046 (N_3046,In_399,In_1145);
nor U3047 (N_3047,In_1917,In_1873);
nor U3048 (N_3048,In_92,In_664);
nor U3049 (N_3049,In_1279,In_1766);
nor U3050 (N_3050,In_2079,In_24);
or U3051 (N_3051,In_700,In_181);
nand U3052 (N_3052,In_82,In_1051);
and U3053 (N_3053,In_1170,In_1332);
nor U3054 (N_3054,In_2224,In_1180);
or U3055 (N_3055,In_1987,In_1401);
and U3056 (N_3056,In_927,In_1539);
xnor U3057 (N_3057,In_751,In_771);
nor U3058 (N_3058,In_1401,In_1404);
and U3059 (N_3059,In_1004,In_2309);
xnor U3060 (N_3060,In_1930,In_1243);
nand U3061 (N_3061,In_1353,In_1491);
nor U3062 (N_3062,In_189,In_1823);
or U3063 (N_3063,In_1046,In_2142);
or U3064 (N_3064,In_2271,In_1995);
xnor U3065 (N_3065,In_576,In_394);
or U3066 (N_3066,In_1710,In_614);
or U3067 (N_3067,In_2131,In_1764);
and U3068 (N_3068,In_1721,In_2007);
nor U3069 (N_3069,In_448,In_1283);
nand U3070 (N_3070,In_1236,In_687);
nor U3071 (N_3071,In_804,In_1439);
nand U3072 (N_3072,In_246,In_2096);
nand U3073 (N_3073,In_974,In_836);
nor U3074 (N_3074,In_1629,In_353);
and U3075 (N_3075,In_1198,In_1319);
or U3076 (N_3076,In_347,In_709);
nand U3077 (N_3077,In_1559,In_2367);
or U3078 (N_3078,In_413,In_1672);
nand U3079 (N_3079,In_602,In_1062);
nor U3080 (N_3080,In_1539,In_276);
xnor U3081 (N_3081,In_2352,In_322);
or U3082 (N_3082,In_2370,In_1017);
nor U3083 (N_3083,In_839,In_2076);
and U3084 (N_3084,In_693,In_2083);
and U3085 (N_3085,In_1909,In_1968);
nor U3086 (N_3086,In_1973,In_1995);
and U3087 (N_3087,In_589,In_1874);
nand U3088 (N_3088,In_1460,In_1900);
nand U3089 (N_3089,In_1120,In_1338);
or U3090 (N_3090,In_592,In_2324);
nor U3091 (N_3091,In_2201,In_1227);
and U3092 (N_3092,In_975,In_764);
nor U3093 (N_3093,In_262,In_777);
nor U3094 (N_3094,In_76,In_1411);
nor U3095 (N_3095,In_1897,In_2180);
nor U3096 (N_3096,In_241,In_1155);
nor U3097 (N_3097,In_2004,In_25);
nand U3098 (N_3098,In_2491,In_1652);
or U3099 (N_3099,In_896,In_1536);
and U3100 (N_3100,In_1734,In_1202);
or U3101 (N_3101,In_2489,In_1445);
or U3102 (N_3102,In_287,In_1202);
nand U3103 (N_3103,In_642,In_1179);
xnor U3104 (N_3104,In_2094,In_386);
and U3105 (N_3105,In_732,In_494);
or U3106 (N_3106,In_795,In_2354);
nand U3107 (N_3107,In_1592,In_1156);
nand U3108 (N_3108,In_1956,In_532);
nand U3109 (N_3109,In_1738,In_543);
xor U3110 (N_3110,In_1778,In_1800);
nor U3111 (N_3111,In_2054,In_351);
nor U3112 (N_3112,In_1782,In_960);
nor U3113 (N_3113,In_719,In_135);
nand U3114 (N_3114,In_447,In_2394);
nand U3115 (N_3115,In_976,In_1037);
and U3116 (N_3116,In_152,In_1804);
nor U3117 (N_3117,In_2399,In_179);
and U3118 (N_3118,In_1065,In_2166);
and U3119 (N_3119,In_1931,In_962);
nor U3120 (N_3120,In_992,In_2124);
or U3121 (N_3121,In_2480,In_98);
or U3122 (N_3122,In_2416,In_2388);
xnor U3123 (N_3123,In_1502,In_41);
nor U3124 (N_3124,In_1826,In_624);
or U3125 (N_3125,In_865,In_2293);
or U3126 (N_3126,In_247,In_1673);
nand U3127 (N_3127,In_985,In_1227);
nor U3128 (N_3128,In_317,In_985);
or U3129 (N_3129,In_1477,In_873);
nand U3130 (N_3130,In_2111,In_1985);
nand U3131 (N_3131,In_1254,In_1029);
nor U3132 (N_3132,In_2304,In_1290);
or U3133 (N_3133,In_1676,In_2433);
or U3134 (N_3134,In_1349,In_1880);
xor U3135 (N_3135,In_2248,In_2007);
nand U3136 (N_3136,In_762,In_1906);
nor U3137 (N_3137,In_1531,In_462);
xor U3138 (N_3138,In_351,In_271);
and U3139 (N_3139,In_373,In_1720);
nor U3140 (N_3140,In_2043,In_2095);
or U3141 (N_3141,In_1396,In_959);
or U3142 (N_3142,In_677,In_1598);
nand U3143 (N_3143,In_2434,In_1208);
nor U3144 (N_3144,In_1937,In_173);
and U3145 (N_3145,In_1021,In_483);
nor U3146 (N_3146,In_2218,In_195);
nand U3147 (N_3147,In_557,In_1880);
and U3148 (N_3148,In_1691,In_956);
and U3149 (N_3149,In_1425,In_1589);
or U3150 (N_3150,In_1834,In_332);
nand U3151 (N_3151,In_134,In_1902);
or U3152 (N_3152,In_251,In_661);
and U3153 (N_3153,In_1280,In_140);
xor U3154 (N_3154,In_659,In_1288);
or U3155 (N_3155,In_137,In_290);
nand U3156 (N_3156,In_2456,In_222);
and U3157 (N_3157,In_115,In_378);
and U3158 (N_3158,In_1140,In_131);
nand U3159 (N_3159,In_687,In_1271);
nand U3160 (N_3160,In_1300,In_35);
nand U3161 (N_3161,In_498,In_2380);
nor U3162 (N_3162,In_583,In_869);
xnor U3163 (N_3163,In_237,In_1678);
xor U3164 (N_3164,In_99,In_1431);
and U3165 (N_3165,In_1796,In_1308);
or U3166 (N_3166,In_1263,In_1102);
or U3167 (N_3167,In_1465,In_52);
nand U3168 (N_3168,In_1716,In_462);
nor U3169 (N_3169,In_157,In_2057);
nor U3170 (N_3170,In_903,In_1318);
nand U3171 (N_3171,In_467,In_1166);
nor U3172 (N_3172,In_1046,In_1131);
nand U3173 (N_3173,In_656,In_1663);
xor U3174 (N_3174,In_1845,In_63);
nand U3175 (N_3175,In_694,In_1618);
nand U3176 (N_3176,In_602,In_2131);
nor U3177 (N_3177,In_1229,In_1757);
xor U3178 (N_3178,In_2348,In_1239);
or U3179 (N_3179,In_2175,In_184);
nor U3180 (N_3180,In_1437,In_714);
or U3181 (N_3181,In_2417,In_1868);
nand U3182 (N_3182,In_259,In_1611);
nor U3183 (N_3183,In_1313,In_285);
and U3184 (N_3184,In_1506,In_1692);
xor U3185 (N_3185,In_1643,In_2124);
and U3186 (N_3186,In_2100,In_1066);
nor U3187 (N_3187,In_309,In_2346);
nand U3188 (N_3188,In_788,In_55);
nand U3189 (N_3189,In_994,In_2023);
and U3190 (N_3190,In_1968,In_1610);
or U3191 (N_3191,In_1487,In_1787);
and U3192 (N_3192,In_1921,In_2378);
and U3193 (N_3193,In_1183,In_1728);
or U3194 (N_3194,In_1751,In_1016);
xor U3195 (N_3195,In_404,In_226);
xor U3196 (N_3196,In_213,In_632);
or U3197 (N_3197,In_1962,In_474);
and U3198 (N_3198,In_595,In_2413);
or U3199 (N_3199,In_1123,In_1155);
nor U3200 (N_3200,In_700,In_1589);
xnor U3201 (N_3201,In_1843,In_2288);
nand U3202 (N_3202,In_1214,In_1097);
or U3203 (N_3203,In_1619,In_2014);
or U3204 (N_3204,In_2337,In_2059);
nand U3205 (N_3205,In_469,In_1439);
xnor U3206 (N_3206,In_2350,In_574);
nor U3207 (N_3207,In_1586,In_1450);
nand U3208 (N_3208,In_350,In_1535);
or U3209 (N_3209,In_1033,In_751);
nand U3210 (N_3210,In_1046,In_707);
and U3211 (N_3211,In_1865,In_290);
or U3212 (N_3212,In_1222,In_2308);
and U3213 (N_3213,In_1151,In_583);
xor U3214 (N_3214,In_1261,In_725);
nand U3215 (N_3215,In_1826,In_1397);
nor U3216 (N_3216,In_799,In_1847);
nor U3217 (N_3217,In_765,In_985);
nor U3218 (N_3218,In_576,In_1608);
or U3219 (N_3219,In_60,In_2399);
nand U3220 (N_3220,In_80,In_1157);
nor U3221 (N_3221,In_988,In_720);
or U3222 (N_3222,In_2413,In_2432);
or U3223 (N_3223,In_584,In_730);
nor U3224 (N_3224,In_1350,In_2139);
and U3225 (N_3225,In_2377,In_1186);
nand U3226 (N_3226,In_821,In_38);
and U3227 (N_3227,In_702,In_1573);
xor U3228 (N_3228,In_1961,In_2383);
nand U3229 (N_3229,In_2435,In_1726);
xnor U3230 (N_3230,In_1782,In_2052);
xor U3231 (N_3231,In_1095,In_642);
or U3232 (N_3232,In_552,In_1358);
and U3233 (N_3233,In_1966,In_1994);
nor U3234 (N_3234,In_1875,In_32);
nand U3235 (N_3235,In_1587,In_2254);
nor U3236 (N_3236,In_1309,In_473);
nand U3237 (N_3237,In_947,In_1246);
nor U3238 (N_3238,In_1417,In_1323);
and U3239 (N_3239,In_462,In_2295);
nand U3240 (N_3240,In_1378,In_2378);
nand U3241 (N_3241,In_2047,In_132);
and U3242 (N_3242,In_760,In_2446);
nor U3243 (N_3243,In_2306,In_502);
nor U3244 (N_3244,In_1068,In_458);
or U3245 (N_3245,In_302,In_2420);
and U3246 (N_3246,In_2451,In_2322);
nor U3247 (N_3247,In_1319,In_730);
nand U3248 (N_3248,In_1827,In_976);
and U3249 (N_3249,In_159,In_1049);
nand U3250 (N_3250,In_139,In_677);
xnor U3251 (N_3251,In_1661,In_1563);
or U3252 (N_3252,In_534,In_2497);
nor U3253 (N_3253,In_613,In_786);
nand U3254 (N_3254,In_2031,In_499);
or U3255 (N_3255,In_883,In_102);
nand U3256 (N_3256,In_1910,In_458);
or U3257 (N_3257,In_1988,In_1350);
or U3258 (N_3258,In_1742,In_1993);
nand U3259 (N_3259,In_440,In_1608);
or U3260 (N_3260,In_1321,In_831);
and U3261 (N_3261,In_1516,In_983);
or U3262 (N_3262,In_1743,In_147);
or U3263 (N_3263,In_1993,In_2423);
and U3264 (N_3264,In_896,In_634);
and U3265 (N_3265,In_275,In_1071);
and U3266 (N_3266,In_2409,In_2349);
xnor U3267 (N_3267,In_87,In_52);
nand U3268 (N_3268,In_1994,In_1709);
nor U3269 (N_3269,In_1842,In_233);
nand U3270 (N_3270,In_1622,In_221);
or U3271 (N_3271,In_1693,In_20);
xor U3272 (N_3272,In_2196,In_783);
and U3273 (N_3273,In_2186,In_644);
xor U3274 (N_3274,In_712,In_876);
or U3275 (N_3275,In_1032,In_2165);
nor U3276 (N_3276,In_1283,In_1324);
nand U3277 (N_3277,In_1479,In_502);
nor U3278 (N_3278,In_1506,In_763);
nor U3279 (N_3279,In_1119,In_6);
xnor U3280 (N_3280,In_936,In_437);
and U3281 (N_3281,In_2257,In_621);
nand U3282 (N_3282,In_109,In_2248);
or U3283 (N_3283,In_976,In_1458);
nand U3284 (N_3284,In_1874,In_236);
nand U3285 (N_3285,In_179,In_878);
nand U3286 (N_3286,In_2267,In_1850);
and U3287 (N_3287,In_1311,In_2138);
nor U3288 (N_3288,In_686,In_1276);
nand U3289 (N_3289,In_383,In_2199);
nand U3290 (N_3290,In_950,In_3);
nand U3291 (N_3291,In_2397,In_844);
and U3292 (N_3292,In_607,In_244);
nand U3293 (N_3293,In_192,In_326);
nor U3294 (N_3294,In_2434,In_348);
nor U3295 (N_3295,In_1637,In_2066);
or U3296 (N_3296,In_389,In_195);
or U3297 (N_3297,In_1522,In_164);
and U3298 (N_3298,In_870,In_254);
and U3299 (N_3299,In_1551,In_287);
and U3300 (N_3300,In_643,In_541);
nor U3301 (N_3301,In_2085,In_1851);
or U3302 (N_3302,In_1561,In_788);
xor U3303 (N_3303,In_1099,In_1357);
nor U3304 (N_3304,In_94,In_1765);
nand U3305 (N_3305,In_1681,In_1445);
and U3306 (N_3306,In_1410,In_1816);
or U3307 (N_3307,In_1949,In_56);
or U3308 (N_3308,In_1643,In_1798);
or U3309 (N_3309,In_991,In_529);
or U3310 (N_3310,In_1415,In_1018);
and U3311 (N_3311,In_1066,In_837);
nor U3312 (N_3312,In_78,In_1348);
xnor U3313 (N_3313,In_1371,In_549);
or U3314 (N_3314,In_1958,In_866);
and U3315 (N_3315,In_1578,In_1660);
nand U3316 (N_3316,In_2495,In_933);
nor U3317 (N_3317,In_1323,In_346);
xor U3318 (N_3318,In_2118,In_825);
nand U3319 (N_3319,In_1300,In_281);
and U3320 (N_3320,In_1896,In_2467);
nand U3321 (N_3321,In_1206,In_1560);
or U3322 (N_3322,In_614,In_307);
nand U3323 (N_3323,In_1537,In_2471);
nor U3324 (N_3324,In_1568,In_629);
nor U3325 (N_3325,In_1539,In_2422);
xnor U3326 (N_3326,In_2156,In_1104);
nor U3327 (N_3327,In_1369,In_381);
nand U3328 (N_3328,In_2367,In_2010);
xor U3329 (N_3329,In_2327,In_551);
nor U3330 (N_3330,In_1910,In_1790);
or U3331 (N_3331,In_832,In_711);
nand U3332 (N_3332,In_2289,In_1483);
and U3333 (N_3333,In_813,In_626);
nor U3334 (N_3334,In_1021,In_1101);
nand U3335 (N_3335,In_2484,In_311);
or U3336 (N_3336,In_891,In_2275);
and U3337 (N_3337,In_692,In_1595);
nor U3338 (N_3338,In_680,In_1229);
or U3339 (N_3339,In_1681,In_1734);
nor U3340 (N_3340,In_299,In_88);
xor U3341 (N_3341,In_771,In_2019);
and U3342 (N_3342,In_1533,In_937);
nor U3343 (N_3343,In_1728,In_1949);
xor U3344 (N_3344,In_837,In_966);
nand U3345 (N_3345,In_1164,In_1433);
and U3346 (N_3346,In_1109,In_499);
and U3347 (N_3347,In_1462,In_1991);
nor U3348 (N_3348,In_604,In_1904);
and U3349 (N_3349,In_1729,In_522);
or U3350 (N_3350,In_1365,In_1887);
nor U3351 (N_3351,In_1733,In_273);
nand U3352 (N_3352,In_1503,In_2474);
nor U3353 (N_3353,In_265,In_1003);
nand U3354 (N_3354,In_2199,In_2201);
nor U3355 (N_3355,In_1270,In_1192);
xor U3356 (N_3356,In_126,In_981);
and U3357 (N_3357,In_1956,In_548);
nand U3358 (N_3358,In_1485,In_346);
nand U3359 (N_3359,In_2124,In_1111);
and U3360 (N_3360,In_724,In_2233);
or U3361 (N_3361,In_1236,In_561);
or U3362 (N_3362,In_1224,In_721);
nor U3363 (N_3363,In_413,In_54);
xor U3364 (N_3364,In_1534,In_269);
and U3365 (N_3365,In_1827,In_1523);
nor U3366 (N_3366,In_1802,In_1276);
and U3367 (N_3367,In_801,In_2335);
and U3368 (N_3368,In_1662,In_1241);
nand U3369 (N_3369,In_1426,In_727);
or U3370 (N_3370,In_1797,In_1416);
xnor U3371 (N_3371,In_1888,In_1348);
and U3372 (N_3372,In_2198,In_783);
nor U3373 (N_3373,In_2227,In_1776);
or U3374 (N_3374,In_293,In_780);
nor U3375 (N_3375,In_262,In_759);
nand U3376 (N_3376,In_44,In_441);
nor U3377 (N_3377,In_86,In_245);
or U3378 (N_3378,In_1627,In_1034);
nor U3379 (N_3379,In_1222,In_1760);
nor U3380 (N_3380,In_1347,In_1901);
and U3381 (N_3381,In_1742,In_486);
nor U3382 (N_3382,In_655,In_626);
nand U3383 (N_3383,In_1012,In_858);
nand U3384 (N_3384,In_1651,In_778);
or U3385 (N_3385,In_322,In_1914);
and U3386 (N_3386,In_47,In_1134);
or U3387 (N_3387,In_892,In_131);
or U3388 (N_3388,In_1307,In_1457);
and U3389 (N_3389,In_10,In_837);
nor U3390 (N_3390,In_533,In_1315);
and U3391 (N_3391,In_2424,In_1820);
nor U3392 (N_3392,In_1114,In_1826);
and U3393 (N_3393,In_1338,In_1380);
and U3394 (N_3394,In_911,In_820);
nand U3395 (N_3395,In_943,In_1619);
nor U3396 (N_3396,In_547,In_2131);
nor U3397 (N_3397,In_2413,In_1511);
and U3398 (N_3398,In_1532,In_957);
or U3399 (N_3399,In_2313,In_1046);
and U3400 (N_3400,In_178,In_406);
and U3401 (N_3401,In_1467,In_1154);
xnor U3402 (N_3402,In_144,In_129);
nor U3403 (N_3403,In_1474,In_1699);
nor U3404 (N_3404,In_533,In_781);
nor U3405 (N_3405,In_2091,In_2163);
or U3406 (N_3406,In_2221,In_1821);
nor U3407 (N_3407,In_1468,In_1986);
xor U3408 (N_3408,In_1726,In_362);
and U3409 (N_3409,In_227,In_1698);
nand U3410 (N_3410,In_149,In_2076);
nor U3411 (N_3411,In_1926,In_484);
and U3412 (N_3412,In_135,In_80);
nor U3413 (N_3413,In_405,In_2081);
and U3414 (N_3414,In_174,In_245);
nor U3415 (N_3415,In_1911,In_9);
and U3416 (N_3416,In_1138,In_645);
or U3417 (N_3417,In_1999,In_2095);
nand U3418 (N_3418,In_747,In_517);
nand U3419 (N_3419,In_534,In_1676);
and U3420 (N_3420,In_2062,In_2499);
xnor U3421 (N_3421,In_1824,In_1144);
and U3422 (N_3422,In_141,In_1512);
nor U3423 (N_3423,In_1381,In_547);
nand U3424 (N_3424,In_330,In_1246);
or U3425 (N_3425,In_654,In_151);
nand U3426 (N_3426,In_392,In_856);
nand U3427 (N_3427,In_1823,In_2445);
nor U3428 (N_3428,In_198,In_941);
or U3429 (N_3429,In_1451,In_50);
xor U3430 (N_3430,In_796,In_2233);
nand U3431 (N_3431,In_287,In_917);
xnor U3432 (N_3432,In_1426,In_435);
xor U3433 (N_3433,In_321,In_2035);
nand U3434 (N_3434,In_1247,In_979);
nand U3435 (N_3435,In_706,In_1857);
or U3436 (N_3436,In_1014,In_2315);
or U3437 (N_3437,In_1220,In_668);
xor U3438 (N_3438,In_1332,In_1217);
xor U3439 (N_3439,In_1825,In_1257);
and U3440 (N_3440,In_1159,In_290);
nor U3441 (N_3441,In_853,In_2492);
nand U3442 (N_3442,In_848,In_1920);
nor U3443 (N_3443,In_1715,In_791);
or U3444 (N_3444,In_744,In_1641);
and U3445 (N_3445,In_1266,In_301);
nand U3446 (N_3446,In_2398,In_643);
nand U3447 (N_3447,In_853,In_1108);
nand U3448 (N_3448,In_2242,In_426);
nand U3449 (N_3449,In_1681,In_412);
or U3450 (N_3450,In_971,In_1015);
nand U3451 (N_3451,In_906,In_1763);
or U3452 (N_3452,In_721,In_438);
xnor U3453 (N_3453,In_1475,In_1585);
and U3454 (N_3454,In_1021,In_2008);
nand U3455 (N_3455,In_730,In_2409);
and U3456 (N_3456,In_838,In_1196);
or U3457 (N_3457,In_1293,In_852);
nor U3458 (N_3458,In_1960,In_2046);
nor U3459 (N_3459,In_1020,In_1820);
nor U3460 (N_3460,In_97,In_1786);
nor U3461 (N_3461,In_1018,In_412);
or U3462 (N_3462,In_782,In_1303);
or U3463 (N_3463,In_920,In_1448);
nand U3464 (N_3464,In_1568,In_929);
or U3465 (N_3465,In_1162,In_778);
and U3466 (N_3466,In_1197,In_1321);
nand U3467 (N_3467,In_2364,In_2386);
xnor U3468 (N_3468,In_264,In_502);
nor U3469 (N_3469,In_1089,In_1845);
and U3470 (N_3470,In_2222,In_1215);
and U3471 (N_3471,In_611,In_1574);
and U3472 (N_3472,In_637,In_583);
and U3473 (N_3473,In_2306,In_2325);
nand U3474 (N_3474,In_2153,In_1780);
nor U3475 (N_3475,In_944,In_1415);
nand U3476 (N_3476,In_2268,In_1970);
or U3477 (N_3477,In_260,In_279);
nor U3478 (N_3478,In_560,In_2124);
or U3479 (N_3479,In_2492,In_170);
and U3480 (N_3480,In_284,In_471);
xor U3481 (N_3481,In_2424,In_1406);
nor U3482 (N_3482,In_2110,In_301);
nand U3483 (N_3483,In_1604,In_2295);
nand U3484 (N_3484,In_163,In_2448);
nand U3485 (N_3485,In_66,In_2200);
or U3486 (N_3486,In_609,In_1330);
or U3487 (N_3487,In_182,In_1241);
or U3488 (N_3488,In_5,In_2441);
or U3489 (N_3489,In_1506,In_2013);
and U3490 (N_3490,In_2344,In_386);
and U3491 (N_3491,In_1719,In_786);
and U3492 (N_3492,In_793,In_2114);
and U3493 (N_3493,In_700,In_371);
nor U3494 (N_3494,In_212,In_2429);
nand U3495 (N_3495,In_539,In_699);
or U3496 (N_3496,In_763,In_942);
nand U3497 (N_3497,In_1613,In_1132);
or U3498 (N_3498,In_2054,In_1726);
nor U3499 (N_3499,In_122,In_604);
xnor U3500 (N_3500,In_621,In_1089);
and U3501 (N_3501,In_1741,In_43);
or U3502 (N_3502,In_1354,In_2441);
or U3503 (N_3503,In_98,In_2400);
or U3504 (N_3504,In_1376,In_2388);
nand U3505 (N_3505,In_165,In_1199);
and U3506 (N_3506,In_540,In_1822);
nand U3507 (N_3507,In_873,In_2217);
nand U3508 (N_3508,In_2296,In_1729);
or U3509 (N_3509,In_1567,In_2075);
nor U3510 (N_3510,In_1475,In_469);
nand U3511 (N_3511,In_1959,In_457);
and U3512 (N_3512,In_461,In_2193);
xor U3513 (N_3513,In_1072,In_14);
or U3514 (N_3514,In_1391,In_63);
and U3515 (N_3515,In_536,In_1315);
and U3516 (N_3516,In_1050,In_347);
and U3517 (N_3517,In_2299,In_1118);
and U3518 (N_3518,In_1534,In_1406);
or U3519 (N_3519,In_1798,In_323);
and U3520 (N_3520,In_2252,In_1238);
or U3521 (N_3521,In_1684,In_2116);
nor U3522 (N_3522,In_2014,In_926);
and U3523 (N_3523,In_35,In_2154);
or U3524 (N_3524,In_1085,In_78);
nor U3525 (N_3525,In_2004,In_737);
and U3526 (N_3526,In_296,In_2016);
xor U3527 (N_3527,In_1152,In_1374);
nand U3528 (N_3528,In_1260,In_1500);
nand U3529 (N_3529,In_1230,In_817);
or U3530 (N_3530,In_1723,In_1734);
or U3531 (N_3531,In_362,In_2459);
nand U3532 (N_3532,In_1779,In_2406);
xor U3533 (N_3533,In_1667,In_114);
or U3534 (N_3534,In_925,In_485);
or U3535 (N_3535,In_1308,In_389);
or U3536 (N_3536,In_1397,In_130);
and U3537 (N_3537,In_624,In_699);
nand U3538 (N_3538,In_1831,In_1981);
or U3539 (N_3539,In_2222,In_65);
or U3540 (N_3540,In_1281,In_2397);
nand U3541 (N_3541,In_779,In_235);
nor U3542 (N_3542,In_689,In_987);
xor U3543 (N_3543,In_1878,In_2125);
and U3544 (N_3544,In_1130,In_931);
nor U3545 (N_3545,In_1941,In_117);
nor U3546 (N_3546,In_1266,In_2165);
or U3547 (N_3547,In_2080,In_2139);
nand U3548 (N_3548,In_1969,In_994);
nor U3549 (N_3549,In_138,In_1040);
nor U3550 (N_3550,In_545,In_793);
xnor U3551 (N_3551,In_1575,In_133);
nand U3552 (N_3552,In_2006,In_1306);
nand U3553 (N_3553,In_309,In_1101);
nor U3554 (N_3554,In_1923,In_550);
nand U3555 (N_3555,In_800,In_1403);
or U3556 (N_3556,In_1930,In_1849);
nor U3557 (N_3557,In_2316,In_1805);
or U3558 (N_3558,In_2316,In_1861);
xnor U3559 (N_3559,In_1214,In_109);
or U3560 (N_3560,In_2116,In_1637);
xnor U3561 (N_3561,In_783,In_1084);
xor U3562 (N_3562,In_1629,In_2423);
and U3563 (N_3563,In_575,In_2431);
or U3564 (N_3564,In_2340,In_703);
nand U3565 (N_3565,In_543,In_293);
nand U3566 (N_3566,In_1122,In_930);
or U3567 (N_3567,In_1386,In_1226);
nand U3568 (N_3568,In_2068,In_2200);
and U3569 (N_3569,In_48,In_1697);
or U3570 (N_3570,In_663,In_531);
nor U3571 (N_3571,In_1231,In_2174);
xnor U3572 (N_3572,In_2188,In_2171);
or U3573 (N_3573,In_895,In_1571);
or U3574 (N_3574,In_1942,In_190);
and U3575 (N_3575,In_2095,In_1263);
xnor U3576 (N_3576,In_938,In_1746);
or U3577 (N_3577,In_1930,In_519);
xor U3578 (N_3578,In_1564,In_1055);
nor U3579 (N_3579,In_1302,In_2321);
nor U3580 (N_3580,In_284,In_2371);
or U3581 (N_3581,In_2427,In_1485);
nor U3582 (N_3582,In_734,In_166);
nand U3583 (N_3583,In_2101,In_2265);
and U3584 (N_3584,In_1324,In_2245);
nor U3585 (N_3585,In_844,In_183);
and U3586 (N_3586,In_1904,In_2109);
xor U3587 (N_3587,In_392,In_2145);
or U3588 (N_3588,In_50,In_1670);
nor U3589 (N_3589,In_2113,In_1917);
nand U3590 (N_3590,In_2088,In_1102);
and U3591 (N_3591,In_1628,In_155);
nand U3592 (N_3592,In_1492,In_1555);
or U3593 (N_3593,In_425,In_1241);
and U3594 (N_3594,In_567,In_777);
or U3595 (N_3595,In_600,In_1198);
or U3596 (N_3596,In_1833,In_2078);
or U3597 (N_3597,In_2049,In_206);
nand U3598 (N_3598,In_717,In_142);
or U3599 (N_3599,In_1809,In_1076);
nand U3600 (N_3600,In_694,In_632);
or U3601 (N_3601,In_520,In_1355);
nor U3602 (N_3602,In_250,In_1137);
and U3603 (N_3603,In_743,In_2029);
xnor U3604 (N_3604,In_683,In_1489);
xor U3605 (N_3605,In_1701,In_919);
nand U3606 (N_3606,In_717,In_117);
nor U3607 (N_3607,In_1331,In_1891);
or U3608 (N_3608,In_1176,In_1444);
nand U3609 (N_3609,In_1109,In_572);
nand U3610 (N_3610,In_1109,In_975);
or U3611 (N_3611,In_2292,In_1922);
nor U3612 (N_3612,In_1148,In_729);
or U3613 (N_3613,In_980,In_695);
or U3614 (N_3614,In_147,In_1309);
nand U3615 (N_3615,In_861,In_262);
and U3616 (N_3616,In_1259,In_2250);
and U3617 (N_3617,In_1914,In_2416);
nand U3618 (N_3618,In_158,In_463);
nand U3619 (N_3619,In_278,In_1281);
nor U3620 (N_3620,In_1717,In_1481);
and U3621 (N_3621,In_1548,In_793);
nor U3622 (N_3622,In_906,In_1229);
nor U3623 (N_3623,In_1920,In_709);
or U3624 (N_3624,In_91,In_1713);
or U3625 (N_3625,In_998,In_189);
nand U3626 (N_3626,In_728,In_421);
and U3627 (N_3627,In_709,In_692);
xnor U3628 (N_3628,In_1852,In_1467);
and U3629 (N_3629,In_892,In_886);
or U3630 (N_3630,In_649,In_1202);
and U3631 (N_3631,In_92,In_1899);
xnor U3632 (N_3632,In_2087,In_1221);
or U3633 (N_3633,In_2068,In_2100);
nand U3634 (N_3634,In_293,In_342);
and U3635 (N_3635,In_553,In_1689);
and U3636 (N_3636,In_2490,In_583);
and U3637 (N_3637,In_2471,In_1086);
or U3638 (N_3638,In_1434,In_125);
xnor U3639 (N_3639,In_1412,In_1308);
or U3640 (N_3640,In_2189,In_673);
or U3641 (N_3641,In_2150,In_1484);
nand U3642 (N_3642,In_2080,In_446);
nor U3643 (N_3643,In_715,In_1137);
nor U3644 (N_3644,In_1484,In_2222);
or U3645 (N_3645,In_1080,In_1790);
nor U3646 (N_3646,In_2152,In_2307);
or U3647 (N_3647,In_402,In_846);
and U3648 (N_3648,In_2363,In_1880);
nor U3649 (N_3649,In_1951,In_615);
or U3650 (N_3650,In_1374,In_1196);
nor U3651 (N_3651,In_595,In_886);
nand U3652 (N_3652,In_1456,In_1032);
nand U3653 (N_3653,In_252,In_1477);
xnor U3654 (N_3654,In_459,In_1788);
nor U3655 (N_3655,In_596,In_1186);
nor U3656 (N_3656,In_1306,In_1262);
or U3657 (N_3657,In_1231,In_1028);
and U3658 (N_3658,In_1953,In_761);
nand U3659 (N_3659,In_1228,In_1935);
nor U3660 (N_3660,In_1353,In_44);
and U3661 (N_3661,In_1845,In_273);
nor U3662 (N_3662,In_2104,In_1131);
nor U3663 (N_3663,In_712,In_1710);
or U3664 (N_3664,In_881,In_260);
and U3665 (N_3665,In_2152,In_2221);
nand U3666 (N_3666,In_489,In_989);
and U3667 (N_3667,In_754,In_679);
nor U3668 (N_3668,In_393,In_1784);
and U3669 (N_3669,In_164,In_1174);
nor U3670 (N_3670,In_1416,In_1433);
and U3671 (N_3671,In_1111,In_422);
and U3672 (N_3672,In_2265,In_2349);
nand U3673 (N_3673,In_2139,In_2470);
or U3674 (N_3674,In_1094,In_1447);
or U3675 (N_3675,In_2245,In_1884);
or U3676 (N_3676,In_215,In_1765);
and U3677 (N_3677,In_1923,In_306);
nand U3678 (N_3678,In_385,In_2015);
nand U3679 (N_3679,In_2133,In_666);
or U3680 (N_3680,In_1576,In_762);
xnor U3681 (N_3681,In_1111,In_1145);
nor U3682 (N_3682,In_1760,In_2214);
nor U3683 (N_3683,In_1815,In_1504);
xor U3684 (N_3684,In_2058,In_1858);
and U3685 (N_3685,In_809,In_1121);
and U3686 (N_3686,In_2387,In_982);
nor U3687 (N_3687,In_2326,In_329);
nand U3688 (N_3688,In_517,In_865);
and U3689 (N_3689,In_1817,In_517);
and U3690 (N_3690,In_21,In_2135);
and U3691 (N_3691,In_1324,In_2290);
or U3692 (N_3692,In_76,In_1304);
nor U3693 (N_3693,In_2380,In_589);
nand U3694 (N_3694,In_878,In_974);
and U3695 (N_3695,In_330,In_1771);
and U3696 (N_3696,In_578,In_280);
nand U3697 (N_3697,In_1471,In_471);
and U3698 (N_3698,In_2354,In_1304);
and U3699 (N_3699,In_2022,In_524);
nand U3700 (N_3700,In_1880,In_328);
nand U3701 (N_3701,In_1148,In_1961);
nor U3702 (N_3702,In_2327,In_397);
and U3703 (N_3703,In_1564,In_903);
and U3704 (N_3704,In_248,In_180);
xor U3705 (N_3705,In_223,In_1500);
or U3706 (N_3706,In_1198,In_1911);
and U3707 (N_3707,In_2378,In_1582);
nand U3708 (N_3708,In_442,In_2013);
or U3709 (N_3709,In_1810,In_510);
and U3710 (N_3710,In_1135,In_915);
and U3711 (N_3711,In_1528,In_1698);
and U3712 (N_3712,In_2238,In_974);
xor U3713 (N_3713,In_1247,In_1693);
nor U3714 (N_3714,In_1604,In_625);
and U3715 (N_3715,In_2350,In_649);
nand U3716 (N_3716,In_2489,In_2148);
and U3717 (N_3717,In_485,In_1501);
nor U3718 (N_3718,In_89,In_1343);
nand U3719 (N_3719,In_1268,In_1059);
xnor U3720 (N_3720,In_1545,In_1343);
or U3721 (N_3721,In_1066,In_2206);
nand U3722 (N_3722,In_2009,In_88);
nand U3723 (N_3723,In_1693,In_363);
and U3724 (N_3724,In_515,In_2049);
xor U3725 (N_3725,In_4,In_1246);
nor U3726 (N_3726,In_1838,In_1193);
or U3727 (N_3727,In_2207,In_1651);
nor U3728 (N_3728,In_1968,In_1681);
nor U3729 (N_3729,In_2488,In_1128);
or U3730 (N_3730,In_803,In_859);
nand U3731 (N_3731,In_1704,In_24);
and U3732 (N_3732,In_732,In_215);
or U3733 (N_3733,In_2109,In_1334);
or U3734 (N_3734,In_1926,In_467);
and U3735 (N_3735,In_1966,In_1027);
nand U3736 (N_3736,In_1140,In_1551);
and U3737 (N_3737,In_166,In_1052);
nor U3738 (N_3738,In_774,In_2197);
or U3739 (N_3739,In_1390,In_1049);
nor U3740 (N_3740,In_1390,In_2347);
nor U3741 (N_3741,In_1378,In_56);
nor U3742 (N_3742,In_396,In_1178);
nand U3743 (N_3743,In_2250,In_1841);
and U3744 (N_3744,In_2066,In_228);
nor U3745 (N_3745,In_1529,In_1037);
nor U3746 (N_3746,In_1311,In_2133);
nand U3747 (N_3747,In_1784,In_748);
nor U3748 (N_3748,In_82,In_1919);
and U3749 (N_3749,In_1289,In_1855);
nor U3750 (N_3750,In_636,In_1312);
and U3751 (N_3751,In_2319,In_1188);
and U3752 (N_3752,In_1774,In_1877);
nand U3753 (N_3753,In_863,In_11);
and U3754 (N_3754,In_806,In_441);
nor U3755 (N_3755,In_220,In_1616);
and U3756 (N_3756,In_80,In_1011);
nor U3757 (N_3757,In_1184,In_90);
xnor U3758 (N_3758,In_526,In_1390);
nand U3759 (N_3759,In_1528,In_1434);
or U3760 (N_3760,In_1109,In_323);
nand U3761 (N_3761,In_2179,In_1004);
or U3762 (N_3762,In_951,In_1054);
nand U3763 (N_3763,In_688,In_1428);
nand U3764 (N_3764,In_1739,In_2378);
nor U3765 (N_3765,In_561,In_364);
nand U3766 (N_3766,In_1590,In_1279);
nor U3767 (N_3767,In_562,In_206);
or U3768 (N_3768,In_1766,In_696);
and U3769 (N_3769,In_1788,In_816);
or U3770 (N_3770,In_2163,In_1483);
and U3771 (N_3771,In_1561,In_2384);
and U3772 (N_3772,In_679,In_2168);
nor U3773 (N_3773,In_417,In_2492);
and U3774 (N_3774,In_1217,In_319);
nand U3775 (N_3775,In_2491,In_337);
and U3776 (N_3776,In_892,In_979);
or U3777 (N_3777,In_1130,In_2203);
and U3778 (N_3778,In_1601,In_285);
and U3779 (N_3779,In_1044,In_1493);
and U3780 (N_3780,In_1841,In_406);
nand U3781 (N_3781,In_1827,In_302);
or U3782 (N_3782,In_231,In_47);
or U3783 (N_3783,In_2247,In_1194);
or U3784 (N_3784,In_66,In_2155);
and U3785 (N_3785,In_905,In_182);
or U3786 (N_3786,In_2248,In_2114);
nor U3787 (N_3787,In_245,In_54);
and U3788 (N_3788,In_1781,In_963);
nor U3789 (N_3789,In_926,In_709);
nor U3790 (N_3790,In_1092,In_1407);
and U3791 (N_3791,In_252,In_2354);
and U3792 (N_3792,In_1289,In_245);
xor U3793 (N_3793,In_2056,In_768);
or U3794 (N_3794,In_581,In_700);
and U3795 (N_3795,In_305,In_1181);
nor U3796 (N_3796,In_840,In_2279);
xnor U3797 (N_3797,In_1626,In_992);
and U3798 (N_3798,In_482,In_2469);
or U3799 (N_3799,In_1880,In_2462);
nor U3800 (N_3800,In_990,In_992);
nor U3801 (N_3801,In_1708,In_1376);
nor U3802 (N_3802,In_1435,In_1799);
xnor U3803 (N_3803,In_996,In_2058);
nand U3804 (N_3804,In_2262,In_1474);
nor U3805 (N_3805,In_1916,In_547);
nand U3806 (N_3806,In_1760,In_833);
and U3807 (N_3807,In_2028,In_14);
or U3808 (N_3808,In_96,In_1593);
nand U3809 (N_3809,In_1740,In_257);
or U3810 (N_3810,In_574,In_137);
nor U3811 (N_3811,In_115,In_99);
nand U3812 (N_3812,In_959,In_610);
and U3813 (N_3813,In_632,In_2375);
xnor U3814 (N_3814,In_555,In_2433);
nor U3815 (N_3815,In_1396,In_1757);
and U3816 (N_3816,In_766,In_1089);
nor U3817 (N_3817,In_1987,In_789);
or U3818 (N_3818,In_266,In_555);
nor U3819 (N_3819,In_2291,In_2290);
nor U3820 (N_3820,In_2150,In_1244);
xnor U3821 (N_3821,In_2438,In_1923);
nor U3822 (N_3822,In_337,In_619);
nand U3823 (N_3823,In_436,In_2075);
and U3824 (N_3824,In_478,In_1148);
or U3825 (N_3825,In_1190,In_1054);
nor U3826 (N_3826,In_1869,In_784);
nand U3827 (N_3827,In_2183,In_1374);
and U3828 (N_3828,In_1203,In_391);
nand U3829 (N_3829,In_635,In_783);
and U3830 (N_3830,In_294,In_257);
or U3831 (N_3831,In_985,In_148);
and U3832 (N_3832,In_830,In_1772);
xnor U3833 (N_3833,In_1480,In_797);
nand U3834 (N_3834,In_315,In_16);
xor U3835 (N_3835,In_192,In_1680);
nor U3836 (N_3836,In_1923,In_179);
nand U3837 (N_3837,In_2355,In_2150);
and U3838 (N_3838,In_1361,In_1457);
or U3839 (N_3839,In_1836,In_240);
or U3840 (N_3840,In_2149,In_1033);
or U3841 (N_3841,In_260,In_1918);
or U3842 (N_3842,In_1326,In_1105);
or U3843 (N_3843,In_476,In_819);
nand U3844 (N_3844,In_1849,In_1814);
or U3845 (N_3845,In_553,In_113);
or U3846 (N_3846,In_1310,In_1092);
nor U3847 (N_3847,In_2355,In_2064);
xor U3848 (N_3848,In_1927,In_36);
nor U3849 (N_3849,In_1607,In_868);
and U3850 (N_3850,In_870,In_444);
and U3851 (N_3851,In_2352,In_1289);
xnor U3852 (N_3852,In_1526,In_1521);
and U3853 (N_3853,In_1465,In_708);
and U3854 (N_3854,In_2133,In_1194);
xnor U3855 (N_3855,In_376,In_2271);
nand U3856 (N_3856,In_1982,In_2466);
nand U3857 (N_3857,In_166,In_14);
nor U3858 (N_3858,In_2430,In_1656);
nor U3859 (N_3859,In_849,In_322);
nand U3860 (N_3860,In_2086,In_143);
or U3861 (N_3861,In_1578,In_716);
nand U3862 (N_3862,In_286,In_1492);
nor U3863 (N_3863,In_1553,In_2218);
xor U3864 (N_3864,In_991,In_678);
and U3865 (N_3865,In_1989,In_1587);
or U3866 (N_3866,In_2301,In_2239);
nor U3867 (N_3867,In_2462,In_1889);
nand U3868 (N_3868,In_1142,In_821);
xnor U3869 (N_3869,In_1494,In_708);
or U3870 (N_3870,In_719,In_500);
and U3871 (N_3871,In_1192,In_2337);
or U3872 (N_3872,In_1804,In_253);
nor U3873 (N_3873,In_1351,In_1281);
nand U3874 (N_3874,In_1995,In_793);
nor U3875 (N_3875,In_1586,In_950);
and U3876 (N_3876,In_1249,In_504);
or U3877 (N_3877,In_1017,In_586);
and U3878 (N_3878,In_432,In_480);
xnor U3879 (N_3879,In_1788,In_2236);
nor U3880 (N_3880,In_591,In_781);
nor U3881 (N_3881,In_486,In_142);
nand U3882 (N_3882,In_1870,In_2173);
and U3883 (N_3883,In_2390,In_1769);
or U3884 (N_3884,In_222,In_1789);
and U3885 (N_3885,In_833,In_857);
and U3886 (N_3886,In_1481,In_1272);
nor U3887 (N_3887,In_2096,In_346);
and U3888 (N_3888,In_524,In_1488);
and U3889 (N_3889,In_295,In_1474);
nor U3890 (N_3890,In_1571,In_82);
nand U3891 (N_3891,In_1329,In_799);
nand U3892 (N_3892,In_2012,In_650);
or U3893 (N_3893,In_672,In_749);
or U3894 (N_3894,In_1887,In_481);
or U3895 (N_3895,In_827,In_1637);
nor U3896 (N_3896,In_2378,In_2258);
xnor U3897 (N_3897,In_213,In_728);
or U3898 (N_3898,In_36,In_745);
nand U3899 (N_3899,In_2483,In_1423);
nand U3900 (N_3900,In_115,In_319);
and U3901 (N_3901,In_1044,In_944);
nor U3902 (N_3902,In_2197,In_54);
xor U3903 (N_3903,In_614,In_277);
xnor U3904 (N_3904,In_582,In_1702);
or U3905 (N_3905,In_863,In_664);
nor U3906 (N_3906,In_442,In_1011);
nand U3907 (N_3907,In_404,In_460);
and U3908 (N_3908,In_696,In_1399);
and U3909 (N_3909,In_2291,In_1832);
nor U3910 (N_3910,In_50,In_1982);
xor U3911 (N_3911,In_394,In_965);
nor U3912 (N_3912,In_42,In_2028);
nor U3913 (N_3913,In_1653,In_1475);
or U3914 (N_3914,In_2360,In_743);
and U3915 (N_3915,In_763,In_45);
and U3916 (N_3916,In_2287,In_1777);
or U3917 (N_3917,In_747,In_1410);
and U3918 (N_3918,In_1914,In_1433);
and U3919 (N_3919,In_1678,In_1508);
nand U3920 (N_3920,In_772,In_2306);
nand U3921 (N_3921,In_1619,In_1813);
or U3922 (N_3922,In_677,In_1167);
xor U3923 (N_3923,In_140,In_1456);
nand U3924 (N_3924,In_34,In_379);
nand U3925 (N_3925,In_964,In_998);
nand U3926 (N_3926,In_2330,In_364);
xor U3927 (N_3927,In_1843,In_1039);
and U3928 (N_3928,In_4,In_485);
and U3929 (N_3929,In_1773,In_147);
and U3930 (N_3930,In_1898,In_728);
or U3931 (N_3931,In_2473,In_1991);
or U3932 (N_3932,In_685,In_1445);
and U3933 (N_3933,In_2018,In_1023);
and U3934 (N_3934,In_211,In_1886);
or U3935 (N_3935,In_429,In_877);
nand U3936 (N_3936,In_894,In_1208);
or U3937 (N_3937,In_249,In_1273);
and U3938 (N_3938,In_2456,In_564);
and U3939 (N_3939,In_2176,In_163);
or U3940 (N_3940,In_1724,In_2215);
and U3941 (N_3941,In_2228,In_262);
nor U3942 (N_3942,In_2108,In_1476);
nand U3943 (N_3943,In_2425,In_2495);
nor U3944 (N_3944,In_16,In_293);
nor U3945 (N_3945,In_346,In_1722);
nor U3946 (N_3946,In_428,In_1081);
or U3947 (N_3947,In_2371,In_1979);
xor U3948 (N_3948,In_2486,In_1326);
and U3949 (N_3949,In_1822,In_630);
or U3950 (N_3950,In_1389,In_1235);
or U3951 (N_3951,In_1620,In_1246);
and U3952 (N_3952,In_1469,In_2280);
or U3953 (N_3953,In_1554,In_1489);
or U3954 (N_3954,In_459,In_77);
nand U3955 (N_3955,In_744,In_2336);
xnor U3956 (N_3956,In_1978,In_683);
or U3957 (N_3957,In_970,In_1755);
or U3958 (N_3958,In_752,In_946);
or U3959 (N_3959,In_836,In_298);
nand U3960 (N_3960,In_1206,In_1114);
nor U3961 (N_3961,In_2111,In_1618);
xor U3962 (N_3962,In_1195,In_1153);
or U3963 (N_3963,In_433,In_744);
and U3964 (N_3964,In_1041,In_381);
nand U3965 (N_3965,In_1297,In_854);
or U3966 (N_3966,In_762,In_2037);
nor U3967 (N_3967,In_495,In_1080);
nand U3968 (N_3968,In_679,In_2498);
nor U3969 (N_3969,In_106,In_494);
nand U3970 (N_3970,In_70,In_2101);
nand U3971 (N_3971,In_567,In_1830);
nor U3972 (N_3972,In_736,In_218);
nor U3973 (N_3973,In_2171,In_2174);
and U3974 (N_3974,In_1508,In_493);
and U3975 (N_3975,In_808,In_2013);
or U3976 (N_3976,In_306,In_1844);
nand U3977 (N_3977,In_1949,In_2357);
nor U3978 (N_3978,In_312,In_316);
or U3979 (N_3979,In_36,In_1797);
xor U3980 (N_3980,In_1944,In_2288);
and U3981 (N_3981,In_1880,In_2005);
and U3982 (N_3982,In_564,In_2219);
nor U3983 (N_3983,In_641,In_2182);
xnor U3984 (N_3984,In_631,In_2398);
and U3985 (N_3985,In_1059,In_79);
nand U3986 (N_3986,In_2078,In_1982);
nor U3987 (N_3987,In_2185,In_1140);
nor U3988 (N_3988,In_2372,In_959);
nand U3989 (N_3989,In_2088,In_1056);
or U3990 (N_3990,In_2336,In_1738);
and U3991 (N_3991,In_826,In_2227);
nor U3992 (N_3992,In_740,In_1894);
or U3993 (N_3993,In_2078,In_1091);
and U3994 (N_3994,In_961,In_101);
nand U3995 (N_3995,In_1632,In_2489);
nor U3996 (N_3996,In_930,In_1982);
nand U3997 (N_3997,In_717,In_580);
or U3998 (N_3998,In_398,In_1778);
or U3999 (N_3999,In_1505,In_2036);
or U4000 (N_4000,In_1582,In_304);
and U4001 (N_4001,In_1095,In_1942);
and U4002 (N_4002,In_1548,In_217);
and U4003 (N_4003,In_1242,In_29);
xnor U4004 (N_4004,In_2192,In_101);
nand U4005 (N_4005,In_1458,In_2283);
nand U4006 (N_4006,In_509,In_858);
or U4007 (N_4007,In_2224,In_1969);
nor U4008 (N_4008,In_220,In_768);
nand U4009 (N_4009,In_2148,In_138);
or U4010 (N_4010,In_1225,In_2461);
nor U4011 (N_4011,In_1351,In_956);
or U4012 (N_4012,In_281,In_1073);
nand U4013 (N_4013,In_712,In_2489);
nand U4014 (N_4014,In_2481,In_667);
and U4015 (N_4015,In_2138,In_803);
xnor U4016 (N_4016,In_2114,In_810);
and U4017 (N_4017,In_1898,In_1593);
and U4018 (N_4018,In_2281,In_2029);
and U4019 (N_4019,In_1168,In_690);
xnor U4020 (N_4020,In_1107,In_1540);
nand U4021 (N_4021,In_200,In_2090);
nor U4022 (N_4022,In_730,In_610);
or U4023 (N_4023,In_2351,In_1500);
or U4024 (N_4024,In_1804,In_555);
or U4025 (N_4025,In_1436,In_2302);
and U4026 (N_4026,In_2327,In_142);
or U4027 (N_4027,In_1606,In_382);
nand U4028 (N_4028,In_829,In_639);
nand U4029 (N_4029,In_1364,In_440);
nand U4030 (N_4030,In_397,In_653);
xnor U4031 (N_4031,In_119,In_2128);
and U4032 (N_4032,In_270,In_992);
nor U4033 (N_4033,In_418,In_316);
nor U4034 (N_4034,In_1495,In_1510);
or U4035 (N_4035,In_637,In_1307);
and U4036 (N_4036,In_2093,In_1329);
nor U4037 (N_4037,In_1588,In_1102);
nand U4038 (N_4038,In_892,In_1413);
or U4039 (N_4039,In_360,In_590);
and U4040 (N_4040,In_908,In_1951);
and U4041 (N_4041,In_1232,In_1900);
nor U4042 (N_4042,In_1970,In_890);
or U4043 (N_4043,In_932,In_1398);
and U4044 (N_4044,In_1444,In_635);
nand U4045 (N_4045,In_2380,In_366);
or U4046 (N_4046,In_1002,In_1345);
nand U4047 (N_4047,In_2149,In_23);
nor U4048 (N_4048,In_775,In_236);
nor U4049 (N_4049,In_1871,In_2196);
nor U4050 (N_4050,In_789,In_296);
nor U4051 (N_4051,In_1320,In_1291);
xor U4052 (N_4052,In_1734,In_977);
nand U4053 (N_4053,In_1975,In_1882);
and U4054 (N_4054,In_2433,In_1751);
or U4055 (N_4055,In_2470,In_1184);
nand U4056 (N_4056,In_345,In_572);
and U4057 (N_4057,In_2477,In_1177);
xnor U4058 (N_4058,In_1210,In_1381);
xor U4059 (N_4059,In_1130,In_2119);
nand U4060 (N_4060,In_1050,In_2047);
xor U4061 (N_4061,In_432,In_1845);
nand U4062 (N_4062,In_251,In_1048);
nand U4063 (N_4063,In_1956,In_2237);
and U4064 (N_4064,In_27,In_1629);
and U4065 (N_4065,In_670,In_2027);
xor U4066 (N_4066,In_2215,In_1728);
and U4067 (N_4067,In_2416,In_2046);
nand U4068 (N_4068,In_2239,In_2238);
xor U4069 (N_4069,In_500,In_1373);
nand U4070 (N_4070,In_868,In_19);
and U4071 (N_4071,In_1268,In_1310);
nand U4072 (N_4072,In_1339,In_356);
and U4073 (N_4073,In_1396,In_2341);
or U4074 (N_4074,In_1982,In_107);
nand U4075 (N_4075,In_1026,In_949);
and U4076 (N_4076,In_1404,In_1731);
nand U4077 (N_4077,In_2062,In_1523);
nor U4078 (N_4078,In_611,In_2203);
nand U4079 (N_4079,In_796,In_736);
or U4080 (N_4080,In_2170,In_2436);
xnor U4081 (N_4081,In_998,In_1778);
nand U4082 (N_4082,In_601,In_1229);
nor U4083 (N_4083,In_1671,In_64);
nor U4084 (N_4084,In_1993,In_102);
and U4085 (N_4085,In_2283,In_1717);
nand U4086 (N_4086,In_526,In_159);
xnor U4087 (N_4087,In_442,In_1631);
nand U4088 (N_4088,In_2408,In_176);
or U4089 (N_4089,In_2312,In_2314);
or U4090 (N_4090,In_916,In_2259);
nor U4091 (N_4091,In_648,In_827);
nand U4092 (N_4092,In_552,In_2346);
nand U4093 (N_4093,In_1440,In_540);
nand U4094 (N_4094,In_1216,In_1905);
nand U4095 (N_4095,In_488,In_413);
nor U4096 (N_4096,In_1428,In_492);
nand U4097 (N_4097,In_1573,In_2452);
nand U4098 (N_4098,In_1596,In_96);
or U4099 (N_4099,In_1371,In_2076);
and U4100 (N_4100,In_811,In_166);
or U4101 (N_4101,In_1578,In_209);
xor U4102 (N_4102,In_2233,In_69);
and U4103 (N_4103,In_1326,In_2237);
and U4104 (N_4104,In_797,In_1492);
and U4105 (N_4105,In_2154,In_735);
or U4106 (N_4106,In_1447,In_1397);
and U4107 (N_4107,In_1500,In_559);
nor U4108 (N_4108,In_2269,In_1369);
and U4109 (N_4109,In_675,In_509);
nand U4110 (N_4110,In_89,In_1445);
nand U4111 (N_4111,In_2016,In_1836);
xor U4112 (N_4112,In_1203,In_2418);
xnor U4113 (N_4113,In_959,In_1082);
and U4114 (N_4114,In_1708,In_2350);
nand U4115 (N_4115,In_1394,In_848);
or U4116 (N_4116,In_2356,In_1782);
or U4117 (N_4117,In_2489,In_2318);
nand U4118 (N_4118,In_1440,In_1252);
or U4119 (N_4119,In_2472,In_422);
or U4120 (N_4120,In_2441,In_56);
nor U4121 (N_4121,In_1719,In_1991);
and U4122 (N_4122,In_366,In_1938);
nand U4123 (N_4123,In_2053,In_1796);
and U4124 (N_4124,In_958,In_1025);
and U4125 (N_4125,In_2188,In_587);
and U4126 (N_4126,In_404,In_1973);
nor U4127 (N_4127,In_768,In_1625);
or U4128 (N_4128,In_1492,In_2037);
and U4129 (N_4129,In_683,In_2010);
nand U4130 (N_4130,In_630,In_1980);
and U4131 (N_4131,In_2188,In_1001);
and U4132 (N_4132,In_1135,In_1844);
and U4133 (N_4133,In_2261,In_994);
xor U4134 (N_4134,In_1861,In_1070);
nand U4135 (N_4135,In_2435,In_1222);
nand U4136 (N_4136,In_160,In_1260);
or U4137 (N_4137,In_1525,In_842);
nand U4138 (N_4138,In_415,In_1350);
nor U4139 (N_4139,In_2211,In_1951);
and U4140 (N_4140,In_1395,In_1097);
or U4141 (N_4141,In_2407,In_1989);
nor U4142 (N_4142,In_718,In_640);
xnor U4143 (N_4143,In_1558,In_1008);
nand U4144 (N_4144,In_2460,In_2214);
nor U4145 (N_4145,In_1277,In_1903);
xor U4146 (N_4146,In_439,In_1760);
xnor U4147 (N_4147,In_1712,In_1809);
or U4148 (N_4148,In_294,In_1090);
nor U4149 (N_4149,In_594,In_790);
nor U4150 (N_4150,In_2076,In_796);
xor U4151 (N_4151,In_2324,In_2062);
nand U4152 (N_4152,In_2368,In_1908);
and U4153 (N_4153,In_1842,In_711);
and U4154 (N_4154,In_2400,In_15);
or U4155 (N_4155,In_131,In_629);
nor U4156 (N_4156,In_1109,In_901);
xnor U4157 (N_4157,In_246,In_237);
nor U4158 (N_4158,In_2386,In_463);
nand U4159 (N_4159,In_1578,In_1738);
nand U4160 (N_4160,In_2384,In_1551);
and U4161 (N_4161,In_1805,In_1636);
xnor U4162 (N_4162,In_2314,In_331);
and U4163 (N_4163,In_1615,In_1532);
and U4164 (N_4164,In_581,In_1127);
nand U4165 (N_4165,In_77,In_359);
nand U4166 (N_4166,In_2120,In_2432);
nand U4167 (N_4167,In_137,In_922);
nor U4168 (N_4168,In_2062,In_30);
or U4169 (N_4169,In_2338,In_1853);
and U4170 (N_4170,In_2127,In_1349);
nand U4171 (N_4171,In_351,In_1965);
xor U4172 (N_4172,In_130,In_2436);
or U4173 (N_4173,In_304,In_1749);
or U4174 (N_4174,In_544,In_2216);
nand U4175 (N_4175,In_2168,In_854);
or U4176 (N_4176,In_1510,In_1054);
nand U4177 (N_4177,In_1248,In_1389);
nand U4178 (N_4178,In_1814,In_1696);
or U4179 (N_4179,In_1129,In_1639);
nand U4180 (N_4180,In_1678,In_1637);
or U4181 (N_4181,In_1286,In_2276);
or U4182 (N_4182,In_1221,In_1484);
and U4183 (N_4183,In_725,In_1802);
nor U4184 (N_4184,In_723,In_439);
and U4185 (N_4185,In_605,In_1986);
and U4186 (N_4186,In_1636,In_1448);
nand U4187 (N_4187,In_1059,In_215);
nand U4188 (N_4188,In_519,In_378);
and U4189 (N_4189,In_1083,In_1044);
and U4190 (N_4190,In_659,In_2088);
nor U4191 (N_4191,In_196,In_416);
nand U4192 (N_4192,In_189,In_2238);
or U4193 (N_4193,In_2263,In_1436);
and U4194 (N_4194,In_1474,In_1135);
nand U4195 (N_4195,In_344,In_522);
or U4196 (N_4196,In_2003,In_805);
nor U4197 (N_4197,In_819,In_353);
nor U4198 (N_4198,In_1498,In_2312);
and U4199 (N_4199,In_413,In_1422);
xor U4200 (N_4200,In_1268,In_2064);
or U4201 (N_4201,In_121,In_1723);
or U4202 (N_4202,In_1670,In_801);
or U4203 (N_4203,In_481,In_1274);
or U4204 (N_4204,In_1122,In_371);
nor U4205 (N_4205,In_1559,In_282);
or U4206 (N_4206,In_1372,In_478);
nand U4207 (N_4207,In_76,In_2174);
nand U4208 (N_4208,In_1345,In_1850);
xnor U4209 (N_4209,In_1707,In_1077);
or U4210 (N_4210,In_605,In_715);
nor U4211 (N_4211,In_2331,In_1493);
or U4212 (N_4212,In_1847,In_2099);
xor U4213 (N_4213,In_1173,In_1475);
nand U4214 (N_4214,In_1674,In_1749);
xor U4215 (N_4215,In_2475,In_280);
nor U4216 (N_4216,In_1295,In_684);
nor U4217 (N_4217,In_211,In_131);
xor U4218 (N_4218,In_190,In_1440);
and U4219 (N_4219,In_2156,In_2282);
xor U4220 (N_4220,In_2236,In_396);
or U4221 (N_4221,In_254,In_1755);
xor U4222 (N_4222,In_2314,In_2332);
nand U4223 (N_4223,In_1553,In_158);
nand U4224 (N_4224,In_1316,In_903);
and U4225 (N_4225,In_2312,In_1103);
nor U4226 (N_4226,In_2472,In_1234);
nand U4227 (N_4227,In_757,In_2209);
and U4228 (N_4228,In_2275,In_1650);
or U4229 (N_4229,In_1781,In_857);
or U4230 (N_4230,In_2340,In_666);
and U4231 (N_4231,In_584,In_1407);
nor U4232 (N_4232,In_836,In_2462);
and U4233 (N_4233,In_687,In_1807);
or U4234 (N_4234,In_2411,In_2309);
nand U4235 (N_4235,In_1508,In_1971);
or U4236 (N_4236,In_865,In_1858);
nand U4237 (N_4237,In_1759,In_938);
nor U4238 (N_4238,In_2138,In_1759);
or U4239 (N_4239,In_1259,In_321);
and U4240 (N_4240,In_380,In_102);
xnor U4241 (N_4241,In_1679,In_1500);
or U4242 (N_4242,In_907,In_2449);
xor U4243 (N_4243,In_569,In_2125);
and U4244 (N_4244,In_1571,In_2194);
nand U4245 (N_4245,In_954,In_645);
and U4246 (N_4246,In_127,In_447);
nor U4247 (N_4247,In_1519,In_2097);
xnor U4248 (N_4248,In_385,In_1659);
xnor U4249 (N_4249,In_2199,In_397);
nor U4250 (N_4250,In_1524,In_227);
and U4251 (N_4251,In_1880,In_545);
or U4252 (N_4252,In_2051,In_755);
or U4253 (N_4253,In_255,In_2351);
nor U4254 (N_4254,In_2439,In_2430);
or U4255 (N_4255,In_579,In_2443);
xor U4256 (N_4256,In_2233,In_1667);
nor U4257 (N_4257,In_540,In_2079);
and U4258 (N_4258,In_550,In_270);
nand U4259 (N_4259,In_2171,In_560);
and U4260 (N_4260,In_2158,In_1288);
nor U4261 (N_4261,In_937,In_1373);
nand U4262 (N_4262,In_1085,In_1928);
nor U4263 (N_4263,In_153,In_2115);
or U4264 (N_4264,In_1511,In_104);
and U4265 (N_4265,In_368,In_1537);
xor U4266 (N_4266,In_1613,In_746);
nand U4267 (N_4267,In_237,In_1600);
nor U4268 (N_4268,In_2373,In_241);
nor U4269 (N_4269,In_1612,In_2257);
nor U4270 (N_4270,In_458,In_2258);
nand U4271 (N_4271,In_1579,In_2268);
nand U4272 (N_4272,In_1722,In_2383);
and U4273 (N_4273,In_1138,In_1944);
nor U4274 (N_4274,In_2179,In_976);
and U4275 (N_4275,In_243,In_597);
and U4276 (N_4276,In_352,In_2408);
and U4277 (N_4277,In_2482,In_466);
and U4278 (N_4278,In_657,In_1826);
or U4279 (N_4279,In_1889,In_1879);
nand U4280 (N_4280,In_1745,In_1648);
xnor U4281 (N_4281,In_2391,In_2121);
nor U4282 (N_4282,In_1996,In_1050);
and U4283 (N_4283,In_2157,In_1045);
nand U4284 (N_4284,In_405,In_987);
nor U4285 (N_4285,In_2178,In_797);
or U4286 (N_4286,In_992,In_527);
or U4287 (N_4287,In_1436,In_1116);
nor U4288 (N_4288,In_1343,In_2195);
nor U4289 (N_4289,In_2004,In_343);
and U4290 (N_4290,In_1303,In_1812);
nor U4291 (N_4291,In_1660,In_2394);
nand U4292 (N_4292,In_2290,In_1831);
xor U4293 (N_4293,In_1952,In_2413);
and U4294 (N_4294,In_1263,In_1453);
nor U4295 (N_4295,In_141,In_2080);
or U4296 (N_4296,In_1038,In_2410);
nor U4297 (N_4297,In_1264,In_2265);
nor U4298 (N_4298,In_1814,In_2490);
or U4299 (N_4299,In_474,In_1294);
nand U4300 (N_4300,In_1883,In_1247);
or U4301 (N_4301,In_2093,In_90);
and U4302 (N_4302,In_2225,In_1153);
nand U4303 (N_4303,In_1041,In_1379);
or U4304 (N_4304,In_2267,In_901);
xor U4305 (N_4305,In_865,In_1336);
nand U4306 (N_4306,In_416,In_2171);
xor U4307 (N_4307,In_1978,In_47);
nand U4308 (N_4308,In_135,In_1950);
xor U4309 (N_4309,In_1462,In_2053);
nand U4310 (N_4310,In_3,In_138);
nor U4311 (N_4311,In_472,In_325);
nor U4312 (N_4312,In_281,In_774);
xnor U4313 (N_4313,In_1138,In_547);
nor U4314 (N_4314,In_180,In_2119);
nor U4315 (N_4315,In_1812,In_2185);
nor U4316 (N_4316,In_246,In_2464);
and U4317 (N_4317,In_232,In_1478);
nor U4318 (N_4318,In_1082,In_2017);
and U4319 (N_4319,In_67,In_1721);
nand U4320 (N_4320,In_648,In_108);
xnor U4321 (N_4321,In_1205,In_1589);
and U4322 (N_4322,In_2210,In_645);
and U4323 (N_4323,In_57,In_218);
xor U4324 (N_4324,In_1139,In_474);
or U4325 (N_4325,In_1338,In_577);
nor U4326 (N_4326,In_412,In_2085);
nor U4327 (N_4327,In_272,In_1043);
nand U4328 (N_4328,In_1949,In_1977);
nand U4329 (N_4329,In_31,In_688);
nor U4330 (N_4330,In_2019,In_2448);
nand U4331 (N_4331,In_2436,In_2409);
and U4332 (N_4332,In_1770,In_369);
xnor U4333 (N_4333,In_1994,In_2409);
nand U4334 (N_4334,In_292,In_525);
nand U4335 (N_4335,In_370,In_239);
and U4336 (N_4336,In_37,In_4);
nor U4337 (N_4337,In_968,In_2272);
and U4338 (N_4338,In_304,In_1713);
or U4339 (N_4339,In_1959,In_458);
or U4340 (N_4340,In_718,In_1125);
and U4341 (N_4341,In_1490,In_2002);
and U4342 (N_4342,In_2026,In_874);
nor U4343 (N_4343,In_2334,In_763);
or U4344 (N_4344,In_1708,In_2192);
or U4345 (N_4345,In_210,In_1666);
nor U4346 (N_4346,In_956,In_591);
nand U4347 (N_4347,In_612,In_2004);
nand U4348 (N_4348,In_2445,In_1757);
nor U4349 (N_4349,In_841,In_2155);
and U4350 (N_4350,In_2107,In_280);
nand U4351 (N_4351,In_1907,In_2158);
or U4352 (N_4352,In_410,In_2106);
or U4353 (N_4353,In_74,In_1284);
nor U4354 (N_4354,In_562,In_2111);
and U4355 (N_4355,In_773,In_847);
nor U4356 (N_4356,In_1356,In_1197);
nor U4357 (N_4357,In_799,In_1278);
xor U4358 (N_4358,In_2105,In_632);
nor U4359 (N_4359,In_579,In_2293);
nor U4360 (N_4360,In_1012,In_1990);
and U4361 (N_4361,In_1373,In_251);
and U4362 (N_4362,In_1569,In_540);
or U4363 (N_4363,In_401,In_2442);
and U4364 (N_4364,In_875,In_2374);
nor U4365 (N_4365,In_557,In_2073);
nand U4366 (N_4366,In_742,In_1095);
or U4367 (N_4367,In_1973,In_1166);
nand U4368 (N_4368,In_2093,In_338);
and U4369 (N_4369,In_2216,In_1281);
nand U4370 (N_4370,In_800,In_2104);
nand U4371 (N_4371,In_2062,In_1414);
and U4372 (N_4372,In_2197,In_164);
nand U4373 (N_4373,In_2145,In_804);
xnor U4374 (N_4374,In_2100,In_1233);
and U4375 (N_4375,In_214,In_934);
or U4376 (N_4376,In_1601,In_1576);
nor U4377 (N_4377,In_1266,In_454);
nand U4378 (N_4378,In_1868,In_144);
or U4379 (N_4379,In_2098,In_1722);
or U4380 (N_4380,In_2232,In_1750);
nand U4381 (N_4381,In_1098,In_1099);
nand U4382 (N_4382,In_1640,In_178);
or U4383 (N_4383,In_815,In_1996);
or U4384 (N_4384,In_1360,In_1325);
or U4385 (N_4385,In_1592,In_1481);
or U4386 (N_4386,In_1728,In_821);
or U4387 (N_4387,In_1666,In_915);
nor U4388 (N_4388,In_331,In_1528);
and U4389 (N_4389,In_1675,In_601);
and U4390 (N_4390,In_1613,In_2001);
or U4391 (N_4391,In_255,In_2122);
nor U4392 (N_4392,In_2233,In_104);
or U4393 (N_4393,In_237,In_1399);
xnor U4394 (N_4394,In_2444,In_2104);
or U4395 (N_4395,In_656,In_790);
nor U4396 (N_4396,In_135,In_2316);
xnor U4397 (N_4397,In_1854,In_1449);
and U4398 (N_4398,In_2097,In_1562);
nand U4399 (N_4399,In_139,In_1866);
nand U4400 (N_4400,In_441,In_1353);
nor U4401 (N_4401,In_2017,In_1137);
nor U4402 (N_4402,In_6,In_1614);
nor U4403 (N_4403,In_2345,In_849);
nor U4404 (N_4404,In_1179,In_1886);
nand U4405 (N_4405,In_1611,In_1388);
nor U4406 (N_4406,In_1630,In_2381);
or U4407 (N_4407,In_2023,In_2488);
nand U4408 (N_4408,In_1368,In_2181);
nand U4409 (N_4409,In_306,In_727);
nor U4410 (N_4410,In_2135,In_1548);
and U4411 (N_4411,In_1648,In_1904);
and U4412 (N_4412,In_941,In_1940);
or U4413 (N_4413,In_2156,In_595);
nand U4414 (N_4414,In_2103,In_987);
and U4415 (N_4415,In_1171,In_1861);
xor U4416 (N_4416,In_174,In_1508);
or U4417 (N_4417,In_2207,In_1055);
and U4418 (N_4418,In_769,In_761);
or U4419 (N_4419,In_2033,In_781);
and U4420 (N_4420,In_1229,In_2199);
or U4421 (N_4421,In_1748,In_1978);
nand U4422 (N_4422,In_2332,In_640);
nor U4423 (N_4423,In_722,In_1494);
nor U4424 (N_4424,In_613,In_52);
nor U4425 (N_4425,In_1032,In_1520);
xnor U4426 (N_4426,In_1646,In_1597);
and U4427 (N_4427,In_680,In_413);
or U4428 (N_4428,In_200,In_834);
nor U4429 (N_4429,In_264,In_398);
nor U4430 (N_4430,In_105,In_607);
nand U4431 (N_4431,In_248,In_1178);
nand U4432 (N_4432,In_463,In_126);
nor U4433 (N_4433,In_2123,In_374);
or U4434 (N_4434,In_732,In_299);
xnor U4435 (N_4435,In_1493,In_386);
xnor U4436 (N_4436,In_1775,In_1869);
or U4437 (N_4437,In_341,In_1776);
and U4438 (N_4438,In_2262,In_1721);
and U4439 (N_4439,In_1393,In_1332);
nor U4440 (N_4440,In_735,In_2170);
xor U4441 (N_4441,In_129,In_84);
or U4442 (N_4442,In_1610,In_2225);
and U4443 (N_4443,In_2468,In_468);
nor U4444 (N_4444,In_625,In_2270);
xnor U4445 (N_4445,In_345,In_268);
nand U4446 (N_4446,In_588,In_1956);
nor U4447 (N_4447,In_1022,In_599);
and U4448 (N_4448,In_473,In_925);
nor U4449 (N_4449,In_2167,In_1757);
nor U4450 (N_4450,In_2425,In_798);
nand U4451 (N_4451,In_2321,In_573);
xnor U4452 (N_4452,In_2223,In_149);
nand U4453 (N_4453,In_1922,In_980);
nand U4454 (N_4454,In_2185,In_1980);
nor U4455 (N_4455,In_1749,In_1519);
nand U4456 (N_4456,In_901,In_2060);
nand U4457 (N_4457,In_606,In_1072);
nor U4458 (N_4458,In_2229,In_2401);
or U4459 (N_4459,In_1634,In_1998);
or U4460 (N_4460,In_1709,In_885);
and U4461 (N_4461,In_729,In_717);
or U4462 (N_4462,In_1551,In_263);
and U4463 (N_4463,In_2379,In_74);
nor U4464 (N_4464,In_334,In_577);
or U4465 (N_4465,In_1209,In_694);
xnor U4466 (N_4466,In_1143,In_1269);
or U4467 (N_4467,In_1264,In_1791);
and U4468 (N_4468,In_820,In_1804);
and U4469 (N_4469,In_1104,In_997);
nand U4470 (N_4470,In_324,In_2393);
xor U4471 (N_4471,In_1481,In_1268);
nand U4472 (N_4472,In_151,In_1383);
nand U4473 (N_4473,In_2091,In_2028);
and U4474 (N_4474,In_1835,In_1904);
or U4475 (N_4475,In_322,In_2305);
nor U4476 (N_4476,In_1650,In_2107);
and U4477 (N_4477,In_155,In_1637);
nand U4478 (N_4478,In_2380,In_981);
and U4479 (N_4479,In_112,In_1379);
or U4480 (N_4480,In_899,In_1560);
nor U4481 (N_4481,In_1427,In_1000);
xor U4482 (N_4482,In_494,In_980);
or U4483 (N_4483,In_548,In_2313);
nand U4484 (N_4484,In_1724,In_339);
nand U4485 (N_4485,In_619,In_201);
nand U4486 (N_4486,In_1186,In_1899);
nand U4487 (N_4487,In_975,In_1716);
nand U4488 (N_4488,In_1447,In_1819);
or U4489 (N_4489,In_184,In_2233);
and U4490 (N_4490,In_2405,In_1134);
and U4491 (N_4491,In_282,In_847);
nand U4492 (N_4492,In_510,In_1967);
or U4493 (N_4493,In_1618,In_0);
or U4494 (N_4494,In_25,In_788);
nor U4495 (N_4495,In_112,In_1757);
nand U4496 (N_4496,In_2067,In_1312);
nand U4497 (N_4497,In_1825,In_1576);
and U4498 (N_4498,In_2448,In_1083);
nor U4499 (N_4499,In_1634,In_885);
or U4500 (N_4500,In_2087,In_1704);
or U4501 (N_4501,In_1987,In_2422);
and U4502 (N_4502,In_1531,In_1548);
nand U4503 (N_4503,In_1074,In_1573);
nor U4504 (N_4504,In_150,In_430);
nor U4505 (N_4505,In_2292,In_1699);
and U4506 (N_4506,In_2005,In_508);
or U4507 (N_4507,In_2484,In_1195);
or U4508 (N_4508,In_982,In_40);
or U4509 (N_4509,In_28,In_126);
nand U4510 (N_4510,In_1208,In_700);
nand U4511 (N_4511,In_1885,In_1546);
nor U4512 (N_4512,In_908,In_2050);
nand U4513 (N_4513,In_1401,In_1792);
nand U4514 (N_4514,In_1736,In_2076);
or U4515 (N_4515,In_1930,In_969);
nand U4516 (N_4516,In_1162,In_1657);
nor U4517 (N_4517,In_2464,In_1346);
xnor U4518 (N_4518,In_1593,In_1628);
or U4519 (N_4519,In_1731,In_125);
and U4520 (N_4520,In_217,In_132);
nand U4521 (N_4521,In_482,In_734);
or U4522 (N_4522,In_1410,In_2035);
nor U4523 (N_4523,In_2378,In_1534);
or U4524 (N_4524,In_1077,In_2277);
and U4525 (N_4525,In_1260,In_2412);
nor U4526 (N_4526,In_2160,In_2272);
xnor U4527 (N_4527,In_2062,In_1927);
or U4528 (N_4528,In_1099,In_2388);
nor U4529 (N_4529,In_1156,In_805);
or U4530 (N_4530,In_2462,In_1330);
or U4531 (N_4531,In_1175,In_1298);
and U4532 (N_4532,In_756,In_1555);
nand U4533 (N_4533,In_1583,In_2241);
and U4534 (N_4534,In_1382,In_27);
xor U4535 (N_4535,In_920,In_269);
nor U4536 (N_4536,In_1797,In_2130);
xor U4537 (N_4537,In_1432,In_1476);
nor U4538 (N_4538,In_2194,In_2439);
or U4539 (N_4539,In_1841,In_1322);
nand U4540 (N_4540,In_2452,In_1118);
and U4541 (N_4541,In_2355,In_2443);
nand U4542 (N_4542,In_18,In_75);
nand U4543 (N_4543,In_2290,In_1479);
nor U4544 (N_4544,In_1562,In_2153);
nand U4545 (N_4545,In_926,In_2182);
or U4546 (N_4546,In_1334,In_2442);
or U4547 (N_4547,In_455,In_947);
nand U4548 (N_4548,In_685,In_1178);
or U4549 (N_4549,In_1196,In_266);
and U4550 (N_4550,In_1151,In_2106);
and U4551 (N_4551,In_2281,In_1392);
nor U4552 (N_4552,In_1245,In_391);
and U4553 (N_4553,In_1310,In_1351);
nor U4554 (N_4554,In_2154,In_1731);
nor U4555 (N_4555,In_2272,In_269);
nor U4556 (N_4556,In_1150,In_1657);
and U4557 (N_4557,In_603,In_1171);
xnor U4558 (N_4558,In_401,In_1771);
nor U4559 (N_4559,In_2233,In_1434);
and U4560 (N_4560,In_914,In_1924);
and U4561 (N_4561,In_2193,In_1977);
nand U4562 (N_4562,In_1419,In_617);
and U4563 (N_4563,In_2165,In_2241);
and U4564 (N_4564,In_14,In_1702);
or U4565 (N_4565,In_1883,In_759);
xor U4566 (N_4566,In_159,In_1501);
and U4567 (N_4567,In_1519,In_2112);
or U4568 (N_4568,In_819,In_1630);
and U4569 (N_4569,In_672,In_2119);
nand U4570 (N_4570,In_1154,In_801);
or U4571 (N_4571,In_1108,In_1482);
or U4572 (N_4572,In_2487,In_1534);
nand U4573 (N_4573,In_993,In_1207);
xor U4574 (N_4574,In_1741,In_1898);
or U4575 (N_4575,In_1724,In_1009);
and U4576 (N_4576,In_507,In_190);
or U4577 (N_4577,In_2119,In_1872);
nand U4578 (N_4578,In_701,In_2139);
nor U4579 (N_4579,In_365,In_1463);
nor U4580 (N_4580,In_650,In_150);
xor U4581 (N_4581,In_736,In_193);
and U4582 (N_4582,In_727,In_2031);
or U4583 (N_4583,In_1457,In_669);
nor U4584 (N_4584,In_725,In_1710);
and U4585 (N_4585,In_1433,In_2427);
xnor U4586 (N_4586,In_36,In_2447);
nor U4587 (N_4587,In_928,In_2441);
nand U4588 (N_4588,In_1732,In_554);
and U4589 (N_4589,In_470,In_2218);
xnor U4590 (N_4590,In_1155,In_333);
and U4591 (N_4591,In_124,In_1314);
and U4592 (N_4592,In_1595,In_1314);
xnor U4593 (N_4593,In_2366,In_2097);
nor U4594 (N_4594,In_999,In_401);
nand U4595 (N_4595,In_418,In_2317);
nor U4596 (N_4596,In_934,In_1120);
xnor U4597 (N_4597,In_56,In_2043);
xor U4598 (N_4598,In_781,In_2329);
nand U4599 (N_4599,In_357,In_2165);
xor U4600 (N_4600,In_1353,In_278);
nand U4601 (N_4601,In_496,In_558);
and U4602 (N_4602,In_1436,In_879);
or U4603 (N_4603,In_2062,In_2090);
xnor U4604 (N_4604,In_722,In_1202);
nor U4605 (N_4605,In_46,In_1720);
nor U4606 (N_4606,In_1479,In_1496);
and U4607 (N_4607,In_1879,In_1193);
or U4608 (N_4608,In_968,In_146);
nand U4609 (N_4609,In_1125,In_1275);
or U4610 (N_4610,In_793,In_1790);
and U4611 (N_4611,In_1844,In_953);
and U4612 (N_4612,In_1707,In_1612);
and U4613 (N_4613,In_722,In_672);
or U4614 (N_4614,In_825,In_2269);
and U4615 (N_4615,In_409,In_576);
or U4616 (N_4616,In_1564,In_802);
and U4617 (N_4617,In_663,In_2242);
nand U4618 (N_4618,In_546,In_2418);
nand U4619 (N_4619,In_301,In_1839);
nand U4620 (N_4620,In_346,In_2391);
or U4621 (N_4621,In_193,In_713);
and U4622 (N_4622,In_105,In_2120);
nand U4623 (N_4623,In_403,In_22);
nor U4624 (N_4624,In_1735,In_391);
and U4625 (N_4625,In_1146,In_318);
xnor U4626 (N_4626,In_433,In_1601);
and U4627 (N_4627,In_2008,In_2162);
nand U4628 (N_4628,In_1080,In_283);
nand U4629 (N_4629,In_2042,In_2456);
and U4630 (N_4630,In_2307,In_953);
or U4631 (N_4631,In_692,In_752);
xnor U4632 (N_4632,In_1723,In_2299);
or U4633 (N_4633,In_562,In_16);
xnor U4634 (N_4634,In_10,In_1861);
nor U4635 (N_4635,In_2220,In_1375);
or U4636 (N_4636,In_1119,In_2176);
nor U4637 (N_4637,In_2113,In_682);
and U4638 (N_4638,In_587,In_529);
nor U4639 (N_4639,In_2020,In_524);
or U4640 (N_4640,In_1632,In_749);
and U4641 (N_4641,In_2306,In_1146);
xor U4642 (N_4642,In_1825,In_1902);
and U4643 (N_4643,In_1840,In_1282);
nand U4644 (N_4644,In_673,In_1253);
nor U4645 (N_4645,In_2396,In_1754);
nand U4646 (N_4646,In_2077,In_1821);
or U4647 (N_4647,In_1632,In_1577);
or U4648 (N_4648,In_603,In_1766);
and U4649 (N_4649,In_1354,In_1691);
and U4650 (N_4650,In_443,In_2397);
or U4651 (N_4651,In_2216,In_42);
xnor U4652 (N_4652,In_66,In_2234);
nand U4653 (N_4653,In_1289,In_2112);
and U4654 (N_4654,In_2200,In_1344);
and U4655 (N_4655,In_780,In_2085);
nand U4656 (N_4656,In_97,In_1984);
xnor U4657 (N_4657,In_78,In_1565);
and U4658 (N_4658,In_183,In_141);
or U4659 (N_4659,In_2220,In_1173);
nand U4660 (N_4660,In_1918,In_2461);
or U4661 (N_4661,In_1378,In_1868);
nand U4662 (N_4662,In_2482,In_161);
nor U4663 (N_4663,In_2271,In_1552);
and U4664 (N_4664,In_1313,In_862);
nor U4665 (N_4665,In_2017,In_1209);
nand U4666 (N_4666,In_1463,In_1841);
and U4667 (N_4667,In_2383,In_1586);
xnor U4668 (N_4668,In_1269,In_925);
nand U4669 (N_4669,In_2031,In_1307);
and U4670 (N_4670,In_422,In_935);
nor U4671 (N_4671,In_1627,In_2254);
nor U4672 (N_4672,In_1356,In_1553);
nor U4673 (N_4673,In_167,In_288);
nor U4674 (N_4674,In_17,In_861);
nand U4675 (N_4675,In_2009,In_15);
or U4676 (N_4676,In_36,In_1149);
nand U4677 (N_4677,In_1844,In_1181);
nor U4678 (N_4678,In_2127,In_3);
and U4679 (N_4679,In_1295,In_852);
nor U4680 (N_4680,In_3,In_2225);
nor U4681 (N_4681,In_651,In_422);
xor U4682 (N_4682,In_1583,In_448);
or U4683 (N_4683,In_1662,In_1207);
nor U4684 (N_4684,In_273,In_1587);
nor U4685 (N_4685,In_1422,In_877);
nand U4686 (N_4686,In_1501,In_1365);
xor U4687 (N_4687,In_1332,In_2281);
nand U4688 (N_4688,In_174,In_1080);
nor U4689 (N_4689,In_1517,In_810);
nand U4690 (N_4690,In_2364,In_1894);
nor U4691 (N_4691,In_779,In_392);
and U4692 (N_4692,In_1480,In_182);
nand U4693 (N_4693,In_327,In_294);
xor U4694 (N_4694,In_1558,In_468);
or U4695 (N_4695,In_2181,In_1475);
and U4696 (N_4696,In_1157,In_2234);
or U4697 (N_4697,In_119,In_1357);
and U4698 (N_4698,In_1597,In_350);
or U4699 (N_4699,In_145,In_2162);
and U4700 (N_4700,In_1451,In_2432);
nand U4701 (N_4701,In_2260,In_926);
or U4702 (N_4702,In_1172,In_306);
nor U4703 (N_4703,In_256,In_1896);
nand U4704 (N_4704,In_1420,In_2104);
or U4705 (N_4705,In_1767,In_902);
nor U4706 (N_4706,In_1371,In_1310);
nor U4707 (N_4707,In_491,In_2110);
nor U4708 (N_4708,In_2428,In_316);
and U4709 (N_4709,In_2045,In_2001);
and U4710 (N_4710,In_1916,In_636);
nand U4711 (N_4711,In_2215,In_932);
or U4712 (N_4712,In_637,In_1531);
or U4713 (N_4713,In_1158,In_310);
nand U4714 (N_4714,In_190,In_1589);
nand U4715 (N_4715,In_407,In_699);
nor U4716 (N_4716,In_1611,In_703);
nor U4717 (N_4717,In_1166,In_1690);
nor U4718 (N_4718,In_1674,In_1138);
or U4719 (N_4719,In_2325,In_1153);
xnor U4720 (N_4720,In_532,In_872);
or U4721 (N_4721,In_1674,In_2287);
nor U4722 (N_4722,In_146,In_977);
nor U4723 (N_4723,In_1353,In_1656);
nand U4724 (N_4724,In_1341,In_867);
nand U4725 (N_4725,In_102,In_284);
nand U4726 (N_4726,In_1325,In_1709);
nor U4727 (N_4727,In_2369,In_2040);
or U4728 (N_4728,In_1667,In_1480);
or U4729 (N_4729,In_332,In_1725);
nor U4730 (N_4730,In_1883,In_2004);
nor U4731 (N_4731,In_139,In_830);
nand U4732 (N_4732,In_1052,In_1565);
or U4733 (N_4733,In_615,In_1953);
or U4734 (N_4734,In_504,In_160);
nand U4735 (N_4735,In_2041,In_1216);
or U4736 (N_4736,In_365,In_1663);
or U4737 (N_4737,In_644,In_2174);
nor U4738 (N_4738,In_870,In_37);
or U4739 (N_4739,In_1391,In_1155);
and U4740 (N_4740,In_775,In_746);
nor U4741 (N_4741,In_1738,In_118);
or U4742 (N_4742,In_1180,In_1155);
and U4743 (N_4743,In_673,In_1825);
nor U4744 (N_4744,In_1190,In_1222);
xnor U4745 (N_4745,In_1420,In_379);
or U4746 (N_4746,In_1623,In_3);
or U4747 (N_4747,In_1605,In_1540);
nor U4748 (N_4748,In_1013,In_1986);
nor U4749 (N_4749,In_1329,In_156);
and U4750 (N_4750,In_595,In_63);
nor U4751 (N_4751,In_275,In_999);
nor U4752 (N_4752,In_1678,In_2103);
and U4753 (N_4753,In_1535,In_499);
nand U4754 (N_4754,In_1403,In_1159);
and U4755 (N_4755,In_618,In_2393);
or U4756 (N_4756,In_1910,In_1294);
nor U4757 (N_4757,In_2229,In_1293);
nor U4758 (N_4758,In_431,In_342);
nor U4759 (N_4759,In_898,In_2390);
nand U4760 (N_4760,In_2314,In_2046);
or U4761 (N_4761,In_1802,In_512);
or U4762 (N_4762,In_987,In_1331);
nand U4763 (N_4763,In_1420,In_727);
or U4764 (N_4764,In_1902,In_1635);
xnor U4765 (N_4765,In_784,In_915);
or U4766 (N_4766,In_1006,In_1795);
or U4767 (N_4767,In_1552,In_242);
or U4768 (N_4768,In_570,In_1669);
and U4769 (N_4769,In_1451,In_582);
nand U4770 (N_4770,In_1811,In_868);
xor U4771 (N_4771,In_2410,In_2369);
or U4772 (N_4772,In_1807,In_1301);
or U4773 (N_4773,In_1874,In_1568);
nand U4774 (N_4774,In_1767,In_1808);
nor U4775 (N_4775,In_2150,In_1769);
or U4776 (N_4776,In_1506,In_243);
or U4777 (N_4777,In_898,In_1833);
nor U4778 (N_4778,In_2042,In_523);
and U4779 (N_4779,In_254,In_2074);
and U4780 (N_4780,In_1474,In_2070);
nor U4781 (N_4781,In_1433,In_1488);
or U4782 (N_4782,In_1568,In_289);
nor U4783 (N_4783,In_1191,In_870);
or U4784 (N_4784,In_2094,In_854);
nor U4785 (N_4785,In_551,In_453);
or U4786 (N_4786,In_694,In_619);
nor U4787 (N_4787,In_1564,In_1632);
or U4788 (N_4788,In_1110,In_1697);
xnor U4789 (N_4789,In_2313,In_1180);
and U4790 (N_4790,In_1818,In_1081);
or U4791 (N_4791,In_1177,In_2480);
xor U4792 (N_4792,In_759,In_1321);
and U4793 (N_4793,In_1603,In_1827);
nor U4794 (N_4794,In_2140,In_1627);
or U4795 (N_4795,In_635,In_1835);
and U4796 (N_4796,In_1280,In_773);
and U4797 (N_4797,In_492,In_1426);
or U4798 (N_4798,In_2180,In_1533);
and U4799 (N_4799,In_104,In_158);
nor U4800 (N_4800,In_60,In_2023);
xnor U4801 (N_4801,In_1185,In_1622);
xor U4802 (N_4802,In_2258,In_1509);
xor U4803 (N_4803,In_2142,In_1397);
nand U4804 (N_4804,In_999,In_1226);
nor U4805 (N_4805,In_2307,In_1253);
nor U4806 (N_4806,In_2479,In_2282);
nor U4807 (N_4807,In_1528,In_970);
or U4808 (N_4808,In_791,In_1650);
or U4809 (N_4809,In_1859,In_543);
and U4810 (N_4810,In_1358,In_1641);
and U4811 (N_4811,In_469,In_1813);
nand U4812 (N_4812,In_1473,In_36);
nand U4813 (N_4813,In_2241,In_2180);
and U4814 (N_4814,In_146,In_2346);
and U4815 (N_4815,In_615,In_1783);
nor U4816 (N_4816,In_795,In_161);
nand U4817 (N_4817,In_1705,In_1560);
nand U4818 (N_4818,In_258,In_1756);
and U4819 (N_4819,In_126,In_365);
or U4820 (N_4820,In_1858,In_2037);
and U4821 (N_4821,In_2177,In_163);
nor U4822 (N_4822,In_1180,In_252);
and U4823 (N_4823,In_2037,In_1674);
and U4824 (N_4824,In_1422,In_595);
or U4825 (N_4825,In_507,In_1858);
or U4826 (N_4826,In_2253,In_1852);
or U4827 (N_4827,In_2328,In_1032);
or U4828 (N_4828,In_140,In_270);
nor U4829 (N_4829,In_1930,In_1207);
or U4830 (N_4830,In_43,In_808);
xnor U4831 (N_4831,In_815,In_1827);
nand U4832 (N_4832,In_270,In_742);
nand U4833 (N_4833,In_1135,In_2320);
xor U4834 (N_4834,In_1069,In_795);
and U4835 (N_4835,In_2032,In_959);
xnor U4836 (N_4836,In_1869,In_2152);
nor U4837 (N_4837,In_760,In_956);
xnor U4838 (N_4838,In_930,In_2212);
nand U4839 (N_4839,In_368,In_371);
and U4840 (N_4840,In_2230,In_596);
nor U4841 (N_4841,In_853,In_2232);
nor U4842 (N_4842,In_2222,In_216);
nand U4843 (N_4843,In_759,In_2416);
or U4844 (N_4844,In_2234,In_722);
and U4845 (N_4845,In_771,In_1207);
nand U4846 (N_4846,In_2023,In_1939);
or U4847 (N_4847,In_1336,In_1891);
nand U4848 (N_4848,In_1319,In_930);
or U4849 (N_4849,In_2240,In_171);
and U4850 (N_4850,In_2491,In_589);
and U4851 (N_4851,In_2344,In_1017);
nand U4852 (N_4852,In_2156,In_182);
nand U4853 (N_4853,In_213,In_589);
xnor U4854 (N_4854,In_1069,In_2434);
nor U4855 (N_4855,In_907,In_648);
and U4856 (N_4856,In_2277,In_2247);
nor U4857 (N_4857,In_1504,In_497);
nor U4858 (N_4858,In_411,In_1289);
nor U4859 (N_4859,In_2046,In_667);
xnor U4860 (N_4860,In_1854,In_2229);
or U4861 (N_4861,In_1380,In_2370);
nor U4862 (N_4862,In_162,In_307);
nor U4863 (N_4863,In_7,In_2150);
or U4864 (N_4864,In_692,In_173);
or U4865 (N_4865,In_317,In_930);
or U4866 (N_4866,In_1468,In_860);
or U4867 (N_4867,In_554,In_978);
and U4868 (N_4868,In_1898,In_2200);
or U4869 (N_4869,In_505,In_1926);
or U4870 (N_4870,In_307,In_1735);
and U4871 (N_4871,In_2483,In_1049);
nor U4872 (N_4872,In_1173,In_1403);
nor U4873 (N_4873,In_1804,In_1383);
and U4874 (N_4874,In_644,In_1011);
or U4875 (N_4875,In_833,In_372);
nand U4876 (N_4876,In_1413,In_1827);
and U4877 (N_4877,In_197,In_440);
and U4878 (N_4878,In_1495,In_2214);
or U4879 (N_4879,In_1978,In_75);
or U4880 (N_4880,In_639,In_1318);
and U4881 (N_4881,In_667,In_1759);
and U4882 (N_4882,In_2228,In_1112);
nor U4883 (N_4883,In_1474,In_1000);
nor U4884 (N_4884,In_2442,In_532);
or U4885 (N_4885,In_1351,In_1913);
nand U4886 (N_4886,In_956,In_1315);
or U4887 (N_4887,In_2410,In_2476);
nand U4888 (N_4888,In_501,In_1821);
nand U4889 (N_4889,In_133,In_359);
or U4890 (N_4890,In_539,In_1092);
nor U4891 (N_4891,In_1863,In_734);
nor U4892 (N_4892,In_426,In_2492);
and U4893 (N_4893,In_255,In_963);
and U4894 (N_4894,In_555,In_1119);
nor U4895 (N_4895,In_1190,In_1753);
or U4896 (N_4896,In_62,In_1356);
or U4897 (N_4897,In_2256,In_217);
or U4898 (N_4898,In_143,In_964);
and U4899 (N_4899,In_2397,In_1359);
and U4900 (N_4900,In_405,In_1345);
and U4901 (N_4901,In_2326,In_277);
and U4902 (N_4902,In_1180,In_89);
or U4903 (N_4903,In_234,In_2419);
or U4904 (N_4904,In_1498,In_2473);
nand U4905 (N_4905,In_2280,In_1108);
or U4906 (N_4906,In_2082,In_1114);
and U4907 (N_4907,In_200,In_2289);
and U4908 (N_4908,In_1687,In_2194);
or U4909 (N_4909,In_546,In_2074);
and U4910 (N_4910,In_64,In_903);
nor U4911 (N_4911,In_2292,In_285);
or U4912 (N_4912,In_1735,In_1213);
nand U4913 (N_4913,In_1949,In_1348);
and U4914 (N_4914,In_1247,In_1729);
nor U4915 (N_4915,In_2286,In_1437);
nand U4916 (N_4916,In_1387,In_755);
nor U4917 (N_4917,In_1532,In_729);
nand U4918 (N_4918,In_1252,In_735);
or U4919 (N_4919,In_412,In_1281);
nand U4920 (N_4920,In_1473,In_1292);
nand U4921 (N_4921,In_806,In_1317);
nand U4922 (N_4922,In_1696,In_1029);
nand U4923 (N_4923,In_2258,In_894);
nand U4924 (N_4924,In_828,In_1029);
and U4925 (N_4925,In_1210,In_752);
nor U4926 (N_4926,In_1314,In_1630);
or U4927 (N_4927,In_1722,In_1133);
nor U4928 (N_4928,In_611,In_2316);
xor U4929 (N_4929,In_2433,In_2265);
nor U4930 (N_4930,In_1215,In_2163);
and U4931 (N_4931,In_649,In_1213);
nor U4932 (N_4932,In_611,In_1504);
or U4933 (N_4933,In_1548,In_633);
nor U4934 (N_4934,In_1043,In_1784);
and U4935 (N_4935,In_1765,In_721);
nand U4936 (N_4936,In_1616,In_533);
and U4937 (N_4937,In_2209,In_1450);
and U4938 (N_4938,In_1393,In_84);
nand U4939 (N_4939,In_2155,In_1133);
or U4940 (N_4940,In_95,In_841);
and U4941 (N_4941,In_1632,In_2288);
and U4942 (N_4942,In_1607,In_1119);
xor U4943 (N_4943,In_256,In_1148);
and U4944 (N_4944,In_441,In_637);
or U4945 (N_4945,In_457,In_2264);
nor U4946 (N_4946,In_481,In_415);
nand U4947 (N_4947,In_2255,In_1067);
xnor U4948 (N_4948,In_1914,In_1444);
nor U4949 (N_4949,In_2288,In_864);
or U4950 (N_4950,In_888,In_2271);
and U4951 (N_4951,In_1913,In_583);
nor U4952 (N_4952,In_2349,In_265);
and U4953 (N_4953,In_669,In_1120);
xor U4954 (N_4954,In_115,In_2363);
nor U4955 (N_4955,In_93,In_2102);
xnor U4956 (N_4956,In_516,In_1720);
nor U4957 (N_4957,In_359,In_1388);
or U4958 (N_4958,In_646,In_1174);
nor U4959 (N_4959,In_1718,In_557);
nor U4960 (N_4960,In_2465,In_1231);
nand U4961 (N_4961,In_1971,In_206);
nand U4962 (N_4962,In_688,In_432);
and U4963 (N_4963,In_311,In_406);
xor U4964 (N_4964,In_980,In_1498);
and U4965 (N_4965,In_162,In_922);
nor U4966 (N_4966,In_492,In_1029);
or U4967 (N_4967,In_625,In_428);
or U4968 (N_4968,In_2421,In_869);
or U4969 (N_4969,In_2,In_1628);
and U4970 (N_4970,In_1393,In_988);
or U4971 (N_4971,In_1553,In_45);
nand U4972 (N_4972,In_116,In_1833);
or U4973 (N_4973,In_645,In_2040);
nand U4974 (N_4974,In_2272,In_2384);
nor U4975 (N_4975,In_740,In_1043);
or U4976 (N_4976,In_2198,In_1091);
nor U4977 (N_4977,In_2417,In_1791);
or U4978 (N_4978,In_830,In_291);
or U4979 (N_4979,In_677,In_1991);
nor U4980 (N_4980,In_268,In_926);
xnor U4981 (N_4981,In_232,In_992);
or U4982 (N_4982,In_619,In_406);
nor U4983 (N_4983,In_1305,In_1088);
nand U4984 (N_4984,In_286,In_762);
nand U4985 (N_4985,In_931,In_306);
nor U4986 (N_4986,In_1427,In_1351);
or U4987 (N_4987,In_1904,In_1546);
and U4988 (N_4988,In_1541,In_2097);
or U4989 (N_4989,In_1518,In_2049);
nor U4990 (N_4990,In_2491,In_477);
nand U4991 (N_4991,In_2338,In_1897);
nor U4992 (N_4992,In_2304,In_1903);
nor U4993 (N_4993,In_1336,In_1557);
nor U4994 (N_4994,In_1860,In_2472);
nor U4995 (N_4995,In_974,In_268);
and U4996 (N_4996,In_1370,In_157);
xnor U4997 (N_4997,In_81,In_1927);
or U4998 (N_4998,In_2183,In_801);
and U4999 (N_4999,In_1887,In_363);
nand U5000 (N_5000,N_858,N_3409);
and U5001 (N_5001,N_2660,N_1248);
xor U5002 (N_5002,N_2049,N_554);
nand U5003 (N_5003,N_3074,N_3188);
xnor U5004 (N_5004,N_4855,N_624);
nand U5005 (N_5005,N_4303,N_1487);
and U5006 (N_5006,N_1637,N_2921);
nand U5007 (N_5007,N_1472,N_3938);
and U5008 (N_5008,N_1474,N_598);
xnor U5009 (N_5009,N_36,N_1754);
nor U5010 (N_5010,N_1595,N_2973);
nor U5011 (N_5011,N_2007,N_844);
nor U5012 (N_5012,N_4581,N_1062);
nand U5013 (N_5013,N_1651,N_4053);
nand U5014 (N_5014,N_1049,N_2335);
nand U5015 (N_5015,N_4722,N_927);
xnor U5016 (N_5016,N_2106,N_3854);
and U5017 (N_5017,N_34,N_1163);
nor U5018 (N_5018,N_3113,N_1841);
nand U5019 (N_5019,N_342,N_2438);
nand U5020 (N_5020,N_3819,N_1438);
and U5021 (N_5021,N_1981,N_2277);
and U5022 (N_5022,N_2704,N_4791);
and U5023 (N_5023,N_4258,N_1698);
nor U5024 (N_5024,N_4655,N_782);
or U5025 (N_5025,N_1796,N_509);
nand U5026 (N_5026,N_1645,N_1385);
xor U5027 (N_5027,N_2554,N_815);
or U5028 (N_5028,N_4294,N_703);
nand U5029 (N_5029,N_1358,N_744);
xor U5030 (N_5030,N_3443,N_1910);
or U5031 (N_5031,N_2748,N_787);
nor U5032 (N_5032,N_3024,N_4533);
and U5033 (N_5033,N_3086,N_4556);
xnor U5034 (N_5034,N_2800,N_3355);
nand U5035 (N_5035,N_1809,N_4668);
or U5036 (N_5036,N_2528,N_3628);
and U5037 (N_5037,N_3407,N_4492);
and U5038 (N_5038,N_3633,N_1074);
nand U5039 (N_5039,N_3745,N_4026);
and U5040 (N_5040,N_4198,N_347);
nor U5041 (N_5041,N_4142,N_834);
or U5042 (N_5042,N_154,N_1011);
or U5043 (N_5043,N_3866,N_3822);
nand U5044 (N_5044,N_4285,N_281);
or U5045 (N_5045,N_1235,N_1236);
or U5046 (N_5046,N_2046,N_3444);
or U5047 (N_5047,N_2126,N_1260);
nor U5048 (N_5048,N_1334,N_2994);
nand U5049 (N_5049,N_5,N_100);
and U5050 (N_5050,N_4852,N_2239);
and U5051 (N_5051,N_3458,N_2926);
xor U5052 (N_5052,N_3011,N_3582);
or U5053 (N_5053,N_2038,N_293);
nand U5054 (N_5054,N_2874,N_1047);
nor U5055 (N_5055,N_4460,N_141);
nor U5056 (N_5056,N_2111,N_1804);
nor U5057 (N_5057,N_1045,N_560);
and U5058 (N_5058,N_4279,N_264);
or U5059 (N_5059,N_2726,N_4520);
xor U5060 (N_5060,N_1097,N_947);
or U5061 (N_5061,N_2405,N_2589);
xnor U5062 (N_5062,N_4642,N_898);
nor U5063 (N_5063,N_571,N_2386);
nand U5064 (N_5064,N_1723,N_3305);
and U5065 (N_5065,N_1722,N_1530);
nor U5066 (N_5066,N_2911,N_4506);
or U5067 (N_5067,N_2464,N_2556);
and U5068 (N_5068,N_3619,N_47);
nor U5069 (N_5069,N_2840,N_2207);
nor U5070 (N_5070,N_2352,N_4212);
nor U5071 (N_5071,N_3876,N_3008);
or U5072 (N_5072,N_1737,N_1437);
nand U5073 (N_5073,N_2297,N_4792);
or U5074 (N_5074,N_1565,N_2646);
and U5075 (N_5075,N_1513,N_2847);
or U5076 (N_5076,N_1345,N_4023);
nor U5077 (N_5077,N_3667,N_4169);
nor U5078 (N_5078,N_2068,N_3816);
xnor U5079 (N_5079,N_3429,N_1276);
nand U5080 (N_5080,N_1324,N_970);
and U5081 (N_5081,N_3194,N_3940);
nand U5082 (N_5082,N_2922,N_4085);
and U5083 (N_5083,N_4180,N_1375);
nor U5084 (N_5084,N_1293,N_4172);
nand U5085 (N_5085,N_3851,N_1112);
or U5086 (N_5086,N_612,N_4171);
and U5087 (N_5087,N_308,N_106);
and U5088 (N_5088,N_3980,N_303);
nor U5089 (N_5089,N_345,N_4341);
or U5090 (N_5090,N_1557,N_1263);
nor U5091 (N_5091,N_2624,N_4761);
and U5092 (N_5092,N_658,N_258);
and U5093 (N_5093,N_2951,N_4548);
and U5094 (N_5094,N_3336,N_3702);
and U5095 (N_5095,N_3416,N_177);
nand U5096 (N_5096,N_586,N_4297);
and U5097 (N_5097,N_1707,N_2032);
and U5098 (N_5098,N_300,N_826);
nor U5099 (N_5099,N_3119,N_2446);
nand U5100 (N_5100,N_2059,N_1328);
and U5101 (N_5101,N_3029,N_164);
nor U5102 (N_5102,N_3027,N_3560);
nand U5103 (N_5103,N_2070,N_1653);
nor U5104 (N_5104,N_896,N_3123);
nand U5105 (N_5105,N_55,N_1745);
and U5106 (N_5106,N_1610,N_3857);
nor U5107 (N_5107,N_3034,N_488);
nor U5108 (N_5108,N_1633,N_1411);
nand U5109 (N_5109,N_965,N_1904);
and U5110 (N_5110,N_3133,N_3030);
nor U5111 (N_5111,N_1788,N_3732);
nand U5112 (N_5112,N_2853,N_2146);
or U5113 (N_5113,N_182,N_939);
or U5114 (N_5114,N_1543,N_3558);
and U5115 (N_5115,N_3922,N_1216);
and U5116 (N_5116,N_1784,N_2750);
nand U5117 (N_5117,N_865,N_4406);
nand U5118 (N_5118,N_3430,N_3406);
and U5119 (N_5119,N_2166,N_552);
nand U5120 (N_5120,N_1744,N_4921);
or U5121 (N_5121,N_2003,N_1226);
or U5122 (N_5122,N_2429,N_203);
nor U5123 (N_5123,N_4249,N_2550);
nand U5124 (N_5124,N_2783,N_1980);
nand U5125 (N_5125,N_1848,N_3057);
or U5126 (N_5126,N_2863,N_4778);
nand U5127 (N_5127,N_3920,N_2320);
nor U5128 (N_5128,N_731,N_4827);
nand U5129 (N_5129,N_4537,N_1685);
and U5130 (N_5130,N_827,N_4076);
or U5131 (N_5131,N_4199,N_87);
nand U5132 (N_5132,N_2671,N_4344);
nor U5133 (N_5133,N_3629,N_3672);
or U5134 (N_5134,N_1446,N_775);
nor U5135 (N_5135,N_2423,N_3110);
nand U5136 (N_5136,N_1355,N_3686);
xor U5137 (N_5137,N_3427,N_1902);
or U5138 (N_5138,N_325,N_1329);
or U5139 (N_5139,N_1435,N_1059);
nor U5140 (N_5140,N_1982,N_2005);
nor U5141 (N_5141,N_804,N_4321);
and U5142 (N_5142,N_4715,N_3346);
or U5143 (N_5143,N_272,N_692);
and U5144 (N_5144,N_2017,N_2823);
and U5145 (N_5145,N_3002,N_3928);
nor U5146 (N_5146,N_1708,N_2889);
nand U5147 (N_5147,N_2494,N_3679);
and U5148 (N_5148,N_4898,N_656);
xor U5149 (N_5149,N_1673,N_4122);
nand U5150 (N_5150,N_3743,N_1410);
and U5151 (N_5151,N_2174,N_2736);
nor U5152 (N_5152,N_4652,N_3186);
or U5153 (N_5153,N_1457,N_44);
and U5154 (N_5154,N_3697,N_1903);
or U5155 (N_5155,N_1132,N_4110);
nor U5156 (N_5156,N_4283,N_3567);
and U5157 (N_5157,N_298,N_1793);
nand U5158 (N_5158,N_1413,N_2340);
or U5159 (N_5159,N_1022,N_2522);
and U5160 (N_5160,N_4699,N_4476);
or U5161 (N_5161,N_242,N_3576);
or U5162 (N_5162,N_4989,N_3946);
and U5163 (N_5163,N_4416,N_950);
and U5164 (N_5164,N_3303,N_1999);
xor U5165 (N_5165,N_536,N_160);
nor U5166 (N_5166,N_3019,N_3983);
or U5167 (N_5167,N_3933,N_2377);
nand U5168 (N_5168,N_2398,N_565);
nor U5169 (N_5169,N_2380,N_486);
nand U5170 (N_5170,N_1890,N_4578);
or U5171 (N_5171,N_1976,N_3124);
nand U5172 (N_5172,N_4500,N_3972);
nor U5173 (N_5173,N_1277,N_1232);
and U5174 (N_5174,N_247,N_4762);
or U5175 (N_5175,N_3712,N_4600);
nor U5176 (N_5176,N_4557,N_3256);
or U5177 (N_5177,N_4884,N_2856);
xnor U5178 (N_5178,N_1171,N_1986);
xnor U5179 (N_5179,N_3053,N_2989);
nand U5180 (N_5180,N_4790,N_1766);
nor U5181 (N_5181,N_3596,N_4307);
and U5182 (N_5182,N_4413,N_4339);
nand U5183 (N_5183,N_2453,N_2520);
or U5184 (N_5184,N_1210,N_3442);
xnor U5185 (N_5185,N_4112,N_1196);
nand U5186 (N_5186,N_2093,N_4608);
nand U5187 (N_5187,N_3175,N_4851);
nor U5188 (N_5188,N_3840,N_3991);
xnor U5189 (N_5189,N_482,N_2591);
nor U5190 (N_5190,N_367,N_2403);
nor U5191 (N_5191,N_3696,N_2728);
nor U5192 (N_5192,N_2455,N_3206);
or U5193 (N_5193,N_3422,N_1702);
nor U5194 (N_5194,N_1073,N_3916);
or U5195 (N_5195,N_3321,N_2312);
nor U5196 (N_5196,N_3635,N_2581);
xnor U5197 (N_5197,N_103,N_2640);
and U5198 (N_5198,N_3097,N_3795);
or U5199 (N_5199,N_3222,N_4562);
nor U5200 (N_5200,N_1183,N_4982);
nand U5201 (N_5201,N_4874,N_3117);
and U5202 (N_5202,N_3494,N_4645);
nand U5203 (N_5203,N_3967,N_3420);
or U5204 (N_5204,N_3032,N_954);
nand U5205 (N_5205,N_2721,N_1063);
nand U5206 (N_5206,N_1013,N_189);
nor U5207 (N_5207,N_1170,N_3881);
nor U5208 (N_5208,N_4255,N_1190);
and U5209 (N_5209,N_4767,N_3936);
and U5210 (N_5210,N_1310,N_4358);
nand U5211 (N_5211,N_3258,N_2545);
and U5212 (N_5212,N_246,N_4496);
or U5213 (N_5213,N_136,N_314);
xnor U5214 (N_5214,N_1089,N_3168);
and U5215 (N_5215,N_3826,N_2997);
and U5216 (N_5216,N_2127,N_2546);
nor U5217 (N_5217,N_94,N_3814);
xor U5218 (N_5218,N_4411,N_2001);
xnor U5219 (N_5219,N_4310,N_309);
and U5220 (N_5220,N_3181,N_3156);
and U5221 (N_5221,N_842,N_4695);
nand U5222 (N_5222,N_3921,N_3036);
and U5223 (N_5223,N_4241,N_4676);
nor U5224 (N_5224,N_640,N_631);
and U5225 (N_5225,N_2406,N_831);
nand U5226 (N_5226,N_4649,N_3863);
or U5227 (N_5227,N_4003,N_3050);
nand U5228 (N_5228,N_4019,N_4809);
and U5229 (N_5229,N_3246,N_1879);
nand U5230 (N_5230,N_3620,N_1179);
and U5231 (N_5231,N_4661,N_376);
nor U5232 (N_5232,N_4326,N_2339);
xor U5233 (N_5233,N_2898,N_2828);
or U5234 (N_5234,N_3411,N_4766);
nand U5235 (N_5235,N_2244,N_550);
nand U5236 (N_5236,N_3875,N_1211);
and U5237 (N_5237,N_415,N_3077);
nor U5238 (N_5238,N_3451,N_162);
nor U5239 (N_5239,N_2037,N_3387);
xor U5240 (N_5240,N_3600,N_3711);
nor U5241 (N_5241,N_4129,N_193);
nand U5242 (N_5242,N_283,N_248);
xor U5243 (N_5243,N_1193,N_1761);
nor U5244 (N_5244,N_1096,N_2670);
nor U5245 (N_5245,N_1587,N_820);
nor U5246 (N_5246,N_419,N_1729);
xnor U5247 (N_5247,N_1835,N_3249);
nor U5248 (N_5248,N_546,N_4997);
nor U5249 (N_5249,N_3102,N_2759);
or U5250 (N_5250,N_448,N_2971);
nand U5251 (N_5251,N_2950,N_772);
xor U5252 (N_5252,N_3959,N_4049);
and U5253 (N_5253,N_1325,N_3661);
and U5254 (N_5254,N_3884,N_2516);
or U5255 (N_5255,N_1770,N_4013);
and U5256 (N_5256,N_4860,N_1116);
and U5257 (N_5257,N_2098,N_2855);
or U5258 (N_5258,N_287,N_4032);
xnor U5259 (N_5259,N_3380,N_3196);
xnor U5260 (N_5260,N_778,N_1775);
xor U5261 (N_5261,N_99,N_3170);
or U5262 (N_5262,N_1718,N_1528);
and U5263 (N_5263,N_2145,N_2211);
and U5264 (N_5264,N_1883,N_1522);
or U5265 (N_5265,N_2932,N_2618);
or U5266 (N_5266,N_17,N_3939);
xnor U5267 (N_5267,N_369,N_4619);
nor U5268 (N_5268,N_2753,N_4765);
and U5269 (N_5269,N_1174,N_4945);
nor U5270 (N_5270,N_1612,N_405);
nand U5271 (N_5271,N_79,N_3401);
nor U5272 (N_5272,N_2283,N_1396);
xor U5273 (N_5273,N_3997,N_4984);
or U5274 (N_5274,N_3758,N_1317);
and U5275 (N_5275,N_1735,N_2892);
xnor U5276 (N_5276,N_1387,N_2956);
nand U5277 (N_5277,N_3561,N_4218);
and U5278 (N_5278,N_1495,N_3051);
nor U5279 (N_5279,N_1621,N_1878);
nor U5280 (N_5280,N_1647,N_3219);
and U5281 (N_5281,N_4682,N_2777);
or U5282 (N_5282,N_3631,N_4304);
nor U5283 (N_5283,N_3621,N_540);
and U5284 (N_5284,N_1273,N_1639);
or U5285 (N_5285,N_1608,N_1948);
nor U5286 (N_5286,N_4916,N_2521);
nor U5287 (N_5287,N_3289,N_2472);
and U5288 (N_5288,N_1582,N_3512);
and U5289 (N_5289,N_1379,N_1778);
nor U5290 (N_5290,N_3926,N_3426);
or U5291 (N_5291,N_291,N_4208);
or U5292 (N_5292,N_3211,N_4813);
nand U5293 (N_5293,N_2611,N_873);
and U5294 (N_5294,N_1929,N_3052);
or U5295 (N_5295,N_3499,N_4173);
and U5296 (N_5296,N_4717,N_62);
nor U5297 (N_5297,N_2101,N_3423);
or U5298 (N_5298,N_1613,N_1868);
and U5299 (N_5299,N_4434,N_2462);
or U5300 (N_5300,N_1831,N_3045);
xor U5301 (N_5301,N_1360,N_3271);
or U5302 (N_5302,N_2980,N_1627);
or U5303 (N_5303,N_4130,N_2171);
or U5304 (N_5304,N_3383,N_4861);
and U5305 (N_5305,N_1882,N_2848);
and U5306 (N_5306,N_3329,N_697);
nor U5307 (N_5307,N_3167,N_503);
and U5308 (N_5308,N_1794,N_758);
or U5309 (N_5309,N_757,N_523);
nand U5310 (N_5310,N_654,N_297);
xor U5311 (N_5311,N_2397,N_3389);
nor U5312 (N_5312,N_400,N_4305);
and U5313 (N_5313,N_4237,N_2129);
and U5314 (N_5314,N_3569,N_531);
and U5315 (N_5315,N_988,N_74);
nand U5316 (N_5316,N_4958,N_1314);
or U5317 (N_5317,N_3463,N_784);
nand U5318 (N_5318,N_1025,N_2292);
and U5319 (N_5319,N_2231,N_2158);
xor U5320 (N_5320,N_4463,N_905);
nand U5321 (N_5321,N_3166,N_3970);
and U5322 (N_5322,N_903,N_4473);
xor U5323 (N_5323,N_4196,N_1222);
or U5324 (N_5324,N_2715,N_4215);
and U5325 (N_5325,N_296,N_401);
xor U5326 (N_5326,N_1463,N_1007);
or U5327 (N_5327,N_2480,N_2587);
nand U5328 (N_5328,N_3134,N_877);
and U5329 (N_5329,N_2843,N_4482);
and U5330 (N_5330,N_3975,N_4074);
nor U5331 (N_5331,N_4610,N_1044);
nand U5332 (N_5332,N_2103,N_4170);
nor U5333 (N_5333,N_4585,N_746);
and U5334 (N_5334,N_2476,N_1580);
nor U5335 (N_5335,N_4651,N_1800);
nand U5336 (N_5336,N_2755,N_535);
and U5337 (N_5337,N_157,N_3604);
and U5338 (N_5338,N_4001,N_3799);
nand U5339 (N_5339,N_2580,N_2267);
nand U5340 (N_5340,N_2746,N_2458);
or U5341 (N_5341,N_919,N_1065);
and U5342 (N_5342,N_4477,N_1665);
nand U5343 (N_5343,N_2809,N_4856);
nand U5344 (N_5344,N_1019,N_4389);
or U5345 (N_5345,N_3751,N_4746);
and U5346 (N_5346,N_3112,N_3136);
and U5347 (N_5347,N_390,N_4786);
and U5348 (N_5348,N_3578,N_1947);
or U5349 (N_5349,N_191,N_3588);
xor U5350 (N_5350,N_2224,N_2383);
or U5351 (N_5351,N_4664,N_3727);
nor U5352 (N_5352,N_3931,N_64);
nand U5353 (N_5353,N_1266,N_1023);
nand U5354 (N_5354,N_1806,N_590);
nor U5355 (N_5355,N_262,N_649);
nor U5356 (N_5356,N_1040,N_4186);
nor U5357 (N_5357,N_3292,N_1875);
or U5358 (N_5358,N_4103,N_2667);
nand U5359 (N_5359,N_1675,N_3436);
nand U5360 (N_5360,N_2302,N_852);
nand U5361 (N_5361,N_974,N_2372);
nand U5362 (N_5362,N_3138,N_2165);
and U5363 (N_5363,N_4667,N_33);
nand U5364 (N_5364,N_3634,N_4366);
nor U5365 (N_5365,N_3551,N_284);
or U5366 (N_5366,N_2474,N_1897);
nor U5367 (N_5367,N_622,N_2949);
nor U5368 (N_5368,N_3058,N_1041);
nor U5369 (N_5369,N_326,N_3068);
nor U5370 (N_5370,N_4734,N_2953);
nand U5371 (N_5371,N_3664,N_102);
nand U5372 (N_5372,N_112,N_4216);
and U5373 (N_5373,N_2531,N_3116);
and U5374 (N_5374,N_4634,N_2459);
nor U5375 (N_5375,N_993,N_3202);
nor U5376 (N_5376,N_558,N_1414);
and U5377 (N_5377,N_4227,N_739);
or U5378 (N_5378,N_3475,N_492);
nor U5379 (N_5379,N_4947,N_639);
and U5380 (N_5380,N_4771,N_2693);
and U5381 (N_5381,N_3753,N_159);
or U5382 (N_5382,N_1491,N_3941);
nand U5383 (N_5383,N_742,N_904);
xor U5384 (N_5384,N_1838,N_4516);
nand U5385 (N_5385,N_4336,N_457);
or U5386 (N_5386,N_4685,N_3948);
nor U5387 (N_5387,N_578,N_4690);
nand U5388 (N_5388,N_1867,N_2815);
or U5389 (N_5389,N_851,N_319);
nand U5390 (N_5390,N_674,N_4333);
or U5391 (N_5391,N_257,N_104);
or U5392 (N_5392,N_1241,N_375);
or U5393 (N_5393,N_2529,N_4329);
or U5394 (N_5394,N_4257,N_3744);
and U5395 (N_5395,N_3597,N_3900);
nor U5396 (N_5396,N_3747,N_3267);
and U5397 (N_5397,N_124,N_4331);
or U5398 (N_5398,N_548,N_2904);
or U5399 (N_5399,N_4663,N_3049);
or U5400 (N_5400,N_3693,N_4864);
and U5401 (N_5401,N_3522,N_4374);
nand U5402 (N_5402,N_698,N_1483);
and U5403 (N_5403,N_123,N_4932);
and U5404 (N_5404,N_539,N_1120);
or U5405 (N_5405,N_3844,N_866);
nor U5406 (N_5406,N_3198,N_179);
nand U5407 (N_5407,N_765,N_1807);
nor U5408 (N_5408,N_295,N_4179);
xor U5409 (N_5409,N_4881,N_1819);
nand U5410 (N_5410,N_2349,N_994);
and U5411 (N_5411,N_1768,N_2191);
nand U5412 (N_5412,N_3284,N_440);
nor U5413 (N_5413,N_4816,N_3377);
nor U5414 (N_5414,N_2388,N_3091);
and U5415 (N_5415,N_1336,N_1450);
nor U5416 (N_5416,N_4299,N_679);
or U5417 (N_5417,N_153,N_4880);
and U5418 (N_5418,N_3710,N_3956);
xor U5419 (N_5419,N_251,N_1787);
and U5420 (N_5420,N_4168,N_4252);
or U5421 (N_5421,N_1346,N_4461);
nor U5422 (N_5422,N_3668,N_1257);
and U5423 (N_5423,N_1155,N_4393);
or U5424 (N_5424,N_556,N_3683);
xnor U5425 (N_5425,N_3784,N_4700);
nand U5426 (N_5426,N_4638,N_1760);
and U5427 (N_5427,N_4143,N_173);
and U5428 (N_5428,N_2159,N_3467);
and U5429 (N_5429,N_661,N_3071);
and U5430 (N_5430,N_1080,N_4472);
nand U5431 (N_5431,N_270,N_691);
and U5432 (N_5432,N_4347,N_2699);
and U5433 (N_5433,N_797,N_813);
nor U5434 (N_5434,N_2967,N_1180);
nand U5435 (N_5435,N_3352,N_3491);
and U5436 (N_5436,N_4902,N_884);
and U5437 (N_5437,N_3418,N_3590);
or U5438 (N_5438,N_3237,N_3856);
or U5439 (N_5439,N_1123,N_525);
nand U5440 (N_5440,N_341,N_4993);
and U5441 (N_5441,N_4005,N_645);
and U5442 (N_5442,N_4917,N_585);
nor U5443 (N_5443,N_4770,N_56);
or U5444 (N_5444,N_1989,N_3520);
or U5445 (N_5445,N_4798,N_1365);
nor U5446 (N_5446,N_690,N_1240);
nor U5447 (N_5447,N_2974,N_2078);
nand U5448 (N_5448,N_4821,N_1111);
or U5449 (N_5449,N_4099,N_1270);
or U5450 (N_5450,N_3660,N_3290);
or U5451 (N_5451,N_3268,N_1181);
or U5452 (N_5452,N_437,N_1469);
and U5453 (N_5453,N_4590,N_943);
nand U5454 (N_5454,N_1602,N_4095);
or U5455 (N_5455,N_613,N_4543);
nand U5456 (N_5456,N_625,N_3031);
nor U5457 (N_5457,N_1326,N_1519);
nor U5458 (N_5458,N_2601,N_4203);
or U5459 (N_5459,N_1547,N_2826);
or U5460 (N_5460,N_1606,N_515);
or U5461 (N_5461,N_427,N_1710);
or U5462 (N_5462,N_3085,N_763);
nand U5463 (N_5463,N_290,N_1777);
nand U5464 (N_5464,N_1197,N_901);
and U5465 (N_5465,N_1477,N_2389);
nor U5466 (N_5466,N_4245,N_2381);
or U5467 (N_5467,N_4635,N_2912);
nand U5468 (N_5468,N_1367,N_2551);
or U5469 (N_5469,N_1577,N_2557);
nor U5470 (N_5470,N_961,N_412);
or U5471 (N_5471,N_3216,N_3534);
or U5472 (N_5472,N_987,N_1660);
nor U5473 (N_5473,N_4487,N_4390);
or U5474 (N_5474,N_2197,N_4637);
or U5475 (N_5475,N_2117,N_3824);
or U5476 (N_5476,N_4814,N_2831);
xnor U5477 (N_5477,N_1889,N_1916);
nand U5478 (N_5478,N_2758,N_3915);
xor U5479 (N_5479,N_4614,N_3332);
nand U5480 (N_5480,N_1337,N_4991);
nand U5481 (N_5481,N_3090,N_1009);
or U5482 (N_5482,N_2636,N_4574);
nor U5483 (N_5483,N_610,N_522);
or U5484 (N_5484,N_150,N_2797);
or U5485 (N_5485,N_3677,N_3195);
xnor U5486 (N_5486,N_3248,N_791);
or U5487 (N_5487,N_2719,N_328);
or U5488 (N_5488,N_2121,N_879);
or U5489 (N_5489,N_2865,N_3073);
xor U5490 (N_5490,N_1238,N_1117);
nand U5491 (N_5491,N_2366,N_3811);
nand U5492 (N_5492,N_4157,N_2247);
nor U5493 (N_5493,N_2844,N_1896);
nor U5494 (N_5494,N_3266,N_549);
nor U5495 (N_5495,N_2504,N_3888);
nand U5496 (N_5496,N_10,N_4938);
or U5497 (N_5497,N_4862,N_1713);
and U5498 (N_5498,N_4131,N_1465);
nor U5499 (N_5499,N_2401,N_2642);
nor U5500 (N_5500,N_1296,N_2113);
nor U5501 (N_5501,N_3366,N_2326);
nand U5502 (N_5502,N_3337,N_1998);
and U5503 (N_5503,N_3233,N_4034);
and U5504 (N_5504,N_3793,N_696);
and U5505 (N_5505,N_256,N_3963);
and U5506 (N_5506,N_2270,N_1227);
nor U5507 (N_5507,N_2257,N_3836);
or U5508 (N_5508,N_4153,N_632);
nand U5509 (N_5509,N_2437,N_1185);
or U5510 (N_5510,N_921,N_1578);
nor U5511 (N_5511,N_1506,N_3670);
nand U5512 (N_5512,N_4037,N_498);
nand U5513 (N_5513,N_2527,N_4288);
xnor U5514 (N_5514,N_2610,N_3402);
and U5515 (N_5515,N_1844,N_2345);
or U5516 (N_5516,N_1,N_3379);
or U5517 (N_5517,N_3911,N_2220);
and U5518 (N_5518,N_27,N_642);
and U5519 (N_5519,N_2631,N_2764);
or U5520 (N_5520,N_471,N_2234);
nand U5521 (N_5521,N_2680,N_3858);
nor U5522 (N_5522,N_1318,N_641);
and U5523 (N_5523,N_2333,N_4156);
xor U5524 (N_5524,N_420,N_705);
and U5525 (N_5525,N_1348,N_3974);
or U5526 (N_5526,N_2138,N_95);
nor U5527 (N_5527,N_4913,N_4704);
or U5528 (N_5528,N_2762,N_992);
nand U5529 (N_5529,N_6,N_4750);
nor U5530 (N_5530,N_2996,N_1301);
nand U5531 (N_5531,N_676,N_2594);
nor U5532 (N_5532,N_4259,N_1458);
nand U5533 (N_5533,N_1656,N_2722);
and U5534 (N_5534,N_1706,N_4755);
and U5535 (N_5535,N_2788,N_2050);
nor U5536 (N_5536,N_1699,N_1849);
or U5537 (N_5537,N_767,N_469);
nand U5538 (N_5538,N_1940,N_4627);
nor U5539 (N_5539,N_1489,N_213);
or U5540 (N_5540,N_3934,N_1812);
or U5541 (N_5541,N_4918,N_4004);
nor U5542 (N_5542,N_860,N_2724);
xor U5543 (N_5543,N_1644,N_2433);
or U5544 (N_5544,N_2269,N_4698);
or U5545 (N_5545,N_4731,N_2771);
and U5546 (N_5546,N_4973,N_931);
or U5547 (N_5547,N_3657,N_4857);
xnor U5548 (N_5548,N_4568,N_3954);
nand U5549 (N_5549,N_647,N_2254);
xnor U5550 (N_5550,N_2278,N_180);
nor U5551 (N_5551,N_2714,N_3791);
and U5552 (N_5552,N_3557,N_4597);
nand U5553 (N_5553,N_908,N_1290);
nor U5554 (N_5554,N_1175,N_4739);
nand U5555 (N_5555,N_4485,N_2463);
nand U5556 (N_5556,N_2524,N_2408);
and U5557 (N_5557,N_2261,N_2296);
nand U5558 (N_5558,N_1148,N_2947);
or U5559 (N_5559,N_2782,N_874);
nand U5560 (N_5560,N_2955,N_2478);
nand U5561 (N_5561,N_2088,N_3262);
nand U5562 (N_5562,N_2779,N_4885);
or U5563 (N_5563,N_311,N_3253);
nand U5564 (N_5564,N_2605,N_3080);
and U5565 (N_5565,N_1035,N_4483);
xor U5566 (N_5566,N_606,N_3918);
nor U5567 (N_5567,N_1021,N_847);
nor U5568 (N_5568,N_1709,N_186);
xnor U5569 (N_5569,N_3584,N_3470);
and U5570 (N_5570,N_2639,N_4486);
nand U5571 (N_5571,N_4323,N_3438);
nor U5572 (N_5572,N_1462,N_544);
xor U5573 (N_5573,N_185,N_3809);
xor U5574 (N_5574,N_2004,N_669);
or U5575 (N_5575,N_4193,N_2440);
nand U5576 (N_5576,N_1188,N_1281);
nand U5577 (N_5577,N_3472,N_893);
and U5578 (N_5578,N_86,N_85);
nor U5579 (N_5579,N_1927,N_2732);
nand U5580 (N_5580,N_2065,N_1884);
or U5581 (N_5581,N_3681,N_2658);
nand U5582 (N_5582,N_4164,N_840);
or U5583 (N_5583,N_4542,N_1072);
nand U5584 (N_5584,N_1319,N_2313);
nand U5585 (N_5585,N_1847,N_4956);
or U5586 (N_5586,N_4963,N_3391);
or U5587 (N_5587,N_4449,N_2124);
and U5588 (N_5588,N_3001,N_3322);
nand U5589 (N_5589,N_3006,N_4536);
nor U5590 (N_5590,N_438,N_3501);
xor U5591 (N_5591,N_1730,N_1850);
xnor U5592 (N_5592,N_4035,N_2569);
nand U5593 (N_5593,N_557,N_4671);
or U5594 (N_5594,N_1140,N_4426);
xor U5595 (N_5595,N_4760,N_2081);
and U5596 (N_5596,N_288,N_829);
or U5597 (N_5597,N_4365,N_2583);
nand U5598 (N_5598,N_211,N_2334);
or U5599 (N_5599,N_1368,N_3126);
nor U5600 (N_5600,N_1481,N_1027);
nor U5601 (N_5601,N_3500,N_1246);
or U5602 (N_5602,N_559,N_2873);
nand U5603 (N_5603,N_951,N_3552);
nand U5604 (N_5604,N_1341,N_3505);
and U5605 (N_5605,N_4233,N_3384);
nand U5606 (N_5606,N_4117,N_2567);
or U5607 (N_5607,N_475,N_2725);
nand U5608 (N_5608,N_66,N_3804);
nand U5609 (N_5609,N_3174,N_3218);
nand U5610 (N_5610,N_811,N_2303);
and U5611 (N_5611,N_1876,N_2519);
and U5612 (N_5612,N_43,N_433);
or U5613 (N_5613,N_4818,N_11);
nor U5614 (N_5614,N_479,N_307);
and U5615 (N_5615,N_1558,N_4301);
nand U5616 (N_5616,N_1593,N_1624);
nand U5617 (N_5617,N_3944,N_3742);
and U5618 (N_5618,N_2275,N_4148);
and U5619 (N_5619,N_2432,N_2087);
nor U5620 (N_5620,N_3827,N_3526);
or U5621 (N_5621,N_856,N_3238);
or U5622 (N_5622,N_3725,N_4281);
nand U5623 (N_5623,N_2284,N_1563);
nor U5624 (N_5624,N_4908,N_3328);
nor U5625 (N_5625,N_686,N_3356);
nor U5626 (N_5626,N_4191,N_2883);
nor U5627 (N_5627,N_4381,N_3414);
xnor U5628 (N_5628,N_3445,N_953);
and U5629 (N_5629,N_4751,N_4296);
and U5630 (N_5630,N_2535,N_1299);
nor U5631 (N_5631,N_1338,N_4371);
nor U5632 (N_5632,N_2744,N_2887);
and U5633 (N_5633,N_1993,N_1416);
and U5634 (N_5634,N_3013,N_3432);
xnor U5635 (N_5635,N_1460,N_3154);
nor U5636 (N_5636,N_3078,N_1030);
or U5637 (N_5637,N_317,N_609);
nor U5638 (N_5638,N_51,N_2448);
nand U5639 (N_5639,N_4563,N_1084);
nor U5640 (N_5640,N_4395,N_4988);
xor U5641 (N_5641,N_3987,N_2582);
nand U5642 (N_5642,N_3771,N_2016);
and U5643 (N_5643,N_1344,N_4546);
or U5644 (N_5644,N_3986,N_603);
xor U5645 (N_5645,N_2014,N_2192);
nor U5646 (N_5646,N_4182,N_483);
and U5647 (N_5647,N_3288,N_2707);
nand U5648 (N_5648,N_2492,N_1259);
or U5649 (N_5649,N_4720,N_1204);
or U5650 (N_5650,N_3368,N_1974);
nor U5651 (N_5651,N_1134,N_3606);
or U5652 (N_5652,N_81,N_3208);
and U5653 (N_5653,N_3848,N_2170);
nand U5654 (N_5654,N_839,N_3227);
and U5655 (N_5655,N_1031,N_3792);
or U5656 (N_5656,N_1058,N_3680);
and U5657 (N_5657,N_2882,N_4996);
or U5658 (N_5658,N_4123,N_218);
and U5659 (N_5659,N_1623,N_199);
xnor U5660 (N_5660,N_3439,N_1198);
nor U5661 (N_5661,N_1725,N_2559);
or U5662 (N_5662,N_4205,N_3563);
nor U5663 (N_5663,N_1938,N_3917);
nor U5664 (N_5664,N_465,N_777);
or U5665 (N_5665,N_1905,N_428);
and U5666 (N_5666,N_72,N_4120);
and U5667 (N_5667,N_3594,N_430);
nor U5668 (N_5668,N_2128,N_4726);
xnor U5669 (N_5669,N_1100,N_2487);
or U5670 (N_5670,N_2295,N_621);
nand U5671 (N_5671,N_962,N_241);
or U5672 (N_5672,N_1664,N_4363);
nor U5673 (N_5673,N_4111,N_3838);
nor U5674 (N_5674,N_4446,N_2354);
nor U5675 (N_5675,N_4146,N_2225);
xor U5676 (N_5676,N_1803,N_1631);
and U5677 (N_5677,N_714,N_3644);
and U5678 (N_5678,N_2315,N_633);
nor U5679 (N_5679,N_1694,N_89);
xor U5680 (N_5680,N_2272,N_1743);
or U5681 (N_5681,N_198,N_4501);
xor U5682 (N_5682,N_2252,N_232);
nor U5683 (N_5683,N_4504,N_2052);
nor U5684 (N_5684,N_386,N_196);
or U5685 (N_5685,N_1560,N_1894);
nand U5686 (N_5686,N_434,N_3232);
nor U5687 (N_5687,N_4105,N_1880);
nand U5688 (N_5688,N_899,N_3957);
nor U5689 (N_5689,N_3287,N_3626);
and U5690 (N_5690,N_887,N_3291);
nor U5691 (N_5691,N_1321,N_2045);
nor U5692 (N_5692,N_4998,N_3473);
or U5693 (N_5693,N_4269,N_260);
xnor U5694 (N_5694,N_3285,N_4702);
or U5695 (N_5695,N_212,N_1165);
and U5696 (N_5696,N_510,N_2365);
nand U5697 (N_5697,N_1567,N_2977);
nor U5698 (N_5698,N_2813,N_1795);
and U5699 (N_5699,N_766,N_2204);
and U5700 (N_5700,N_4630,N_4625);
nor U5701 (N_5701,N_4260,N_728);
or U5702 (N_5702,N_355,N_3755);
nor U5703 (N_5703,N_1106,N_2214);
nand U5704 (N_5704,N_1680,N_781);
nand U5705 (N_5705,N_512,N_143);
or U5706 (N_5706,N_1421,N_3641);
nor U5707 (N_5707,N_1842,N_1160);
nand U5708 (N_5708,N_1042,N_1827);
and U5709 (N_5709,N_1516,N_3889);
or U5710 (N_5710,N_4980,N_46);
xnor U5711 (N_5711,N_4050,N_3525);
or U5712 (N_5712,N_4825,N_2035);
nor U5713 (N_5713,N_237,N_1690);
nand U5714 (N_5714,N_209,N_3550);
nand U5715 (N_5715,N_2473,N_3158);
and U5716 (N_5716,N_330,N_938);
nand U5717 (N_5717,N_280,N_920);
or U5718 (N_5718,N_591,N_3541);
nand U5719 (N_5719,N_285,N_4960);
or U5720 (N_5720,N_137,N_1086);
nor U5721 (N_5721,N_1946,N_1893);
nor U5722 (N_5722,N_2307,N_4189);
and U5723 (N_5723,N_4274,N_1378);
nand U5724 (N_5724,N_1217,N_1810);
or U5725 (N_5725,N_1088,N_4797);
xor U5726 (N_5726,N_1311,N_1525);
nand U5727 (N_5727,N_3200,N_4894);
and U5728 (N_5728,N_339,N_1415);
nand U5729 (N_5729,N_269,N_2903);
nand U5730 (N_5730,N_671,N_3782);
nor U5731 (N_5731,N_4733,N_2511);
nand U5732 (N_5732,N_4706,N_4470);
nor U5733 (N_5733,N_477,N_3638);
or U5734 (N_5734,N_1350,N_1607);
and U5735 (N_5735,N_4666,N_1915);
nor U5736 (N_5736,N_3270,N_3184);
or U5737 (N_5737,N_4452,N_505);
or U5738 (N_5738,N_1366,N_2573);
or U5739 (N_5739,N_3437,N_1178);
xor U5740 (N_5740,N_4839,N_730);
or U5741 (N_5741,N_4896,N_4058);
nor U5742 (N_5742,N_3878,N_4566);
nor U5743 (N_5743,N_1629,N_823);
and U5744 (N_5744,N_3599,N_1101);
nand U5745 (N_5745,N_3130,N_35);
or U5746 (N_5746,N_1546,N_4879);
xor U5747 (N_5747,N_63,N_4589);
xor U5748 (N_5748,N_2891,N_655);
and U5749 (N_5749,N_602,N_4789);
and U5750 (N_5750,N_1388,N_4787);
xnor U5751 (N_5751,N_2899,N_2375);
or U5752 (N_5752,N_3038,N_3545);
nor U5753 (N_5753,N_720,N_2766);
and U5754 (N_5754,N_1461,N_1967);
or U5755 (N_5755,N_3100,N_984);
or U5756 (N_5756,N_2051,N_4235);
nand U5757 (N_5757,N_3966,N_377);
or U5758 (N_5758,N_4280,N_4838);
nor U5759 (N_5759,N_4910,N_737);
xor U5760 (N_5760,N_4223,N_2177);
nand U5761 (N_5761,N_2264,N_3351);
nand U5762 (N_5762,N_4712,N_2651);
or U5763 (N_5763,N_4386,N_1298);
nand U5764 (N_5764,N_3129,N_4137);
and U5765 (N_5765,N_4745,N_2493);
or U5766 (N_5766,N_4815,N_4519);
or U5767 (N_5767,N_1026,N_3004);
and U5768 (N_5768,N_4622,N_2854);
nand U5769 (N_5769,N_3257,N_4442);
or U5770 (N_5770,N_1256,N_2125);
or U5771 (N_5771,N_4409,N_2697);
and U5772 (N_5772,N_3450,N_680);
nand U5773 (N_5773,N_3675,N_2217);
or U5774 (N_5774,N_2615,N_4774);
or U5775 (N_5775,N_2652,N_1245);
and U5776 (N_5776,N_4886,N_3964);
nor U5777 (N_5777,N_215,N_2028);
nand U5778 (N_5778,N_1510,N_316);
nor U5779 (N_5779,N_4540,N_2906);
and U5780 (N_5780,N_2560,N_1369);
and U5781 (N_5781,N_4802,N_1959);
and U5782 (N_5782,N_2930,N_1340);
xor U5783 (N_5783,N_2905,N_2555);
and U5784 (N_5784,N_4757,N_1970);
and U5785 (N_5785,N_4854,N_71);
xnor U5786 (N_5786,N_2394,N_1550);
or U5787 (N_5787,N_4041,N_4271);
nand U5788 (N_5788,N_3935,N_4201);
or U5789 (N_5789,N_406,N_3513);
or U5790 (N_5790,N_4410,N_4686);
and U5791 (N_5791,N_2650,N_1092);
nor U5792 (N_5792,N_3201,N_4125);
xor U5793 (N_5793,N_2399,N_545);
and U5794 (N_5794,N_4840,N_534);
and U5795 (N_5795,N_3978,N_4660);
nor U5796 (N_5796,N_2970,N_3831);
nor U5797 (N_5797,N_4541,N_2767);
xor U5798 (N_5798,N_1268,N_4957);
xor U5799 (N_5799,N_693,N_1774);
nand U5800 (N_5800,N_2328,N_1555);
or U5801 (N_5801,N_2357,N_4348);
nand U5802 (N_5802,N_1147,N_2230);
and U5803 (N_5803,N_2628,N_3490);
and U5804 (N_5804,N_4607,N_4006);
and U5805 (N_5805,N_4783,N_2663);
or U5806 (N_5806,N_4448,N_2201);
nand U5807 (N_5807,N_2233,N_2626);
or U5808 (N_5808,N_630,N_2890);
and U5809 (N_5809,N_2851,N_4009);
or U5810 (N_5810,N_2570,N_3028);
or U5811 (N_5811,N_3165,N_4396);
nor U5812 (N_5812,N_3605,N_4054);
nor U5813 (N_5813,N_1828,N_1056);
or U5814 (N_5814,N_2179,N_2888);
or U5815 (N_5815,N_701,N_2530);
nand U5816 (N_5816,N_2752,N_3082);
and U5817 (N_5817,N_1275,N_1408);
and U5818 (N_5818,N_1207,N_1284);
nand U5819 (N_5819,N_3846,N_395);
nor U5820 (N_5820,N_2937,N_4665);
or U5821 (N_5821,N_1561,N_3242);
nand U5822 (N_5822,N_4939,N_1315);
nor U5823 (N_5823,N_4972,N_2358);
and U5824 (N_5824,N_2833,N_3283);
and U5825 (N_5825,N_4822,N_702);
and U5826 (N_5826,N_3717,N_4843);
or U5827 (N_5827,N_4401,N_952);
nor U5828 (N_5828,N_918,N_2859);
nand U5829 (N_5829,N_2180,N_2213);
xnor U5830 (N_5830,N_2666,N_4990);
nor U5831 (N_5831,N_4992,N_688);
nor U5832 (N_5832,N_1957,N_4232);
nor U5833 (N_5833,N_4376,N_3101);
nor U5834 (N_5834,N_4335,N_568);
or U5835 (N_5835,N_2327,N_426);
xor U5836 (N_5836,N_3255,N_895);
nand U5837 (N_5837,N_1224,N_1493);
and U5838 (N_5838,N_3805,N_1802);
nand U5839 (N_5839,N_1242,N_4421);
xnor U5840 (N_5840,N_4458,N_4656);
xor U5841 (N_5841,N_4983,N_3235);
or U5842 (N_5842,N_1843,N_3497);
nor U5843 (N_5843,N_1184,N_4222);
nor U5844 (N_5844,N_1670,N_2008);
nor U5845 (N_5845,N_2316,N_384);
nor U5846 (N_5846,N_4639,N_3359);
and U5847 (N_5847,N_244,N_2260);
and U5848 (N_5848,N_1430,N_4673);
nand U5849 (N_5849,N_4805,N_1750);
or U5850 (N_5850,N_1853,N_2139);
nand U5851 (N_5851,N_3904,N_3025);
and U5852 (N_5852,N_733,N_2781);
nor U5853 (N_5853,N_4159,N_49);
or U5854 (N_5854,N_3141,N_1356);
nor U5855 (N_5855,N_1576,N_1650);
and U5856 (N_5856,N_2107,N_3988);
or U5857 (N_5857,N_2376,N_599);
nor U5858 (N_5858,N_2481,N_805);
nand U5859 (N_5859,N_3122,N_3345);
and U5860 (N_5860,N_3056,N_4200);
or U5861 (N_5861,N_4844,N_1395);
xor U5862 (N_5862,N_3842,N_3930);
nand U5863 (N_5863,N_4718,N_1984);
and U5864 (N_5864,N_2141,N_3221);
and U5865 (N_5865,N_2701,N_4756);
and U5866 (N_5866,N_3774,N_4924);
or U5867 (N_5867,N_91,N_4007);
nor U5868 (N_5868,N_1130,N_4832);
xnor U5869 (N_5869,N_2568,N_793);
nor U5870 (N_5870,N_3883,N_790);
nor U5871 (N_5871,N_4969,N_4708);
or U5872 (N_5872,N_707,N_455);
nor U5873 (N_5873,N_2643,N_2803);
xnor U5874 (N_5874,N_1603,N_1601);
or U5875 (N_5875,N_2747,N_82);
nor U5876 (N_5876,N_3976,N_2935);
xor U5877 (N_5877,N_1267,N_2999);
or U5878 (N_5878,N_60,N_2308);
nand U5879 (N_5879,N_1467,N_4437);
and U5880 (N_5880,N_2209,N_3554);
nand U5881 (N_5881,N_4535,N_2413);
nand U5882 (N_5882,N_1076,N_2858);
nor U5883 (N_5883,N_1055,N_1816);
nor U5884 (N_5884,N_1452,N_2805);
or U5885 (N_5885,N_254,N_313);
nor U5886 (N_5886,N_399,N_760);
nand U5887 (N_5887,N_4162,N_449);
nor U5888 (N_5888,N_4465,N_1444);
nand U5889 (N_5889,N_4829,N_249);
nand U5890 (N_5890,N_955,N_678);
xor U5891 (N_5891,N_1655,N_1852);
or U5892 (N_5892,N_3642,N_4728);
and U5893 (N_5893,N_3813,N_1090);
nand U5894 (N_5894,N_3610,N_2544);
nor U5895 (N_5895,N_1724,N_3548);
or U5896 (N_5896,N_2547,N_1705);
nand U5897 (N_5897,N_2468,N_3733);
and U5898 (N_5898,N_2227,N_3396);
nor U5899 (N_5899,N_4826,N_2015);
or U5900 (N_5900,N_306,N_4210);
nor U5901 (N_5901,N_1652,N_416);
or U5902 (N_5902,N_1202,N_282);
nor U5903 (N_5903,N_853,N_808);
and U5904 (N_5904,N_1762,N_4278);
and U5905 (N_5905,N_634,N_1825);
nor U5906 (N_5906,N_3135,N_2538);
nand U5907 (N_5907,N_4048,N_422);
and U5908 (N_5908,N_1973,N_3347);
nor U5909 (N_5909,N_2827,N_841);
nor U5910 (N_5910,N_2677,N_3225);
nor U5911 (N_5911,N_2069,N_2665);
xor U5912 (N_5912,N_3764,N_3757);
nand U5913 (N_5913,N_4197,N_1870);
and U5914 (N_5914,N_2259,N_414);
and U5915 (N_5915,N_4711,N_2893);
or U5916 (N_5916,N_2109,N_1785);
nand U5917 (N_5917,N_729,N_2995);
nand U5918 (N_5918,N_1083,N_3254);
and U5919 (N_5919,N_197,N_1873);
nand U5920 (N_5920,N_594,N_3955);
nand U5921 (N_5921,N_2543,N_907);
nand U5922 (N_5922,N_4735,N_1081);
and U5923 (N_5923,N_1711,N_1343);
xnor U5924 (N_5924,N_4265,N_0);
or U5925 (N_5925,N_4422,N_2802);
and U5926 (N_5926,N_1417,N_1162);
or U5927 (N_5927,N_2806,N_4388);
and U5928 (N_5928,N_3455,N_155);
nand U5929 (N_5929,N_3798,N_301);
xnor U5930 (N_5930,N_128,N_2318);
or U5931 (N_5931,N_3182,N_2410);
xor U5932 (N_5932,N_233,N_4582);
xor U5933 (N_5933,N_1028,N_3808);
and U5934 (N_5934,N_4941,N_900);
and U5935 (N_5935,N_3482,N_3736);
nand U5936 (N_5936,N_513,N_3796);
or U5937 (N_5937,N_370,N_3752);
nor U5938 (N_5938,N_4432,N_2499);
or U5939 (N_5939,N_3010,N_4318);
nand U5940 (N_5940,N_2627,N_2536);
nand U5941 (N_5941,N_1922,N_1630);
and U5942 (N_5942,N_4641,N_2563);
or U5943 (N_5943,N_3177,N_3962);
nor U5944 (N_5944,N_2884,N_3115);
and U5945 (N_5945,N_4555,N_431);
and U5946 (N_5946,N_1158,N_2729);
or U5947 (N_5947,N_1394,N_2731);
and U5948 (N_5948,N_614,N_116);
or U5949 (N_5949,N_1553,N_3949);
nor U5950 (N_5950,N_3183,N_378);
nand U5951 (N_5951,N_1046,N_2202);
nor U5952 (N_5952,N_738,N_1594);
or U5953 (N_5953,N_1118,N_3453);
or U5954 (N_5954,N_3327,N_2790);
or U5955 (N_5955,N_4572,N_561);
and U5956 (N_5956,N_2424,N_354);
and U5957 (N_5957,N_1888,N_3229);
xor U5958 (N_5958,N_4583,N_4097);
nand U5959 (N_5959,N_4440,N_2488);
and U5960 (N_5960,N_3731,N_1149);
or U5961 (N_5961,N_2864,N_4353);
xor U5962 (N_5962,N_3425,N_2894);
nor U5963 (N_5963,N_3690,N_1913);
xor U5964 (N_5964,N_3121,N_2501);
and U5965 (N_5965,N_456,N_3595);
nand U5966 (N_5966,N_704,N_28);
nand U5967 (N_5967,N_1863,N_2082);
and U5968 (N_5968,N_1574,N_3251);
and U5969 (N_5969,N_2449,N_1006);
nor U5970 (N_5970,N_273,N_3273);
or U5971 (N_5971,N_1468,N_111);
nand U5972 (N_5972,N_4643,N_3719);
nor U5973 (N_5973,N_2657,N_4077);
nand U5974 (N_5974,N_933,N_759);
and U5975 (N_5975,N_2723,N_2835);
nand U5976 (N_5976,N_2872,N_4515);
nor U5977 (N_5977,N_364,N_1018);
xor U5978 (N_5978,N_646,N_476);
or U5979 (N_5979,N_2607,N_1562);
nand U5980 (N_5980,N_4466,N_481);
nor U5981 (N_5981,N_3413,N_3107);
nor U5982 (N_5982,N_4907,N_4441);
xor U5983 (N_5983,N_562,N_4357);
or U5984 (N_5984,N_2915,N_25);
nand U5985 (N_5985,N_3643,N_487);
nand U5986 (N_5986,N_4769,N_1128);
nand U5987 (N_5987,N_3531,N_3701);
xnor U5988 (N_5988,N_2143,N_734);
nor U5989 (N_5989,N_2635,N_1808);
or U5990 (N_5990,N_2745,N_2978);
or U5991 (N_5991,N_2625,N_2164);
or U5992 (N_5992,N_4251,N_350);
or U5993 (N_5993,N_770,N_1497);
or U5994 (N_5994,N_2910,N_2871);
xnor U5995 (N_5995,N_4763,N_1676);
nand U5996 (N_5996,N_208,N_1390);
and U5997 (N_5997,N_3652,N_4306);
nand U5998 (N_5998,N_3803,N_3689);
or U5999 (N_5999,N_1790,N_3585);
and U6000 (N_6000,N_2434,N_239);
and U6001 (N_6001,N_1071,N_4290);
or U6002 (N_6002,N_3245,N_3761);
and U6003 (N_6003,N_3378,N_3022);
and U6004 (N_6004,N_1033,N_2206);
nand U6005 (N_6005,N_4311,N_3493);
nand U6006 (N_6006,N_4847,N_2154);
and U6007 (N_6007,N_1249,N_1626);
nor U6008 (N_6008,N_2656,N_1518);
or U6009 (N_6009,N_2285,N_2710);
or U6010 (N_6010,N_4202,N_4526);
nand U6011 (N_6011,N_2925,N_2485);
and U6012 (N_6012,N_4190,N_4324);
and U6013 (N_6013,N_1403,N_2599);
nand U6014 (N_6014,N_3220,N_1538);
nor U6015 (N_6015,N_524,N_806);
nand U6016 (N_6016,N_2024,N_677);
and U6017 (N_6017,N_3990,N_1440);
xor U6018 (N_6018,N_255,N_1466);
nor U6019 (N_6019,N_1524,N_3947);
nor U6020 (N_6020,N_4067,N_148);
nor U6021 (N_6021,N_2218,N_447);
or U6022 (N_6022,N_2976,N_2703);
xnor U6023 (N_6023,N_50,N_1500);
nor U6024 (N_6024,N_221,N_2265);
nand U6025 (N_6025,N_3958,N_423);
nand U6026 (N_6026,N_3197,N_3320);
or U6027 (N_6027,N_4768,N_127);
nand U6028 (N_6028,N_3790,N_3880);
and U6029 (N_6029,N_4887,N_2392);
nor U6030 (N_6030,N_3054,N_4571);
and U6031 (N_6031,N_4433,N_4184);
nor U6032 (N_6032,N_333,N_4273);
nor U6033 (N_6033,N_1811,N_2713);
and U6034 (N_6034,N_3277,N_2644);
and U6035 (N_6035,N_576,N_1886);
or U6036 (N_6036,N_3874,N_225);
and U6037 (N_6037,N_547,N_114);
and U6038 (N_6038,N_1866,N_2393);
or U6039 (N_6039,N_2541,N_995);
nand U6040 (N_6040,N_3766,N_2857);
nand U6041 (N_6041,N_1434,N_3017);
nor U6042 (N_6042,N_1782,N_57);
and U6043 (N_6043,N_4033,N_2115);
nand U6044 (N_6044,N_4749,N_4616);
nor U6045 (N_6045,N_1721,N_2431);
or U6046 (N_6046,N_2181,N_3981);
and U6047 (N_6047,N_1380,N_3787);
and U6048 (N_6048,N_4253,N_1054);
xor U6049 (N_6049,N_2048,N_3312);
or U6050 (N_6050,N_4419,N_3);
and U6051 (N_6051,N_3137,N_1590);
and U6052 (N_6052,N_2092,N_3820);
nor U6053 (N_6053,N_3269,N_1895);
and U6054 (N_6054,N_4497,N_2990);
or U6055 (N_6055,N_583,N_724);
nor U6056 (N_6056,N_999,N_1978);
nor U6057 (N_6057,N_3353,N_1931);
nor U6058 (N_6058,N_13,N_2592);
nand U6059 (N_6059,N_2355,N_648);
nor U6060 (N_6060,N_3924,N_3523);
xor U6061 (N_6061,N_3713,N_1282);
or U6062 (N_6062,N_3370,N_1159);
or U6063 (N_6063,N_664,N_4378);
or U6064 (N_6064,N_4705,N_1381);
or U6065 (N_6065,N_1936,N_4895);
or U6066 (N_6066,N_3330,N_4490);
and U6067 (N_6067,N_4207,N_3397);
or U6068 (N_6068,N_1928,N_4338);
nand U6069 (N_6069,N_721,N_1944);
and U6070 (N_6070,N_3779,N_1901);
or U6071 (N_6071,N_4412,N_480);
nor U6072 (N_6072,N_4970,N_3412);
nor U6073 (N_6073,N_3908,N_1996);
or U6074 (N_6074,N_1303,N_4560);
xnor U6075 (N_6075,N_1549,N_2294);
and U6076 (N_6076,N_2867,N_3549);
or U6077 (N_6077,N_4263,N_139);
and U6078 (N_6078,N_2373,N_2205);
nor U6079 (N_6079,N_445,N_444);
nor U6080 (N_6080,N_3150,N_1133);
and U6081 (N_6081,N_750,N_252);
xnor U6082 (N_6082,N_3040,N_4534);
and U6083 (N_6083,N_2338,N_3297);
or U6084 (N_6084,N_940,N_4987);
or U6085 (N_6085,N_726,N_4282);
or U6086 (N_6086,N_380,N_336);
nand U6087 (N_6087,N_3786,N_1858);
nand U6088 (N_6088,N_4246,N_4104);
nor U6089 (N_6089,N_774,N_880);
nor U6090 (N_6090,N_2168,N_2185);
or U6091 (N_6091,N_563,N_2927);
or U6092 (N_6092,N_3705,N_3602);
xor U6093 (N_6093,N_843,N_2391);
or U6094 (N_6094,N_4491,N_3203);
nand U6095 (N_6095,N_2768,N_4906);
or U6096 (N_6096,N_4662,N_3763);
nor U6097 (N_6097,N_668,N_618);
nand U6098 (N_6098,N_3464,N_3519);
or U6099 (N_6099,N_3466,N_22);
nand U6100 (N_6100,N_1300,N_4359);
nand U6101 (N_6101,N_675,N_4);
nand U6102 (N_6102,N_4867,N_1017);
nor U6103 (N_6103,N_4644,N_528);
nor U6104 (N_6104,N_491,N_4510);
nor U6105 (N_6105,N_3363,N_2679);
or U6106 (N_6106,N_4377,N_2288);
nand U6107 (N_6107,N_3655,N_1376);
xor U6108 (N_6108,N_2010,N_4484);
or U6109 (N_6109,N_4633,N_3897);
nand U6110 (N_6110,N_2832,N_4971);
nor U6111 (N_6111,N_2498,N_2241);
nor U6112 (N_6112,N_2176,N_1189);
or U6113 (N_6113,N_4059,N_538);
nor U6114 (N_6114,N_3394,N_3419);
and U6115 (N_6115,N_859,N_181);
nand U6116 (N_6116,N_1714,N_1921);
and U6117 (N_6117,N_1749,N_2513);
nand U6118 (N_6118,N_1129,N_1584);
nor U6119 (N_6119,N_3640,N_601);
or U6120 (N_6120,N_2153,N_4055);
xor U6121 (N_6121,N_3835,N_1252);
nand U6122 (N_6122,N_3083,N_1269);
nor U6123 (N_6123,N_1508,N_2346);
nor U6124 (N_6124,N_786,N_4408);
nand U6125 (N_6125,N_727,N_2609);
nand U6126 (N_6126,N_1671,N_4926);
nand U6127 (N_6127,N_2984,N_236);
nor U6128 (N_6128,N_4592,N_176);
nand U6129 (N_6129,N_2600,N_4738);
or U6130 (N_6130,N_543,N_776);
or U6131 (N_6131,N_1667,N_1570);
and U6132 (N_6132,N_59,N_1214);
nand U6133 (N_6133,N_327,N_3171);
and U6134 (N_6134,N_885,N_67);
and U6135 (N_6135,N_2425,N_243);
and U6136 (N_6136,N_3060,N_2691);
and U6137 (N_6137,N_4512,N_1034);
xnor U6138 (N_6138,N_1320,N_3446);
or U6139 (N_6139,N_4599,N_3617);
or U6140 (N_6140,N_861,N_3785);
nor U6141 (N_6141,N_2271,N_2071);
nand U6142 (N_6142,N_3319,N_58);
or U6143 (N_6143,N_985,N_3492);
or U6144 (N_6144,N_2824,N_651);
and U6145 (N_6145,N_2810,N_2688);
nand U6146 (N_6146,N_3503,N_1053);
xor U6147 (N_6147,N_660,N_1384);
or U6148 (N_6148,N_2299,N_4611);
and U6149 (N_6149,N_1920,N_659);
nor U6150 (N_6150,N_2040,N_1684);
and U6151 (N_6151,N_2928,N_3906);
xnor U6152 (N_6152,N_122,N_332);
or U6153 (N_6153,N_3362,N_39);
nand U6154 (N_6154,N_3506,N_4382);
xnor U6155 (N_6155,N_3340,N_2445);
or U6156 (N_6156,N_3872,N_2118);
or U6157 (N_6157,N_4084,N_725);
nor U6158 (N_6158,N_4391,N_2939);
and U6159 (N_6159,N_527,N_519);
and U6160 (N_6160,N_2332,N_1291);
nor U6161 (N_6161,N_3794,N_52);
and U6162 (N_6162,N_4462,N_3344);
nor U6163 (N_6163,N_1925,N_1194);
nand U6164 (N_6164,N_3887,N_1914);
nor U6165 (N_6165,N_1305,N_3913);
or U6166 (N_6166,N_4415,N_4803);
nor U6167 (N_6167,N_4943,N_2085);
nand U6168 (N_6168,N_567,N_1727);
or U6169 (N_6169,N_835,N_2532);
nor U6170 (N_6170,N_3684,N_3815);
nor U6171 (N_6171,N_4870,N_1288);
nor U6172 (N_6172,N_2741,N_1526);
nand U6173 (N_6173,N_2490,N_2378);
nand U6174 (N_6174,N_3937,N_2616);
xor U6175 (N_6175,N_4545,N_1122);
nor U6176 (N_6176,N_3647,N_3511);
nor U6177 (N_6177,N_4594,N_2298);
nand U6178 (N_6178,N_906,N_1898);
or U6179 (N_6179,N_4725,N_3861);
and U6180 (N_6180,N_3265,N_1509);
nand U6181 (N_6181,N_2022,N_3063);
and U6182 (N_6182,N_1119,N_1051);
or U6183 (N_6183,N_3261,N_4370);
nand U6184 (N_6184,N_2161,N_121);
nor U6185 (N_6185,N_3326,N_4425);
nor U6186 (N_6186,N_3995,N_4397);
nor U6187 (N_6187,N_161,N_2036);
and U6188 (N_6188,N_3867,N_1751);
nand U6189 (N_6189,N_2221,N_3295);
or U6190 (N_6190,N_935,N_3390);
and U6191 (N_6191,N_4275,N_1666);
nand U6192 (N_6192,N_2960,N_1107);
or U6193 (N_6193,N_76,N_2102);
nor U6194 (N_6194,N_1154,N_3873);
nand U6195 (N_6195,N_566,N_4312);
or U6196 (N_6196,N_4935,N_409);
nor U6197 (N_6197,N_2620,N_4453);
xor U6198 (N_6198,N_2861,N_981);
nand U6199 (N_6199,N_1223,N_2770);
and U6200 (N_6200,N_4595,N_2018);
nand U6201 (N_6201,N_1769,N_3770);
or U6202 (N_6202,N_1668,N_4498);
nand U6203 (N_6203,N_3839,N_4954);
nand U6204 (N_6204,N_1681,N_413);
nor U6205 (N_6205,N_3003,N_4262);
and U6206 (N_6206,N_2360,N_2842);
nor U6207 (N_6207,N_4132,N_4352);
and U6208 (N_6208,N_1349,N_3613);
nor U6209 (N_6209,N_2743,N_917);
or U6210 (N_6210,N_689,N_3555);
nor U6211 (N_6211,N_684,N_2456);
nand U6212 (N_6212,N_2095,N_3817);
nor U6213 (N_6213,N_533,N_105);
or U6214 (N_6214,N_3694,N_3176);
nor U6215 (N_6215,N_68,N_4567);
nor U6216 (N_6216,N_40,N_478);
nand U6217 (N_6217,N_2785,N_2287);
nand U6218 (N_6218,N_2948,N_2331);
or U6219 (N_6219,N_4604,N_494);
and U6220 (N_6220,N_719,N_32);
nand U6221 (N_6221,N_3833,N_4384);
nor U6222 (N_6222,N_4247,N_2268);
or U6223 (N_6223,N_4865,N_3299);
and U6224 (N_6224,N_946,N_4772);
or U6225 (N_6225,N_4025,N_2041);
nand U6226 (N_6226,N_132,N_2194);
nor U6227 (N_6227,N_3658,N_4584);
nor U6228 (N_6228,N_4101,N_222);
nand U6229 (N_6229,N_3035,N_504);
xor U6230 (N_6230,N_2451,N_214);
and U6231 (N_6231,N_846,N_142);
nand U6232 (N_6232,N_1199,N_588);
nor U6233 (N_6233,N_816,N_234);
nor U6234 (N_6234,N_1772,N_4051);
and U6235 (N_6235,N_2226,N_4603);
and U6236 (N_6236,N_2420,N_3544);
nand U6237 (N_6237,N_892,N_223);
nand U6238 (N_6238,N_518,N_3304);
nand U6239 (N_6239,N_2675,N_2875);
xnor U6240 (N_6240,N_989,N_3120);
nor U6241 (N_6241,N_4740,N_3853);
and U6242 (N_6242,N_4944,N_3301);
or U6243 (N_6243,N_1869,N_1114);
and U6244 (N_6244,N_4060,N_3611);
or U6245 (N_6245,N_3315,N_3350);
nor U6246 (N_6246,N_1264,N_188);
nand U6247 (N_6247,N_3149,N_3892);
and U6248 (N_6248,N_3151,N_4481);
and U6249 (N_6249,N_4979,N_854);
nand U6250 (N_6250,N_1539,N_4475);
or U6251 (N_6251,N_18,N_3272);
nand U6252 (N_6252,N_3890,N_2820);
nand U6253 (N_6253,N_1877,N_635);
nor U6254 (N_6254,N_2484,N_2940);
nand U6255 (N_6255,N_1164,N_732);
nor U6256 (N_6256,N_2711,N_3568);
nand U6257 (N_6257,N_4691,N_1370);
xnor U6258 (N_6258,N_3324,N_526);
nand U6259 (N_6259,N_3537,N_3064);
nor U6260 (N_6260,N_3476,N_3228);
nor U6261 (N_6261,N_1036,N_1364);
or U6262 (N_6262,N_1121,N_3951);
nand U6263 (N_6263,N_2457,N_3012);
or U6264 (N_6264,N_3373,N_1597);
nor U6265 (N_6265,N_4428,N_3859);
or U6266 (N_6266,N_2902,N_1616);
nand U6267 (N_6267,N_4707,N_4513);
or U6268 (N_6268,N_1393,N_1649);
or U6269 (N_6269,N_2060,N_3532);
nand U6270 (N_6270,N_2183,N_2336);
nand U6271 (N_6271,N_1950,N_1686);
nor U6272 (N_6272,N_2664,N_4220);
nor U6273 (N_6273,N_338,N_2602);
xor U6274 (N_6274,N_97,N_265);
and U6275 (N_6275,N_2959,N_1231);
or U6276 (N_6276,N_3207,N_4373);
or U6277 (N_6277,N_1482,N_387);
and U6278 (N_6278,N_1427,N_3066);
nor U6279 (N_6279,N_4836,N_388);
or U6280 (N_6280,N_1103,N_4807);
or U6281 (N_6281,N_4624,N_3308);
nor U6282 (N_6282,N_4659,N_807);
and U6283 (N_6283,N_3388,N_3616);
xor U6284 (N_6284,N_4593,N_3231);
or U6285 (N_6285,N_2941,N_1564);
nor U6286 (N_6286,N_809,N_3448);
or U6287 (N_6287,N_2495,N_261);
nor U6288 (N_6288,N_1475,N_3518);
nor U6289 (N_6289,N_3737,N_4309);
and U6290 (N_6290,N_4646,N_2523);
xor U6291 (N_6291,N_4729,N_2822);
or U6292 (N_6292,N_975,N_1377);
nor U6293 (N_6293,N_1739,N_3855);
and U6294 (N_6294,N_4136,N_1401);
nor U6295 (N_6295,N_1992,N_2526);
and U6296 (N_6296,N_1934,N_3932);
xnor U6297 (N_6297,N_2416,N_4591);
xor U6298 (N_6298,N_1704,N_175);
nand U6299 (N_6299,N_2235,N_1459);
or U6300 (N_6300,N_1503,N_2369);
or U6301 (N_6301,N_3612,N_286);
xor U6302 (N_6302,N_4334,N_323);
nor U6303 (N_6303,N_2341,N_2775);
and U6304 (N_6304,N_2913,N_340);
or U6305 (N_6305,N_913,N_1228);
or U6306 (N_6306,N_499,N_4454);
or U6307 (N_6307,N_2598,N_553);
nand U6308 (N_6308,N_4863,N_2962);
nor U6309 (N_6309,N_2020,N_3673);
nor U6310 (N_6310,N_3046,N_1741);
nor U6311 (N_6311,N_2415,N_402);
and U6312 (N_6312,N_3618,N_2730);
or U6313 (N_6313,N_4243,N_2137);
or U6314 (N_6314,N_65,N_3603);
or U6315 (N_6315,N_1642,N_2030);
nor U6316 (N_6316,N_2132,N_3741);
and U6317 (N_6317,N_956,N_3447);
nor U6318 (N_6318,N_183,N_4356);
and U6319 (N_6319,N_4028,N_949);
and U6320 (N_6320,N_4909,N_1496);
nand U6321 (N_6321,N_3274,N_700);
or U6322 (N_6322,N_3160,N_863);
or U6323 (N_6323,N_3424,N_3193);
xor U6324 (N_6324,N_53,N_4276);
or U6325 (N_6325,N_3260,N_1306);
or U6326 (N_6326,N_410,N_4126);
nor U6327 (N_6327,N_1692,N_2190);
xnor U6328 (N_6328,N_4234,N_4152);
or U6329 (N_6329,N_857,N_4061);
xor U6330 (N_6330,N_3783,N_2896);
or U6331 (N_6331,N_2593,N_747);
nand U6332 (N_6332,N_1618,N_2700);
or U6333 (N_6333,N_592,N_2825);
nor U6334 (N_6334,N_451,N_3636);
nand U6335 (N_6335,N_4030,N_1150);
xnor U6336 (N_6336,N_334,N_4889);
xor U6337 (N_6337,N_4100,N_3147);
nor U6338 (N_6338,N_1638,N_910);
nand U6339 (N_6339,N_2054,N_3800);
and U6340 (N_6340,N_202,N_1443);
nand U6341 (N_6341,N_2791,N_21);
nand U6342 (N_6342,N_302,N_541);
nor U6343 (N_6343,N_4576,N_2619);
nor U6344 (N_6344,N_329,N_3527);
nor U6345 (N_6345,N_4211,N_3325);
nor U6346 (N_6346,N_383,N_238);
or U6347 (N_6347,N_1254,N_1429);
nand U6348 (N_6348,N_3044,N_2908);
nand U6349 (N_6349,N_1731,N_577);
xnor U6350 (N_6350,N_38,N_4464);
or U6351 (N_6351,N_1586,N_876);
xor U6352 (N_6352,N_2566,N_1486);
or U6353 (N_6353,N_220,N_977);
nand U6354 (N_6354,N_497,N_2025);
and U6355 (N_6355,N_2505,N_2807);
or U6356 (N_6356,N_4781,N_3339);
and U6357 (N_6357,N_1715,N_3185);
and U6358 (N_6358,N_3923,N_2692);
or U6359 (N_6359,N_936,N_4457);
nor U6360 (N_6360,N_4286,N_2662);
nor U6361 (N_6361,N_2786,N_1641);
nand U6362 (N_6362,N_156,N_3417);
and U6363 (N_6363,N_991,N_2739);
and U6364 (N_6364,N_2136,N_1405);
or U6365 (N_6365,N_4689,N_3692);
nand U6366 (N_6366,N_2880,N_580);
and U6367 (N_6367,N_2773,N_3656);
nand U6368 (N_6368,N_1332,N_4965);
nand U6369 (N_6369,N_3234,N_360);
and U6370 (N_6370,N_187,N_1383);
nor U6371 (N_6371,N_2178,N_2042);
nand U6372 (N_6372,N_4163,N_1470);
or U6373 (N_6373,N_2981,N_2062);
nor U6374 (N_6374,N_3704,N_3143);
or U6375 (N_6375,N_3695,N_1732);
nor U6376 (N_6376,N_3317,N_1309);
xnor U6377 (N_6377,N_374,N_2150);
nor U6378 (N_6378,N_90,N_521);
and U6379 (N_6379,N_3333,N_4617);
nor U6380 (N_6380,N_3089,N_2549);
nand U6381 (N_6381,N_3372,N_3023);
or U6382 (N_6382,N_542,N_4091);
and U6383 (N_6383,N_4147,N_2525);
nor U6384 (N_6384,N_3776,N_4029);
or U6385 (N_6385,N_2441,N_4764);
xnor U6386 (N_6386,N_1425,N_3488);
or U6387 (N_6387,N_1095,N_2027);
nor U6388 (N_6388,N_3236,N_2281);
and U6389 (N_6389,N_1447,N_267);
nand U6390 (N_6390,N_2595,N_1203);
and U6391 (N_6391,N_1420,N_998);
nand U6392 (N_6392,N_1507,N_2160);
nand U6393 (N_6393,N_748,N_2119);
nor U6394 (N_6394,N_1200,N_2966);
and U6395 (N_6395,N_3769,N_718);
xor U6396 (N_6396,N_3172,N_2716);
xnor U6397 (N_6397,N_3832,N_20);
nor U6398 (N_6398,N_4647,N_3801);
and U6399 (N_6399,N_2837,N_3070);
and U6400 (N_6400,N_3998,N_2253);
nand U6401 (N_6401,N_2512,N_1104);
and U6402 (N_6402,N_4113,N_3180);
and U6403 (N_6403,N_4517,N_4444);
or U6404 (N_6404,N_2852,N_3486);
or U6405 (N_6405,N_2669,N_4342);
nand U6406 (N_6406,N_3896,N_976);
or U6407 (N_6407,N_4086,N_3106);
or U6408 (N_6408,N_3825,N_2698);
nand U6409 (N_6409,N_4811,N_1533);
nand U6410 (N_6410,N_574,N_948);
nor U6411 (N_6411,N_3259,N_670);
nand U6412 (N_6412,N_2157,N_2110);
nor U6413 (N_6413,N_2661,N_4758);
or U6414 (N_6414,N_2575,N_2706);
or U6415 (N_6415,N_628,N_3639);
and U6416 (N_6416,N_2885,N_4052);
and U6417 (N_6417,N_1995,N_3128);
nor U6418 (N_6418,N_4387,N_2798);
nor U6419 (N_6419,N_3777,N_1823);
nor U6420 (N_6420,N_1569,N_3461);
nor U6421 (N_6421,N_611,N_1908);
nand U6422 (N_6422,N_2648,N_2361);
nand U6423 (N_6423,N_3105,N_349);
xnor U6424 (N_6424,N_305,N_2672);
or U6425 (N_6425,N_4601,N_1442);
or U6426 (N_6426,N_1734,N_1137);
or U6427 (N_6427,N_530,N_1068);
nor U6428 (N_6428,N_3169,N_1043);
nand U6429 (N_6429,N_2021,N_1488);
nand U6430 (N_6430,N_3885,N_3666);
or U6431 (N_6431,N_263,N_2702);
or U6432 (N_6432,N_4628,N_2649);
xor U6433 (N_6433,N_3398,N_4443);
or U6434 (N_6434,N_4447,N_1881);
nand U6435 (N_6435,N_2614,N_3108);
nor U6436 (N_6436,N_4812,N_2503);
nor U6437 (N_6437,N_3374,N_4436);
or U6438 (N_6438,N_1449,N_1824);
and U6439 (N_6439,N_424,N_2237);
nor U6440 (N_6440,N_3263,N_452);
nor U6441 (N_6441,N_1016,N_1274);
or U6442 (N_6442,N_2849,N_2804);
nor U6443 (N_6443,N_1361,N_3903);
nor U6444 (N_6444,N_717,N_3540);
and U6445 (N_6445,N_4124,N_694);
or U6446 (N_6446,N_4069,N_800);
nand U6447 (N_6447,N_1131,N_979);
or U6448 (N_6448,N_3140,N_3781);
and U6449 (N_6449,N_2836,N_4149);
or U6450 (N_6450,N_2131,N_4903);
nand U6451 (N_6451,N_4605,N_2687);
nor U6452 (N_6452,N_4891,N_4626);
or U6453 (N_6453,N_2152,N_4531);
xnor U6454 (N_6454,N_1478,N_1397);
and U6455 (N_6455,N_4905,N_37);
nor U6456 (N_6456,N_4876,N_4530);
and U6457 (N_6457,N_113,N_2632);
nor U6458 (N_6458,N_1874,N_1887);
nor U6459 (N_6459,N_1672,N_1144);
nor U6460 (N_6460,N_1529,N_2811);
nor U6461 (N_6461,N_365,N_1779);
xor U6462 (N_6462,N_4547,N_502);
and U6463 (N_6463,N_2623,N_4018);
xnor U6464 (N_6464,N_2982,N_1255);
or U6465 (N_6465,N_2907,N_4904);
or U6466 (N_6466,N_1661,N_429);
or U6467 (N_6467,N_1728,N_472);
and U6468 (N_6468,N_385,N_2212);
xor U6469 (N_6469,N_3361,N_1335);
nand U6470 (N_6470,N_3369,N_170);
xnor U6471 (N_6471,N_3671,N_743);
and U6472 (N_6472,N_3730,N_1674);
xor U6473 (N_6473,N_3069,N_1247);
and U6474 (N_6474,N_845,N_3609);
or U6475 (N_6475,N_226,N_569);
and U6476 (N_6476,N_4355,N_3076);
nand U6477 (N_6477,N_2056,N_2238);
or U6478 (N_6478,N_1924,N_881);
nand U6479 (N_6479,N_75,N_353);
or U6480 (N_6480,N_924,N_466);
nor U6481 (N_6481,N_3627,N_3546);
xnor U6482 (N_6482,N_3517,N_4031);
or U6483 (N_6483,N_3275,N_30);
nand U6484 (N_6484,N_2878,N_460);
nor U6485 (N_6485,N_2765,N_2466);
nor U6486 (N_6486,N_959,N_3614);
xor U6487 (N_6487,N_1531,N_2838);
and U6488 (N_6488,N_836,N_4340);
nand U6489 (N_6489,N_4950,N_3925);
nor U6490 (N_6490,N_4090,N_3484);
and U6491 (N_6491,N_1609,N_2066);
nor U6492 (N_6492,N_926,N_4165);
nor U6493 (N_6493,N_1422,N_982);
nand U6494 (N_6494,N_2428,N_1789);
and U6495 (N_6495,N_2578,N_4094);
nand U6496 (N_6496,N_2506,N_171);
nand U6497 (N_6497,N_663,N_986);
nor U6498 (N_6498,N_146,N_2407);
nor U6499 (N_6499,N_960,N_2571);
or U6500 (N_6500,N_4808,N_4849);
nor U6501 (N_6501,N_4151,N_4002);
and U6502 (N_6502,N_277,N_362);
and U6503 (N_6503,N_564,N_4912);
or U6504 (N_6504,N_3485,N_3164);
nor U6505 (N_6505,N_2869,N_2439);
and U6506 (N_6506,N_4658,N_3688);
and U6507 (N_6507,N_2368,N_432);
and U6508 (N_6508,N_2208,N_712);
nand U6509 (N_6509,N_3734,N_1746);
nor U6510 (N_6510,N_2841,N_268);
xor U6511 (N_6511,N_441,N_888);
nor U6512 (N_6512,N_1719,N_4952);
xnor U6513 (N_6513,N_2816,N_135);
nor U6514 (N_6514,N_2076,N_3909);
xnor U6515 (N_6515,N_666,N_2047);
nand U6516 (N_6516,N_764,N_4552);
nor U6517 (N_6517,N_983,N_4872);
or U6518 (N_6518,N_2850,N_4489);
and U6519 (N_6519,N_4561,N_2236);
and U6520 (N_6520,N_1253,N_133);
nand U6521 (N_6521,N_4804,N_3759);
or U6522 (N_6522,N_2964,N_166);
nor U6523 (N_6523,N_1471,N_1759);
nor U6524 (N_6524,N_425,N_1177);
and U6525 (N_6525,N_3043,N_1127);
nand U6526 (N_6526,N_745,N_3132);
xnor U6527 (N_6527,N_3571,N_2266);
nor U6528 (N_6528,N_4040,N_2104);
nand U6529 (N_6529,N_761,N_818);
and U6530 (N_6530,N_1125,N_803);
xor U6531 (N_6531,N_4175,N_1105);
nor U6532 (N_6532,N_3968,N_4518);
and U6533 (N_6533,N_1142,N_1559);
and U6534 (N_6534,N_4213,N_2923);
or U6535 (N_6535,N_138,N_4511);
or U6536 (N_6536,N_1292,N_3316);
xor U6537 (N_6537,N_2251,N_3341);
nand U6538 (N_6538,N_4933,N_101);
or U6539 (N_6539,N_4785,N_2696);
nand U6540 (N_6540,N_484,N_1689);
and U6541 (N_6541,N_131,N_2819);
and U6542 (N_6542,N_864,N_2839);
nor U6543 (N_6543,N_1433,N_1826);
nand U6544 (N_6544,N_3037,N_4846);
and U6545 (N_6545,N_4036,N_2282);
xor U6546 (N_6546,N_2879,N_4360);
or U6547 (N_6547,N_366,N_3215);
nand U6548 (N_6548,N_4385,N_192);
and U6549 (N_6549,N_4527,N_459);
nand U6550 (N_6550,N_3516,N_883);
nand U6551 (N_6551,N_2367,N_1786);
nor U6552 (N_6552,N_822,N_1965);
xnor U6553 (N_6553,N_4532,N_194);
nand U6554 (N_6554,N_4474,N_3300);
or U6555 (N_6555,N_4883,N_2641);
or U6556 (N_6556,N_2311,N_3026);
nor U6557 (N_6557,N_4092,N_224);
and U6558 (N_6558,N_4493,N_4010);
nand U6559 (N_6559,N_2634,N_2189);
nand U6560 (N_6560,N_4139,N_1703);
and U6561 (N_6561,N_4343,N_2742);
or U6562 (N_6562,N_381,N_2784);
nand U6563 (N_6563,N_1233,N_2140);
nor U6564 (N_6564,N_118,N_1070);
xor U6565 (N_6565,N_1733,N_4748);
nand U6566 (N_6566,N_344,N_2756);
xor U6567 (N_6567,N_4929,N_4868);
nand U6568 (N_6568,N_517,N_1012);
nand U6569 (N_6569,N_1079,N_31);
xor U6570 (N_6570,N_1620,N_2830);
or U6571 (N_6571,N_4621,N_3279);
or U6572 (N_6572,N_3148,N_1327);
or U6573 (N_6573,N_709,N_1599);
nor U6574 (N_6574,N_2475,N_2796);
nand U6575 (N_6575,N_1077,N_1899);
nand U6576 (N_6576,N_1094,N_4308);
or U6577 (N_6577,N_749,N_3965);
nor U6578 (N_6578,N_2936,N_3371);
xor U6579 (N_6579,N_3653,N_3021);
nor U6580 (N_6580,N_4743,N_3586);
or U6581 (N_6581,N_358,N_869);
or U6582 (N_6582,N_2653,N_2868);
and U6583 (N_6583,N_1820,N_1840);
and U6584 (N_6584,N_3191,N_2659);
xnor U6585 (N_6585,N_4674,N_3738);
and U6586 (N_6586,N_4062,N_98);
nand U6587 (N_6587,N_723,N_1261);
and U6588 (N_6588,N_3929,N_496);
and U6589 (N_6589,N_2914,N_1726);
and U6590 (N_6590,N_1061,N_1700);
nand U6591 (N_6591,N_4317,N_4688);
or U6592 (N_6592,N_2304,N_2043);
nand U6593 (N_6593,N_1926,N_4796);
and U6594 (N_6594,N_1135,N_1373);
xor U6595 (N_6595,N_117,N_3772);
or U6596 (N_6596,N_2943,N_331);
and U6597 (N_6597,N_24,N_3294);
and U6598 (N_6598,N_4160,N_1008);
or U6599 (N_6599,N_3163,N_1537);
nor U6600 (N_6600,N_3159,N_4072);
nor U6601 (N_6601,N_1353,N_4853);
and U6602 (N_6602,N_41,N_3767);
nor U6603 (N_6603,N_4116,N_3375);
nor U6604 (N_6604,N_2359,N_2749);
or U6605 (N_6605,N_838,N_4372);
nor U6606 (N_6606,N_3296,N_474);
nand U6607 (N_6607,N_3645,N_4858);
or U6608 (N_6608,N_4837,N_1658);
nor U6609 (N_6609,N_1278,N_1585);
and U6610 (N_6610,N_4882,N_1514);
nor U6611 (N_6611,N_3365,N_3349);
nand U6612 (N_6612,N_4580,N_4261);
and U6613 (N_6613,N_3721,N_2780);
or U6614 (N_6614,N_716,N_3598);
nor U6615 (N_6615,N_2245,N_2647);
or U6616 (N_6616,N_4964,N_151);
and U6617 (N_6617,N_4256,N_1136);
nor U6618 (N_6618,N_1935,N_2727);
xnor U6619 (N_6619,N_1968,N_4505);
nor U6620 (N_6620,N_1456,N_2576);
nand U6621 (N_6621,N_490,N_1919);
nand U6622 (N_6622,N_3927,N_1657);
nor U6623 (N_6623,N_4820,N_1872);
or U6624 (N_6624,N_4351,N_4732);
nand U6625 (N_6625,N_4330,N_3474);
or U6626 (N_6626,N_184,N_4400);
nand U6627 (N_6627,N_3376,N_1832);
nand U6628 (N_6628,N_4609,N_4773);
nor U6629 (N_6629,N_2289,N_167);
nand U6630 (N_6630,N_4228,N_890);
nor U6631 (N_6631,N_657,N_2156);
and U6632 (N_6632,N_3740,N_1818);
and U6633 (N_6633,N_1987,N_3131);
or U6634 (N_6634,N_4579,N_1152);
xor U6635 (N_6635,N_2633,N_1854);
nor U6636 (N_6636,N_1679,N_1682);
nor U6637 (N_6637,N_4598,N_3243);
nor U6638 (N_6638,N_3849,N_3410);
or U6639 (N_6639,N_3624,N_3061);
and U6640 (N_6640,N_2983,N_2002);
nor U6641 (N_6641,N_2674,N_2552);
or U6642 (N_6642,N_537,N_4230);
and U6643 (N_6643,N_2182,N_753);
xor U6644 (N_6644,N_2099,N_4495);
or U6645 (N_6645,N_4719,N_608);
nor U6646 (N_6646,N_404,N_4158);
nor U6647 (N_6647,N_1691,N_4565);
and U6648 (N_6648,N_2735,N_4133);
and U6649 (N_6649,N_2258,N_2712);
or U6650 (N_6650,N_4670,N_4612);
nand U6651 (N_6651,N_2467,N_393);
nand U6652 (N_6652,N_1109,N_755);
xor U6653 (N_6653,N_3434,N_507);
xor U6654 (N_6654,N_3479,N_626);
and U6655 (N_6655,N_4066,N_867);
nand U6656 (N_6656,N_695,N_2579);
xnor U6657 (N_6657,N_205,N_1330);
or U6658 (N_6658,N_4430,N_1956);
and U6659 (N_6659,N_4291,N_4368);
nor U6660 (N_6660,N_3905,N_485);
xor U6661 (N_6661,N_964,N_4287);
nor U6662 (N_6662,N_3580,N_229);
and U6663 (N_6663,N_3700,N_3364);
and U6664 (N_6664,N_2933,N_699);
nand U6665 (N_6665,N_3864,N_3821);
nand U6666 (N_6666,N_925,N_1801);
or U6667 (N_6667,N_4523,N_3095);
xnor U6668 (N_6668,N_3392,N_3481);
and U6669 (N_6669,N_1157,N_3118);
nor U6670 (N_6670,N_2044,N_4586);
or U6671 (N_6671,N_922,N_1082);
xnor U6672 (N_6672,N_615,N_2992);
or U6673 (N_6673,N_1971,N_3706);
nor U6674 (N_6674,N_1424,N_4068);
xnor U6675 (N_6675,N_2353,N_2829);
and U6676 (N_6676,N_3632,N_575);
xnor U6677 (N_6677,N_2187,N_120);
nor U6678 (N_6678,N_3648,N_1991);
nor U6679 (N_6679,N_3762,N_2945);
nand U6680 (N_6680,N_201,N_2860);
and U6681 (N_6681,N_1272,N_3103);
nor U6682 (N_6682,N_1357,N_2695);
nor U6683 (N_6683,N_4936,N_4544);
xnor U6684 (N_6684,N_819,N_4239);
or U6685 (N_6685,N_312,N_149);
and U6686 (N_6686,N_3487,N_1830);
nor U6687 (N_6687,N_1052,N_638);
nand U6688 (N_6688,N_3901,N_4976);
nor U6689 (N_6689,N_1402,N_2073);
nand U6690 (N_6690,N_1219,N_363);
xor U6691 (N_6691,N_4456,N_4684);
xnor U6692 (N_6692,N_1575,N_130);
nand U6693 (N_6693,N_3583,N_3593);
and U6694 (N_6694,N_3205,N_417);
xor U6695 (N_6695,N_2684,N_1622);
nor U6696 (N_6696,N_3907,N_4915);
nor U6697 (N_6697,N_2577,N_3528);
or U6698 (N_6698,N_2023,N_3309);
and U6699 (N_6699,N_2167,N_3144);
nor U6700 (N_6700,N_555,N_1544);
or U6701 (N_6701,N_1108,N_4899);
or U6702 (N_6702,N_2586,N_2300);
nor U6703 (N_6703,N_411,N_3072);
or U6704 (N_6704,N_1540,N_824);
and U6705 (N_6705,N_3161,N_1918);
or U6706 (N_6706,N_2079,N_4451);
or U6707 (N_6707,N_3099,N_3020);
or U6708 (N_6708,N_1640,N_4345);
and U6709 (N_6709,N_1523,N_3943);
and U6710 (N_6710,N_45,N_1307);
xor U6711 (N_6711,N_930,N_1900);
and U6712 (N_6712,N_2203,N_1738);
nand U6713 (N_6713,N_1339,N_3404);
and U6714 (N_6714,N_1453,N_4955);
nand U6715 (N_6715,N_2091,N_802);
or U6716 (N_6716,N_3252,N_3217);
xnor U6717 (N_6717,N_1592,N_8);
nand U6718 (N_6718,N_4657,N_3812);
nand U6719 (N_6719,N_4640,N_1736);
or U6720 (N_6720,N_2363,N_593);
nand U6721 (N_6721,N_636,N_911);
or U6722 (N_6722,N_4779,N_3687);
nand U6723 (N_6723,N_1696,N_3950);
or U6724 (N_6724,N_2931,N_442);
or U6725 (N_6725,N_168,N_4314);
nor U6726 (N_6726,N_1432,N_3678);
nand U6727 (N_6727,N_3698,N_463);
nand U6728 (N_6728,N_828,N_2876);
nor U6729 (N_6729,N_681,N_4959);
and U6730 (N_6730,N_3104,N_2029);
or U6731 (N_6731,N_1143,N_1287);
nor U6732 (N_6732,N_1556,N_3042);
xor U6733 (N_6733,N_1860,N_2305);
and U6734 (N_6734,N_2337,N_1480);
nand U6735 (N_6735,N_1085,N_2778);
or U6736 (N_6736,N_4940,N_2216);
nand U6737 (N_6737,N_2916,N_4514);
xor U6738 (N_6738,N_1697,N_4934);
or U6739 (N_6739,N_1372,N_3087);
and U6740 (N_6740,N_4925,N_2542);
nor U6741 (N_6741,N_453,N_4866);
and U6742 (N_6742,N_2184,N_1634);
nand U6743 (N_6743,N_4529,N_4587);
or U6744 (N_6744,N_4575,N_1780);
xnor U6745 (N_6745,N_1763,N_4127);
nor U6746 (N_6746,N_4427,N_3067);
xor U6747 (N_6747,N_4300,N_1262);
and U6748 (N_6748,N_1773,N_172);
nand U6749 (N_6749,N_3264,N_3662);
nand U6750 (N_6750,N_4450,N_4873);
xnor U6751 (N_6751,N_4044,N_1548);
nor U6752 (N_6752,N_1990,N_4414);
nor U6753 (N_6753,N_1911,N_1939);
xor U6754 (N_6754,N_2301,N_4354);
and U6755 (N_6755,N_1445,N_1909);
and U6756 (N_6756,N_3084,N_2929);
nand U6757 (N_6757,N_4842,N_3240);
and U6758 (N_6758,N_4892,N_3860);
nand U6759 (N_6759,N_582,N_1115);
nand U6760 (N_6760,N_3837,N_2243);
or U6761 (N_6761,N_1983,N_2496);
nand U6762 (N_6762,N_1473,N_3535);
and U6763 (N_6763,N_163,N_3313);
nor U6764 (N_6764,N_1182,N_4623);
or U6765 (N_6765,N_1961,N_169);
xnor U6766 (N_6766,N_1250,N_3199);
xnor U6767 (N_6767,N_2162,N_3187);
nor U6768 (N_6768,N_3898,N_4399);
and U6769 (N_6769,N_3179,N_1221);
nand U6770 (N_6770,N_3454,N_4801);
or U6771 (N_6771,N_2074,N_1966);
and U6772 (N_6772,N_1797,N_3850);
xnor U6773 (N_6773,N_4776,N_3173);
nand U6774 (N_6774,N_506,N_3714);
nand U6775 (N_6775,N_3802,N_3754);
nand U6776 (N_6776,N_4268,N_1351);
xor U6777 (N_6777,N_4369,N_2794);
nor U6778 (N_6778,N_2895,N_3230);
nand U6779 (N_6779,N_4697,N_3335);
and U6780 (N_6780,N_1955,N_7);
nor U6781 (N_6781,N_2033,N_2963);
xnor U6782 (N_6782,N_2382,N_107);
and U6783 (N_6783,N_1669,N_2011);
and U6784 (N_6784,N_3723,N_3239);
or U6785 (N_6785,N_3469,N_4919);
nand U6786 (N_6786,N_468,N_216);
and U6787 (N_6787,N_1294,N_2274);
nor U6788 (N_6788,N_1964,N_2900);
nor U6789 (N_6789,N_4692,N_276);
nor U6790 (N_6790,N_398,N_914);
nor U6791 (N_6791,N_4248,N_2263);
nor U6792 (N_6792,N_932,N_1740);
nand U6793 (N_6793,N_4948,N_662);
nor U6794 (N_6794,N_2229,N_4242);
xnor U6795 (N_6795,N_126,N_4316);
xor U6796 (N_6796,N_650,N_4949);
or U6797 (N_6797,N_4696,N_4744);
nor U6798 (N_6798,N_3059,N_2116);
or U6799 (N_6799,N_4439,N_644);
nand U6800 (N_6800,N_3868,N_4349);
nand U6801 (N_6801,N_2919,N_1145);
and U6802 (N_6802,N_125,N_3994);
nor U6803 (N_6803,N_2329,N_3845);
nand U6804 (N_6804,N_2514,N_2310);
nand U6805 (N_6805,N_2681,N_1975);
nand U6806 (N_6806,N_4038,N_3495);
and U6807 (N_6807,N_2491,N_1605);
or U6808 (N_6808,N_4753,N_941);
or U6809 (N_6809,N_3247,N_3979);
or U6810 (N_6810,N_2120,N_3209);
and U6811 (N_6811,N_4678,N_1419);
and U6812 (N_6812,N_3088,N_1436);
or U6813 (N_6813,N_3592,N_3226);
and U6814 (N_6814,N_833,N_589);
nand U6815 (N_6815,N_1906,N_1941);
or U6816 (N_6816,N_1814,N_2881);
nor U6817 (N_6817,N_3559,N_2590);
nand U6818 (N_6818,N_1716,N_1962);
xor U6819 (N_6819,N_1359,N_3910);
or U6820 (N_6820,N_2097,N_373);
or U6821 (N_6821,N_3608,N_1839);
xnor U6822 (N_6822,N_771,N_4859);
nand U6823 (N_6823,N_1333,N_357);
nand U6824 (N_6824,N_1494,N_796);
xnor U6825 (N_6825,N_4494,N_3079);
and U6826 (N_6826,N_3722,N_2515);
and U6827 (N_6827,N_4588,N_2565);
and U6828 (N_6828,N_3047,N_4021);
xnor U6829 (N_6829,N_4150,N_4057);
nor U6830 (N_6830,N_2561,N_821);
xnor U6831 (N_6831,N_3405,N_1566);
and U6832 (N_6832,N_4503,N_1752);
nor U6833 (N_6833,N_1102,N_2322);
nand U6834 (N_6834,N_1407,N_957);
and U6835 (N_6835,N_4819,N_3870);
and U6836 (N_6836,N_392,N_2718);
nor U6837 (N_6837,N_1907,N_1091);
nand U6838 (N_6838,N_92,N_119);
xor U6839 (N_6839,N_4554,N_3460);
and U6840 (N_6840,N_605,N_3062);
xor U6841 (N_6841,N_2053,N_4841);
nor U6842 (N_6842,N_3162,N_3382);
nand U6843 (N_6843,N_3823,N_3573);
or U6844 (N_6844,N_4701,N_4974);
or U6845 (N_6845,N_2387,N_3539);
or U6846 (N_6846,N_3311,N_4680);
xnor U6847 (N_6847,N_1280,N_3607);
nand U6848 (N_6848,N_3307,N_1323);
nand U6849 (N_6849,N_2533,N_2362);
and U6850 (N_6850,N_1943,N_3982);
and U6851 (N_6851,N_1168,N_3478);
nand U6852 (N_6852,N_4528,N_2009);
and U6853 (N_6853,N_2222,N_1234);
nand U6854 (N_6854,N_1399,N_271);
or U6855 (N_6855,N_915,N_310);
or U6856 (N_6856,N_3708,N_3869);
and U6857 (N_6857,N_2112,N_2787);
nor U6858 (N_6858,N_4946,N_3852);
and U6859 (N_6859,N_3715,N_945);
nand U6860 (N_6860,N_4145,N_3192);
nand U6861 (N_6861,N_3735,N_2603);
nor U6862 (N_6862,N_1972,N_2286);
and U6863 (N_6863,N_1717,N_871);
xor U6864 (N_6864,N_4710,N_968);
nand U6865 (N_6865,N_2961,N_1271);
xnor U6866 (N_6866,N_1067,N_2946);
and U6867 (N_6867,N_1186,N_4468);
and U6868 (N_6868,N_1050,N_3650);
nor U6869 (N_6869,N_4736,N_4995);
or U6870 (N_6870,N_3882,N_652);
or U6871 (N_6871,N_4098,N_3589);
nor U6872 (N_6872,N_4115,N_4206);
or U6873 (N_6873,N_3456,N_408);
nor U6874 (N_6874,N_207,N_1215);
xor U6875 (N_6875,N_1834,N_2100);
and U6876 (N_6876,N_473,N_3189);
nor U6877 (N_6877,N_206,N_368);
and U6878 (N_6878,N_2414,N_850);
or U6879 (N_6879,N_1504,N_3989);
and U6880 (N_6880,N_4424,N_4901);
nor U6881 (N_6881,N_4250,N_1598);
nand U6882 (N_6882,N_4975,N_3709);
xor U6883 (N_6883,N_2452,N_4911);
nand U6884 (N_6884,N_2134,N_1205);
xnor U6885 (N_6885,N_4418,N_470);
or U6886 (N_6886,N_2799,N_653);
nand U6887 (N_6887,N_3457,N_3400);
nand U6888 (N_6888,N_2314,N_4890);
and U6889 (N_6889,N_584,N_1492);
xnor U6890 (N_6890,N_2421,N_61);
nor U6891 (N_6891,N_3562,N_3862);
or U6892 (N_6892,N_2169,N_1000);
nor U6893 (N_6893,N_3081,N_2606);
xnor U6894 (N_6894,N_351,N_1756);
nand U6895 (N_6895,N_1952,N_2866);
nor U6896 (N_6896,N_2013,N_1099);
nor U6897 (N_6897,N_462,N_1374);
nor U6898 (N_6898,N_4226,N_3984);
and U6899 (N_6899,N_2678,N_3039);
and U6900 (N_6900,N_3993,N_912);
and U6901 (N_6901,N_1362,N_4392);
and U6902 (N_6902,N_2055,N_4799);
or U6903 (N_6903,N_3756,N_4254);
or U6904 (N_6904,N_2920,N_1851);
nor U6905 (N_6905,N_1001,N_1078);
nand U6906 (N_6906,N_3415,N_2862);
or U6907 (N_6907,N_889,N_3536);
nand U6908 (N_6908,N_1821,N_1124);
nor U6909 (N_6909,N_4109,N_783);
and U6910 (N_6910,N_516,N_4106);
and U6911 (N_6911,N_762,N_1662);
nor U6912 (N_6912,N_3094,N_958);
nand U6913 (N_6913,N_706,N_1297);
nand U6914 (N_6914,N_830,N_4008);
and U6915 (N_6915,N_210,N_3343);
or U6916 (N_6916,N_219,N_923);
nand U6917 (N_6917,N_2709,N_4264);
nand U6918 (N_6918,N_235,N_1520);
or U6919 (N_6919,N_4293,N_3992);
or U6920 (N_6920,N_4108,N_4875);
or U6921 (N_6921,N_4488,N_1517);
and U6922 (N_6922,N_1153,N_4968);
nor U6923 (N_6923,N_2348,N_928);
and U6924 (N_6924,N_279,N_321);
and U6925 (N_6925,N_3178,N_1951);
nand U6926 (N_6926,N_2979,N_673);
and U6927 (N_6927,N_3865,N_2877);
and U6928 (N_6928,N_493,N_1316);
nand U6929 (N_6929,N_1342,N_973);
and U6930 (N_6930,N_1138,N_4042);
and U6931 (N_6931,N_292,N_2454);
xor U6932 (N_6932,N_2371,N_1862);
or U6933 (N_6933,N_356,N_2186);
nand U6934 (N_6934,N_4022,N_274);
or U6935 (N_6935,N_2471,N_4632);
nor U6936 (N_6936,N_4648,N_3775);
and U6937 (N_6937,N_1166,N_1521);
or U6938 (N_6938,N_3489,N_1169);
nor U6939 (N_6939,N_1923,N_2019);
or U6940 (N_6940,N_1815,N_2486);
nor U6941 (N_6941,N_1747,N_2061);
nand U6942 (N_6942,N_4267,N_4631);
nand U6943 (N_6943,N_4167,N_2094);
nand U6944 (N_6944,N_1371,N_2924);
and U6945 (N_6945,N_500,N_1015);
or U6946 (N_6946,N_2834,N_4194);
or U6947 (N_6947,N_4405,N_4231);
nand U6948 (N_6948,N_937,N_768);
or U6949 (N_6949,N_604,N_3306);
nand U6950 (N_6950,N_3459,N_4478);
nand U6951 (N_6951,N_253,N_1600);
and U6952 (N_6952,N_2083,N_4780);
and U6953 (N_6953,N_1404,N_2395);
nand U6954 (N_6954,N_3899,N_1302);
or U6955 (N_6955,N_3408,N_2279);
and U6956 (N_6956,N_3646,N_4155);
nor U6957 (N_6957,N_619,N_2517);
nand U6958 (N_6958,N_967,N_3281);
xnor U6959 (N_6959,N_4236,N_4174);
or U6960 (N_6960,N_3386,N_2350);
xor U6961 (N_6961,N_3428,N_3729);
nand U6962 (N_6962,N_3298,N_4747);
nor U6963 (N_6963,N_1643,N_2342);
or U6964 (N_6964,N_1693,N_4830);
nand U6965 (N_6965,N_1833,N_1037);
nor U6966 (N_6966,N_4178,N_1426);
and U6967 (N_6967,N_1663,N_2705);
nand U6968 (N_6968,N_2250,N_2356);
or U6969 (N_6969,N_2846,N_3919);
nand U6970 (N_6970,N_4292,N_3435);
nand U6971 (N_6971,N_2988,N_3572);
or U6972 (N_6972,N_3314,N_4073);
nor U6973 (N_6973,N_4119,N_3016);
nor U6974 (N_6974,N_4362,N_4777);
or U6975 (N_6975,N_1846,N_3912);
nor U6976 (N_6976,N_4431,N_2155);
or U6977 (N_6977,N_2763,N_352);
or U6978 (N_6978,N_3999,N_4845);
and U6979 (N_6979,N_756,N_2255);
and U6980 (N_6980,N_3480,N_343);
xor U6981 (N_6981,N_2938,N_230);
or U6982 (N_6982,N_855,N_1541);
xor U6983 (N_6983,N_4942,N_4553);
xor U6984 (N_6984,N_397,N_454);
nand U6985 (N_6985,N_2958,N_4089);
nor U6986 (N_6986,N_2364,N_620);
or U6987 (N_6987,N_1392,N_2934);
nand U6988 (N_6988,N_1505,N_1511);
nand U6989 (N_6989,N_1243,N_3556);
nand U6990 (N_6990,N_4045,N_2172);
nand U6991 (N_6991,N_1791,N_4011);
xor U6992 (N_6992,N_1441,N_2482);
nand U6993 (N_6993,N_2685,N_4154);
nor U6994 (N_6994,N_371,N_2760);
and U6995 (N_6995,N_3524,N_1146);
nand U6996 (N_6996,N_4380,N_2774);
or U6997 (N_6997,N_93,N_4093);
nor U6998 (N_6998,N_2351,N_174);
nand U6999 (N_6999,N_1552,N_3797);
and U7000 (N_7000,N_2789,N_4654);
nor U7001 (N_7001,N_3142,N_1695);
xnor U7002 (N_7002,N_2418,N_4114);
and U7003 (N_7003,N_3765,N_4166);
nand U7004 (N_7004,N_1765,N_3515);
and U7005 (N_7005,N_3788,N_1836);
xor U7006 (N_7006,N_4118,N_304);
nand U7007 (N_7007,N_3622,N_1010);
and U7008 (N_7008,N_3847,N_3748);
and U7009 (N_7009,N_4810,N_2886);
nor U7010 (N_7010,N_2072,N_1212);
and U7011 (N_7011,N_245,N_83);
nand U7012 (N_7012,N_2309,N_2676);
and U7013 (N_7013,N_1632,N_514);
or U7014 (N_7014,N_1589,N_532);
and U7015 (N_7015,N_1251,N_3691);
and U7016 (N_7016,N_751,N_779);
nand U7017 (N_7017,N_4914,N_29);
or U7018 (N_7018,N_4833,N_1829);
nand U7019 (N_7019,N_1448,N_4752);
xor U7020 (N_7020,N_3780,N_458);
nor U7021 (N_7021,N_1382,N_1572);
or U7022 (N_7022,N_3098,N_322);
nor U7023 (N_7023,N_4549,N_4313);
or U7024 (N_7024,N_1864,N_1363);
nor U7025 (N_7025,N_3676,N_4999);
nor U7026 (N_7026,N_4204,N_1614);
xnor U7027 (N_7027,N_4302,N_2151);
or U7028 (N_7028,N_346,N_897);
nand U7029 (N_7029,N_944,N_1209);
nor U7030 (N_7030,N_1156,N_1813);
or U7031 (N_7031,N_4070,N_886);
or U7032 (N_7032,N_3914,N_4459);
or U7033 (N_7033,N_1892,N_96);
or U7034 (N_7034,N_1942,N_4679);
nor U7035 (N_7035,N_1113,N_266);
nand U7036 (N_7036,N_3570,N_2249);
and U7037 (N_7037,N_3726,N_3591);
nor U7038 (N_7038,N_3969,N_2293);
or U7039 (N_7039,N_1225,N_382);
or U7040 (N_7040,N_2063,N_2198);
nor U7041 (N_7041,N_4618,N_627);
and U7042 (N_7042,N_4083,N_4183);
or U7043 (N_7043,N_4985,N_2985);
or U7044 (N_7044,N_4824,N_685);
nand U7045 (N_7045,N_2443,N_418);
nand U7046 (N_7046,N_4266,N_581);
and U7047 (N_7047,N_4081,N_4602);
nor U7048 (N_7048,N_1213,N_2944);
and U7049 (N_7049,N_741,N_2248);
and U7050 (N_7050,N_4015,N_337);
or U7051 (N_7051,N_1075,N_1817);
nor U7052 (N_7052,N_2509,N_1464);
and U7053 (N_7053,N_4559,N_3746);
and U7054 (N_7054,N_3718,N_4000);
or U7055 (N_7055,N_4047,N_4046);
or U7056 (N_7056,N_3750,N_3310);
nand U7057 (N_7057,N_4724,N_3471);
xor U7058 (N_7058,N_4502,N_2039);
nor U7059 (N_7059,N_2444,N_2757);
xnor U7060 (N_7060,N_1002,N_3280);
nor U7061 (N_7061,N_795,N_4521);
or U7062 (N_7062,N_2057,N_1960);
nand U7063 (N_7063,N_4850,N_2683);
nor U7064 (N_7064,N_972,N_2682);
nor U7065 (N_7065,N_4509,N_2108);
nand U7066 (N_7066,N_3960,N_1126);
nand U7067 (N_7067,N_990,N_4192);
nor U7068 (N_7068,N_3773,N_1020);
nand U7069 (N_7069,N_966,N_4043);
nand U7070 (N_7070,N_1499,N_882);
nand U7071 (N_7071,N_1932,N_3096);
nand U7072 (N_7072,N_3048,N_3157);
xor U7073 (N_7073,N_2772,N_969);
and U7074 (N_7074,N_1206,N_3553);
or U7075 (N_7075,N_48,N_4923);
and U7076 (N_7076,N_1861,N_421);
or U7077 (N_7077,N_4928,N_2064);
and U7078 (N_7078,N_4289,N_2422);
and U7079 (N_7079,N_2500,N_4877);
or U7080 (N_7080,N_1412,N_1167);
nand U7081 (N_7081,N_4404,N_2497);
nand U7082 (N_7082,N_2870,N_1571);
nand U7083 (N_7083,N_3575,N_4471);
xor U7084 (N_7084,N_3367,N_2954);
nand U7085 (N_7085,N_4650,N_1431);
or U7086 (N_7086,N_3973,N_2075);
nand U7087 (N_7087,N_372,N_587);
or U7088 (N_7088,N_3625,N_4742);
and U7089 (N_7089,N_1678,N_2720);
nor U7090 (N_7090,N_3953,N_1753);
and U7091 (N_7091,N_4469,N_2612);
nand U7092 (N_7092,N_3465,N_2769);
nor U7093 (N_7093,N_1687,N_1398);
and U7094 (N_7094,N_3542,N_637);
nor U7095 (N_7095,N_4238,N_2510);
or U7096 (N_7096,N_2330,N_4878);
nand U7097 (N_7097,N_4141,N_4848);
nor U7098 (N_7098,N_2290,N_2122);
or U7099 (N_7099,N_2694,N_3015);
nand U7100 (N_7100,N_3153,N_2400);
and U7101 (N_7101,N_3577,N_359);
nor U7102 (N_7102,N_3348,N_315);
xnor U7103 (N_7103,N_3961,N_3977);
xnor U7104 (N_7104,N_3114,N_1933);
and U7105 (N_7105,N_2306,N_2572);
nand U7106 (N_7106,N_278,N_396);
and U7107 (N_7107,N_4455,N_617);
nand U7108 (N_7108,N_769,N_3125);
and U7109 (N_7109,N_1579,N_3498);
nor U7110 (N_7110,N_1237,N_2477);
xor U7111 (N_7111,N_3996,N_2689);
nand U7112 (N_7112,N_4063,N_3468);
or U7113 (N_7113,N_1501,N_4079);
and U7114 (N_7114,N_3533,N_711);
nor U7115 (N_7115,N_2617,N_1191);
xor U7116 (N_7116,N_2585,N_2942);
or U7117 (N_7117,N_3623,N_2219);
or U7118 (N_7118,N_2738,N_4937);
nor U7119 (N_7119,N_2562,N_4508);
nand U7120 (N_7120,N_69,N_4187);
or U7121 (N_7121,N_2534,N_2384);
or U7122 (N_7122,N_595,N_3778);
xnor U7123 (N_7123,N_3334,N_4977);
nor U7124 (N_7124,N_2814,N_3538);
and U7125 (N_7125,N_320,N_3041);
nor U7126 (N_7126,N_4741,N_144);
nand U7127 (N_7127,N_1857,N_814);
nand U7128 (N_7128,N_3139,N_3818);
nor U7129 (N_7129,N_2645,N_4834);
and U7130 (N_7130,N_4244,N_794);
nor U7131 (N_7131,N_1720,N_2149);
or U7132 (N_7132,N_672,N_3357);
nand U7133 (N_7133,N_4800,N_1798);
nand U7134 (N_7134,N_1596,N_894);
or U7135 (N_7135,N_1048,N_4327);
xor U7136 (N_7136,N_1837,N_2737);
or U7137 (N_7137,N_4056,N_70);
nor U7138 (N_7138,N_2479,N_4714);
nand U7139 (N_7139,N_2690,N_4017);
nor U7140 (N_7140,N_4499,N_1799);
and U7141 (N_7141,N_4606,N_596);
nor U7142 (N_7142,N_4078,N_4014);
or U7143 (N_7143,N_1066,N_4027);
nand U7144 (N_7144,N_2123,N_2751);
or U7145 (N_7145,N_2708,N_2795);
and U7146 (N_7146,N_394,N_1805);
or U7147 (N_7147,N_996,N_3665);
or U7148 (N_7148,N_1871,N_1093);
and U7149 (N_7149,N_4978,N_4088);
nand U7150 (N_7150,N_1591,N_2686);
and U7151 (N_7151,N_3507,N_4806);
nand U7152 (N_7152,N_3381,N_1313);
and U7153 (N_7153,N_868,N_4823);
nand U7154 (N_7154,N_1917,N_2733);
and U7155 (N_7155,N_1024,N_2597);
nor U7156 (N_7156,N_3005,N_2465);
nor U7157 (N_7157,N_1161,N_4835);
nand U7158 (N_7158,N_4020,N_2574);
nand U7159 (N_7159,N_997,N_832);
or U7160 (N_7160,N_1912,N_4284);
nor U7161 (N_7161,N_4138,N_2317);
nor U7162 (N_7162,N_4687,N_4445);
or U7163 (N_7163,N_115,N_1611);
nor U7164 (N_7164,N_616,N_195);
or U7165 (N_7165,N_4550,N_4930);
and U7166 (N_7166,N_785,N_1757);
and U7167 (N_7167,N_3496,N_3360);
and U7168 (N_7168,N_4564,N_1304);
xor U7169 (N_7169,N_3433,N_1648);
and U7170 (N_7170,N_2613,N_1244);
or U7171 (N_7171,N_1485,N_2991);
or U7172 (N_7172,N_1289,N_4927);
or U7173 (N_7173,N_4423,N_1683);
and U7174 (N_7174,N_108,N_1792);
or U7175 (N_7175,N_1654,N_3212);
nand U7176 (N_7176,N_4716,N_2034);
nor U7177 (N_7177,N_1771,N_2442);
and U7178 (N_7178,N_2654,N_2436);
or U7179 (N_7179,N_4573,N_1352);
nor U7180 (N_7180,N_3510,N_129);
nand U7181 (N_7181,N_324,N_3543);
nand U7182 (N_7182,N_3075,N_3716);
nand U7183 (N_7183,N_3009,N_4831);
nor U7184 (N_7184,N_607,N_2096);
and U7185 (N_7185,N_2483,N_2734);
or U7186 (N_7186,N_1230,N_3055);
or U7187 (N_7187,N_1439,N_464);
nor U7188 (N_7188,N_2975,N_4102);
nor U7189 (N_7189,N_1677,N_110);
nor U7190 (N_7190,N_3651,N_299);
or U7191 (N_7191,N_2130,N_2540);
xor U7192 (N_7192,N_501,N_752);
nor U7193 (N_7193,N_2817,N_2801);
and U7194 (N_7194,N_3581,N_1625);
or U7195 (N_7195,N_227,N_3728);
nand U7196 (N_7196,N_2084,N_446);
nor U7197 (N_7197,N_2604,N_4795);
or U7198 (N_7198,N_1822,N_4177);
nand U7199 (N_7199,N_2558,N_4967);
nor U7200 (N_7200,N_4788,N_2965);
or U7201 (N_7201,N_2379,N_1659);
xnor U7202 (N_7202,N_3574,N_403);
or U7203 (N_7203,N_2972,N_3749);
nor U7204 (N_7204,N_2058,N_4754);
and U7205 (N_7205,N_1004,N_1937);
and U7206 (N_7206,N_3276,N_1391);
nand U7207 (N_7207,N_4272,N_391);
or U7208 (N_7208,N_3529,N_2993);
xor U7209 (N_7209,N_4270,N_2193);
nand U7210 (N_7210,N_2909,N_600);
nor U7211 (N_7211,N_529,N_862);
nand U7212 (N_7212,N_2417,N_3615);
xor U7213 (N_7213,N_4551,N_4694);
nor U7214 (N_7214,N_1172,N_4107);
or U7215 (N_7215,N_4681,N_1347);
and U7216 (N_7216,N_2419,N_178);
and U7217 (N_7217,N_773,N_1490);
or U7218 (N_7218,N_240,N_2630);
and U7219 (N_7219,N_4315,N_2280);
xor U7220 (N_7220,N_4480,N_1997);
and U7221 (N_7221,N_1098,N_4981);
nand U7222 (N_7222,N_4524,N_1418);
or U7223 (N_7223,N_3895,N_4417);
nor U7224 (N_7224,N_4429,N_1958);
nor U7225 (N_7225,N_3871,N_4071);
nor U7226 (N_7226,N_335,N_3127);
nor U7227 (N_7227,N_3452,N_4087);
nand U7228 (N_7228,N_3354,N_4675);
nor U7229 (N_7229,N_4615,N_3521);
and U7230 (N_7230,N_1038,N_2321);
nor U7231 (N_7231,N_909,N_735);
nor U7232 (N_7232,N_1865,N_2596);
and U7233 (N_7233,N_1454,N_1985);
or U7234 (N_7234,N_3807,N_2450);
nor U7235 (N_7235,N_1069,N_3155);
xor U7236 (N_7236,N_4539,N_2969);
or U7237 (N_7237,N_4319,N_2901);
and U7238 (N_7238,N_2347,N_2385);
and U7239 (N_7239,N_4569,N_4782);
and U7240 (N_7240,N_26,N_4775);
nor U7241 (N_7241,N_4931,N_2195);
and U7242 (N_7242,N_23,N_4727);
and U7243 (N_7243,N_14,N_1322);
or U7244 (N_7244,N_3477,N_4209);
or U7245 (N_7245,N_929,N_4161);
and U7246 (N_7246,N_4435,N_1635);
nand U7247 (N_7247,N_2548,N_3891);
or U7248 (N_7248,N_3111,N_4195);
nand U7249 (N_7249,N_4229,N_3282);
and U7250 (N_7250,N_3564,N_2276);
nand U7251 (N_7251,N_4721,N_520);
and U7252 (N_7252,N_54,N_190);
and U7253 (N_7253,N_2006,N_1573);
and U7254 (N_7254,N_1029,N_4039);
or U7255 (N_7255,N_4794,N_837);
and U7256 (N_7256,N_4337,N_4298);
nand U7257 (N_7257,N_1515,N_4065);
or U7258 (N_7258,N_2114,N_3331);
xor U7259 (N_7259,N_4570,N_3241);
or U7260 (N_7260,N_1141,N_2210);
and U7261 (N_7261,N_450,N_3395);
nor U7262 (N_7262,N_872,N_2323);
xnor U7263 (N_7263,N_3385,N_4082);
nand U7264 (N_7264,N_4224,N_147);
nand U7265 (N_7265,N_4364,N_3952);
and U7266 (N_7266,N_461,N_3109);
or U7267 (N_7267,N_3659,N_3244);
nand U7268 (N_7268,N_934,N_4709);
and U7269 (N_7269,N_2147,N_4295);
nand U7270 (N_7270,N_3204,N_3828);
nor U7271 (N_7271,N_3768,N_12);
nand U7272 (N_7272,N_294,N_2897);
and U7273 (N_7273,N_4951,N_1512);
and U7274 (N_7274,N_4375,N_3318);
nand U7275 (N_7275,N_4817,N_2390);
nor U7276 (N_7276,N_551,N_2142);
and U7277 (N_7277,N_4075,N_3789);
nor U7278 (N_7278,N_4525,N_2952);
and U7279 (N_7279,N_4784,N_3707);
and U7280 (N_7280,N_1742,N_1855);
and U7281 (N_7281,N_2325,N_140);
nand U7282 (N_7282,N_2242,N_3674);
xnor U7283 (N_7283,N_2402,N_439);
xnor U7284 (N_7284,N_4325,N_3843);
nand U7285 (N_7285,N_4672,N_2175);
and U7286 (N_7286,N_1688,N_4869);
nor U7287 (N_7287,N_1498,N_4713);
or U7288 (N_7288,N_3152,N_4636);
and U7289 (N_7289,N_902,N_16);
nand U7290 (N_7290,N_4128,N_19);
xor U7291 (N_7291,N_4723,N_2427);
nand U7292 (N_7292,N_3092,N_1581);
or U7293 (N_7293,N_1389,N_4064);
or U7294 (N_7294,N_4240,N_3830);
or U7295 (N_7295,N_2622,N_3579);
or U7296 (N_7296,N_1712,N_798);
or U7297 (N_7297,N_849,N_228);
or U7298 (N_7298,N_1536,N_495);
nor U7299 (N_7299,N_825,N_2246);
nand U7300 (N_7300,N_2821,N_3654);
nor U7301 (N_7301,N_4629,N_715);
and U7302 (N_7302,N_1885,N_3703);
and U7303 (N_7303,N_3000,N_4900);
and U7304 (N_7304,N_3669,N_687);
nand U7305 (N_7305,N_80,N_2026);
nor U7306 (N_7306,N_4737,N_3033);
xor U7307 (N_7307,N_942,N_3145);
xor U7308 (N_7308,N_3302,N_3879);
and U7309 (N_7309,N_597,N_573);
nand U7310 (N_7310,N_1354,N_3323);
xnor U7311 (N_7311,N_623,N_4144);
or U7312 (N_7312,N_3509,N_2717);
nand U7313 (N_7313,N_2344,N_1308);
and U7314 (N_7314,N_2324,N_2655);
nand U7315 (N_7315,N_1954,N_754);
xnor U7316 (N_7316,N_2067,N_1781);
or U7317 (N_7317,N_2144,N_3007);
or U7318 (N_7318,N_1534,N_2163);
nand U7319 (N_7319,N_1758,N_1409);
or U7320 (N_7320,N_1192,N_2262);
or U7321 (N_7321,N_2588,N_2968);
xnor U7322 (N_7322,N_1551,N_3431);
xor U7323 (N_7323,N_158,N_318);
nor U7324 (N_7324,N_579,N_963);
nand U7325 (N_7325,N_1554,N_3250);
nor U7326 (N_7326,N_1295,N_2319);
nand U7327 (N_7327,N_3760,N_2343);
nand U7328 (N_7328,N_1110,N_2089);
and U7329 (N_7329,N_875,N_3806);
nand U7330 (N_7330,N_1988,N_2518);
nor U7331 (N_7331,N_2374,N_2761);
nor U7332 (N_7332,N_4217,N_2987);
or U7333 (N_7333,N_2000,N_1845);
nor U7334 (N_7334,N_2370,N_2776);
nand U7335 (N_7335,N_2240,N_165);
nor U7336 (N_7336,N_3065,N_1891);
nor U7337 (N_7337,N_2539,N_3985);
and U7338 (N_7338,N_3440,N_2200);
nand U7339 (N_7339,N_4683,N_2668);
xnor U7340 (N_7340,N_2173,N_3547);
nor U7341 (N_7341,N_4438,N_1285);
nor U7342 (N_7342,N_4080,N_713);
and U7343 (N_7343,N_801,N_2196);
or U7344 (N_7344,N_2818,N_2077);
and U7345 (N_7345,N_4221,N_1279);
nor U7346 (N_7346,N_4522,N_3601);
and U7347 (N_7347,N_2998,N_2489);
and U7348 (N_7348,N_870,N_467);
or U7349 (N_7349,N_1239,N_1476);
and U7350 (N_7350,N_3893,N_4828);
nand U7351 (N_7351,N_1265,N_3342);
or U7352 (N_7352,N_361,N_4407);
and U7353 (N_7353,N_4383,N_443);
nand U7354 (N_7354,N_1428,N_2537);
and U7355 (N_7355,N_2917,N_3508);
nor U7356 (N_7356,N_3441,N_4479);
nand U7357 (N_7357,N_3886,N_4350);
or U7358 (N_7358,N_3566,N_2412);
xnor U7359 (N_7359,N_1208,N_4793);
and U7360 (N_7360,N_1527,N_1979);
nor U7361 (N_7361,N_4181,N_643);
nand U7362 (N_7362,N_848,N_980);
and U7363 (N_7363,N_1139,N_916);
nor U7364 (N_7364,N_3587,N_217);
xor U7365 (N_7365,N_4140,N_3449);
and U7366 (N_7366,N_348,N_710);
or U7367 (N_7367,N_1176,N_3514);
and U7368 (N_7368,N_780,N_4966);
or U7369 (N_7369,N_379,N_740);
nor U7370 (N_7370,N_1187,N_1173);
nor U7371 (N_7371,N_1005,N_4185);
nand U7372 (N_7372,N_1542,N_4703);
xnor U7373 (N_7373,N_3637,N_436);
nor U7374 (N_7374,N_3663,N_2845);
or U7375 (N_7375,N_2228,N_4961);
and U7376 (N_7376,N_77,N_2223);
nand U7377 (N_7377,N_4225,N_4398);
and U7378 (N_7378,N_4420,N_1312);
and U7379 (N_7379,N_3942,N_2090);
and U7380 (N_7380,N_4012,N_4219);
nand U7381 (N_7381,N_1451,N_3210);
nor U7382 (N_7382,N_1003,N_2135);
nor U7383 (N_7383,N_3739,N_9);
nor U7384 (N_7384,N_3630,N_4920);
nand U7385 (N_7385,N_4577,N_1535);
nand U7386 (N_7386,N_789,N_3223);
nand U7387 (N_7387,N_2553,N_3214);
nor U7388 (N_7388,N_511,N_3877);
xnor U7389 (N_7389,N_4096,N_1014);
xnor U7390 (N_7390,N_3213,N_4693);
xnor U7391 (N_7391,N_204,N_1636);
nor U7392 (N_7392,N_4922,N_2986);
or U7393 (N_7393,N_1039,N_1032);
and U7394 (N_7394,N_2754,N_1617);
and U7395 (N_7395,N_722,N_4653);
or U7396 (N_7396,N_4134,N_1764);
or U7397 (N_7397,N_250,N_4403);
xor U7398 (N_7398,N_2808,N_2957);
or U7399 (N_7399,N_3293,N_4188);
or U7400 (N_7400,N_667,N_152);
nor U7401 (N_7401,N_2584,N_1977);
nand U7402 (N_7402,N_1963,N_3945);
and U7403 (N_7403,N_1386,N_4024);
or U7404 (N_7404,N_4538,N_2435);
and U7405 (N_7405,N_1151,N_3014);
or U7406 (N_7406,N_200,N_2740);
nand U7407 (N_7407,N_1455,N_683);
nand U7408 (N_7408,N_2508,N_572);
or U7409 (N_7409,N_259,N_15);
nor U7410 (N_7410,N_3834,N_736);
nor U7411 (N_7411,N_1406,N_407);
or U7412 (N_7412,N_2564,N_4277);
or U7413 (N_7413,N_3971,N_231);
or U7414 (N_7414,N_971,N_4322);
nand U7415 (N_7415,N_1258,N_1619);
nor U7416 (N_7416,N_1615,N_2608);
and U7417 (N_7417,N_629,N_4986);
or U7418 (N_7418,N_134,N_3720);
and U7419 (N_7419,N_4328,N_2629);
and U7420 (N_7420,N_4759,N_3421);
or U7421 (N_7421,N_1479,N_3403);
nand U7422 (N_7422,N_508,N_4730);
or U7423 (N_7423,N_145,N_4613);
xnor U7424 (N_7424,N_1331,N_1748);
or U7425 (N_7425,N_1229,N_1423);
and U7426 (N_7426,N_42,N_4176);
nor U7427 (N_7427,N_665,N_489);
and U7428 (N_7428,N_1568,N_878);
nand U7429 (N_7429,N_3399,N_2);
nand U7430 (N_7430,N_1502,N_1945);
and U7431 (N_7431,N_2460,N_3530);
or U7432 (N_7432,N_1701,N_2430);
and U7433 (N_7433,N_3841,N_3462);
and U7434 (N_7434,N_1060,N_4394);
or U7435 (N_7435,N_1220,N_3894);
nor U7436 (N_7436,N_1057,N_1484);
and U7437 (N_7437,N_4346,N_682);
nand U7438 (N_7438,N_3190,N_1588);
nand U7439 (N_7439,N_4669,N_2148);
xor U7440 (N_7440,N_1583,N_3902);
nand U7441 (N_7441,N_1767,N_1286);
and U7442 (N_7442,N_4893,N_2918);
or U7443 (N_7443,N_812,N_4332);
and U7444 (N_7444,N_2086,N_1545);
nand U7445 (N_7445,N_73,N_3286);
nand U7446 (N_7446,N_2793,N_4467);
nor U7447 (N_7447,N_1646,N_570);
nand U7448 (N_7448,N_1628,N_3093);
nor U7449 (N_7449,N_1218,N_2502);
nor U7450 (N_7450,N_2188,N_2199);
and U7451 (N_7451,N_3565,N_2012);
nor U7452 (N_7452,N_3338,N_2637);
or U7453 (N_7453,N_3699,N_3502);
and U7454 (N_7454,N_817,N_792);
nand U7455 (N_7455,N_2638,N_3278);
and U7456 (N_7456,N_1064,N_4888);
or U7457 (N_7457,N_978,N_1994);
nor U7458 (N_7458,N_3358,N_275);
and U7459 (N_7459,N_1604,N_4871);
nor U7460 (N_7460,N_2256,N_1783);
nor U7461 (N_7461,N_2080,N_1969);
nor U7462 (N_7462,N_4016,N_1087);
nor U7463 (N_7463,N_1953,N_708);
nand U7464 (N_7464,N_3393,N_3810);
and U7465 (N_7465,N_2673,N_2273);
nor U7466 (N_7466,N_2470,N_4596);
and U7467 (N_7467,N_788,N_3649);
or U7468 (N_7468,N_2291,N_1283);
or U7469 (N_7469,N_4214,N_1532);
or U7470 (N_7470,N_2031,N_3829);
or U7471 (N_7471,N_4135,N_799);
nand U7472 (N_7472,N_4367,N_78);
or U7473 (N_7473,N_1755,N_3685);
and U7474 (N_7474,N_4677,N_4897);
or U7475 (N_7475,N_3724,N_109);
nor U7476 (N_7476,N_2404,N_1195);
nor U7477 (N_7477,N_84,N_3146);
nor U7478 (N_7478,N_3504,N_891);
nand U7479 (N_7479,N_2105,N_1776);
or U7480 (N_7480,N_1856,N_2133);
and U7481 (N_7481,N_4121,N_2461);
or U7482 (N_7482,N_4953,N_2812);
nor U7483 (N_7483,N_1400,N_4994);
or U7484 (N_7484,N_2507,N_810);
and U7485 (N_7485,N_2215,N_2792);
nand U7486 (N_7486,N_1201,N_2411);
nor U7487 (N_7487,N_4558,N_1859);
nor U7488 (N_7488,N_3682,N_2469);
or U7489 (N_7489,N_2232,N_1930);
nand U7490 (N_7490,N_389,N_2426);
and U7491 (N_7491,N_435,N_4507);
xor U7492 (N_7492,N_4320,N_2396);
and U7493 (N_7493,N_2409,N_3018);
or U7494 (N_7494,N_1949,N_4361);
nor U7495 (N_7495,N_4620,N_4962);
nand U7496 (N_7496,N_3224,N_4402);
and U7497 (N_7497,N_4379,N_88);
or U7498 (N_7498,N_3483,N_289);
nor U7499 (N_7499,N_2447,N_2621);
or U7500 (N_7500,N_3920,N_2553);
or U7501 (N_7501,N_4775,N_3045);
nand U7502 (N_7502,N_2064,N_583);
nand U7503 (N_7503,N_3632,N_3343);
nand U7504 (N_7504,N_63,N_1079);
nand U7505 (N_7505,N_484,N_522);
nor U7506 (N_7506,N_3059,N_3948);
xnor U7507 (N_7507,N_857,N_3971);
nand U7508 (N_7508,N_1720,N_2774);
nand U7509 (N_7509,N_3739,N_3040);
nand U7510 (N_7510,N_3260,N_1952);
nand U7511 (N_7511,N_208,N_348);
xor U7512 (N_7512,N_4394,N_683);
and U7513 (N_7513,N_1568,N_2189);
xnor U7514 (N_7514,N_4728,N_4856);
nor U7515 (N_7515,N_2906,N_2579);
nor U7516 (N_7516,N_3815,N_3698);
nor U7517 (N_7517,N_570,N_4828);
nor U7518 (N_7518,N_3865,N_2506);
nor U7519 (N_7519,N_492,N_3462);
or U7520 (N_7520,N_1014,N_1906);
or U7521 (N_7521,N_1622,N_115);
nand U7522 (N_7522,N_2550,N_4383);
nor U7523 (N_7523,N_3792,N_972);
or U7524 (N_7524,N_3229,N_83);
nand U7525 (N_7525,N_1145,N_920);
xnor U7526 (N_7526,N_1618,N_3213);
and U7527 (N_7527,N_201,N_1881);
nand U7528 (N_7528,N_1921,N_4468);
nand U7529 (N_7529,N_1270,N_906);
nand U7530 (N_7530,N_2588,N_3907);
and U7531 (N_7531,N_1173,N_4381);
nand U7532 (N_7532,N_3144,N_1481);
nand U7533 (N_7533,N_2749,N_2091);
and U7534 (N_7534,N_3181,N_4355);
xnor U7535 (N_7535,N_3825,N_4207);
and U7536 (N_7536,N_3568,N_3808);
nor U7537 (N_7537,N_2829,N_3606);
or U7538 (N_7538,N_1506,N_309);
or U7539 (N_7539,N_2897,N_652);
nand U7540 (N_7540,N_2743,N_2377);
nand U7541 (N_7541,N_3094,N_1977);
nand U7542 (N_7542,N_1980,N_3838);
xnor U7543 (N_7543,N_510,N_4257);
or U7544 (N_7544,N_4779,N_1067);
and U7545 (N_7545,N_2367,N_3610);
and U7546 (N_7546,N_2256,N_882);
nand U7547 (N_7547,N_4933,N_963);
nor U7548 (N_7548,N_2777,N_4680);
and U7549 (N_7549,N_1941,N_3898);
nor U7550 (N_7550,N_91,N_3450);
or U7551 (N_7551,N_828,N_1995);
nor U7552 (N_7552,N_1064,N_4281);
and U7553 (N_7553,N_4955,N_2250);
nor U7554 (N_7554,N_4444,N_3134);
nor U7555 (N_7555,N_1296,N_686);
nor U7556 (N_7556,N_1797,N_1431);
nor U7557 (N_7557,N_4933,N_725);
or U7558 (N_7558,N_4733,N_869);
and U7559 (N_7559,N_4740,N_3256);
or U7560 (N_7560,N_4210,N_3512);
nand U7561 (N_7561,N_2610,N_572);
nand U7562 (N_7562,N_4314,N_2060);
and U7563 (N_7563,N_4807,N_4897);
or U7564 (N_7564,N_458,N_2874);
xnor U7565 (N_7565,N_363,N_4535);
nand U7566 (N_7566,N_2628,N_2402);
nand U7567 (N_7567,N_3869,N_656);
or U7568 (N_7568,N_1513,N_3064);
nor U7569 (N_7569,N_3823,N_1252);
nand U7570 (N_7570,N_4288,N_3457);
xnor U7571 (N_7571,N_1757,N_22);
nor U7572 (N_7572,N_3023,N_1230);
and U7573 (N_7573,N_3522,N_1857);
and U7574 (N_7574,N_254,N_1613);
nor U7575 (N_7575,N_2626,N_2870);
nor U7576 (N_7576,N_4951,N_2212);
or U7577 (N_7577,N_1875,N_2425);
or U7578 (N_7578,N_4352,N_3945);
and U7579 (N_7579,N_3303,N_3239);
nor U7580 (N_7580,N_1359,N_4284);
xor U7581 (N_7581,N_4599,N_969);
or U7582 (N_7582,N_175,N_3424);
and U7583 (N_7583,N_2838,N_4618);
or U7584 (N_7584,N_243,N_2719);
nand U7585 (N_7585,N_297,N_4136);
nand U7586 (N_7586,N_333,N_2040);
nand U7587 (N_7587,N_4518,N_1550);
or U7588 (N_7588,N_1914,N_781);
nor U7589 (N_7589,N_4923,N_203);
xor U7590 (N_7590,N_4115,N_205);
and U7591 (N_7591,N_4812,N_3681);
nand U7592 (N_7592,N_4924,N_2703);
or U7593 (N_7593,N_4870,N_4789);
or U7594 (N_7594,N_4085,N_927);
nand U7595 (N_7595,N_1767,N_4051);
xnor U7596 (N_7596,N_124,N_3299);
or U7597 (N_7597,N_415,N_3361);
xor U7598 (N_7598,N_1719,N_4036);
nor U7599 (N_7599,N_3477,N_1726);
and U7600 (N_7600,N_187,N_4596);
nor U7601 (N_7601,N_128,N_3143);
nand U7602 (N_7602,N_730,N_2880);
and U7603 (N_7603,N_1711,N_3170);
nand U7604 (N_7604,N_1605,N_4595);
nand U7605 (N_7605,N_4253,N_1221);
nand U7606 (N_7606,N_863,N_431);
nand U7607 (N_7607,N_3178,N_2492);
or U7608 (N_7608,N_1975,N_4441);
nor U7609 (N_7609,N_856,N_596);
or U7610 (N_7610,N_640,N_235);
nand U7611 (N_7611,N_28,N_278);
nor U7612 (N_7612,N_4886,N_4354);
or U7613 (N_7613,N_3490,N_3962);
and U7614 (N_7614,N_905,N_2348);
nor U7615 (N_7615,N_1372,N_4595);
and U7616 (N_7616,N_161,N_3767);
nor U7617 (N_7617,N_3801,N_2320);
and U7618 (N_7618,N_1365,N_2510);
and U7619 (N_7619,N_2066,N_1946);
xor U7620 (N_7620,N_1146,N_1676);
xor U7621 (N_7621,N_1213,N_4523);
or U7622 (N_7622,N_1586,N_893);
and U7623 (N_7623,N_2452,N_4489);
or U7624 (N_7624,N_2622,N_3502);
nand U7625 (N_7625,N_402,N_4549);
nand U7626 (N_7626,N_4924,N_1479);
xor U7627 (N_7627,N_1836,N_1549);
nor U7628 (N_7628,N_3347,N_4428);
nand U7629 (N_7629,N_1207,N_1644);
and U7630 (N_7630,N_2601,N_4558);
nor U7631 (N_7631,N_4185,N_370);
nor U7632 (N_7632,N_1200,N_2506);
or U7633 (N_7633,N_4733,N_3893);
nand U7634 (N_7634,N_4198,N_4997);
nand U7635 (N_7635,N_4601,N_2078);
and U7636 (N_7636,N_582,N_3375);
or U7637 (N_7637,N_1227,N_4785);
xor U7638 (N_7638,N_4314,N_4986);
nor U7639 (N_7639,N_4338,N_1324);
xnor U7640 (N_7640,N_4017,N_4316);
and U7641 (N_7641,N_1325,N_1674);
or U7642 (N_7642,N_4501,N_1507);
nor U7643 (N_7643,N_4864,N_2942);
and U7644 (N_7644,N_4079,N_116);
nor U7645 (N_7645,N_2561,N_2724);
nor U7646 (N_7646,N_1108,N_1132);
nor U7647 (N_7647,N_3041,N_3015);
nor U7648 (N_7648,N_1474,N_310);
and U7649 (N_7649,N_3513,N_3212);
and U7650 (N_7650,N_574,N_1691);
nor U7651 (N_7651,N_2539,N_2744);
or U7652 (N_7652,N_3824,N_2842);
or U7653 (N_7653,N_2427,N_1899);
and U7654 (N_7654,N_1039,N_4568);
and U7655 (N_7655,N_4118,N_3398);
nand U7656 (N_7656,N_3592,N_4964);
xnor U7657 (N_7657,N_3113,N_4561);
or U7658 (N_7658,N_10,N_4436);
nand U7659 (N_7659,N_606,N_693);
or U7660 (N_7660,N_3279,N_4132);
and U7661 (N_7661,N_2129,N_4532);
or U7662 (N_7662,N_82,N_3454);
or U7663 (N_7663,N_2178,N_4369);
and U7664 (N_7664,N_4410,N_3493);
nor U7665 (N_7665,N_2193,N_4346);
nand U7666 (N_7666,N_4195,N_2229);
and U7667 (N_7667,N_3656,N_1991);
and U7668 (N_7668,N_4011,N_2377);
and U7669 (N_7669,N_857,N_548);
and U7670 (N_7670,N_4709,N_4833);
and U7671 (N_7671,N_4838,N_4614);
nand U7672 (N_7672,N_4154,N_4551);
nand U7673 (N_7673,N_1751,N_1115);
xor U7674 (N_7674,N_1530,N_412);
or U7675 (N_7675,N_2463,N_175);
nor U7676 (N_7676,N_2469,N_4053);
nand U7677 (N_7677,N_4883,N_4652);
and U7678 (N_7678,N_1047,N_3136);
and U7679 (N_7679,N_1606,N_3212);
xor U7680 (N_7680,N_1395,N_1410);
xnor U7681 (N_7681,N_4956,N_2190);
xnor U7682 (N_7682,N_3591,N_4380);
nand U7683 (N_7683,N_2863,N_945);
nand U7684 (N_7684,N_1283,N_852);
nor U7685 (N_7685,N_1914,N_1948);
and U7686 (N_7686,N_1691,N_3947);
or U7687 (N_7687,N_3805,N_819);
or U7688 (N_7688,N_4615,N_4826);
and U7689 (N_7689,N_1187,N_88);
or U7690 (N_7690,N_3172,N_3587);
and U7691 (N_7691,N_1555,N_344);
and U7692 (N_7692,N_1431,N_1625);
nand U7693 (N_7693,N_3656,N_3974);
nor U7694 (N_7694,N_4711,N_1619);
or U7695 (N_7695,N_2576,N_3665);
xor U7696 (N_7696,N_2711,N_518);
xor U7697 (N_7697,N_62,N_690);
nand U7698 (N_7698,N_2830,N_823);
nor U7699 (N_7699,N_543,N_994);
nand U7700 (N_7700,N_706,N_2229);
xor U7701 (N_7701,N_1498,N_771);
and U7702 (N_7702,N_2862,N_4269);
xor U7703 (N_7703,N_704,N_521);
or U7704 (N_7704,N_2861,N_4447);
and U7705 (N_7705,N_438,N_4139);
nor U7706 (N_7706,N_4190,N_2745);
or U7707 (N_7707,N_3806,N_878);
or U7708 (N_7708,N_4189,N_2640);
and U7709 (N_7709,N_1657,N_776);
and U7710 (N_7710,N_964,N_2964);
nand U7711 (N_7711,N_697,N_1034);
nor U7712 (N_7712,N_4927,N_3681);
or U7713 (N_7713,N_2355,N_2353);
or U7714 (N_7714,N_4934,N_4700);
xor U7715 (N_7715,N_3034,N_4434);
nand U7716 (N_7716,N_629,N_501);
nand U7717 (N_7717,N_3228,N_1964);
or U7718 (N_7718,N_4429,N_1853);
or U7719 (N_7719,N_1449,N_1916);
nand U7720 (N_7720,N_3472,N_359);
nand U7721 (N_7721,N_577,N_2322);
or U7722 (N_7722,N_2719,N_3834);
nand U7723 (N_7723,N_1172,N_2822);
and U7724 (N_7724,N_1005,N_1158);
nand U7725 (N_7725,N_1208,N_1481);
nor U7726 (N_7726,N_1654,N_2162);
nand U7727 (N_7727,N_4981,N_878);
and U7728 (N_7728,N_174,N_2789);
nand U7729 (N_7729,N_4692,N_4547);
xnor U7730 (N_7730,N_2329,N_2209);
or U7731 (N_7731,N_4926,N_3077);
or U7732 (N_7732,N_2890,N_2112);
or U7733 (N_7733,N_3706,N_573);
or U7734 (N_7734,N_4529,N_3209);
nand U7735 (N_7735,N_3871,N_1519);
or U7736 (N_7736,N_4676,N_4997);
and U7737 (N_7737,N_2666,N_946);
or U7738 (N_7738,N_75,N_2970);
xnor U7739 (N_7739,N_3544,N_4499);
nor U7740 (N_7740,N_1442,N_737);
xor U7741 (N_7741,N_175,N_4979);
nor U7742 (N_7742,N_3317,N_2420);
and U7743 (N_7743,N_4991,N_1522);
or U7744 (N_7744,N_3570,N_4415);
nor U7745 (N_7745,N_1490,N_2725);
nand U7746 (N_7746,N_790,N_4954);
xor U7747 (N_7747,N_3127,N_3724);
or U7748 (N_7748,N_3593,N_3292);
xnor U7749 (N_7749,N_3798,N_724);
or U7750 (N_7750,N_1987,N_1978);
or U7751 (N_7751,N_1309,N_3135);
nor U7752 (N_7752,N_917,N_3731);
or U7753 (N_7753,N_1166,N_4542);
or U7754 (N_7754,N_4456,N_3442);
nor U7755 (N_7755,N_4060,N_1234);
or U7756 (N_7756,N_185,N_1984);
nor U7757 (N_7757,N_1251,N_3858);
nor U7758 (N_7758,N_3658,N_2508);
nand U7759 (N_7759,N_1630,N_398);
or U7760 (N_7760,N_1869,N_4191);
nor U7761 (N_7761,N_660,N_4187);
nor U7762 (N_7762,N_2747,N_1788);
nand U7763 (N_7763,N_4357,N_4882);
or U7764 (N_7764,N_1031,N_4147);
or U7765 (N_7765,N_957,N_1406);
nor U7766 (N_7766,N_1840,N_1910);
or U7767 (N_7767,N_4251,N_4576);
nor U7768 (N_7768,N_3253,N_2225);
nand U7769 (N_7769,N_544,N_2448);
xnor U7770 (N_7770,N_1387,N_1172);
or U7771 (N_7771,N_4501,N_2408);
and U7772 (N_7772,N_3786,N_3857);
xnor U7773 (N_7773,N_4943,N_1925);
nor U7774 (N_7774,N_4320,N_4584);
nor U7775 (N_7775,N_4799,N_3471);
and U7776 (N_7776,N_2995,N_1042);
or U7777 (N_7777,N_2463,N_66);
xnor U7778 (N_7778,N_1722,N_4470);
nand U7779 (N_7779,N_676,N_777);
and U7780 (N_7780,N_3666,N_2038);
and U7781 (N_7781,N_3833,N_1196);
nor U7782 (N_7782,N_1555,N_3374);
nor U7783 (N_7783,N_3411,N_4713);
or U7784 (N_7784,N_1816,N_3721);
or U7785 (N_7785,N_893,N_3374);
nor U7786 (N_7786,N_4188,N_320);
nor U7787 (N_7787,N_2100,N_2059);
and U7788 (N_7788,N_4317,N_878);
and U7789 (N_7789,N_4288,N_908);
nand U7790 (N_7790,N_3533,N_1077);
nor U7791 (N_7791,N_968,N_3709);
nand U7792 (N_7792,N_4430,N_667);
or U7793 (N_7793,N_1265,N_4790);
nand U7794 (N_7794,N_320,N_3800);
and U7795 (N_7795,N_3315,N_4949);
nand U7796 (N_7796,N_668,N_4656);
or U7797 (N_7797,N_871,N_2596);
and U7798 (N_7798,N_413,N_2256);
nand U7799 (N_7799,N_1376,N_1358);
xnor U7800 (N_7800,N_1197,N_781);
and U7801 (N_7801,N_3398,N_4154);
xor U7802 (N_7802,N_397,N_2913);
nand U7803 (N_7803,N_2622,N_3878);
or U7804 (N_7804,N_4762,N_3403);
and U7805 (N_7805,N_1402,N_4971);
nor U7806 (N_7806,N_1420,N_3112);
nand U7807 (N_7807,N_1085,N_2892);
or U7808 (N_7808,N_264,N_4006);
or U7809 (N_7809,N_4739,N_2335);
or U7810 (N_7810,N_4534,N_797);
nor U7811 (N_7811,N_2607,N_4564);
nand U7812 (N_7812,N_3778,N_4048);
and U7813 (N_7813,N_1485,N_2603);
nor U7814 (N_7814,N_2138,N_4578);
and U7815 (N_7815,N_1635,N_219);
and U7816 (N_7816,N_4090,N_2307);
nand U7817 (N_7817,N_3492,N_4746);
nor U7818 (N_7818,N_1464,N_3216);
and U7819 (N_7819,N_2372,N_1951);
or U7820 (N_7820,N_167,N_1879);
nor U7821 (N_7821,N_2019,N_2416);
nand U7822 (N_7822,N_1876,N_2025);
nor U7823 (N_7823,N_1099,N_2191);
xnor U7824 (N_7824,N_2031,N_3284);
or U7825 (N_7825,N_30,N_3862);
and U7826 (N_7826,N_231,N_81);
nor U7827 (N_7827,N_1573,N_4748);
and U7828 (N_7828,N_702,N_3801);
nand U7829 (N_7829,N_4685,N_4583);
or U7830 (N_7830,N_2910,N_3867);
nor U7831 (N_7831,N_4916,N_1623);
nand U7832 (N_7832,N_2426,N_1059);
nor U7833 (N_7833,N_4690,N_3542);
nor U7834 (N_7834,N_755,N_1969);
and U7835 (N_7835,N_4792,N_1366);
nor U7836 (N_7836,N_3809,N_1512);
xor U7837 (N_7837,N_3772,N_2383);
or U7838 (N_7838,N_4222,N_4127);
xnor U7839 (N_7839,N_1540,N_344);
nor U7840 (N_7840,N_3364,N_3122);
and U7841 (N_7841,N_1662,N_4880);
or U7842 (N_7842,N_1555,N_3552);
nand U7843 (N_7843,N_854,N_4452);
or U7844 (N_7844,N_564,N_2105);
and U7845 (N_7845,N_3469,N_3978);
nor U7846 (N_7846,N_2302,N_784);
nor U7847 (N_7847,N_4775,N_3864);
nor U7848 (N_7848,N_1525,N_2511);
or U7849 (N_7849,N_4899,N_4980);
nand U7850 (N_7850,N_685,N_687);
nand U7851 (N_7851,N_3287,N_702);
nand U7852 (N_7852,N_208,N_3654);
nand U7853 (N_7853,N_1091,N_2556);
or U7854 (N_7854,N_3330,N_3787);
or U7855 (N_7855,N_1001,N_1618);
nand U7856 (N_7856,N_2445,N_2294);
or U7857 (N_7857,N_4118,N_3056);
and U7858 (N_7858,N_594,N_2013);
and U7859 (N_7859,N_2079,N_4591);
nand U7860 (N_7860,N_3327,N_2908);
nand U7861 (N_7861,N_3900,N_2338);
or U7862 (N_7862,N_1039,N_4210);
nand U7863 (N_7863,N_1900,N_1390);
nand U7864 (N_7864,N_3199,N_3920);
nor U7865 (N_7865,N_3781,N_3823);
nor U7866 (N_7866,N_361,N_899);
and U7867 (N_7867,N_3730,N_2301);
and U7868 (N_7868,N_264,N_35);
or U7869 (N_7869,N_3323,N_1778);
nor U7870 (N_7870,N_885,N_3882);
nand U7871 (N_7871,N_4421,N_3301);
nand U7872 (N_7872,N_4579,N_1986);
and U7873 (N_7873,N_2520,N_147);
or U7874 (N_7874,N_1370,N_4875);
and U7875 (N_7875,N_2983,N_1928);
and U7876 (N_7876,N_3869,N_924);
and U7877 (N_7877,N_1287,N_1739);
nor U7878 (N_7878,N_3714,N_752);
nor U7879 (N_7879,N_3932,N_4415);
xor U7880 (N_7880,N_4570,N_3695);
or U7881 (N_7881,N_1446,N_2452);
nor U7882 (N_7882,N_4598,N_3446);
nor U7883 (N_7883,N_3784,N_3314);
or U7884 (N_7884,N_4123,N_2200);
nor U7885 (N_7885,N_1692,N_2066);
or U7886 (N_7886,N_450,N_1100);
and U7887 (N_7887,N_1023,N_2074);
nor U7888 (N_7888,N_1579,N_1227);
and U7889 (N_7889,N_3203,N_694);
nor U7890 (N_7890,N_271,N_3809);
nor U7891 (N_7891,N_1952,N_728);
xnor U7892 (N_7892,N_570,N_3936);
xor U7893 (N_7893,N_4871,N_1318);
and U7894 (N_7894,N_2303,N_2014);
or U7895 (N_7895,N_4962,N_1107);
and U7896 (N_7896,N_3951,N_3926);
or U7897 (N_7897,N_3994,N_3507);
and U7898 (N_7898,N_2627,N_3672);
xnor U7899 (N_7899,N_4801,N_4697);
and U7900 (N_7900,N_4996,N_461);
or U7901 (N_7901,N_1179,N_4515);
nor U7902 (N_7902,N_64,N_376);
or U7903 (N_7903,N_1857,N_1891);
xor U7904 (N_7904,N_4736,N_1291);
and U7905 (N_7905,N_3154,N_4356);
or U7906 (N_7906,N_1360,N_1075);
nand U7907 (N_7907,N_1060,N_550);
and U7908 (N_7908,N_1209,N_3258);
nor U7909 (N_7909,N_767,N_2235);
and U7910 (N_7910,N_1606,N_3777);
and U7911 (N_7911,N_4401,N_2733);
xnor U7912 (N_7912,N_319,N_1693);
and U7913 (N_7913,N_323,N_140);
xnor U7914 (N_7914,N_2968,N_1929);
or U7915 (N_7915,N_4325,N_3742);
nor U7916 (N_7916,N_3524,N_4460);
nand U7917 (N_7917,N_2138,N_4243);
nor U7918 (N_7918,N_4250,N_4735);
nand U7919 (N_7919,N_3643,N_897);
nand U7920 (N_7920,N_2432,N_1956);
and U7921 (N_7921,N_4866,N_3606);
nor U7922 (N_7922,N_3322,N_4879);
nand U7923 (N_7923,N_3916,N_1897);
or U7924 (N_7924,N_2447,N_2286);
nand U7925 (N_7925,N_4335,N_2902);
nor U7926 (N_7926,N_2748,N_1875);
nor U7927 (N_7927,N_1959,N_4874);
or U7928 (N_7928,N_4902,N_4766);
xnor U7929 (N_7929,N_2741,N_1386);
nand U7930 (N_7930,N_1828,N_3083);
or U7931 (N_7931,N_3370,N_2682);
or U7932 (N_7932,N_4235,N_1888);
nor U7933 (N_7933,N_1807,N_2887);
and U7934 (N_7934,N_2557,N_3948);
nand U7935 (N_7935,N_4250,N_1522);
xnor U7936 (N_7936,N_3540,N_3205);
and U7937 (N_7937,N_1258,N_1876);
or U7938 (N_7938,N_596,N_350);
or U7939 (N_7939,N_4158,N_4923);
and U7940 (N_7940,N_3358,N_3461);
nor U7941 (N_7941,N_1365,N_2811);
xnor U7942 (N_7942,N_1716,N_634);
xnor U7943 (N_7943,N_1756,N_3815);
or U7944 (N_7944,N_3570,N_4292);
and U7945 (N_7945,N_4339,N_236);
nand U7946 (N_7946,N_2129,N_431);
nand U7947 (N_7947,N_186,N_141);
or U7948 (N_7948,N_3149,N_3663);
nand U7949 (N_7949,N_2675,N_4401);
and U7950 (N_7950,N_3254,N_1760);
nand U7951 (N_7951,N_3475,N_1314);
nor U7952 (N_7952,N_3268,N_4157);
or U7953 (N_7953,N_4396,N_3272);
nor U7954 (N_7954,N_3791,N_412);
and U7955 (N_7955,N_3771,N_875);
or U7956 (N_7956,N_360,N_1491);
nand U7957 (N_7957,N_4742,N_3661);
nor U7958 (N_7958,N_207,N_2231);
nand U7959 (N_7959,N_1173,N_3339);
and U7960 (N_7960,N_1323,N_4082);
nand U7961 (N_7961,N_1795,N_2223);
nand U7962 (N_7962,N_1894,N_4);
xor U7963 (N_7963,N_85,N_3155);
xnor U7964 (N_7964,N_734,N_3985);
or U7965 (N_7965,N_3969,N_1621);
nand U7966 (N_7966,N_2123,N_3295);
xnor U7967 (N_7967,N_2766,N_4624);
or U7968 (N_7968,N_1666,N_3851);
or U7969 (N_7969,N_295,N_3080);
or U7970 (N_7970,N_560,N_2686);
nand U7971 (N_7971,N_2689,N_4037);
nand U7972 (N_7972,N_2625,N_3354);
and U7973 (N_7973,N_2892,N_3939);
and U7974 (N_7974,N_1846,N_4022);
or U7975 (N_7975,N_1983,N_4278);
or U7976 (N_7976,N_2931,N_4804);
nand U7977 (N_7977,N_279,N_3360);
nor U7978 (N_7978,N_1238,N_2610);
nand U7979 (N_7979,N_3882,N_445);
nand U7980 (N_7980,N_2248,N_3145);
nand U7981 (N_7981,N_1791,N_2098);
nand U7982 (N_7982,N_2906,N_1463);
or U7983 (N_7983,N_1444,N_3417);
and U7984 (N_7984,N_4069,N_2868);
nand U7985 (N_7985,N_4385,N_2303);
or U7986 (N_7986,N_1270,N_2249);
nor U7987 (N_7987,N_4453,N_1318);
or U7988 (N_7988,N_1895,N_3133);
and U7989 (N_7989,N_4067,N_1189);
and U7990 (N_7990,N_2294,N_4295);
and U7991 (N_7991,N_1601,N_4972);
nand U7992 (N_7992,N_3717,N_1175);
or U7993 (N_7993,N_1470,N_2242);
nor U7994 (N_7994,N_4958,N_1317);
and U7995 (N_7995,N_1252,N_2580);
nor U7996 (N_7996,N_2034,N_2508);
nand U7997 (N_7997,N_743,N_887);
and U7998 (N_7998,N_511,N_1156);
nand U7999 (N_7999,N_4137,N_3623);
nand U8000 (N_8000,N_1593,N_3347);
or U8001 (N_8001,N_2997,N_149);
nor U8002 (N_8002,N_2163,N_4034);
nor U8003 (N_8003,N_2264,N_4864);
nand U8004 (N_8004,N_2944,N_1568);
and U8005 (N_8005,N_4515,N_460);
and U8006 (N_8006,N_2456,N_116);
nand U8007 (N_8007,N_2490,N_4226);
nor U8008 (N_8008,N_1224,N_248);
nand U8009 (N_8009,N_3448,N_1431);
or U8010 (N_8010,N_2994,N_1981);
nand U8011 (N_8011,N_3892,N_155);
nor U8012 (N_8012,N_4758,N_1684);
nand U8013 (N_8013,N_4969,N_372);
nand U8014 (N_8014,N_2363,N_3337);
nand U8015 (N_8015,N_2304,N_809);
and U8016 (N_8016,N_1424,N_2415);
nand U8017 (N_8017,N_363,N_1764);
nor U8018 (N_8018,N_3669,N_3459);
xor U8019 (N_8019,N_1661,N_2377);
and U8020 (N_8020,N_602,N_2264);
and U8021 (N_8021,N_2344,N_4956);
nand U8022 (N_8022,N_3296,N_380);
or U8023 (N_8023,N_4867,N_4100);
nor U8024 (N_8024,N_3521,N_3176);
and U8025 (N_8025,N_4694,N_32);
or U8026 (N_8026,N_2137,N_3579);
or U8027 (N_8027,N_2880,N_1134);
nand U8028 (N_8028,N_708,N_2311);
nor U8029 (N_8029,N_2499,N_4790);
or U8030 (N_8030,N_3215,N_4480);
nand U8031 (N_8031,N_711,N_1408);
and U8032 (N_8032,N_3352,N_4514);
xnor U8033 (N_8033,N_162,N_2272);
or U8034 (N_8034,N_2458,N_619);
or U8035 (N_8035,N_1019,N_3441);
and U8036 (N_8036,N_2051,N_334);
xnor U8037 (N_8037,N_2480,N_22);
xnor U8038 (N_8038,N_1305,N_1042);
or U8039 (N_8039,N_1462,N_2835);
or U8040 (N_8040,N_2738,N_3308);
xnor U8041 (N_8041,N_4322,N_160);
nand U8042 (N_8042,N_4806,N_4432);
nand U8043 (N_8043,N_3638,N_4114);
or U8044 (N_8044,N_459,N_2387);
nor U8045 (N_8045,N_3209,N_1337);
xnor U8046 (N_8046,N_4104,N_4870);
xnor U8047 (N_8047,N_3536,N_3861);
and U8048 (N_8048,N_1791,N_4268);
and U8049 (N_8049,N_4459,N_256);
nor U8050 (N_8050,N_4004,N_3468);
xnor U8051 (N_8051,N_4881,N_2808);
nand U8052 (N_8052,N_2751,N_3753);
nand U8053 (N_8053,N_651,N_2113);
and U8054 (N_8054,N_4729,N_1320);
nor U8055 (N_8055,N_1957,N_2697);
and U8056 (N_8056,N_4209,N_4046);
and U8057 (N_8057,N_4752,N_1590);
nor U8058 (N_8058,N_1990,N_3420);
and U8059 (N_8059,N_4500,N_1328);
or U8060 (N_8060,N_93,N_4382);
or U8061 (N_8061,N_1532,N_1090);
nand U8062 (N_8062,N_2469,N_3617);
and U8063 (N_8063,N_2525,N_2485);
nand U8064 (N_8064,N_2058,N_3479);
or U8065 (N_8065,N_2370,N_376);
xor U8066 (N_8066,N_1011,N_4826);
nand U8067 (N_8067,N_4860,N_585);
and U8068 (N_8068,N_2335,N_1036);
nor U8069 (N_8069,N_553,N_1840);
nand U8070 (N_8070,N_1266,N_1499);
nor U8071 (N_8071,N_4417,N_1765);
and U8072 (N_8072,N_4613,N_830);
nor U8073 (N_8073,N_3367,N_1861);
nor U8074 (N_8074,N_902,N_4726);
nor U8075 (N_8075,N_1498,N_4630);
or U8076 (N_8076,N_1274,N_3025);
and U8077 (N_8077,N_4517,N_173);
nand U8078 (N_8078,N_1391,N_1084);
nor U8079 (N_8079,N_1989,N_4875);
or U8080 (N_8080,N_2010,N_4932);
or U8081 (N_8081,N_2419,N_2194);
xor U8082 (N_8082,N_4685,N_306);
nor U8083 (N_8083,N_859,N_3654);
nor U8084 (N_8084,N_2838,N_515);
or U8085 (N_8085,N_1949,N_1414);
nor U8086 (N_8086,N_2619,N_4192);
or U8087 (N_8087,N_3235,N_1736);
nand U8088 (N_8088,N_4440,N_4885);
or U8089 (N_8089,N_4877,N_4280);
nor U8090 (N_8090,N_2190,N_2169);
xor U8091 (N_8091,N_3111,N_669);
nor U8092 (N_8092,N_2986,N_3622);
xor U8093 (N_8093,N_2443,N_3606);
or U8094 (N_8094,N_3350,N_1543);
nor U8095 (N_8095,N_1536,N_3173);
nor U8096 (N_8096,N_3674,N_572);
nand U8097 (N_8097,N_3141,N_1106);
nand U8098 (N_8098,N_809,N_4162);
nand U8099 (N_8099,N_3874,N_4543);
or U8100 (N_8100,N_893,N_1806);
and U8101 (N_8101,N_2009,N_1502);
xnor U8102 (N_8102,N_3244,N_4032);
and U8103 (N_8103,N_4099,N_4631);
nand U8104 (N_8104,N_1556,N_3877);
nor U8105 (N_8105,N_3826,N_191);
or U8106 (N_8106,N_1733,N_3386);
nor U8107 (N_8107,N_2426,N_17);
nand U8108 (N_8108,N_4259,N_1114);
nand U8109 (N_8109,N_1195,N_1532);
nor U8110 (N_8110,N_3626,N_641);
and U8111 (N_8111,N_3297,N_2555);
or U8112 (N_8112,N_4793,N_731);
xor U8113 (N_8113,N_3073,N_638);
or U8114 (N_8114,N_2648,N_2443);
or U8115 (N_8115,N_3868,N_2583);
or U8116 (N_8116,N_901,N_187);
nand U8117 (N_8117,N_377,N_881);
nor U8118 (N_8118,N_4257,N_3349);
nand U8119 (N_8119,N_1,N_3965);
nor U8120 (N_8120,N_2279,N_881);
nand U8121 (N_8121,N_2352,N_1458);
and U8122 (N_8122,N_1661,N_3984);
or U8123 (N_8123,N_10,N_587);
nand U8124 (N_8124,N_3170,N_1035);
or U8125 (N_8125,N_4992,N_4457);
nor U8126 (N_8126,N_2300,N_2323);
and U8127 (N_8127,N_1155,N_4569);
or U8128 (N_8128,N_2696,N_1658);
and U8129 (N_8129,N_2357,N_3427);
xor U8130 (N_8130,N_673,N_3786);
or U8131 (N_8131,N_4572,N_2446);
nand U8132 (N_8132,N_4775,N_2683);
or U8133 (N_8133,N_1135,N_1185);
nand U8134 (N_8134,N_1744,N_2135);
nor U8135 (N_8135,N_4887,N_4746);
and U8136 (N_8136,N_3555,N_1326);
nand U8137 (N_8137,N_2909,N_2927);
nor U8138 (N_8138,N_4671,N_2877);
nor U8139 (N_8139,N_1965,N_1998);
nor U8140 (N_8140,N_1323,N_2453);
nor U8141 (N_8141,N_4971,N_4928);
or U8142 (N_8142,N_2645,N_1552);
and U8143 (N_8143,N_750,N_2941);
xor U8144 (N_8144,N_1969,N_4545);
nor U8145 (N_8145,N_2686,N_2696);
nor U8146 (N_8146,N_3309,N_946);
or U8147 (N_8147,N_3248,N_1377);
nand U8148 (N_8148,N_2615,N_2631);
and U8149 (N_8149,N_4001,N_3418);
nand U8150 (N_8150,N_4584,N_1193);
and U8151 (N_8151,N_492,N_433);
and U8152 (N_8152,N_266,N_4922);
nand U8153 (N_8153,N_184,N_2288);
xnor U8154 (N_8154,N_4103,N_1166);
and U8155 (N_8155,N_3490,N_392);
nor U8156 (N_8156,N_4145,N_162);
or U8157 (N_8157,N_2098,N_3642);
nand U8158 (N_8158,N_4213,N_3897);
and U8159 (N_8159,N_1531,N_2801);
xor U8160 (N_8160,N_3045,N_3670);
nor U8161 (N_8161,N_315,N_2431);
nand U8162 (N_8162,N_1704,N_4005);
nand U8163 (N_8163,N_455,N_2575);
or U8164 (N_8164,N_2391,N_407);
nor U8165 (N_8165,N_2652,N_3388);
nand U8166 (N_8166,N_1431,N_4812);
nand U8167 (N_8167,N_3862,N_3217);
nor U8168 (N_8168,N_4591,N_3069);
nor U8169 (N_8169,N_1672,N_3782);
or U8170 (N_8170,N_4204,N_4012);
xnor U8171 (N_8171,N_3504,N_983);
or U8172 (N_8172,N_4116,N_2990);
or U8173 (N_8173,N_2197,N_658);
nor U8174 (N_8174,N_1819,N_362);
nor U8175 (N_8175,N_4083,N_2028);
or U8176 (N_8176,N_809,N_1484);
nand U8177 (N_8177,N_3201,N_3822);
nor U8178 (N_8178,N_2589,N_1527);
xor U8179 (N_8179,N_3851,N_2035);
xor U8180 (N_8180,N_2806,N_1544);
nand U8181 (N_8181,N_267,N_1706);
nand U8182 (N_8182,N_2752,N_134);
and U8183 (N_8183,N_4796,N_2883);
nand U8184 (N_8184,N_568,N_662);
and U8185 (N_8185,N_1048,N_2439);
or U8186 (N_8186,N_2377,N_4405);
and U8187 (N_8187,N_4625,N_1184);
nor U8188 (N_8188,N_1583,N_965);
nor U8189 (N_8189,N_4335,N_1251);
or U8190 (N_8190,N_2868,N_4403);
nor U8191 (N_8191,N_2601,N_1942);
nand U8192 (N_8192,N_138,N_3648);
and U8193 (N_8193,N_146,N_2016);
nor U8194 (N_8194,N_2618,N_1029);
nand U8195 (N_8195,N_814,N_365);
and U8196 (N_8196,N_1002,N_942);
nand U8197 (N_8197,N_2046,N_3037);
and U8198 (N_8198,N_1202,N_3499);
or U8199 (N_8199,N_1701,N_1956);
or U8200 (N_8200,N_3105,N_712);
nor U8201 (N_8201,N_4830,N_3383);
and U8202 (N_8202,N_2369,N_761);
nand U8203 (N_8203,N_4313,N_4187);
nor U8204 (N_8204,N_1923,N_1141);
nor U8205 (N_8205,N_1907,N_389);
or U8206 (N_8206,N_474,N_1325);
or U8207 (N_8207,N_4616,N_508);
and U8208 (N_8208,N_1979,N_4718);
nand U8209 (N_8209,N_2817,N_4206);
nor U8210 (N_8210,N_1578,N_1505);
nor U8211 (N_8211,N_1880,N_4953);
nand U8212 (N_8212,N_828,N_2091);
nand U8213 (N_8213,N_3376,N_1236);
nand U8214 (N_8214,N_3137,N_766);
or U8215 (N_8215,N_3795,N_543);
or U8216 (N_8216,N_4626,N_3284);
nor U8217 (N_8217,N_3125,N_530);
xor U8218 (N_8218,N_4726,N_2917);
and U8219 (N_8219,N_1559,N_1737);
and U8220 (N_8220,N_3227,N_2816);
nor U8221 (N_8221,N_1659,N_260);
nor U8222 (N_8222,N_567,N_505);
or U8223 (N_8223,N_4158,N_3061);
nand U8224 (N_8224,N_2764,N_3431);
nor U8225 (N_8225,N_34,N_4372);
and U8226 (N_8226,N_3268,N_2742);
nor U8227 (N_8227,N_4594,N_4657);
and U8228 (N_8228,N_2826,N_2241);
nor U8229 (N_8229,N_3880,N_2272);
and U8230 (N_8230,N_4398,N_1768);
and U8231 (N_8231,N_508,N_1610);
or U8232 (N_8232,N_4593,N_3276);
nor U8233 (N_8233,N_2791,N_2603);
and U8234 (N_8234,N_427,N_3548);
nor U8235 (N_8235,N_4163,N_2242);
and U8236 (N_8236,N_12,N_1043);
nor U8237 (N_8237,N_4616,N_804);
and U8238 (N_8238,N_4348,N_1726);
and U8239 (N_8239,N_2067,N_2853);
and U8240 (N_8240,N_4293,N_623);
or U8241 (N_8241,N_96,N_2194);
nand U8242 (N_8242,N_3112,N_2738);
and U8243 (N_8243,N_3210,N_4617);
nand U8244 (N_8244,N_2712,N_3059);
nand U8245 (N_8245,N_4434,N_1055);
or U8246 (N_8246,N_4001,N_1485);
nor U8247 (N_8247,N_2648,N_3457);
and U8248 (N_8248,N_2178,N_1471);
nor U8249 (N_8249,N_4791,N_493);
nor U8250 (N_8250,N_1796,N_1150);
and U8251 (N_8251,N_4938,N_1333);
nor U8252 (N_8252,N_4786,N_4733);
or U8253 (N_8253,N_1908,N_3283);
nor U8254 (N_8254,N_1637,N_298);
and U8255 (N_8255,N_4417,N_4500);
or U8256 (N_8256,N_2058,N_858);
nand U8257 (N_8257,N_1920,N_3691);
and U8258 (N_8258,N_1726,N_3834);
nor U8259 (N_8259,N_1135,N_3656);
and U8260 (N_8260,N_1695,N_4813);
xor U8261 (N_8261,N_503,N_249);
nand U8262 (N_8262,N_4849,N_74);
and U8263 (N_8263,N_2907,N_4193);
and U8264 (N_8264,N_710,N_2557);
nor U8265 (N_8265,N_1812,N_3206);
or U8266 (N_8266,N_4370,N_3514);
and U8267 (N_8267,N_806,N_2272);
xnor U8268 (N_8268,N_4734,N_1643);
xnor U8269 (N_8269,N_2820,N_1580);
nand U8270 (N_8270,N_517,N_4411);
and U8271 (N_8271,N_4375,N_276);
and U8272 (N_8272,N_2779,N_3207);
nand U8273 (N_8273,N_229,N_135);
or U8274 (N_8274,N_2830,N_4269);
or U8275 (N_8275,N_3720,N_908);
and U8276 (N_8276,N_2547,N_871);
or U8277 (N_8277,N_4445,N_355);
or U8278 (N_8278,N_2577,N_898);
and U8279 (N_8279,N_4099,N_495);
or U8280 (N_8280,N_483,N_1949);
nor U8281 (N_8281,N_1563,N_3985);
and U8282 (N_8282,N_13,N_2608);
or U8283 (N_8283,N_3775,N_4197);
or U8284 (N_8284,N_1863,N_2571);
nor U8285 (N_8285,N_3256,N_1124);
nand U8286 (N_8286,N_2513,N_4390);
nand U8287 (N_8287,N_2316,N_1703);
nor U8288 (N_8288,N_607,N_3712);
xnor U8289 (N_8289,N_4043,N_3844);
xor U8290 (N_8290,N_3092,N_3194);
and U8291 (N_8291,N_2471,N_39);
nor U8292 (N_8292,N_969,N_1238);
nor U8293 (N_8293,N_3835,N_4220);
nor U8294 (N_8294,N_2639,N_194);
nand U8295 (N_8295,N_2683,N_525);
or U8296 (N_8296,N_336,N_4084);
nand U8297 (N_8297,N_2131,N_2428);
xor U8298 (N_8298,N_1617,N_4521);
nor U8299 (N_8299,N_2011,N_3291);
and U8300 (N_8300,N_643,N_4720);
or U8301 (N_8301,N_1930,N_4449);
and U8302 (N_8302,N_4369,N_3032);
or U8303 (N_8303,N_2186,N_636);
xnor U8304 (N_8304,N_903,N_607);
or U8305 (N_8305,N_3225,N_4875);
or U8306 (N_8306,N_4788,N_1210);
or U8307 (N_8307,N_2733,N_4152);
and U8308 (N_8308,N_3876,N_1637);
nand U8309 (N_8309,N_4870,N_950);
or U8310 (N_8310,N_540,N_4219);
and U8311 (N_8311,N_4547,N_3569);
or U8312 (N_8312,N_1685,N_1360);
nand U8313 (N_8313,N_4647,N_69);
or U8314 (N_8314,N_1145,N_1923);
and U8315 (N_8315,N_4867,N_4194);
or U8316 (N_8316,N_4983,N_3733);
nor U8317 (N_8317,N_3288,N_3888);
nand U8318 (N_8318,N_4616,N_4158);
nand U8319 (N_8319,N_3574,N_4864);
nor U8320 (N_8320,N_4454,N_4074);
nand U8321 (N_8321,N_2551,N_4692);
nor U8322 (N_8322,N_2883,N_2805);
xor U8323 (N_8323,N_3362,N_4886);
nand U8324 (N_8324,N_926,N_753);
nand U8325 (N_8325,N_4760,N_1026);
and U8326 (N_8326,N_2466,N_4672);
or U8327 (N_8327,N_3714,N_80);
nand U8328 (N_8328,N_3970,N_4646);
or U8329 (N_8329,N_1488,N_2523);
or U8330 (N_8330,N_280,N_897);
or U8331 (N_8331,N_3099,N_433);
or U8332 (N_8332,N_4769,N_1647);
or U8333 (N_8333,N_43,N_4867);
xnor U8334 (N_8334,N_3168,N_1338);
nor U8335 (N_8335,N_4552,N_2640);
or U8336 (N_8336,N_3162,N_2221);
nand U8337 (N_8337,N_4941,N_1258);
or U8338 (N_8338,N_467,N_3214);
nand U8339 (N_8339,N_477,N_1733);
or U8340 (N_8340,N_3110,N_3256);
nand U8341 (N_8341,N_4256,N_2992);
or U8342 (N_8342,N_1759,N_46);
nor U8343 (N_8343,N_227,N_147);
and U8344 (N_8344,N_1978,N_4196);
nor U8345 (N_8345,N_698,N_4271);
nand U8346 (N_8346,N_488,N_383);
and U8347 (N_8347,N_4477,N_233);
nor U8348 (N_8348,N_4495,N_1529);
and U8349 (N_8349,N_134,N_2176);
and U8350 (N_8350,N_3105,N_1038);
xnor U8351 (N_8351,N_171,N_2644);
and U8352 (N_8352,N_4143,N_477);
or U8353 (N_8353,N_2483,N_4757);
nand U8354 (N_8354,N_2815,N_4846);
nand U8355 (N_8355,N_874,N_2635);
nand U8356 (N_8356,N_4860,N_3894);
or U8357 (N_8357,N_2424,N_1608);
nand U8358 (N_8358,N_4399,N_2923);
and U8359 (N_8359,N_2959,N_3337);
and U8360 (N_8360,N_1881,N_1050);
and U8361 (N_8361,N_1732,N_4161);
and U8362 (N_8362,N_2335,N_4160);
nand U8363 (N_8363,N_578,N_3410);
xor U8364 (N_8364,N_2383,N_899);
nand U8365 (N_8365,N_3642,N_1132);
nand U8366 (N_8366,N_4229,N_4609);
nor U8367 (N_8367,N_670,N_4518);
or U8368 (N_8368,N_677,N_4489);
or U8369 (N_8369,N_2170,N_2868);
and U8370 (N_8370,N_4825,N_3482);
or U8371 (N_8371,N_3272,N_4705);
nand U8372 (N_8372,N_3167,N_85);
nand U8373 (N_8373,N_1713,N_2392);
and U8374 (N_8374,N_4519,N_2784);
nor U8375 (N_8375,N_3961,N_3690);
and U8376 (N_8376,N_3882,N_56);
nor U8377 (N_8377,N_2172,N_2909);
xnor U8378 (N_8378,N_4211,N_172);
nor U8379 (N_8379,N_2553,N_4872);
nor U8380 (N_8380,N_4824,N_2591);
nand U8381 (N_8381,N_1428,N_1491);
nand U8382 (N_8382,N_1274,N_4365);
and U8383 (N_8383,N_1912,N_4160);
nor U8384 (N_8384,N_3937,N_4009);
and U8385 (N_8385,N_1274,N_2630);
nand U8386 (N_8386,N_1224,N_2197);
nor U8387 (N_8387,N_2659,N_3703);
xnor U8388 (N_8388,N_1729,N_2963);
nor U8389 (N_8389,N_3776,N_2087);
nor U8390 (N_8390,N_1168,N_3140);
nor U8391 (N_8391,N_4693,N_4923);
and U8392 (N_8392,N_2053,N_386);
nand U8393 (N_8393,N_2272,N_2331);
and U8394 (N_8394,N_4538,N_3290);
and U8395 (N_8395,N_2772,N_3846);
and U8396 (N_8396,N_1798,N_818);
and U8397 (N_8397,N_927,N_3197);
xnor U8398 (N_8398,N_3927,N_3801);
or U8399 (N_8399,N_1936,N_2332);
and U8400 (N_8400,N_983,N_3840);
nand U8401 (N_8401,N_3428,N_2077);
nor U8402 (N_8402,N_4374,N_3184);
and U8403 (N_8403,N_2966,N_2055);
nand U8404 (N_8404,N_1442,N_3732);
and U8405 (N_8405,N_939,N_2205);
and U8406 (N_8406,N_1408,N_3960);
or U8407 (N_8407,N_4570,N_3583);
and U8408 (N_8408,N_1323,N_3031);
or U8409 (N_8409,N_962,N_4830);
and U8410 (N_8410,N_851,N_3989);
and U8411 (N_8411,N_4101,N_1789);
nand U8412 (N_8412,N_3758,N_2026);
and U8413 (N_8413,N_2624,N_1403);
or U8414 (N_8414,N_4444,N_3453);
or U8415 (N_8415,N_1889,N_2295);
and U8416 (N_8416,N_3079,N_478);
nor U8417 (N_8417,N_1085,N_960);
or U8418 (N_8418,N_3192,N_4710);
nor U8419 (N_8419,N_2646,N_1230);
or U8420 (N_8420,N_4467,N_1792);
or U8421 (N_8421,N_840,N_3808);
xor U8422 (N_8422,N_98,N_8);
nand U8423 (N_8423,N_3349,N_2003);
nor U8424 (N_8424,N_3709,N_3349);
xor U8425 (N_8425,N_1073,N_344);
nand U8426 (N_8426,N_4819,N_4217);
xor U8427 (N_8427,N_2789,N_3980);
nand U8428 (N_8428,N_2044,N_1709);
or U8429 (N_8429,N_3253,N_1558);
nor U8430 (N_8430,N_3841,N_439);
xnor U8431 (N_8431,N_4255,N_3025);
nor U8432 (N_8432,N_2955,N_174);
nor U8433 (N_8433,N_1665,N_2094);
and U8434 (N_8434,N_2602,N_1538);
nor U8435 (N_8435,N_1012,N_1182);
or U8436 (N_8436,N_4244,N_1895);
nor U8437 (N_8437,N_1973,N_1256);
nand U8438 (N_8438,N_269,N_2634);
or U8439 (N_8439,N_1034,N_1674);
nand U8440 (N_8440,N_628,N_3348);
nor U8441 (N_8441,N_1155,N_1205);
nand U8442 (N_8442,N_1906,N_3129);
nand U8443 (N_8443,N_3021,N_150);
or U8444 (N_8444,N_4623,N_3271);
nand U8445 (N_8445,N_3946,N_3548);
nor U8446 (N_8446,N_1385,N_2822);
xnor U8447 (N_8447,N_229,N_1232);
and U8448 (N_8448,N_4977,N_2717);
nand U8449 (N_8449,N_4348,N_1763);
xnor U8450 (N_8450,N_2619,N_4043);
or U8451 (N_8451,N_4680,N_2897);
and U8452 (N_8452,N_200,N_485);
nand U8453 (N_8453,N_615,N_2470);
and U8454 (N_8454,N_3915,N_850);
and U8455 (N_8455,N_4593,N_308);
nor U8456 (N_8456,N_4409,N_4932);
nor U8457 (N_8457,N_165,N_1083);
nand U8458 (N_8458,N_3488,N_2472);
nand U8459 (N_8459,N_1625,N_2788);
nand U8460 (N_8460,N_4599,N_3375);
nand U8461 (N_8461,N_1316,N_4741);
nor U8462 (N_8462,N_4201,N_1093);
xnor U8463 (N_8463,N_1564,N_4840);
nand U8464 (N_8464,N_2382,N_348);
nand U8465 (N_8465,N_4332,N_3462);
or U8466 (N_8466,N_703,N_1628);
or U8467 (N_8467,N_3522,N_4587);
nand U8468 (N_8468,N_3089,N_215);
nand U8469 (N_8469,N_1047,N_683);
xor U8470 (N_8470,N_2211,N_703);
or U8471 (N_8471,N_2937,N_3873);
and U8472 (N_8472,N_3720,N_3229);
nor U8473 (N_8473,N_3959,N_258);
and U8474 (N_8474,N_2715,N_2832);
and U8475 (N_8475,N_688,N_805);
xor U8476 (N_8476,N_3539,N_310);
nand U8477 (N_8477,N_4239,N_2984);
or U8478 (N_8478,N_2877,N_2070);
or U8479 (N_8479,N_2632,N_1207);
and U8480 (N_8480,N_4014,N_2454);
nand U8481 (N_8481,N_564,N_4796);
nor U8482 (N_8482,N_1310,N_1243);
xor U8483 (N_8483,N_2583,N_636);
or U8484 (N_8484,N_3204,N_1651);
nor U8485 (N_8485,N_221,N_1809);
nand U8486 (N_8486,N_2634,N_4011);
and U8487 (N_8487,N_2245,N_1528);
nor U8488 (N_8488,N_2413,N_1205);
xor U8489 (N_8489,N_3402,N_4935);
xnor U8490 (N_8490,N_180,N_344);
and U8491 (N_8491,N_3964,N_1199);
and U8492 (N_8492,N_3116,N_3579);
nand U8493 (N_8493,N_2650,N_3971);
nand U8494 (N_8494,N_1021,N_927);
nand U8495 (N_8495,N_1798,N_1691);
or U8496 (N_8496,N_2524,N_131);
nand U8497 (N_8497,N_2507,N_4490);
xor U8498 (N_8498,N_3318,N_1697);
nand U8499 (N_8499,N_4907,N_4905);
and U8500 (N_8500,N_4645,N_1658);
xor U8501 (N_8501,N_2285,N_3081);
nand U8502 (N_8502,N_3740,N_657);
nor U8503 (N_8503,N_433,N_4323);
and U8504 (N_8504,N_3406,N_588);
and U8505 (N_8505,N_542,N_526);
nand U8506 (N_8506,N_3207,N_3099);
nand U8507 (N_8507,N_1463,N_408);
or U8508 (N_8508,N_4146,N_3000);
or U8509 (N_8509,N_3254,N_165);
or U8510 (N_8510,N_31,N_4488);
nor U8511 (N_8511,N_4644,N_3478);
or U8512 (N_8512,N_1893,N_4899);
nor U8513 (N_8513,N_336,N_1165);
or U8514 (N_8514,N_562,N_2506);
or U8515 (N_8515,N_1033,N_1802);
and U8516 (N_8516,N_3753,N_2328);
nand U8517 (N_8517,N_4955,N_4768);
nor U8518 (N_8518,N_4254,N_1108);
or U8519 (N_8519,N_2932,N_4355);
nand U8520 (N_8520,N_1293,N_718);
and U8521 (N_8521,N_3060,N_57);
and U8522 (N_8522,N_3146,N_3503);
xnor U8523 (N_8523,N_110,N_1346);
nor U8524 (N_8524,N_4183,N_1259);
nor U8525 (N_8525,N_121,N_4096);
or U8526 (N_8526,N_4493,N_4157);
xnor U8527 (N_8527,N_4819,N_335);
nand U8528 (N_8528,N_3574,N_1788);
or U8529 (N_8529,N_4507,N_3451);
and U8530 (N_8530,N_3162,N_984);
nor U8531 (N_8531,N_4661,N_2363);
and U8532 (N_8532,N_1699,N_538);
xor U8533 (N_8533,N_1677,N_4123);
or U8534 (N_8534,N_3393,N_351);
xnor U8535 (N_8535,N_290,N_3232);
nor U8536 (N_8536,N_1379,N_378);
and U8537 (N_8537,N_2775,N_3493);
and U8538 (N_8538,N_3668,N_4473);
nor U8539 (N_8539,N_350,N_146);
nand U8540 (N_8540,N_2003,N_4047);
nor U8541 (N_8541,N_4734,N_116);
xor U8542 (N_8542,N_2596,N_2826);
nor U8543 (N_8543,N_1917,N_1492);
and U8544 (N_8544,N_1436,N_3002);
xor U8545 (N_8545,N_885,N_1423);
and U8546 (N_8546,N_3299,N_530);
or U8547 (N_8547,N_2106,N_2667);
nand U8548 (N_8548,N_595,N_2789);
and U8549 (N_8549,N_223,N_1827);
or U8550 (N_8550,N_2395,N_2334);
nor U8551 (N_8551,N_2040,N_2011);
and U8552 (N_8552,N_4579,N_1828);
xnor U8553 (N_8553,N_2322,N_4841);
nand U8554 (N_8554,N_3195,N_1204);
and U8555 (N_8555,N_1243,N_1196);
or U8556 (N_8556,N_1136,N_2916);
nor U8557 (N_8557,N_1423,N_4230);
nor U8558 (N_8558,N_3388,N_4371);
xor U8559 (N_8559,N_2663,N_2722);
nand U8560 (N_8560,N_945,N_1565);
nor U8561 (N_8561,N_2493,N_3974);
nand U8562 (N_8562,N_1610,N_3152);
nor U8563 (N_8563,N_1906,N_1716);
and U8564 (N_8564,N_1249,N_1547);
nand U8565 (N_8565,N_3731,N_3649);
and U8566 (N_8566,N_689,N_1516);
nand U8567 (N_8567,N_861,N_1029);
nand U8568 (N_8568,N_3346,N_3455);
or U8569 (N_8569,N_128,N_3066);
and U8570 (N_8570,N_1607,N_1289);
nand U8571 (N_8571,N_2935,N_2747);
and U8572 (N_8572,N_1004,N_2532);
or U8573 (N_8573,N_3874,N_1526);
and U8574 (N_8574,N_4922,N_4115);
xnor U8575 (N_8575,N_959,N_2126);
nor U8576 (N_8576,N_2305,N_4409);
nor U8577 (N_8577,N_4526,N_2868);
or U8578 (N_8578,N_888,N_1476);
or U8579 (N_8579,N_1140,N_4811);
nand U8580 (N_8580,N_1522,N_4998);
or U8581 (N_8581,N_3593,N_4637);
nor U8582 (N_8582,N_814,N_3174);
nor U8583 (N_8583,N_4775,N_4537);
or U8584 (N_8584,N_1966,N_3279);
nand U8585 (N_8585,N_4555,N_196);
or U8586 (N_8586,N_856,N_4225);
xnor U8587 (N_8587,N_1204,N_3552);
and U8588 (N_8588,N_502,N_2105);
nor U8589 (N_8589,N_992,N_4406);
and U8590 (N_8590,N_65,N_2155);
and U8591 (N_8591,N_3135,N_4603);
or U8592 (N_8592,N_3785,N_764);
nand U8593 (N_8593,N_2210,N_467);
nor U8594 (N_8594,N_1303,N_4412);
and U8595 (N_8595,N_242,N_4150);
nor U8596 (N_8596,N_1852,N_3966);
and U8597 (N_8597,N_1355,N_793);
and U8598 (N_8598,N_180,N_2724);
nand U8599 (N_8599,N_2563,N_162);
or U8600 (N_8600,N_3896,N_4986);
and U8601 (N_8601,N_2413,N_3740);
and U8602 (N_8602,N_4517,N_3086);
nor U8603 (N_8603,N_5,N_3140);
and U8604 (N_8604,N_4369,N_4509);
nor U8605 (N_8605,N_3281,N_287);
and U8606 (N_8606,N_1705,N_4295);
nor U8607 (N_8607,N_3777,N_3294);
nor U8608 (N_8608,N_2030,N_3855);
and U8609 (N_8609,N_1225,N_449);
or U8610 (N_8610,N_178,N_1996);
nor U8611 (N_8611,N_2869,N_1014);
or U8612 (N_8612,N_2538,N_3769);
and U8613 (N_8613,N_1378,N_306);
nand U8614 (N_8614,N_3754,N_633);
nand U8615 (N_8615,N_1523,N_2088);
nor U8616 (N_8616,N_1718,N_3531);
or U8617 (N_8617,N_3003,N_1736);
xnor U8618 (N_8618,N_4797,N_11);
and U8619 (N_8619,N_2593,N_3927);
nand U8620 (N_8620,N_4180,N_2001);
nor U8621 (N_8621,N_403,N_721);
or U8622 (N_8622,N_2717,N_3029);
nand U8623 (N_8623,N_1001,N_2955);
xor U8624 (N_8624,N_1976,N_4008);
or U8625 (N_8625,N_3028,N_3717);
nor U8626 (N_8626,N_4892,N_261);
or U8627 (N_8627,N_4918,N_1478);
and U8628 (N_8628,N_2968,N_4461);
or U8629 (N_8629,N_3541,N_4459);
or U8630 (N_8630,N_580,N_1884);
and U8631 (N_8631,N_4097,N_3009);
xnor U8632 (N_8632,N_4498,N_1023);
or U8633 (N_8633,N_1881,N_3252);
or U8634 (N_8634,N_947,N_881);
nand U8635 (N_8635,N_3767,N_1976);
nor U8636 (N_8636,N_3068,N_4245);
or U8637 (N_8637,N_3143,N_654);
and U8638 (N_8638,N_1654,N_1770);
and U8639 (N_8639,N_4979,N_1916);
and U8640 (N_8640,N_1552,N_4529);
nor U8641 (N_8641,N_4881,N_85);
nor U8642 (N_8642,N_3451,N_20);
and U8643 (N_8643,N_2468,N_2928);
nor U8644 (N_8644,N_886,N_17);
nor U8645 (N_8645,N_56,N_3897);
nor U8646 (N_8646,N_1634,N_224);
nor U8647 (N_8647,N_977,N_3529);
nor U8648 (N_8648,N_88,N_2615);
nand U8649 (N_8649,N_2816,N_3512);
or U8650 (N_8650,N_1352,N_2050);
nor U8651 (N_8651,N_339,N_3235);
nand U8652 (N_8652,N_3304,N_1051);
and U8653 (N_8653,N_1316,N_2158);
nand U8654 (N_8654,N_940,N_491);
and U8655 (N_8655,N_176,N_2037);
nand U8656 (N_8656,N_2063,N_1142);
nand U8657 (N_8657,N_2050,N_272);
or U8658 (N_8658,N_32,N_1935);
and U8659 (N_8659,N_1812,N_4325);
or U8660 (N_8660,N_4111,N_1472);
nor U8661 (N_8661,N_618,N_3896);
nor U8662 (N_8662,N_3889,N_2863);
nor U8663 (N_8663,N_102,N_3564);
nand U8664 (N_8664,N_74,N_3820);
nand U8665 (N_8665,N_4770,N_3716);
nor U8666 (N_8666,N_1241,N_3509);
or U8667 (N_8667,N_4805,N_247);
xnor U8668 (N_8668,N_1468,N_2871);
and U8669 (N_8669,N_562,N_2868);
nor U8670 (N_8670,N_756,N_252);
nor U8671 (N_8671,N_4883,N_4935);
nand U8672 (N_8672,N_3735,N_4622);
or U8673 (N_8673,N_2647,N_2961);
nand U8674 (N_8674,N_1390,N_2367);
nand U8675 (N_8675,N_3951,N_371);
nor U8676 (N_8676,N_30,N_674);
and U8677 (N_8677,N_3187,N_4861);
xor U8678 (N_8678,N_310,N_829);
or U8679 (N_8679,N_3803,N_528);
nand U8680 (N_8680,N_3157,N_3131);
nand U8681 (N_8681,N_4621,N_16);
or U8682 (N_8682,N_4871,N_1257);
and U8683 (N_8683,N_2943,N_2409);
and U8684 (N_8684,N_643,N_3515);
nor U8685 (N_8685,N_1964,N_861);
nor U8686 (N_8686,N_4602,N_3377);
and U8687 (N_8687,N_1773,N_4407);
and U8688 (N_8688,N_3495,N_2795);
or U8689 (N_8689,N_1451,N_275);
and U8690 (N_8690,N_1705,N_1789);
nand U8691 (N_8691,N_4720,N_1735);
nor U8692 (N_8692,N_499,N_873);
xnor U8693 (N_8693,N_1789,N_2414);
or U8694 (N_8694,N_3583,N_4697);
nor U8695 (N_8695,N_3416,N_3175);
and U8696 (N_8696,N_4603,N_448);
or U8697 (N_8697,N_45,N_1565);
nand U8698 (N_8698,N_1958,N_4003);
nor U8699 (N_8699,N_4271,N_1614);
nand U8700 (N_8700,N_2201,N_3111);
and U8701 (N_8701,N_4275,N_1538);
and U8702 (N_8702,N_4830,N_960);
nand U8703 (N_8703,N_1698,N_845);
nor U8704 (N_8704,N_3389,N_3360);
or U8705 (N_8705,N_4985,N_2329);
or U8706 (N_8706,N_662,N_1095);
and U8707 (N_8707,N_3688,N_3046);
or U8708 (N_8708,N_2551,N_133);
and U8709 (N_8709,N_3070,N_2100);
nand U8710 (N_8710,N_2488,N_3564);
nor U8711 (N_8711,N_362,N_1623);
nor U8712 (N_8712,N_1189,N_647);
or U8713 (N_8713,N_2291,N_1300);
and U8714 (N_8714,N_3685,N_4831);
xnor U8715 (N_8715,N_4736,N_4504);
nor U8716 (N_8716,N_4100,N_4743);
nand U8717 (N_8717,N_4400,N_3314);
nand U8718 (N_8718,N_4144,N_3740);
nor U8719 (N_8719,N_3344,N_963);
nor U8720 (N_8720,N_1852,N_2168);
or U8721 (N_8721,N_1867,N_2021);
xnor U8722 (N_8722,N_2339,N_720);
nor U8723 (N_8723,N_3331,N_4050);
or U8724 (N_8724,N_91,N_2475);
nand U8725 (N_8725,N_1858,N_4720);
nor U8726 (N_8726,N_540,N_525);
or U8727 (N_8727,N_3137,N_1503);
nand U8728 (N_8728,N_337,N_2184);
nand U8729 (N_8729,N_1883,N_183);
and U8730 (N_8730,N_3168,N_2972);
or U8731 (N_8731,N_2546,N_3982);
nand U8732 (N_8732,N_346,N_1864);
or U8733 (N_8733,N_595,N_1182);
nor U8734 (N_8734,N_4630,N_1821);
and U8735 (N_8735,N_3246,N_4130);
nor U8736 (N_8736,N_3127,N_3832);
nor U8737 (N_8737,N_1334,N_3422);
nor U8738 (N_8738,N_4608,N_1162);
and U8739 (N_8739,N_619,N_2960);
nand U8740 (N_8740,N_1351,N_2109);
nand U8741 (N_8741,N_1004,N_1467);
xnor U8742 (N_8742,N_2877,N_596);
or U8743 (N_8743,N_4083,N_2074);
nand U8744 (N_8744,N_1917,N_504);
or U8745 (N_8745,N_1978,N_3782);
nand U8746 (N_8746,N_503,N_2613);
nand U8747 (N_8747,N_1438,N_984);
xnor U8748 (N_8748,N_336,N_4228);
or U8749 (N_8749,N_4727,N_2363);
nand U8750 (N_8750,N_1276,N_3321);
and U8751 (N_8751,N_3718,N_3757);
or U8752 (N_8752,N_54,N_4161);
nand U8753 (N_8753,N_3145,N_2836);
or U8754 (N_8754,N_81,N_3910);
nand U8755 (N_8755,N_3488,N_4446);
or U8756 (N_8756,N_1255,N_1456);
nand U8757 (N_8757,N_2174,N_433);
nor U8758 (N_8758,N_1370,N_706);
or U8759 (N_8759,N_1275,N_2286);
nand U8760 (N_8760,N_4603,N_157);
or U8761 (N_8761,N_3543,N_3011);
nand U8762 (N_8762,N_725,N_2999);
or U8763 (N_8763,N_474,N_4270);
nand U8764 (N_8764,N_2469,N_4196);
nor U8765 (N_8765,N_1817,N_4017);
and U8766 (N_8766,N_2411,N_1947);
nor U8767 (N_8767,N_2892,N_1640);
nand U8768 (N_8768,N_2888,N_1763);
xnor U8769 (N_8769,N_4701,N_4471);
and U8770 (N_8770,N_2273,N_1891);
nor U8771 (N_8771,N_3661,N_3779);
nor U8772 (N_8772,N_3356,N_4366);
nand U8773 (N_8773,N_3945,N_4502);
and U8774 (N_8774,N_3013,N_3050);
or U8775 (N_8775,N_3214,N_4070);
nand U8776 (N_8776,N_991,N_2865);
and U8777 (N_8777,N_3878,N_4350);
nand U8778 (N_8778,N_762,N_2511);
or U8779 (N_8779,N_1835,N_87);
and U8780 (N_8780,N_3136,N_4566);
nor U8781 (N_8781,N_3905,N_378);
and U8782 (N_8782,N_601,N_205);
and U8783 (N_8783,N_642,N_764);
or U8784 (N_8784,N_4568,N_848);
nand U8785 (N_8785,N_1241,N_4481);
and U8786 (N_8786,N_4073,N_2693);
or U8787 (N_8787,N_2818,N_4318);
nand U8788 (N_8788,N_3282,N_1364);
nand U8789 (N_8789,N_723,N_2063);
nor U8790 (N_8790,N_141,N_4706);
or U8791 (N_8791,N_4549,N_3246);
or U8792 (N_8792,N_1839,N_3505);
nor U8793 (N_8793,N_4413,N_546);
and U8794 (N_8794,N_3773,N_4584);
and U8795 (N_8795,N_2822,N_3053);
xor U8796 (N_8796,N_279,N_770);
or U8797 (N_8797,N_2155,N_930);
nor U8798 (N_8798,N_3386,N_1253);
nand U8799 (N_8799,N_410,N_4025);
nor U8800 (N_8800,N_3695,N_10);
nor U8801 (N_8801,N_2452,N_3362);
nand U8802 (N_8802,N_1754,N_3255);
and U8803 (N_8803,N_2979,N_4490);
nor U8804 (N_8804,N_2696,N_2974);
xor U8805 (N_8805,N_311,N_1010);
or U8806 (N_8806,N_3490,N_2444);
nor U8807 (N_8807,N_257,N_2328);
nor U8808 (N_8808,N_4411,N_3193);
nor U8809 (N_8809,N_4540,N_916);
nand U8810 (N_8810,N_852,N_2868);
and U8811 (N_8811,N_4186,N_929);
nand U8812 (N_8812,N_394,N_3325);
nor U8813 (N_8813,N_165,N_236);
or U8814 (N_8814,N_4174,N_1973);
xor U8815 (N_8815,N_4892,N_686);
nor U8816 (N_8816,N_3237,N_2048);
or U8817 (N_8817,N_1077,N_2791);
nand U8818 (N_8818,N_3588,N_1401);
nand U8819 (N_8819,N_4488,N_2989);
nand U8820 (N_8820,N_4360,N_4130);
nand U8821 (N_8821,N_233,N_347);
or U8822 (N_8822,N_555,N_3008);
or U8823 (N_8823,N_1784,N_3339);
nor U8824 (N_8824,N_4291,N_1370);
or U8825 (N_8825,N_3824,N_1472);
nand U8826 (N_8826,N_1941,N_2140);
and U8827 (N_8827,N_232,N_3135);
nor U8828 (N_8828,N_2291,N_4934);
nor U8829 (N_8829,N_4321,N_2052);
and U8830 (N_8830,N_1645,N_1164);
nor U8831 (N_8831,N_784,N_1278);
nor U8832 (N_8832,N_2190,N_2384);
and U8833 (N_8833,N_2778,N_4224);
and U8834 (N_8834,N_1047,N_1440);
nor U8835 (N_8835,N_4246,N_432);
nor U8836 (N_8836,N_2315,N_4777);
or U8837 (N_8837,N_1154,N_410);
and U8838 (N_8838,N_10,N_1033);
and U8839 (N_8839,N_1267,N_1205);
and U8840 (N_8840,N_515,N_3302);
and U8841 (N_8841,N_2475,N_2982);
nor U8842 (N_8842,N_2762,N_1016);
xnor U8843 (N_8843,N_1764,N_1032);
nand U8844 (N_8844,N_1364,N_1348);
and U8845 (N_8845,N_3590,N_1449);
nor U8846 (N_8846,N_139,N_196);
xor U8847 (N_8847,N_1299,N_2326);
nand U8848 (N_8848,N_13,N_4614);
and U8849 (N_8849,N_3327,N_4767);
or U8850 (N_8850,N_3021,N_3732);
and U8851 (N_8851,N_3235,N_2759);
nor U8852 (N_8852,N_1000,N_4912);
nand U8853 (N_8853,N_4285,N_2278);
xnor U8854 (N_8854,N_3308,N_1022);
or U8855 (N_8855,N_4902,N_4452);
and U8856 (N_8856,N_2041,N_3351);
and U8857 (N_8857,N_3925,N_426);
nand U8858 (N_8858,N_860,N_4568);
nand U8859 (N_8859,N_2891,N_318);
xnor U8860 (N_8860,N_2398,N_733);
or U8861 (N_8861,N_4885,N_1735);
nor U8862 (N_8862,N_4840,N_2444);
or U8863 (N_8863,N_4216,N_3048);
and U8864 (N_8864,N_381,N_2347);
and U8865 (N_8865,N_2284,N_2780);
nor U8866 (N_8866,N_765,N_4737);
or U8867 (N_8867,N_3043,N_2578);
nor U8868 (N_8868,N_3068,N_1564);
nand U8869 (N_8869,N_4383,N_4803);
nor U8870 (N_8870,N_1053,N_3955);
nand U8871 (N_8871,N_1147,N_4828);
or U8872 (N_8872,N_2212,N_1151);
and U8873 (N_8873,N_340,N_972);
xnor U8874 (N_8874,N_2968,N_136);
nor U8875 (N_8875,N_2217,N_4086);
xnor U8876 (N_8876,N_4687,N_4994);
xnor U8877 (N_8877,N_4731,N_111);
xor U8878 (N_8878,N_1484,N_4845);
xnor U8879 (N_8879,N_3019,N_1230);
nand U8880 (N_8880,N_4323,N_3045);
nor U8881 (N_8881,N_3691,N_2153);
nand U8882 (N_8882,N_2099,N_2950);
nand U8883 (N_8883,N_1057,N_1206);
nor U8884 (N_8884,N_2102,N_467);
or U8885 (N_8885,N_3779,N_2313);
and U8886 (N_8886,N_2268,N_2709);
and U8887 (N_8887,N_776,N_1444);
nand U8888 (N_8888,N_4671,N_430);
and U8889 (N_8889,N_27,N_753);
and U8890 (N_8890,N_2538,N_1151);
and U8891 (N_8891,N_1846,N_4405);
nand U8892 (N_8892,N_2421,N_240);
and U8893 (N_8893,N_4603,N_2138);
xnor U8894 (N_8894,N_1827,N_3782);
or U8895 (N_8895,N_4306,N_2147);
and U8896 (N_8896,N_3375,N_2368);
xnor U8897 (N_8897,N_1699,N_2898);
and U8898 (N_8898,N_3585,N_441);
or U8899 (N_8899,N_1524,N_1635);
nand U8900 (N_8900,N_2081,N_2007);
nor U8901 (N_8901,N_2444,N_4073);
and U8902 (N_8902,N_237,N_1901);
nand U8903 (N_8903,N_4094,N_2027);
and U8904 (N_8904,N_2190,N_825);
nand U8905 (N_8905,N_4541,N_1850);
nor U8906 (N_8906,N_2242,N_768);
or U8907 (N_8907,N_3572,N_3207);
nand U8908 (N_8908,N_2101,N_1636);
and U8909 (N_8909,N_2791,N_730);
and U8910 (N_8910,N_576,N_3022);
or U8911 (N_8911,N_4124,N_2976);
nor U8912 (N_8912,N_36,N_1414);
and U8913 (N_8913,N_503,N_990);
nor U8914 (N_8914,N_4950,N_3916);
nand U8915 (N_8915,N_769,N_245);
nand U8916 (N_8916,N_86,N_4903);
xnor U8917 (N_8917,N_3569,N_509);
or U8918 (N_8918,N_422,N_3746);
xnor U8919 (N_8919,N_1875,N_2557);
or U8920 (N_8920,N_1913,N_967);
or U8921 (N_8921,N_517,N_4696);
or U8922 (N_8922,N_744,N_456);
and U8923 (N_8923,N_2612,N_4680);
xor U8924 (N_8924,N_736,N_925);
and U8925 (N_8925,N_1341,N_4400);
nor U8926 (N_8926,N_4735,N_2342);
nand U8927 (N_8927,N_3355,N_759);
nor U8928 (N_8928,N_3272,N_4461);
and U8929 (N_8929,N_2820,N_3005);
or U8930 (N_8930,N_4011,N_2910);
nand U8931 (N_8931,N_2980,N_4600);
or U8932 (N_8932,N_3208,N_3993);
or U8933 (N_8933,N_4838,N_4022);
nand U8934 (N_8934,N_2884,N_2013);
or U8935 (N_8935,N_4116,N_2640);
or U8936 (N_8936,N_2252,N_325);
or U8937 (N_8937,N_1981,N_3945);
xnor U8938 (N_8938,N_888,N_1905);
or U8939 (N_8939,N_2722,N_1871);
nor U8940 (N_8940,N_396,N_39);
nor U8941 (N_8941,N_2344,N_1812);
and U8942 (N_8942,N_1567,N_3038);
nand U8943 (N_8943,N_4814,N_2636);
nand U8944 (N_8944,N_2895,N_175);
and U8945 (N_8945,N_701,N_2127);
or U8946 (N_8946,N_2408,N_2011);
nor U8947 (N_8947,N_2458,N_1880);
nand U8948 (N_8948,N_3568,N_320);
nand U8949 (N_8949,N_1153,N_2527);
nand U8950 (N_8950,N_3645,N_4391);
nand U8951 (N_8951,N_2183,N_1601);
nand U8952 (N_8952,N_4135,N_3746);
or U8953 (N_8953,N_4388,N_1885);
xnor U8954 (N_8954,N_1476,N_3570);
nand U8955 (N_8955,N_3679,N_250);
and U8956 (N_8956,N_2337,N_3865);
nor U8957 (N_8957,N_4769,N_260);
or U8958 (N_8958,N_3704,N_364);
and U8959 (N_8959,N_245,N_90);
xor U8960 (N_8960,N_2861,N_1097);
or U8961 (N_8961,N_1362,N_2218);
xor U8962 (N_8962,N_2152,N_1624);
and U8963 (N_8963,N_619,N_2611);
nor U8964 (N_8964,N_3364,N_3939);
nor U8965 (N_8965,N_723,N_1226);
and U8966 (N_8966,N_2060,N_3502);
and U8967 (N_8967,N_1061,N_1230);
nand U8968 (N_8968,N_1965,N_4458);
and U8969 (N_8969,N_3488,N_259);
nor U8970 (N_8970,N_707,N_2347);
nand U8971 (N_8971,N_993,N_2135);
xnor U8972 (N_8972,N_2926,N_2236);
nand U8973 (N_8973,N_300,N_4546);
nor U8974 (N_8974,N_608,N_2330);
nor U8975 (N_8975,N_2371,N_1066);
nor U8976 (N_8976,N_3502,N_4268);
nor U8977 (N_8977,N_2956,N_4035);
nand U8978 (N_8978,N_1959,N_3235);
xnor U8979 (N_8979,N_2279,N_998);
xor U8980 (N_8980,N_3115,N_381);
nor U8981 (N_8981,N_1290,N_4587);
and U8982 (N_8982,N_4604,N_4453);
and U8983 (N_8983,N_843,N_459);
nand U8984 (N_8984,N_2900,N_2678);
nor U8985 (N_8985,N_3697,N_1020);
or U8986 (N_8986,N_1836,N_17);
or U8987 (N_8987,N_3915,N_329);
nand U8988 (N_8988,N_2871,N_4851);
nor U8989 (N_8989,N_1338,N_2263);
xnor U8990 (N_8990,N_2836,N_3994);
nand U8991 (N_8991,N_784,N_2032);
and U8992 (N_8992,N_2591,N_930);
nor U8993 (N_8993,N_695,N_835);
or U8994 (N_8994,N_4306,N_4895);
nand U8995 (N_8995,N_3943,N_2460);
or U8996 (N_8996,N_735,N_1376);
or U8997 (N_8997,N_4652,N_304);
and U8998 (N_8998,N_1790,N_985);
xor U8999 (N_8999,N_2086,N_3554);
and U9000 (N_9000,N_3184,N_3076);
xor U9001 (N_9001,N_2197,N_1948);
and U9002 (N_9002,N_1132,N_4384);
and U9003 (N_9003,N_804,N_416);
nor U9004 (N_9004,N_153,N_3052);
and U9005 (N_9005,N_886,N_4079);
or U9006 (N_9006,N_3896,N_3170);
xor U9007 (N_9007,N_4750,N_1348);
and U9008 (N_9008,N_3649,N_3856);
or U9009 (N_9009,N_2997,N_533);
and U9010 (N_9010,N_1546,N_4385);
or U9011 (N_9011,N_3254,N_3161);
nor U9012 (N_9012,N_4991,N_587);
and U9013 (N_9013,N_1795,N_193);
and U9014 (N_9014,N_1315,N_1229);
or U9015 (N_9015,N_3389,N_671);
and U9016 (N_9016,N_3475,N_3994);
or U9017 (N_9017,N_810,N_1918);
and U9018 (N_9018,N_535,N_1369);
or U9019 (N_9019,N_743,N_2825);
nor U9020 (N_9020,N_377,N_357);
xnor U9021 (N_9021,N_4693,N_3091);
and U9022 (N_9022,N_4560,N_651);
nor U9023 (N_9023,N_4487,N_1914);
nor U9024 (N_9024,N_3929,N_4220);
nor U9025 (N_9025,N_3397,N_1282);
and U9026 (N_9026,N_2256,N_3344);
nor U9027 (N_9027,N_3455,N_767);
nor U9028 (N_9028,N_4293,N_4246);
nand U9029 (N_9029,N_3800,N_4098);
and U9030 (N_9030,N_847,N_3481);
and U9031 (N_9031,N_148,N_2171);
or U9032 (N_9032,N_2011,N_3193);
and U9033 (N_9033,N_702,N_3530);
and U9034 (N_9034,N_4398,N_2329);
and U9035 (N_9035,N_3568,N_2103);
or U9036 (N_9036,N_150,N_2811);
or U9037 (N_9037,N_4623,N_1044);
and U9038 (N_9038,N_2065,N_505);
or U9039 (N_9039,N_1015,N_1310);
nor U9040 (N_9040,N_3635,N_4575);
nor U9041 (N_9041,N_1366,N_2386);
and U9042 (N_9042,N_2648,N_3958);
nand U9043 (N_9043,N_85,N_3139);
or U9044 (N_9044,N_527,N_4936);
nand U9045 (N_9045,N_934,N_4961);
xnor U9046 (N_9046,N_644,N_1279);
and U9047 (N_9047,N_158,N_2012);
xor U9048 (N_9048,N_4604,N_3920);
xor U9049 (N_9049,N_4412,N_2440);
nand U9050 (N_9050,N_2737,N_212);
and U9051 (N_9051,N_4709,N_2118);
or U9052 (N_9052,N_708,N_3372);
xnor U9053 (N_9053,N_2263,N_2624);
nor U9054 (N_9054,N_2195,N_3832);
xor U9055 (N_9055,N_3356,N_130);
and U9056 (N_9056,N_2021,N_1738);
or U9057 (N_9057,N_4251,N_2624);
nor U9058 (N_9058,N_2377,N_674);
or U9059 (N_9059,N_814,N_3294);
xor U9060 (N_9060,N_2586,N_1945);
or U9061 (N_9061,N_1027,N_2853);
and U9062 (N_9062,N_784,N_3794);
nand U9063 (N_9063,N_2964,N_4656);
and U9064 (N_9064,N_1731,N_4259);
and U9065 (N_9065,N_4994,N_1293);
nor U9066 (N_9066,N_903,N_4287);
nand U9067 (N_9067,N_1046,N_3927);
xor U9068 (N_9068,N_3656,N_3343);
nand U9069 (N_9069,N_1599,N_418);
nand U9070 (N_9070,N_1873,N_3261);
xnor U9071 (N_9071,N_3195,N_1781);
nor U9072 (N_9072,N_2827,N_3722);
xor U9073 (N_9073,N_1712,N_1758);
nor U9074 (N_9074,N_2777,N_3686);
nor U9075 (N_9075,N_3505,N_3401);
nor U9076 (N_9076,N_2087,N_292);
nor U9077 (N_9077,N_1128,N_2359);
and U9078 (N_9078,N_2533,N_3855);
nor U9079 (N_9079,N_2827,N_4312);
or U9080 (N_9080,N_562,N_917);
nor U9081 (N_9081,N_3516,N_1668);
nand U9082 (N_9082,N_3480,N_539);
nor U9083 (N_9083,N_1451,N_3230);
nor U9084 (N_9084,N_3233,N_4271);
or U9085 (N_9085,N_498,N_3304);
and U9086 (N_9086,N_3818,N_2120);
or U9087 (N_9087,N_3246,N_2889);
or U9088 (N_9088,N_3300,N_935);
nor U9089 (N_9089,N_4520,N_277);
or U9090 (N_9090,N_3281,N_3902);
or U9091 (N_9091,N_1652,N_1045);
nand U9092 (N_9092,N_726,N_3458);
and U9093 (N_9093,N_1829,N_4213);
or U9094 (N_9094,N_4972,N_339);
or U9095 (N_9095,N_49,N_4736);
or U9096 (N_9096,N_3720,N_1070);
nor U9097 (N_9097,N_3367,N_1749);
or U9098 (N_9098,N_4200,N_2224);
or U9099 (N_9099,N_868,N_1720);
or U9100 (N_9100,N_1862,N_1191);
xor U9101 (N_9101,N_4584,N_2645);
nor U9102 (N_9102,N_52,N_3037);
or U9103 (N_9103,N_3217,N_4088);
and U9104 (N_9104,N_4670,N_4992);
nor U9105 (N_9105,N_4062,N_3205);
xor U9106 (N_9106,N_551,N_3947);
and U9107 (N_9107,N_913,N_4334);
and U9108 (N_9108,N_317,N_3067);
nor U9109 (N_9109,N_2386,N_4064);
nor U9110 (N_9110,N_4268,N_3092);
or U9111 (N_9111,N_1392,N_3622);
xor U9112 (N_9112,N_793,N_4833);
and U9113 (N_9113,N_2584,N_3004);
nor U9114 (N_9114,N_3550,N_3014);
and U9115 (N_9115,N_2965,N_711);
xnor U9116 (N_9116,N_3631,N_1684);
nor U9117 (N_9117,N_4443,N_4471);
nand U9118 (N_9118,N_889,N_107);
nand U9119 (N_9119,N_4426,N_1034);
or U9120 (N_9120,N_3998,N_4099);
nor U9121 (N_9121,N_480,N_2613);
xnor U9122 (N_9122,N_2635,N_3518);
nand U9123 (N_9123,N_3865,N_2139);
xor U9124 (N_9124,N_433,N_2849);
xor U9125 (N_9125,N_4281,N_3435);
nor U9126 (N_9126,N_3699,N_4753);
or U9127 (N_9127,N_2773,N_2974);
nor U9128 (N_9128,N_464,N_3442);
nand U9129 (N_9129,N_4882,N_3205);
and U9130 (N_9130,N_739,N_4336);
or U9131 (N_9131,N_4541,N_150);
or U9132 (N_9132,N_4084,N_901);
and U9133 (N_9133,N_1010,N_285);
or U9134 (N_9134,N_4644,N_987);
or U9135 (N_9135,N_3787,N_3105);
nor U9136 (N_9136,N_935,N_3199);
or U9137 (N_9137,N_2589,N_2627);
and U9138 (N_9138,N_1093,N_476);
and U9139 (N_9139,N_850,N_4157);
and U9140 (N_9140,N_102,N_3864);
or U9141 (N_9141,N_2095,N_1515);
or U9142 (N_9142,N_4096,N_3183);
nand U9143 (N_9143,N_4417,N_199);
and U9144 (N_9144,N_529,N_4890);
and U9145 (N_9145,N_857,N_3414);
nand U9146 (N_9146,N_2728,N_4250);
nor U9147 (N_9147,N_1035,N_2005);
and U9148 (N_9148,N_1940,N_2703);
nand U9149 (N_9149,N_2816,N_2197);
nand U9150 (N_9150,N_4437,N_3631);
or U9151 (N_9151,N_1919,N_3273);
nor U9152 (N_9152,N_1547,N_2870);
nand U9153 (N_9153,N_1625,N_4499);
nor U9154 (N_9154,N_4191,N_3733);
nor U9155 (N_9155,N_2059,N_2722);
nand U9156 (N_9156,N_2468,N_3779);
and U9157 (N_9157,N_1032,N_2116);
xnor U9158 (N_9158,N_4527,N_2489);
nand U9159 (N_9159,N_1052,N_3369);
nor U9160 (N_9160,N_3609,N_838);
and U9161 (N_9161,N_3143,N_4961);
or U9162 (N_9162,N_3507,N_3911);
nor U9163 (N_9163,N_889,N_315);
nand U9164 (N_9164,N_621,N_3057);
xor U9165 (N_9165,N_4665,N_4086);
xnor U9166 (N_9166,N_2548,N_570);
or U9167 (N_9167,N_747,N_3131);
and U9168 (N_9168,N_4478,N_2700);
xor U9169 (N_9169,N_4568,N_119);
nand U9170 (N_9170,N_590,N_3252);
and U9171 (N_9171,N_2303,N_670);
or U9172 (N_9172,N_4723,N_1689);
or U9173 (N_9173,N_4016,N_4557);
nor U9174 (N_9174,N_2079,N_321);
nor U9175 (N_9175,N_2683,N_3815);
and U9176 (N_9176,N_653,N_4103);
or U9177 (N_9177,N_4317,N_1570);
or U9178 (N_9178,N_3840,N_2600);
nand U9179 (N_9179,N_3798,N_3278);
or U9180 (N_9180,N_1306,N_3610);
and U9181 (N_9181,N_1669,N_4813);
or U9182 (N_9182,N_2593,N_1330);
nand U9183 (N_9183,N_1979,N_61);
nor U9184 (N_9184,N_287,N_613);
nand U9185 (N_9185,N_4925,N_4649);
nand U9186 (N_9186,N_3247,N_3359);
nor U9187 (N_9187,N_3096,N_3900);
or U9188 (N_9188,N_2658,N_199);
nor U9189 (N_9189,N_646,N_3741);
nand U9190 (N_9190,N_1849,N_2653);
nor U9191 (N_9191,N_3290,N_523);
xor U9192 (N_9192,N_4787,N_1055);
nor U9193 (N_9193,N_522,N_3442);
nand U9194 (N_9194,N_2010,N_792);
or U9195 (N_9195,N_3221,N_814);
xor U9196 (N_9196,N_3902,N_2006);
nand U9197 (N_9197,N_55,N_2073);
nor U9198 (N_9198,N_1584,N_4594);
and U9199 (N_9199,N_3259,N_2823);
or U9200 (N_9200,N_2331,N_382);
and U9201 (N_9201,N_1896,N_284);
and U9202 (N_9202,N_1934,N_1647);
and U9203 (N_9203,N_3657,N_1289);
nor U9204 (N_9204,N_1622,N_4507);
or U9205 (N_9205,N_721,N_4346);
or U9206 (N_9206,N_2826,N_2192);
xor U9207 (N_9207,N_617,N_761);
nor U9208 (N_9208,N_1033,N_4923);
and U9209 (N_9209,N_4604,N_2175);
nand U9210 (N_9210,N_2659,N_4663);
or U9211 (N_9211,N_1801,N_2660);
and U9212 (N_9212,N_34,N_1201);
or U9213 (N_9213,N_4613,N_1960);
nor U9214 (N_9214,N_4460,N_1224);
xnor U9215 (N_9215,N_3420,N_4573);
nor U9216 (N_9216,N_3607,N_4321);
nor U9217 (N_9217,N_1724,N_362);
and U9218 (N_9218,N_4262,N_3020);
and U9219 (N_9219,N_3307,N_4467);
or U9220 (N_9220,N_2592,N_4814);
or U9221 (N_9221,N_4458,N_4387);
nand U9222 (N_9222,N_175,N_2112);
or U9223 (N_9223,N_987,N_2550);
xnor U9224 (N_9224,N_3755,N_609);
or U9225 (N_9225,N_2858,N_4293);
or U9226 (N_9226,N_114,N_1984);
nor U9227 (N_9227,N_1502,N_4552);
xnor U9228 (N_9228,N_961,N_3455);
and U9229 (N_9229,N_3765,N_284);
nor U9230 (N_9230,N_2261,N_4389);
nor U9231 (N_9231,N_4034,N_2169);
nand U9232 (N_9232,N_2945,N_160);
nand U9233 (N_9233,N_1586,N_2400);
nand U9234 (N_9234,N_3851,N_499);
nand U9235 (N_9235,N_2109,N_4965);
nor U9236 (N_9236,N_904,N_2704);
or U9237 (N_9237,N_1562,N_2376);
nand U9238 (N_9238,N_4275,N_2506);
nor U9239 (N_9239,N_1557,N_3371);
nor U9240 (N_9240,N_2514,N_1614);
xor U9241 (N_9241,N_3066,N_1355);
nand U9242 (N_9242,N_2755,N_1714);
nand U9243 (N_9243,N_4242,N_3056);
or U9244 (N_9244,N_3573,N_4972);
and U9245 (N_9245,N_2634,N_541);
xnor U9246 (N_9246,N_408,N_3382);
or U9247 (N_9247,N_2344,N_4920);
and U9248 (N_9248,N_1287,N_4381);
nand U9249 (N_9249,N_2311,N_2983);
nor U9250 (N_9250,N_2965,N_943);
and U9251 (N_9251,N_563,N_1927);
or U9252 (N_9252,N_1860,N_2687);
nand U9253 (N_9253,N_3399,N_4442);
nand U9254 (N_9254,N_4975,N_4049);
or U9255 (N_9255,N_686,N_432);
or U9256 (N_9256,N_3480,N_2244);
or U9257 (N_9257,N_2757,N_3623);
nand U9258 (N_9258,N_4434,N_4564);
nand U9259 (N_9259,N_1943,N_346);
or U9260 (N_9260,N_3566,N_3003);
nand U9261 (N_9261,N_3762,N_4560);
nor U9262 (N_9262,N_2838,N_1215);
xnor U9263 (N_9263,N_1271,N_392);
or U9264 (N_9264,N_671,N_4311);
or U9265 (N_9265,N_3986,N_2517);
and U9266 (N_9266,N_4731,N_4901);
or U9267 (N_9267,N_1119,N_1478);
and U9268 (N_9268,N_4218,N_944);
nand U9269 (N_9269,N_3615,N_3035);
nand U9270 (N_9270,N_4891,N_1322);
nor U9271 (N_9271,N_4924,N_1985);
xor U9272 (N_9272,N_746,N_3979);
nand U9273 (N_9273,N_2507,N_1823);
nor U9274 (N_9274,N_3531,N_4370);
or U9275 (N_9275,N_2843,N_2200);
nand U9276 (N_9276,N_4710,N_781);
and U9277 (N_9277,N_1940,N_2107);
or U9278 (N_9278,N_912,N_1318);
nor U9279 (N_9279,N_2314,N_543);
nand U9280 (N_9280,N_4317,N_4213);
nand U9281 (N_9281,N_697,N_1553);
nand U9282 (N_9282,N_3219,N_784);
and U9283 (N_9283,N_3659,N_3937);
or U9284 (N_9284,N_2878,N_1157);
nand U9285 (N_9285,N_3612,N_4694);
and U9286 (N_9286,N_3872,N_1556);
xor U9287 (N_9287,N_4733,N_36);
and U9288 (N_9288,N_3482,N_3071);
and U9289 (N_9289,N_3448,N_2760);
nand U9290 (N_9290,N_514,N_3256);
nor U9291 (N_9291,N_3201,N_4317);
xnor U9292 (N_9292,N_779,N_4537);
nand U9293 (N_9293,N_2839,N_3780);
nor U9294 (N_9294,N_1531,N_4085);
nand U9295 (N_9295,N_4592,N_3455);
xor U9296 (N_9296,N_472,N_572);
xor U9297 (N_9297,N_2916,N_73);
or U9298 (N_9298,N_4993,N_1068);
or U9299 (N_9299,N_4808,N_558);
and U9300 (N_9300,N_2743,N_3805);
and U9301 (N_9301,N_2024,N_56);
xor U9302 (N_9302,N_3196,N_2150);
or U9303 (N_9303,N_38,N_656);
or U9304 (N_9304,N_4006,N_1563);
nor U9305 (N_9305,N_4362,N_1626);
or U9306 (N_9306,N_2353,N_2913);
xor U9307 (N_9307,N_1421,N_555);
nor U9308 (N_9308,N_3909,N_4089);
nor U9309 (N_9309,N_2357,N_582);
xor U9310 (N_9310,N_17,N_2394);
nand U9311 (N_9311,N_4197,N_323);
nand U9312 (N_9312,N_4737,N_4831);
or U9313 (N_9313,N_3762,N_2033);
or U9314 (N_9314,N_1769,N_1815);
nand U9315 (N_9315,N_3674,N_1539);
and U9316 (N_9316,N_1607,N_4963);
or U9317 (N_9317,N_865,N_1509);
xnor U9318 (N_9318,N_1269,N_2093);
nand U9319 (N_9319,N_3219,N_3767);
nand U9320 (N_9320,N_4094,N_4211);
and U9321 (N_9321,N_4987,N_1654);
nor U9322 (N_9322,N_3926,N_1136);
nor U9323 (N_9323,N_1082,N_2994);
and U9324 (N_9324,N_744,N_4528);
and U9325 (N_9325,N_1848,N_2079);
and U9326 (N_9326,N_893,N_2294);
nor U9327 (N_9327,N_143,N_1961);
nor U9328 (N_9328,N_2736,N_401);
nor U9329 (N_9329,N_2704,N_684);
nor U9330 (N_9330,N_3031,N_1960);
or U9331 (N_9331,N_3697,N_985);
nor U9332 (N_9332,N_2722,N_1560);
and U9333 (N_9333,N_808,N_563);
nand U9334 (N_9334,N_3024,N_3248);
or U9335 (N_9335,N_4826,N_936);
and U9336 (N_9336,N_448,N_4862);
or U9337 (N_9337,N_3332,N_4064);
nand U9338 (N_9338,N_3730,N_3841);
xnor U9339 (N_9339,N_4294,N_3820);
nand U9340 (N_9340,N_493,N_2895);
xor U9341 (N_9341,N_2111,N_4473);
nor U9342 (N_9342,N_3597,N_3974);
nand U9343 (N_9343,N_1250,N_3795);
nand U9344 (N_9344,N_3939,N_2730);
or U9345 (N_9345,N_455,N_4068);
nand U9346 (N_9346,N_3706,N_3896);
nor U9347 (N_9347,N_1544,N_3663);
and U9348 (N_9348,N_1490,N_4836);
or U9349 (N_9349,N_4743,N_2086);
or U9350 (N_9350,N_4977,N_759);
and U9351 (N_9351,N_3548,N_4511);
xnor U9352 (N_9352,N_595,N_110);
and U9353 (N_9353,N_4649,N_3719);
and U9354 (N_9354,N_4981,N_4872);
and U9355 (N_9355,N_4828,N_1847);
nor U9356 (N_9356,N_3008,N_4152);
or U9357 (N_9357,N_48,N_1759);
nand U9358 (N_9358,N_1246,N_1095);
xnor U9359 (N_9359,N_1935,N_4873);
and U9360 (N_9360,N_4153,N_4834);
nor U9361 (N_9361,N_3142,N_3419);
nor U9362 (N_9362,N_4224,N_2345);
nor U9363 (N_9363,N_3500,N_4727);
or U9364 (N_9364,N_264,N_1966);
xnor U9365 (N_9365,N_3443,N_3525);
and U9366 (N_9366,N_320,N_1498);
nor U9367 (N_9367,N_1152,N_4189);
xnor U9368 (N_9368,N_44,N_2292);
nand U9369 (N_9369,N_2096,N_3379);
and U9370 (N_9370,N_4610,N_795);
nor U9371 (N_9371,N_3877,N_3917);
or U9372 (N_9372,N_4689,N_3872);
nor U9373 (N_9373,N_4680,N_2972);
xnor U9374 (N_9374,N_742,N_721);
nor U9375 (N_9375,N_1848,N_2594);
nand U9376 (N_9376,N_2878,N_2448);
and U9377 (N_9377,N_2819,N_1573);
and U9378 (N_9378,N_773,N_181);
and U9379 (N_9379,N_1239,N_4671);
and U9380 (N_9380,N_456,N_4365);
nand U9381 (N_9381,N_4857,N_2754);
nand U9382 (N_9382,N_4814,N_4378);
nand U9383 (N_9383,N_1530,N_1143);
nor U9384 (N_9384,N_4766,N_3070);
and U9385 (N_9385,N_3356,N_2044);
or U9386 (N_9386,N_2533,N_3051);
xor U9387 (N_9387,N_620,N_1890);
nand U9388 (N_9388,N_2001,N_3574);
nand U9389 (N_9389,N_3374,N_3640);
nor U9390 (N_9390,N_786,N_4592);
and U9391 (N_9391,N_1960,N_1191);
and U9392 (N_9392,N_4060,N_3309);
or U9393 (N_9393,N_4329,N_2010);
and U9394 (N_9394,N_702,N_4263);
and U9395 (N_9395,N_1968,N_3584);
nor U9396 (N_9396,N_4751,N_1864);
or U9397 (N_9397,N_2976,N_1564);
nand U9398 (N_9398,N_178,N_256);
or U9399 (N_9399,N_4391,N_1228);
and U9400 (N_9400,N_4949,N_3018);
nand U9401 (N_9401,N_567,N_4041);
xnor U9402 (N_9402,N_1022,N_3018);
nand U9403 (N_9403,N_4718,N_828);
xor U9404 (N_9404,N_1733,N_1090);
nand U9405 (N_9405,N_3023,N_1226);
and U9406 (N_9406,N_4058,N_2704);
nor U9407 (N_9407,N_1578,N_3536);
or U9408 (N_9408,N_4735,N_2010);
xnor U9409 (N_9409,N_2503,N_1094);
and U9410 (N_9410,N_4046,N_2947);
xnor U9411 (N_9411,N_2379,N_3706);
nor U9412 (N_9412,N_371,N_3233);
xnor U9413 (N_9413,N_2590,N_3216);
or U9414 (N_9414,N_586,N_3347);
nand U9415 (N_9415,N_3426,N_2073);
or U9416 (N_9416,N_1116,N_1948);
and U9417 (N_9417,N_4599,N_2420);
and U9418 (N_9418,N_626,N_3648);
nor U9419 (N_9419,N_158,N_670);
and U9420 (N_9420,N_3949,N_837);
nand U9421 (N_9421,N_2795,N_2589);
nor U9422 (N_9422,N_3275,N_3304);
and U9423 (N_9423,N_37,N_241);
xnor U9424 (N_9424,N_4515,N_1253);
or U9425 (N_9425,N_3808,N_981);
or U9426 (N_9426,N_2690,N_3327);
nand U9427 (N_9427,N_802,N_2998);
and U9428 (N_9428,N_455,N_1440);
or U9429 (N_9429,N_4946,N_245);
or U9430 (N_9430,N_876,N_1051);
nand U9431 (N_9431,N_3762,N_1356);
nand U9432 (N_9432,N_3137,N_3711);
and U9433 (N_9433,N_3412,N_17);
nor U9434 (N_9434,N_796,N_987);
or U9435 (N_9435,N_3007,N_2199);
nor U9436 (N_9436,N_3180,N_764);
xor U9437 (N_9437,N_467,N_1459);
xnor U9438 (N_9438,N_4053,N_3099);
or U9439 (N_9439,N_4281,N_2546);
or U9440 (N_9440,N_1469,N_4480);
and U9441 (N_9441,N_4320,N_4952);
nor U9442 (N_9442,N_2304,N_1284);
and U9443 (N_9443,N_2980,N_2243);
or U9444 (N_9444,N_2717,N_938);
nand U9445 (N_9445,N_1226,N_1779);
or U9446 (N_9446,N_4560,N_1281);
nand U9447 (N_9447,N_3287,N_238);
nor U9448 (N_9448,N_1529,N_4556);
and U9449 (N_9449,N_93,N_2510);
or U9450 (N_9450,N_1575,N_754);
and U9451 (N_9451,N_598,N_2338);
nor U9452 (N_9452,N_4217,N_3361);
and U9453 (N_9453,N_4461,N_2390);
or U9454 (N_9454,N_1233,N_3115);
and U9455 (N_9455,N_572,N_155);
or U9456 (N_9456,N_1288,N_329);
nor U9457 (N_9457,N_307,N_2357);
nor U9458 (N_9458,N_1252,N_2461);
or U9459 (N_9459,N_1752,N_4628);
and U9460 (N_9460,N_130,N_4399);
nand U9461 (N_9461,N_3630,N_82);
nand U9462 (N_9462,N_1447,N_798);
xor U9463 (N_9463,N_1373,N_2232);
xor U9464 (N_9464,N_1603,N_4234);
nor U9465 (N_9465,N_3571,N_635);
nand U9466 (N_9466,N_4069,N_4099);
or U9467 (N_9467,N_4525,N_4018);
nand U9468 (N_9468,N_312,N_1384);
nor U9469 (N_9469,N_2294,N_2905);
and U9470 (N_9470,N_3048,N_2846);
and U9471 (N_9471,N_4898,N_2286);
or U9472 (N_9472,N_1652,N_4013);
or U9473 (N_9473,N_2010,N_77);
or U9474 (N_9474,N_2300,N_2784);
nor U9475 (N_9475,N_1880,N_845);
nor U9476 (N_9476,N_1739,N_1744);
nand U9477 (N_9477,N_1375,N_949);
nand U9478 (N_9478,N_978,N_827);
nor U9479 (N_9479,N_848,N_2153);
or U9480 (N_9480,N_1943,N_147);
nand U9481 (N_9481,N_237,N_2610);
or U9482 (N_9482,N_2036,N_2728);
xor U9483 (N_9483,N_2702,N_3107);
or U9484 (N_9484,N_2331,N_4749);
nor U9485 (N_9485,N_2173,N_4798);
nand U9486 (N_9486,N_816,N_1121);
and U9487 (N_9487,N_3127,N_912);
and U9488 (N_9488,N_812,N_2868);
or U9489 (N_9489,N_4942,N_4438);
nand U9490 (N_9490,N_1867,N_4270);
or U9491 (N_9491,N_1564,N_3449);
nand U9492 (N_9492,N_1195,N_1574);
and U9493 (N_9493,N_3686,N_4205);
nand U9494 (N_9494,N_2761,N_3512);
nor U9495 (N_9495,N_571,N_4699);
xnor U9496 (N_9496,N_3857,N_4480);
or U9497 (N_9497,N_705,N_4244);
nand U9498 (N_9498,N_2464,N_2355);
or U9499 (N_9499,N_2288,N_4162);
nor U9500 (N_9500,N_1825,N_413);
nor U9501 (N_9501,N_2206,N_661);
nor U9502 (N_9502,N_699,N_3835);
and U9503 (N_9503,N_4056,N_1653);
or U9504 (N_9504,N_2879,N_1096);
nand U9505 (N_9505,N_1507,N_4217);
and U9506 (N_9506,N_91,N_4076);
xnor U9507 (N_9507,N_3312,N_3294);
xor U9508 (N_9508,N_1657,N_640);
nand U9509 (N_9509,N_4806,N_779);
and U9510 (N_9510,N_586,N_3816);
and U9511 (N_9511,N_4053,N_3990);
nor U9512 (N_9512,N_1655,N_2312);
nand U9513 (N_9513,N_486,N_610);
nand U9514 (N_9514,N_1253,N_4128);
and U9515 (N_9515,N_2098,N_2090);
nor U9516 (N_9516,N_1076,N_4468);
nand U9517 (N_9517,N_610,N_2926);
xnor U9518 (N_9518,N_73,N_4319);
or U9519 (N_9519,N_2780,N_4507);
and U9520 (N_9520,N_374,N_52);
nand U9521 (N_9521,N_2139,N_4740);
or U9522 (N_9522,N_3729,N_3152);
nor U9523 (N_9523,N_3030,N_2843);
nor U9524 (N_9524,N_1191,N_2199);
or U9525 (N_9525,N_1565,N_803);
xnor U9526 (N_9526,N_614,N_517);
or U9527 (N_9527,N_4240,N_4986);
nor U9528 (N_9528,N_2603,N_868);
and U9529 (N_9529,N_60,N_1273);
and U9530 (N_9530,N_4809,N_4710);
and U9531 (N_9531,N_439,N_1868);
or U9532 (N_9532,N_2913,N_4076);
and U9533 (N_9533,N_935,N_849);
or U9534 (N_9534,N_1903,N_924);
nand U9535 (N_9535,N_2211,N_2565);
nand U9536 (N_9536,N_2,N_16);
nor U9537 (N_9537,N_1912,N_3182);
and U9538 (N_9538,N_1177,N_1110);
nor U9539 (N_9539,N_475,N_196);
and U9540 (N_9540,N_2126,N_4374);
nor U9541 (N_9541,N_1591,N_4017);
nor U9542 (N_9542,N_1341,N_1731);
and U9543 (N_9543,N_2265,N_3883);
and U9544 (N_9544,N_4438,N_2137);
nor U9545 (N_9545,N_926,N_4331);
nor U9546 (N_9546,N_3840,N_1322);
nand U9547 (N_9547,N_2099,N_4063);
nor U9548 (N_9548,N_2361,N_2890);
and U9549 (N_9549,N_3767,N_2082);
and U9550 (N_9550,N_2893,N_4868);
xor U9551 (N_9551,N_1686,N_2785);
and U9552 (N_9552,N_1660,N_4868);
or U9553 (N_9553,N_3266,N_4717);
or U9554 (N_9554,N_2499,N_3331);
or U9555 (N_9555,N_4391,N_2608);
and U9556 (N_9556,N_1476,N_534);
or U9557 (N_9557,N_684,N_3282);
nand U9558 (N_9558,N_3894,N_2447);
and U9559 (N_9559,N_4856,N_1503);
nor U9560 (N_9560,N_3424,N_1755);
nor U9561 (N_9561,N_4142,N_2632);
and U9562 (N_9562,N_475,N_264);
nand U9563 (N_9563,N_4600,N_185);
nor U9564 (N_9564,N_3719,N_2237);
nor U9565 (N_9565,N_1451,N_1639);
or U9566 (N_9566,N_3499,N_1990);
nor U9567 (N_9567,N_2868,N_2672);
nand U9568 (N_9568,N_1801,N_2760);
nand U9569 (N_9569,N_3872,N_3065);
nand U9570 (N_9570,N_3114,N_2216);
or U9571 (N_9571,N_2113,N_3782);
and U9572 (N_9572,N_448,N_4792);
nor U9573 (N_9573,N_3900,N_2650);
xnor U9574 (N_9574,N_3713,N_4890);
and U9575 (N_9575,N_2176,N_1881);
or U9576 (N_9576,N_3643,N_4408);
nor U9577 (N_9577,N_2486,N_3107);
nor U9578 (N_9578,N_581,N_2731);
or U9579 (N_9579,N_475,N_4803);
xnor U9580 (N_9580,N_351,N_2479);
or U9581 (N_9581,N_930,N_3039);
or U9582 (N_9582,N_1907,N_1193);
nor U9583 (N_9583,N_2606,N_2061);
xor U9584 (N_9584,N_391,N_472);
xor U9585 (N_9585,N_773,N_4296);
nor U9586 (N_9586,N_3016,N_1166);
xnor U9587 (N_9587,N_2192,N_810);
or U9588 (N_9588,N_1176,N_3771);
or U9589 (N_9589,N_1468,N_673);
or U9590 (N_9590,N_3917,N_351);
nor U9591 (N_9591,N_3953,N_2616);
or U9592 (N_9592,N_4727,N_4855);
xnor U9593 (N_9593,N_2444,N_4201);
nand U9594 (N_9594,N_2701,N_3414);
nor U9595 (N_9595,N_1803,N_3178);
and U9596 (N_9596,N_3298,N_4556);
xnor U9597 (N_9597,N_4748,N_2179);
and U9598 (N_9598,N_3479,N_149);
nor U9599 (N_9599,N_3567,N_2722);
and U9600 (N_9600,N_1991,N_4294);
or U9601 (N_9601,N_2261,N_3464);
and U9602 (N_9602,N_870,N_3274);
or U9603 (N_9603,N_1296,N_4288);
and U9604 (N_9604,N_3237,N_528);
and U9605 (N_9605,N_4885,N_4804);
and U9606 (N_9606,N_3182,N_2762);
and U9607 (N_9607,N_1788,N_700);
or U9608 (N_9608,N_458,N_2715);
or U9609 (N_9609,N_2775,N_2836);
nand U9610 (N_9610,N_2020,N_3521);
xor U9611 (N_9611,N_3551,N_2705);
nor U9612 (N_9612,N_2327,N_4001);
nor U9613 (N_9613,N_2041,N_3460);
and U9614 (N_9614,N_1182,N_1664);
nor U9615 (N_9615,N_2481,N_4625);
nor U9616 (N_9616,N_54,N_2418);
or U9617 (N_9617,N_325,N_4723);
nor U9618 (N_9618,N_2914,N_1310);
nand U9619 (N_9619,N_2413,N_4831);
and U9620 (N_9620,N_2540,N_2599);
or U9621 (N_9621,N_2557,N_3024);
and U9622 (N_9622,N_4134,N_4376);
nand U9623 (N_9623,N_3484,N_394);
and U9624 (N_9624,N_3756,N_451);
nand U9625 (N_9625,N_4317,N_2528);
nand U9626 (N_9626,N_2518,N_2864);
xnor U9627 (N_9627,N_328,N_2431);
nand U9628 (N_9628,N_4723,N_3926);
and U9629 (N_9629,N_1534,N_4023);
or U9630 (N_9630,N_4191,N_2182);
xor U9631 (N_9631,N_1213,N_4040);
nand U9632 (N_9632,N_1718,N_3276);
and U9633 (N_9633,N_108,N_4520);
nor U9634 (N_9634,N_2924,N_1811);
nor U9635 (N_9635,N_1504,N_285);
nand U9636 (N_9636,N_4115,N_2274);
or U9637 (N_9637,N_4800,N_231);
and U9638 (N_9638,N_3082,N_1267);
and U9639 (N_9639,N_3467,N_3474);
nand U9640 (N_9640,N_3983,N_2253);
or U9641 (N_9641,N_1729,N_2594);
or U9642 (N_9642,N_4643,N_216);
nor U9643 (N_9643,N_317,N_276);
and U9644 (N_9644,N_799,N_340);
and U9645 (N_9645,N_1150,N_4931);
nand U9646 (N_9646,N_3833,N_1117);
xnor U9647 (N_9647,N_4513,N_2204);
or U9648 (N_9648,N_3165,N_1064);
and U9649 (N_9649,N_1085,N_731);
and U9650 (N_9650,N_4418,N_1948);
nand U9651 (N_9651,N_2953,N_538);
and U9652 (N_9652,N_1535,N_1878);
and U9653 (N_9653,N_2802,N_3739);
or U9654 (N_9654,N_2649,N_508);
xor U9655 (N_9655,N_3544,N_2111);
nor U9656 (N_9656,N_3081,N_210);
or U9657 (N_9657,N_3991,N_2765);
or U9658 (N_9658,N_2632,N_2450);
nor U9659 (N_9659,N_3209,N_2458);
nand U9660 (N_9660,N_880,N_4519);
and U9661 (N_9661,N_351,N_15);
or U9662 (N_9662,N_3027,N_3032);
and U9663 (N_9663,N_4847,N_806);
or U9664 (N_9664,N_2919,N_381);
nand U9665 (N_9665,N_4845,N_4530);
and U9666 (N_9666,N_1511,N_4895);
nand U9667 (N_9667,N_1137,N_893);
nand U9668 (N_9668,N_2824,N_2375);
and U9669 (N_9669,N_170,N_2000);
nor U9670 (N_9670,N_2226,N_3608);
and U9671 (N_9671,N_649,N_4220);
nor U9672 (N_9672,N_2198,N_3218);
nand U9673 (N_9673,N_3375,N_1747);
nand U9674 (N_9674,N_2135,N_1040);
nand U9675 (N_9675,N_3965,N_1877);
xor U9676 (N_9676,N_1760,N_4625);
xnor U9677 (N_9677,N_434,N_3513);
xnor U9678 (N_9678,N_1530,N_3994);
nand U9679 (N_9679,N_3736,N_1314);
or U9680 (N_9680,N_1025,N_2430);
or U9681 (N_9681,N_805,N_3943);
nand U9682 (N_9682,N_3243,N_3641);
nor U9683 (N_9683,N_1306,N_3872);
xnor U9684 (N_9684,N_1206,N_2264);
xor U9685 (N_9685,N_2184,N_4354);
xnor U9686 (N_9686,N_3372,N_2798);
nor U9687 (N_9687,N_458,N_4191);
nand U9688 (N_9688,N_1422,N_643);
or U9689 (N_9689,N_4696,N_1868);
nand U9690 (N_9690,N_1121,N_2352);
and U9691 (N_9691,N_1996,N_161);
nor U9692 (N_9692,N_927,N_1596);
xnor U9693 (N_9693,N_152,N_3264);
and U9694 (N_9694,N_1039,N_3246);
nand U9695 (N_9695,N_757,N_4946);
nor U9696 (N_9696,N_984,N_4395);
or U9697 (N_9697,N_4399,N_1786);
nand U9698 (N_9698,N_1760,N_3001);
nor U9699 (N_9699,N_3943,N_4282);
nand U9700 (N_9700,N_2490,N_533);
or U9701 (N_9701,N_3054,N_4128);
xor U9702 (N_9702,N_3014,N_2131);
xnor U9703 (N_9703,N_4867,N_1602);
or U9704 (N_9704,N_2893,N_1308);
xor U9705 (N_9705,N_432,N_4915);
or U9706 (N_9706,N_2901,N_376);
and U9707 (N_9707,N_4109,N_4691);
or U9708 (N_9708,N_2912,N_3846);
and U9709 (N_9709,N_26,N_3445);
or U9710 (N_9710,N_653,N_2310);
and U9711 (N_9711,N_4988,N_481);
xor U9712 (N_9712,N_3334,N_1444);
nor U9713 (N_9713,N_136,N_2339);
nand U9714 (N_9714,N_4023,N_4632);
xnor U9715 (N_9715,N_784,N_4397);
or U9716 (N_9716,N_3745,N_4802);
nand U9717 (N_9717,N_4989,N_3017);
nand U9718 (N_9718,N_1960,N_1096);
nor U9719 (N_9719,N_1778,N_150);
or U9720 (N_9720,N_645,N_4707);
xor U9721 (N_9721,N_2508,N_1220);
nand U9722 (N_9722,N_3921,N_3140);
and U9723 (N_9723,N_1936,N_4536);
nand U9724 (N_9724,N_2289,N_1007);
or U9725 (N_9725,N_3148,N_4625);
or U9726 (N_9726,N_2993,N_4588);
nor U9727 (N_9727,N_2111,N_2426);
and U9728 (N_9728,N_1992,N_4014);
nor U9729 (N_9729,N_1934,N_1672);
or U9730 (N_9730,N_3511,N_1868);
xor U9731 (N_9731,N_1013,N_2666);
nor U9732 (N_9732,N_1773,N_437);
nor U9733 (N_9733,N_4972,N_2896);
and U9734 (N_9734,N_4075,N_1261);
and U9735 (N_9735,N_502,N_3193);
nand U9736 (N_9736,N_2356,N_1542);
and U9737 (N_9737,N_1884,N_256);
nand U9738 (N_9738,N_1963,N_3888);
or U9739 (N_9739,N_1988,N_1174);
nor U9740 (N_9740,N_3331,N_1638);
and U9741 (N_9741,N_4613,N_3872);
or U9742 (N_9742,N_2193,N_164);
nand U9743 (N_9743,N_4211,N_1474);
xnor U9744 (N_9744,N_333,N_4395);
or U9745 (N_9745,N_2691,N_142);
nor U9746 (N_9746,N_4485,N_1394);
nand U9747 (N_9747,N_130,N_614);
and U9748 (N_9748,N_4344,N_1713);
nand U9749 (N_9749,N_3552,N_4302);
or U9750 (N_9750,N_4095,N_887);
nand U9751 (N_9751,N_1372,N_3239);
or U9752 (N_9752,N_3791,N_858);
nand U9753 (N_9753,N_3165,N_2064);
nand U9754 (N_9754,N_2690,N_1066);
xnor U9755 (N_9755,N_4185,N_527);
nor U9756 (N_9756,N_3393,N_3389);
and U9757 (N_9757,N_2974,N_3565);
and U9758 (N_9758,N_347,N_2859);
nor U9759 (N_9759,N_909,N_4485);
or U9760 (N_9760,N_4730,N_336);
and U9761 (N_9761,N_96,N_4251);
xnor U9762 (N_9762,N_1340,N_123);
nor U9763 (N_9763,N_1692,N_3023);
and U9764 (N_9764,N_3825,N_522);
xor U9765 (N_9765,N_4741,N_3721);
nor U9766 (N_9766,N_3958,N_1015);
and U9767 (N_9767,N_4412,N_2961);
and U9768 (N_9768,N_2671,N_4089);
nor U9769 (N_9769,N_2163,N_3922);
or U9770 (N_9770,N_1740,N_2908);
xnor U9771 (N_9771,N_2495,N_4630);
xor U9772 (N_9772,N_1827,N_2330);
or U9773 (N_9773,N_1066,N_1440);
and U9774 (N_9774,N_1516,N_1881);
or U9775 (N_9775,N_254,N_3369);
or U9776 (N_9776,N_2132,N_2196);
or U9777 (N_9777,N_3505,N_2781);
nor U9778 (N_9778,N_4376,N_2684);
nor U9779 (N_9779,N_1099,N_1096);
nand U9780 (N_9780,N_3284,N_3905);
or U9781 (N_9781,N_189,N_1563);
or U9782 (N_9782,N_1729,N_176);
or U9783 (N_9783,N_4908,N_2255);
and U9784 (N_9784,N_2320,N_4572);
nand U9785 (N_9785,N_4581,N_4141);
or U9786 (N_9786,N_440,N_2641);
nor U9787 (N_9787,N_4974,N_774);
nor U9788 (N_9788,N_2457,N_1893);
nor U9789 (N_9789,N_2712,N_1953);
nand U9790 (N_9790,N_3008,N_849);
nor U9791 (N_9791,N_303,N_1175);
nor U9792 (N_9792,N_3606,N_1608);
or U9793 (N_9793,N_1882,N_2268);
nor U9794 (N_9794,N_986,N_975);
nand U9795 (N_9795,N_748,N_2500);
nand U9796 (N_9796,N_4983,N_784);
nand U9797 (N_9797,N_1417,N_2639);
nor U9798 (N_9798,N_3169,N_4093);
nor U9799 (N_9799,N_2752,N_2906);
and U9800 (N_9800,N_4764,N_4027);
xnor U9801 (N_9801,N_2804,N_2492);
nand U9802 (N_9802,N_2572,N_4150);
and U9803 (N_9803,N_2920,N_3082);
and U9804 (N_9804,N_1346,N_129);
nor U9805 (N_9805,N_2282,N_371);
nand U9806 (N_9806,N_275,N_513);
or U9807 (N_9807,N_3308,N_1918);
nand U9808 (N_9808,N_4160,N_2236);
xnor U9809 (N_9809,N_1296,N_2201);
nand U9810 (N_9810,N_1403,N_3143);
or U9811 (N_9811,N_100,N_2978);
or U9812 (N_9812,N_4440,N_1745);
or U9813 (N_9813,N_3283,N_1916);
and U9814 (N_9814,N_222,N_4104);
nand U9815 (N_9815,N_1726,N_4404);
nor U9816 (N_9816,N_3285,N_2004);
nor U9817 (N_9817,N_4030,N_2202);
nor U9818 (N_9818,N_3621,N_4747);
nor U9819 (N_9819,N_954,N_4227);
nor U9820 (N_9820,N_4038,N_1046);
xor U9821 (N_9821,N_162,N_2140);
and U9822 (N_9822,N_4734,N_2989);
or U9823 (N_9823,N_177,N_2218);
and U9824 (N_9824,N_2594,N_1078);
nand U9825 (N_9825,N_2619,N_2694);
and U9826 (N_9826,N_374,N_3998);
or U9827 (N_9827,N_2265,N_167);
or U9828 (N_9828,N_3591,N_1452);
nor U9829 (N_9829,N_2286,N_726);
or U9830 (N_9830,N_1955,N_4669);
nor U9831 (N_9831,N_2717,N_51);
nand U9832 (N_9832,N_2873,N_3792);
and U9833 (N_9833,N_284,N_3815);
xnor U9834 (N_9834,N_1458,N_1422);
nor U9835 (N_9835,N_1839,N_2165);
and U9836 (N_9836,N_3782,N_3813);
xor U9837 (N_9837,N_3907,N_3381);
nand U9838 (N_9838,N_275,N_521);
xor U9839 (N_9839,N_1339,N_2889);
and U9840 (N_9840,N_4338,N_932);
or U9841 (N_9841,N_960,N_4532);
and U9842 (N_9842,N_4047,N_469);
nand U9843 (N_9843,N_2802,N_3019);
xor U9844 (N_9844,N_1939,N_38);
and U9845 (N_9845,N_3612,N_2185);
or U9846 (N_9846,N_1724,N_916);
nor U9847 (N_9847,N_4712,N_13);
and U9848 (N_9848,N_4078,N_1514);
nand U9849 (N_9849,N_2182,N_4777);
and U9850 (N_9850,N_2801,N_4262);
and U9851 (N_9851,N_1756,N_803);
nand U9852 (N_9852,N_4511,N_3133);
or U9853 (N_9853,N_4594,N_2469);
nand U9854 (N_9854,N_4289,N_4098);
xor U9855 (N_9855,N_3467,N_2979);
nor U9856 (N_9856,N_4305,N_498);
nand U9857 (N_9857,N_492,N_283);
or U9858 (N_9858,N_2970,N_4708);
nand U9859 (N_9859,N_3218,N_1750);
nand U9860 (N_9860,N_664,N_3262);
and U9861 (N_9861,N_1031,N_2484);
or U9862 (N_9862,N_2072,N_4321);
nand U9863 (N_9863,N_578,N_4996);
and U9864 (N_9864,N_4738,N_1975);
nand U9865 (N_9865,N_3141,N_2760);
nor U9866 (N_9866,N_4876,N_4500);
and U9867 (N_9867,N_4044,N_3145);
and U9868 (N_9868,N_4897,N_1458);
nand U9869 (N_9869,N_2997,N_586);
or U9870 (N_9870,N_1612,N_475);
nor U9871 (N_9871,N_4283,N_3251);
and U9872 (N_9872,N_829,N_1599);
nand U9873 (N_9873,N_4974,N_4654);
xnor U9874 (N_9874,N_1763,N_1368);
nand U9875 (N_9875,N_875,N_2312);
nor U9876 (N_9876,N_3885,N_2002);
nor U9877 (N_9877,N_948,N_4718);
nor U9878 (N_9878,N_3384,N_1640);
or U9879 (N_9879,N_1281,N_4137);
and U9880 (N_9880,N_2637,N_1980);
and U9881 (N_9881,N_410,N_3933);
and U9882 (N_9882,N_2242,N_3841);
nor U9883 (N_9883,N_1307,N_3657);
nand U9884 (N_9884,N_3362,N_4658);
nor U9885 (N_9885,N_3956,N_842);
nand U9886 (N_9886,N_806,N_1072);
nand U9887 (N_9887,N_4006,N_194);
nor U9888 (N_9888,N_1376,N_4283);
or U9889 (N_9889,N_4430,N_4096);
nor U9890 (N_9890,N_1158,N_299);
or U9891 (N_9891,N_4635,N_2755);
and U9892 (N_9892,N_917,N_3481);
or U9893 (N_9893,N_279,N_4145);
nand U9894 (N_9894,N_1081,N_3647);
and U9895 (N_9895,N_3229,N_2538);
and U9896 (N_9896,N_3893,N_3153);
or U9897 (N_9897,N_1044,N_2370);
and U9898 (N_9898,N_4802,N_4736);
and U9899 (N_9899,N_1659,N_3881);
nand U9900 (N_9900,N_4553,N_2419);
and U9901 (N_9901,N_1094,N_2027);
nand U9902 (N_9902,N_321,N_3943);
nand U9903 (N_9903,N_2995,N_1963);
nor U9904 (N_9904,N_257,N_4540);
and U9905 (N_9905,N_1058,N_3561);
nor U9906 (N_9906,N_1076,N_4244);
nor U9907 (N_9907,N_4483,N_2826);
xnor U9908 (N_9908,N_4916,N_4577);
nor U9909 (N_9909,N_4530,N_4589);
and U9910 (N_9910,N_1120,N_636);
nand U9911 (N_9911,N_408,N_775);
and U9912 (N_9912,N_2124,N_4839);
nand U9913 (N_9913,N_2483,N_4400);
or U9914 (N_9914,N_4072,N_2021);
nand U9915 (N_9915,N_1940,N_2124);
nand U9916 (N_9916,N_463,N_95);
xor U9917 (N_9917,N_3964,N_3805);
nand U9918 (N_9918,N_4255,N_1663);
xnor U9919 (N_9919,N_1094,N_2242);
nor U9920 (N_9920,N_3593,N_4816);
or U9921 (N_9921,N_4802,N_3541);
nand U9922 (N_9922,N_1068,N_898);
and U9923 (N_9923,N_2567,N_285);
or U9924 (N_9924,N_4715,N_4901);
or U9925 (N_9925,N_3521,N_3657);
or U9926 (N_9926,N_3559,N_4617);
or U9927 (N_9927,N_4830,N_1634);
or U9928 (N_9928,N_2795,N_3302);
or U9929 (N_9929,N_1752,N_1257);
nor U9930 (N_9930,N_3737,N_3345);
nand U9931 (N_9931,N_218,N_3349);
nor U9932 (N_9932,N_745,N_4166);
nor U9933 (N_9933,N_344,N_3894);
nor U9934 (N_9934,N_197,N_579);
or U9935 (N_9935,N_3475,N_622);
and U9936 (N_9936,N_3276,N_2354);
or U9937 (N_9937,N_1409,N_2911);
or U9938 (N_9938,N_217,N_3525);
or U9939 (N_9939,N_527,N_3101);
or U9940 (N_9940,N_2224,N_4316);
xor U9941 (N_9941,N_3688,N_3116);
and U9942 (N_9942,N_3022,N_2457);
nand U9943 (N_9943,N_4282,N_72);
nand U9944 (N_9944,N_3803,N_2471);
nand U9945 (N_9945,N_470,N_1380);
xnor U9946 (N_9946,N_82,N_2969);
nor U9947 (N_9947,N_331,N_3445);
xor U9948 (N_9948,N_612,N_2275);
xnor U9949 (N_9949,N_3010,N_2221);
nand U9950 (N_9950,N_1264,N_3188);
or U9951 (N_9951,N_3911,N_1211);
xnor U9952 (N_9952,N_1860,N_4899);
or U9953 (N_9953,N_1993,N_351);
and U9954 (N_9954,N_1666,N_1782);
nor U9955 (N_9955,N_4538,N_4596);
nor U9956 (N_9956,N_2545,N_1220);
and U9957 (N_9957,N_4094,N_14);
and U9958 (N_9958,N_4387,N_4775);
or U9959 (N_9959,N_764,N_3822);
nand U9960 (N_9960,N_3132,N_3225);
or U9961 (N_9961,N_3429,N_3680);
nor U9962 (N_9962,N_3299,N_4993);
or U9963 (N_9963,N_3868,N_4469);
or U9964 (N_9964,N_1345,N_2655);
nand U9965 (N_9965,N_476,N_4859);
and U9966 (N_9966,N_1170,N_726);
nor U9967 (N_9967,N_1114,N_2500);
or U9968 (N_9968,N_4547,N_785);
nand U9969 (N_9969,N_3475,N_3820);
nor U9970 (N_9970,N_1188,N_458);
nand U9971 (N_9971,N_3419,N_4937);
xnor U9972 (N_9972,N_2555,N_2917);
or U9973 (N_9973,N_4768,N_3616);
nand U9974 (N_9974,N_1328,N_2667);
xnor U9975 (N_9975,N_1250,N_2878);
nor U9976 (N_9976,N_4506,N_4400);
or U9977 (N_9977,N_2264,N_4620);
nor U9978 (N_9978,N_4897,N_694);
or U9979 (N_9979,N_1765,N_1469);
nor U9980 (N_9980,N_3397,N_3200);
xor U9981 (N_9981,N_4845,N_3854);
nand U9982 (N_9982,N_745,N_3669);
or U9983 (N_9983,N_1422,N_3970);
and U9984 (N_9984,N_1986,N_1694);
nor U9985 (N_9985,N_1632,N_4030);
or U9986 (N_9986,N_841,N_4847);
or U9987 (N_9987,N_2220,N_828);
nor U9988 (N_9988,N_4732,N_863);
xnor U9989 (N_9989,N_4834,N_4294);
xnor U9990 (N_9990,N_578,N_745);
nor U9991 (N_9991,N_3387,N_1916);
xor U9992 (N_9992,N_2730,N_3086);
or U9993 (N_9993,N_3836,N_243);
or U9994 (N_9994,N_1083,N_3323);
nand U9995 (N_9995,N_2214,N_3779);
nand U9996 (N_9996,N_4923,N_4286);
or U9997 (N_9997,N_2235,N_3021);
xnor U9998 (N_9998,N_1869,N_2633);
nor U9999 (N_9999,N_3258,N_1387);
nand U10000 (N_10000,N_7863,N_8524);
nand U10001 (N_10001,N_6287,N_9015);
or U10002 (N_10002,N_9475,N_5509);
nor U10003 (N_10003,N_6952,N_9531);
nand U10004 (N_10004,N_9799,N_7486);
or U10005 (N_10005,N_6686,N_7360);
and U10006 (N_10006,N_5834,N_8484);
or U10007 (N_10007,N_9464,N_9256);
xnor U10008 (N_10008,N_8339,N_8024);
or U10009 (N_10009,N_8944,N_9867);
nand U10010 (N_10010,N_9916,N_8340);
and U10011 (N_10011,N_5030,N_9820);
nor U10012 (N_10012,N_8547,N_9018);
or U10013 (N_10013,N_8337,N_8264);
and U10014 (N_10014,N_5308,N_7438);
or U10015 (N_10015,N_8408,N_8834);
or U10016 (N_10016,N_8982,N_8189);
nand U10017 (N_10017,N_6736,N_9051);
xor U10018 (N_10018,N_7504,N_5559);
xor U10019 (N_10019,N_8295,N_9796);
nand U10020 (N_10020,N_5982,N_9486);
and U10021 (N_10021,N_6744,N_8660);
and U10022 (N_10022,N_8810,N_6175);
nand U10023 (N_10023,N_5254,N_8876);
nor U10024 (N_10024,N_8857,N_9188);
nor U10025 (N_10025,N_7700,N_5346);
and U10026 (N_10026,N_9915,N_7988);
or U10027 (N_10027,N_9035,N_5345);
or U10028 (N_10028,N_6578,N_7408);
or U10029 (N_10029,N_5201,N_5879);
and U10030 (N_10030,N_9436,N_8599);
and U10031 (N_10031,N_8055,N_9925);
and U10032 (N_10032,N_6072,N_6332);
nand U10033 (N_10033,N_7778,N_6840);
nand U10034 (N_10034,N_7240,N_7015);
nand U10035 (N_10035,N_5763,N_6319);
or U10036 (N_10036,N_7353,N_6932);
nor U10037 (N_10037,N_8826,N_7218);
and U10038 (N_10038,N_6362,N_7311);
and U10039 (N_10039,N_5418,N_8073);
nor U10040 (N_10040,N_8509,N_5184);
or U10041 (N_10041,N_5284,N_9271);
or U10042 (N_10042,N_6433,N_6328);
nor U10043 (N_10043,N_6834,N_9133);
nand U10044 (N_10044,N_9886,N_8533);
xor U10045 (N_10045,N_8964,N_8867);
nand U10046 (N_10046,N_8182,N_8864);
xor U10047 (N_10047,N_7323,N_9758);
or U10048 (N_10048,N_6029,N_6716);
nand U10049 (N_10049,N_9872,N_9209);
and U10050 (N_10050,N_9408,N_6115);
and U10051 (N_10051,N_5794,N_7586);
nand U10052 (N_10052,N_6698,N_5529);
and U10053 (N_10053,N_9746,N_8743);
xnor U10054 (N_10054,N_8811,N_7362);
and U10055 (N_10055,N_6039,N_5717);
nor U10056 (N_10056,N_6634,N_6585);
or U10057 (N_10057,N_7799,N_5438);
nor U10058 (N_10058,N_7813,N_8054);
nor U10059 (N_10059,N_6277,N_8661);
and U10060 (N_10060,N_8092,N_6633);
nand U10061 (N_10061,N_7435,N_7800);
and U10062 (N_10062,N_5480,N_7202);
or U10063 (N_10063,N_9631,N_7177);
nor U10064 (N_10064,N_5017,N_9666);
and U10065 (N_10065,N_5870,N_9422);
xor U10066 (N_10066,N_9638,N_8248);
and U10067 (N_10067,N_8767,N_8010);
nand U10068 (N_10068,N_7550,N_5640);
and U10069 (N_10069,N_5806,N_6264);
nor U10070 (N_10070,N_6192,N_8332);
nand U10071 (N_10071,N_6389,N_7124);
or U10072 (N_10072,N_5043,N_9564);
nand U10073 (N_10073,N_9870,N_7625);
nor U10074 (N_10074,N_6798,N_9478);
nand U10075 (N_10075,N_6684,N_7477);
or U10076 (N_10076,N_8507,N_5251);
or U10077 (N_10077,N_8620,N_5842);
and U10078 (N_10078,N_8222,N_7050);
nor U10079 (N_10079,N_6385,N_7961);
or U10080 (N_10080,N_9058,N_7642);
and U10081 (N_10081,N_7656,N_6769);
nand U10082 (N_10082,N_8925,N_7650);
xnor U10083 (N_10083,N_6141,N_7102);
or U10084 (N_10084,N_7940,N_8855);
nor U10085 (N_10085,N_8768,N_5570);
or U10086 (N_10086,N_9361,N_5769);
or U10087 (N_10087,N_7298,N_7792);
nor U10088 (N_10088,N_9964,N_9411);
xnor U10089 (N_10089,N_7003,N_6820);
or U10090 (N_10090,N_6282,N_8207);
or U10091 (N_10091,N_6424,N_5857);
nor U10092 (N_10092,N_5174,N_5428);
or U10093 (N_10093,N_7722,N_7972);
or U10094 (N_10094,N_9937,N_9007);
nor U10095 (N_10095,N_7544,N_7502);
nand U10096 (N_10096,N_9332,N_9933);
xor U10097 (N_10097,N_5878,N_9159);
nand U10098 (N_10098,N_8549,N_6823);
and U10099 (N_10099,N_6721,N_9513);
nand U10100 (N_10100,N_9865,N_7578);
nor U10101 (N_10101,N_8276,N_7276);
and U10102 (N_10102,N_5996,N_7838);
and U10103 (N_10103,N_7803,N_9134);
and U10104 (N_10104,N_8459,N_6781);
nor U10105 (N_10105,N_6107,N_9469);
nand U10106 (N_10106,N_7457,N_7583);
nand U10107 (N_10107,N_7216,N_7290);
nor U10108 (N_10108,N_8235,N_8372);
and U10109 (N_10109,N_9982,N_8034);
nand U10110 (N_10110,N_7379,N_6344);
nand U10111 (N_10111,N_9369,N_6213);
nand U10112 (N_10112,N_6479,N_7695);
or U10113 (N_10113,N_6460,N_5257);
nor U10114 (N_10114,N_6811,N_8977);
nor U10115 (N_10115,N_6727,N_7172);
nor U10116 (N_10116,N_5245,N_9935);
nand U10117 (N_10117,N_5215,N_8185);
nand U10118 (N_10118,N_9049,N_5468);
nand U10119 (N_10119,N_7366,N_6281);
and U10120 (N_10120,N_7646,N_6550);
nor U10121 (N_10121,N_7491,N_5984);
nand U10122 (N_10122,N_7345,N_7764);
or U10123 (N_10123,N_7380,N_9519);
nor U10124 (N_10124,N_6041,N_9249);
or U10125 (N_10125,N_8609,N_8036);
nor U10126 (N_10126,N_6379,N_6278);
nand U10127 (N_10127,N_6667,N_5267);
nor U10128 (N_10128,N_7503,N_6280);
nor U10129 (N_10129,N_7356,N_7953);
and U10130 (N_10130,N_7287,N_5786);
nand U10131 (N_10131,N_6937,N_5289);
nand U10132 (N_10132,N_6019,N_7830);
or U10133 (N_10133,N_9538,N_5021);
xnor U10134 (N_10134,N_7051,N_7517);
or U10135 (N_10135,N_6301,N_6742);
nor U10136 (N_10136,N_9731,N_6227);
nand U10137 (N_10137,N_5551,N_6963);
and U10138 (N_10138,N_7652,N_7787);
xor U10139 (N_10139,N_7249,N_6881);
xor U10140 (N_10140,N_9410,N_7350);
nor U10141 (N_10141,N_8851,N_6873);
nor U10142 (N_10142,N_5651,N_5285);
nor U10143 (N_10143,N_8695,N_7344);
xor U10144 (N_10144,N_5507,N_8956);
or U10145 (N_10145,N_5770,N_9741);
nand U10146 (N_10146,N_8902,N_8259);
nand U10147 (N_10147,N_6608,N_6388);
nor U10148 (N_10148,N_8502,N_7014);
and U10149 (N_10149,N_7155,N_9629);
or U10150 (N_10150,N_9177,N_5138);
nor U10151 (N_10151,N_9499,N_7509);
xnor U10152 (N_10152,N_5190,N_7390);
nor U10153 (N_10153,N_9502,N_8909);
and U10154 (N_10154,N_5073,N_8156);
nor U10155 (N_10155,N_5964,N_7377);
nand U10156 (N_10156,N_8359,N_8519);
or U10157 (N_10157,N_8048,N_6659);
nand U10158 (N_10158,N_7531,N_8253);
nand U10159 (N_10159,N_6047,N_6070);
nand U10160 (N_10160,N_6267,N_7569);
or U10161 (N_10161,N_7129,N_6541);
and U10162 (N_10162,N_8541,N_8118);
nand U10163 (N_10163,N_8853,N_6165);
nor U10164 (N_10164,N_8970,N_8001);
and U10165 (N_10165,N_7592,N_7056);
and U10166 (N_10166,N_6642,N_6168);
or U10167 (N_10167,N_7622,N_9019);
and U10168 (N_10168,N_8758,N_8492);
xnor U10169 (N_10169,N_6582,N_6208);
nand U10170 (N_10170,N_8731,N_9505);
and U10171 (N_10171,N_9246,N_9691);
or U10172 (N_10172,N_6569,N_6884);
and U10173 (N_10173,N_5573,N_7682);
nor U10174 (N_10174,N_8070,N_6316);
or U10175 (N_10175,N_9461,N_5130);
nand U10176 (N_10176,N_8446,N_7957);
and U10177 (N_10177,N_8943,N_8198);
nor U10178 (N_10178,N_8984,N_5180);
or U10179 (N_10179,N_5571,N_6290);
or U10180 (N_10180,N_8428,N_6462);
nor U10181 (N_10181,N_5622,N_9186);
nor U10182 (N_10182,N_5682,N_6464);
nand U10183 (N_10183,N_8442,N_7610);
nor U10184 (N_10184,N_9624,N_8421);
nor U10185 (N_10185,N_9041,N_9922);
nand U10186 (N_10186,N_8475,N_7539);
and U10187 (N_10187,N_5916,N_5113);
and U10188 (N_10188,N_5349,N_7798);
nor U10189 (N_10189,N_8949,N_5549);
or U10190 (N_10190,N_7765,N_9802);
nor U10191 (N_10191,N_8701,N_8912);
and U10192 (N_10192,N_8726,N_9111);
and U10193 (N_10193,N_5965,N_8788);
or U10194 (N_10194,N_6522,N_9305);
nand U10195 (N_10195,N_8261,N_5033);
nand U10196 (N_10196,N_5941,N_7186);
nand U10197 (N_10197,N_8184,N_7079);
xnor U10198 (N_10198,N_9273,N_5925);
nand U10199 (N_10199,N_6855,N_6885);
and U10200 (N_10200,N_5329,N_8432);
or U10201 (N_10201,N_9254,N_5676);
and U10202 (N_10202,N_5353,N_6552);
nor U10203 (N_10203,N_7150,N_5635);
or U10204 (N_10204,N_9275,N_6342);
or U10205 (N_10205,N_7779,N_6059);
xor U10206 (N_10206,N_8821,N_8346);
nand U10207 (N_10207,N_7283,N_7042);
nor U10208 (N_10208,N_9244,N_7818);
nor U10209 (N_10209,N_8687,N_7132);
nor U10210 (N_10210,N_9929,N_9043);
or U10211 (N_10211,N_9530,N_5587);
nor U10212 (N_10212,N_9384,N_9658);
nor U10213 (N_10213,N_7244,N_6590);
nor U10214 (N_10214,N_8004,N_5375);
nand U10215 (N_10215,N_9614,N_6745);
nor U10216 (N_10216,N_7157,N_5615);
xor U10217 (N_10217,N_6685,N_9549);
or U10218 (N_10218,N_9036,N_6027);
nand U10219 (N_10219,N_5268,N_7588);
nor U10220 (N_10220,N_5161,N_7512);
nand U10221 (N_10221,N_8969,N_6611);
and U10222 (N_10222,N_6360,N_9783);
or U10223 (N_10223,N_8324,N_7777);
xor U10224 (N_10224,N_8779,N_9226);
xnor U10225 (N_10225,N_9652,N_5880);
and U10226 (N_10226,N_9797,N_6283);
nand U10227 (N_10227,N_5394,N_6321);
nand U10228 (N_10228,N_8848,N_9262);
nand U10229 (N_10229,N_6392,N_6270);
nor U10230 (N_10230,N_5160,N_9554);
and U10231 (N_10231,N_6524,N_6242);
nor U10232 (N_10232,N_8995,N_8501);
nor U10233 (N_10233,N_9492,N_5383);
or U10234 (N_10234,N_5293,N_8503);
nor U10235 (N_10235,N_8735,N_9957);
xnor U10236 (N_10236,N_5080,N_6597);
nand U10237 (N_10237,N_5874,N_7442);
or U10238 (N_10238,N_8476,N_8239);
or U10239 (N_10239,N_6036,N_9034);
nand U10240 (N_10240,N_9642,N_5821);
nor U10241 (N_10241,N_6448,N_5291);
and U10242 (N_10242,N_5337,N_5156);
and U10243 (N_10243,N_6446,N_7995);
nor U10244 (N_10244,N_7144,N_8896);
and U10245 (N_10245,N_5566,N_7549);
or U10246 (N_10246,N_9222,N_6519);
or U10247 (N_10247,N_8763,N_8965);
nand U10248 (N_10248,N_7629,N_6187);
and U10249 (N_10249,N_9374,N_9483);
and U10250 (N_10250,N_6094,N_5176);
nor U10251 (N_10251,N_5679,N_9927);
or U10252 (N_10252,N_9717,N_8742);
nand U10253 (N_10253,N_8143,N_6133);
nand U10254 (N_10254,N_6330,N_5826);
xor U10255 (N_10255,N_9546,N_5825);
nor U10256 (N_10256,N_8579,N_5038);
or U10257 (N_10257,N_5588,N_5482);
and U10258 (N_10258,N_6430,N_7591);
xnor U10259 (N_10259,N_8244,N_6371);
nand U10260 (N_10260,N_8177,N_6688);
xnor U10261 (N_10261,N_8762,N_7872);
and U10262 (N_10262,N_9214,N_6217);
and U10263 (N_10263,N_8534,N_7904);
or U10264 (N_10264,N_6835,N_5844);
or U10265 (N_10265,N_5619,N_8150);
nand U10266 (N_10266,N_6364,N_8319);
or U10267 (N_10267,N_5342,N_8078);
nor U10268 (N_10268,N_7414,N_9328);
or U10269 (N_10269,N_7189,N_8082);
xnor U10270 (N_10270,N_5753,N_9511);
nor U10271 (N_10271,N_9518,N_5934);
or U10272 (N_10272,N_8968,N_7762);
or U10273 (N_10273,N_8570,N_6011);
nor U10274 (N_10274,N_6704,N_7068);
nor U10275 (N_10275,N_8260,N_7984);
nor U10276 (N_10276,N_7483,N_8284);
nand U10277 (N_10277,N_8021,N_5339);
or U10278 (N_10278,N_5528,N_7012);
or U10279 (N_10279,N_5933,N_7378);
xnor U10280 (N_10280,N_6419,N_5417);
or U10281 (N_10281,N_9786,N_5641);
nand U10282 (N_10282,N_8514,N_9683);
nor U10283 (N_10283,N_9515,N_5478);
or U10284 (N_10284,N_8676,N_7288);
and U10285 (N_10285,N_9837,N_7365);
and U10286 (N_10286,N_9924,N_9757);
or U10287 (N_10287,N_8681,N_8387);
nand U10288 (N_10288,N_8472,N_9667);
or U10289 (N_10289,N_8910,N_7420);
or U10290 (N_10290,N_9230,N_8398);
and U10291 (N_10291,N_8338,N_8448);
xnor U10292 (N_10292,N_5690,N_7963);
nand U10293 (N_10293,N_5369,N_8229);
and U10294 (N_10294,N_7690,N_8343);
or U10295 (N_10295,N_6327,N_7309);
and U10296 (N_10296,N_5175,N_6791);
or U10297 (N_10297,N_5382,N_5590);
nand U10298 (N_10298,N_6207,N_6728);
and U10299 (N_10299,N_6712,N_6893);
nor U10300 (N_10300,N_8258,N_5830);
nand U10301 (N_10301,N_9057,N_6390);
nand U10302 (N_10302,N_7923,N_8176);
xor U10303 (N_10303,N_8686,N_5773);
nand U10304 (N_10304,N_9120,N_7825);
or U10305 (N_10305,N_8350,N_8132);
nor U10306 (N_10306,N_9524,N_7370);
and U10307 (N_10307,N_5935,N_8133);
nand U10308 (N_10308,N_9775,N_7201);
nor U10309 (N_10309,N_7008,N_7031);
and U10310 (N_10310,N_6169,N_5315);
and U10311 (N_10311,N_8199,N_5368);
and U10312 (N_10312,N_5592,N_8528);
and U10313 (N_10313,N_5188,N_8022);
nand U10314 (N_10314,N_8617,N_8069);
nor U10315 (N_10315,N_7900,N_8497);
nand U10316 (N_10316,N_9896,N_6476);
nand U10317 (N_10317,N_5716,N_7081);
nor U10318 (N_10318,N_9993,N_6488);
or U10319 (N_10319,N_7870,N_6549);
xnor U10320 (N_10320,N_9286,N_9640);
xor U10321 (N_10321,N_6996,N_7910);
nor U10322 (N_10322,N_8068,N_9711);
and U10323 (N_10323,N_9489,N_8394);
nand U10324 (N_10324,N_9028,N_7460);
nand U10325 (N_10325,N_9815,N_5162);
xnor U10326 (N_10326,N_7243,N_7059);
nor U10327 (N_10327,N_6251,N_8154);
or U10328 (N_10328,N_6012,N_6995);
nand U10329 (N_10329,N_7738,N_7418);
xor U10330 (N_10330,N_9897,N_7396);
and U10331 (N_10331,N_5526,N_6052);
nor U10332 (N_10332,N_6156,N_9462);
and U10333 (N_10333,N_6429,N_5807);
nor U10334 (N_10334,N_5617,N_7901);
and U10335 (N_10335,N_9930,N_6426);
and U10336 (N_10336,N_6773,N_7480);
xor U10337 (N_10337,N_5746,N_7675);
or U10338 (N_10338,N_9413,N_9399);
or U10339 (N_10339,N_5975,N_8088);
nor U10340 (N_10340,N_8685,N_7403);
nor U10341 (N_10341,N_6555,N_8427);
or U10342 (N_10342,N_6225,N_8801);
and U10343 (N_10343,N_7874,N_9782);
or U10344 (N_10344,N_8397,N_7742);
or U10345 (N_10345,N_8066,N_9999);
nor U10346 (N_10346,N_7865,N_7278);
or U10347 (N_10347,N_8254,N_5022);
nand U10348 (N_10348,N_8075,N_6856);
or U10349 (N_10349,N_9107,N_5154);
nor U10350 (N_10350,N_7808,N_6637);
nand U10351 (N_10351,N_6179,N_6400);
or U10352 (N_10352,N_7417,N_9264);
nand U10353 (N_10353,N_6244,N_6195);
and U10354 (N_10354,N_9725,N_7098);
xor U10355 (N_10355,N_5132,N_6037);
nand U10356 (N_10356,N_9781,N_7839);
nor U10357 (N_10357,N_5049,N_6486);
xnor U10358 (N_10358,N_6977,N_8690);
or U10359 (N_10359,N_9849,N_6719);
xor U10360 (N_10360,N_8730,N_6753);
nand U10361 (N_10361,N_9952,N_8736);
and U10362 (N_10362,N_8808,N_8454);
or U10363 (N_10363,N_7727,N_8149);
or U10364 (N_10364,N_6665,N_7116);
nor U10365 (N_10365,N_5993,N_5522);
nor U10366 (N_10366,N_7239,N_6558);
nand U10367 (N_10367,N_8607,N_8757);
nand U10368 (N_10368,N_6897,N_7667);
and U10369 (N_10369,N_5957,N_8100);
nor U10370 (N_10370,N_5700,N_5508);
nand U10371 (N_10371,N_5689,N_9217);
nand U10372 (N_10372,N_9165,N_6553);
and U10373 (N_10373,N_9311,N_6696);
nor U10374 (N_10374,N_8216,N_8228);
or U10375 (N_10375,N_9779,N_5272);
nor U10376 (N_10376,N_5504,N_8613);
and U10377 (N_10377,N_9452,N_6738);
and U10378 (N_10378,N_5663,N_5312);
or U10379 (N_10379,N_7530,N_7536);
nor U10380 (N_10380,N_5462,N_7117);
nor U10381 (N_10381,N_9263,N_8174);
nor U10382 (N_10382,N_7020,N_6074);
or U10383 (N_10383,N_7494,N_9383);
nand U10384 (N_10384,N_7409,N_9045);
or U10385 (N_10385,N_5045,N_7441);
nand U10386 (N_10386,N_5856,N_9054);
nor U10387 (N_10387,N_8847,N_7226);
and U10388 (N_10388,N_7627,N_7782);
or U10389 (N_10389,N_9917,N_8414);
nor U10390 (N_10390,N_7816,N_5466);
or U10391 (N_10391,N_5139,N_9636);
nor U10392 (N_10392,N_6050,N_8085);
nor U10393 (N_10393,N_7598,N_5860);
and U10394 (N_10394,N_8976,N_5929);
nor U10395 (N_10395,N_8854,N_8605);
nand U10396 (N_10396,N_7999,N_7346);
nor U10397 (N_10397,N_5544,N_9071);
and U10398 (N_10398,N_9899,N_6235);
or U10399 (N_10399,N_9176,N_5411);
or U10400 (N_10400,N_7542,N_5359);
nand U10401 (N_10401,N_9685,N_9842);
and U10402 (N_10402,N_5662,N_7316);
nand U10403 (N_10403,N_8094,N_7285);
and U10404 (N_10404,N_6583,N_8702);
xor U10405 (N_10405,N_7703,N_7065);
xnor U10406 (N_10406,N_6949,N_8564);
and U10407 (N_10407,N_6139,N_8275);
xnor U10408 (N_10408,N_9233,N_7585);
nor U10409 (N_10409,N_9920,N_6409);
nand U10410 (N_10410,N_6878,N_5235);
and U10411 (N_10411,N_8866,N_9156);
nor U10412 (N_10412,N_5970,N_9495);
nand U10413 (N_10413,N_6160,N_6702);
or U10414 (N_10414,N_5586,N_5601);
nand U10415 (N_10415,N_9493,N_8148);
nor U10416 (N_10416,N_9889,N_6405);
and U10417 (N_10417,N_8027,N_5674);
nor U10418 (N_10418,N_5968,N_5330);
or U10419 (N_10419,N_9137,N_8355);
and U10420 (N_10420,N_6289,N_6067);
nand U10421 (N_10421,N_8693,N_6166);
and U10422 (N_10422,N_7708,N_6975);
nand U10423 (N_10423,N_9856,N_8850);
nor U10424 (N_10424,N_7720,N_8365);
and U10425 (N_10425,N_5764,N_5388);
nor U10426 (N_10426,N_5789,N_5051);
nand U10427 (N_10427,N_5500,N_7431);
or U10428 (N_10428,N_6147,N_7789);
nand U10429 (N_10429,N_7263,N_7426);
and U10430 (N_10430,N_8265,N_5414);
or U10431 (N_10431,N_8796,N_8578);
xnor U10432 (N_10432,N_5506,N_8106);
nor U10433 (N_10433,N_9845,N_6879);
nand U10434 (N_10434,N_9810,N_6335);
or U10435 (N_10435,N_9155,N_6760);
or U10436 (N_10436,N_6609,N_5638);
and U10437 (N_10437,N_5998,N_7617);
and U10438 (N_10438,N_7935,N_5196);
or U10439 (N_10439,N_8415,N_6323);
nand U10440 (N_10440,N_9963,N_5589);
and U10441 (N_10441,N_6715,N_7686);
or U10442 (N_10442,N_9690,N_7011);
and U10443 (N_10443,N_5492,N_9914);
nand U10444 (N_10444,N_8981,N_9432);
nand U10445 (N_10445,N_9251,N_6620);
nor U10446 (N_10446,N_8941,N_8107);
or U10447 (N_10447,N_6480,N_8733);
nand U10448 (N_10448,N_6313,N_6384);
and U10449 (N_10449,N_6421,N_6625);
or U10450 (N_10450,N_5730,N_7797);
and U10451 (N_10451,N_6383,N_6940);
nand U10452 (N_10452,N_8151,N_9882);
and U10453 (N_10453,N_9807,N_5495);
and U10454 (N_10454,N_6345,N_5863);
nand U10455 (N_10455,N_9995,N_6492);
nand U10456 (N_10456,N_9269,N_6528);
nand U10457 (N_10457,N_6604,N_6030);
nor U10458 (N_10458,N_9737,N_7022);
and U10459 (N_10459,N_6451,N_9871);
nor U10460 (N_10460,N_7982,N_7479);
and U10461 (N_10461,N_9597,N_6116);
nand U10462 (N_10462,N_6422,N_6516);
xor U10463 (N_10463,N_8536,N_9533);
nand U10464 (N_10464,N_7723,N_9127);
nor U10465 (N_10465,N_9138,N_9545);
nand U10466 (N_10466,N_8056,N_7168);
or U10467 (N_10467,N_9829,N_8963);
or U10468 (N_10468,N_8168,N_9894);
or U10469 (N_10469,N_7151,N_6109);
xnor U10470 (N_10470,N_8345,N_8680);
nand U10471 (N_10471,N_5103,N_7925);
or U10472 (N_10472,N_7853,N_6617);
xnor U10473 (N_10473,N_7133,N_6161);
nand U10474 (N_10474,N_6525,N_9303);
nand U10475 (N_10475,N_8918,N_8341);
nand U10476 (N_10476,N_9077,N_5006);
nor U10477 (N_10477,N_7179,N_8431);
nand U10478 (N_10478,N_6456,N_8939);
xnor U10479 (N_10479,N_5241,N_6197);
and U10480 (N_10480,N_9285,N_7987);
nand U10481 (N_10481,N_5403,N_7843);
nor U10482 (N_10482,N_9932,N_9319);
and U10483 (N_10483,N_6567,N_5702);
and U10484 (N_10484,N_5840,N_5486);
or U10485 (N_10485,N_9923,N_9470);
xor U10486 (N_10486,N_5978,N_6485);
xnor U10487 (N_10487,N_7702,N_5936);
nor U10488 (N_10488,N_9552,N_6854);
nor U10489 (N_10489,N_6018,N_8666);
and U10490 (N_10490,N_6145,N_9987);
and U10491 (N_10491,N_9064,N_6586);
nor U10492 (N_10492,N_6089,N_5079);
or U10493 (N_10493,N_8434,N_7579);
and U10494 (N_10494,N_9429,N_6741);
nand U10495 (N_10495,N_7230,N_6357);
or U10496 (N_10496,N_8020,N_7752);
and U10497 (N_10497,N_7891,N_6711);
or U10498 (N_10498,N_9985,N_5032);
nor U10499 (N_10499,N_6477,N_7330);
and U10500 (N_10500,N_8243,N_9123);
nor U10501 (N_10501,N_8167,N_9537);
nand U10502 (N_10502,N_8173,N_5927);
nand U10503 (N_10503,N_6926,N_5944);
and U10504 (N_10504,N_6576,N_8430);
or U10505 (N_10505,N_7694,N_7072);
xnor U10506 (N_10506,N_8957,N_7123);
or U10507 (N_10507,N_8740,N_9003);
nand U10508 (N_10508,N_8749,N_7785);
nand U10509 (N_10509,N_5961,N_8917);
or U10510 (N_10510,N_7104,N_6514);
nor U10511 (N_10511,N_7930,N_9232);
nand U10512 (N_10512,N_5661,N_7898);
or U10513 (N_10513,N_6465,N_9121);
nor U10514 (N_10514,N_7246,N_9444);
nand U10515 (N_10515,N_5275,N_9268);
or U10516 (N_10516,N_7661,N_9850);
nand U10517 (N_10517,N_5081,N_7985);
nand U10518 (N_10518,N_6431,N_7282);
nor U10519 (N_10519,N_5652,N_8436);
nand U10520 (N_10520,N_5818,N_7130);
nand U10521 (N_10521,N_6755,N_9241);
and U10522 (N_10522,N_8009,N_8590);
nor U10523 (N_10523,N_9203,N_9247);
xor U10524 (N_10524,N_7566,N_9231);
xnor U10525 (N_10525,N_5695,N_8232);
nand U10526 (N_10526,N_5599,N_8440);
nor U10527 (N_10527,N_8161,N_7268);
and U10528 (N_10528,N_9736,N_9948);
nor U10529 (N_10529,N_5378,N_6865);
nor U10530 (N_10530,N_8483,N_9401);
or U10531 (N_10531,N_9240,N_6097);
nor U10532 (N_10532,N_8996,N_6310);
nor U10533 (N_10533,N_9888,N_6111);
nor U10534 (N_10534,N_7430,N_6173);
nand U10535 (N_10535,N_6258,N_5243);
nand U10536 (N_10536,N_6750,N_9130);
xor U10537 (N_10537,N_5020,N_7600);
nor U10538 (N_10538,N_5459,N_6177);
nor U10539 (N_10539,N_5814,N_9647);
nand U10540 (N_10540,N_8462,N_5287);
nand U10541 (N_10541,N_9504,N_9853);
nor U10542 (N_10542,N_7521,N_7633);
or U10543 (N_10543,N_7774,N_9713);
nor U10544 (N_10544,N_6518,N_9967);
or U10545 (N_10545,N_9258,N_9664);
and U10546 (N_10546,N_9073,N_8897);
nand U10547 (N_10547,N_5269,N_7302);
or U10548 (N_10548,N_9795,N_9221);
xnor U10549 (N_10549,N_5483,N_7225);
and U10550 (N_10550,N_5451,N_7826);
nor U10551 (N_10551,N_9005,N_6299);
nor U10552 (N_10552,N_6568,N_6325);
xor U10553 (N_10553,N_7207,N_7200);
and U10554 (N_10554,N_6643,N_5340);
nand U10555 (N_10555,N_8437,N_6378);
nand U10556 (N_10556,N_9969,N_8929);
or U10557 (N_10557,N_5782,N_6923);
nor U10558 (N_10558,N_8766,N_8160);
and U10559 (N_10559,N_7562,N_5888);
or U10560 (N_10560,N_8014,N_5246);
and U10561 (N_10561,N_9650,N_6679);
or U10562 (N_10562,N_5109,N_5252);
nand U10563 (N_10563,N_9292,N_8395);
nand U10564 (N_10564,N_9169,N_7547);
and U10565 (N_10565,N_9593,N_6944);
or U10566 (N_10566,N_8400,N_5439);
nor U10567 (N_10567,N_8513,N_9790);
nor U10568 (N_10568,N_5453,N_8256);
and U10569 (N_10569,N_5166,N_9477);
nand U10570 (N_10570,N_8734,N_8494);
nor U10571 (N_10571,N_9378,N_7381);
and U10572 (N_10572,N_8404,N_5708);
or U10573 (N_10573,N_8782,N_8392);
nand U10574 (N_10574,N_9280,N_9874);
and U10575 (N_10575,N_9228,N_5776);
nand U10576 (N_10576,N_6110,N_7847);
or U10577 (N_10577,N_5565,N_9526);
nor U10578 (N_10578,N_7310,N_7715);
nand U10579 (N_10579,N_9097,N_5042);
nor U10580 (N_10580,N_6726,N_7520);
xnor U10581 (N_10581,N_9298,N_9317);
nor U10582 (N_10582,N_6824,N_9668);
and U10583 (N_10583,N_8540,N_7635);
or U10584 (N_10584,N_7804,N_9575);
nand U10585 (N_10585,N_7500,N_5144);
or U10586 (N_10586,N_9581,N_5871);
or U10587 (N_10587,N_5292,N_5406);
xnor U10588 (N_10588,N_9075,N_8347);
xnor U10589 (N_10589,N_5798,N_5598);
nand U10590 (N_10590,N_6122,N_5775);
and U10591 (N_10591,N_9687,N_8269);
and U10592 (N_10592,N_7571,N_7327);
or U10593 (N_10593,N_7584,N_7203);
nor U10594 (N_10594,N_7142,N_9941);
nand U10595 (N_10595,N_7641,N_9027);
nand U10596 (N_10596,N_6697,N_6947);
nor U10597 (N_10597,N_8662,N_9976);
and U10598 (N_10598,N_7010,N_5419);
nor U10599 (N_10599,N_8525,N_5367);
nor U10600 (N_10600,N_5228,N_8606);
or U10601 (N_10601,N_8129,N_5511);
or U10602 (N_10602,N_8111,N_7038);
and U10603 (N_10603,N_7807,N_5833);
and U10604 (N_10604,N_8219,N_9766);
xor U10605 (N_10605,N_8461,N_6226);
and U10606 (N_10606,N_5048,N_5307);
or U10607 (N_10607,N_6482,N_8644);
nor U10608 (N_10608,N_6707,N_5460);
nand U10609 (N_10609,N_9772,N_6123);
or U10610 (N_10610,N_9125,N_5692);
nor U10611 (N_10611,N_6043,N_9416);
nand U10612 (N_10612,N_7689,N_8304);
nor U10613 (N_10613,N_5943,N_7419);
or U10614 (N_10614,N_6209,N_6584);
nand U10615 (N_10615,N_5214,N_7581);
nor U10616 (N_10616,N_5639,N_6709);
or U10617 (N_10617,N_5265,N_8999);
nor U10618 (N_10618,N_7078,N_7555);
nor U10619 (N_10619,N_6619,N_6635);
xor U10620 (N_10620,N_7410,N_5802);
or U10621 (N_10621,N_5634,N_7971);
xor U10622 (N_10622,N_8973,N_8382);
nand U10623 (N_10623,N_9110,N_9335);
nand U10624 (N_10624,N_7358,N_7801);
nand U10625 (N_10625,N_5971,N_8962);
nor U10626 (N_10626,N_9732,N_9627);
nand U10627 (N_10627,N_7447,N_9323);
or U10628 (N_10628,N_9161,N_6513);
nor U10629 (N_10629,N_7678,N_9172);
and U10630 (N_10630,N_7837,N_9544);
nor U10631 (N_10631,N_6414,N_6382);
and U10632 (N_10632,N_7469,N_8558);
nor U10633 (N_10633,N_5686,N_9721);
and U10634 (N_10634,N_6336,N_6381);
nor U10635 (N_10635,N_7574,N_7505);
or U10636 (N_10636,N_7620,N_6628);
nor U10637 (N_10637,N_9083,N_6483);
and U10638 (N_10638,N_9451,N_6565);
nor U10639 (N_10639,N_5318,N_6159);
xnor U10640 (N_10640,N_9858,N_8165);
and U10641 (N_10641,N_8815,N_8930);
nand U10642 (N_10642,N_9639,N_8839);
or U10643 (N_10643,N_9142,N_8527);
nor U10644 (N_10644,N_6554,N_7519);
and U10645 (N_10645,N_5521,N_5656);
or U10646 (N_10646,N_8566,N_6471);
or U10647 (N_10647,N_8648,N_7312);
nand U10648 (N_10648,N_6463,N_8694);
and U10649 (N_10649,N_8268,N_5047);
xor U10650 (N_10650,N_9014,N_7424);
and U10651 (N_10651,N_6681,N_8402);
and U10652 (N_10652,N_9770,N_6563);
and U10653 (N_10653,N_5303,N_5301);
and U10654 (N_10654,N_7304,N_6527);
or U10655 (N_10655,N_9199,N_8664);
xor U10656 (N_10656,N_7856,N_8409);
nand U10657 (N_10657,N_5614,N_9778);
nor U10658 (N_10658,N_9402,N_8357);
xnor U10659 (N_10659,N_5328,N_7744);
nand U10660 (N_10660,N_5488,N_7308);
nand U10661 (N_10661,N_5886,N_9283);
and U10662 (N_10662,N_5644,N_7223);
nand U10663 (N_10663,N_7023,N_8785);
xor U10664 (N_10664,N_7658,N_8732);
nor U10665 (N_10665,N_6228,N_5093);
and U10666 (N_10666,N_6082,N_5013);
nand U10667 (N_10667,N_6042,N_5310);
and U10668 (N_10668,N_7572,N_6777);
or U10669 (N_10669,N_7740,N_9497);
nor U10670 (N_10670,N_5707,N_8250);
nand U10671 (N_10671,N_8146,N_6794);
and U10672 (N_10672,N_6470,N_9836);
nand U10673 (N_10673,N_6454,N_5255);
nor U10674 (N_10674,N_7376,N_8531);
or U10675 (N_10675,N_7590,N_9726);
nand U10676 (N_10676,N_8325,N_9239);
nor U10677 (N_10677,N_8804,N_7508);
nand U10678 (N_10678,N_9122,N_8831);
nor U10679 (N_10679,N_8905,N_7540);
nor U10680 (N_10680,N_6222,N_5364);
and U10681 (N_10681,N_7842,N_8794);
and U10682 (N_10682,N_6091,N_8096);
and U10683 (N_10683,N_5288,N_7432);
or U10684 (N_10684,N_5637,N_7190);
nand U10685 (N_10685,N_8042,N_6804);
and U10686 (N_10686,N_6506,N_5490);
and U10687 (N_10687,N_9739,N_7384);
or U10688 (N_10688,N_8843,N_8725);
or U10689 (N_10689,N_6795,N_5035);
nor U10690 (N_10690,N_9900,N_9106);
or U10691 (N_10691,N_7791,N_8879);
and U10692 (N_10692,N_6980,N_8257);
nand U10693 (N_10693,N_6521,N_7933);
and U10694 (N_10694,N_9341,N_8596);
or U10695 (N_10695,N_8871,N_5758);
nor U10696 (N_10696,N_9587,N_5575);
nor U10697 (N_10697,N_9229,N_9387);
nand U10698 (N_10698,N_8581,N_6532);
or U10699 (N_10699,N_5959,N_5973);
or U10700 (N_10700,N_9662,N_9831);
xnor U10701 (N_10701,N_6761,N_6489);
nand U10702 (N_10702,N_7293,N_6100);
nand U10703 (N_10703,N_7859,N_5891);
nand U10704 (N_10704,N_8712,N_6640);
or U10705 (N_10705,N_9686,N_5606);
and U10706 (N_10706,N_7258,N_6275);
nand U10707 (N_10707,N_5819,N_6880);
nor U10708 (N_10708,N_9032,N_5595);
or U10709 (N_10709,N_5939,N_9541);
or U10710 (N_10710,N_5680,N_8241);
and U10711 (N_10711,N_9825,N_6809);
or U10712 (N_10712,N_8186,N_8420);
and U10713 (N_10713,N_6032,N_9694);
or U10714 (N_10714,N_7554,N_6988);
nor U10715 (N_10715,N_5256,N_6331);
nand U10716 (N_10716,N_9342,N_6857);
nand U10717 (N_10717,N_9816,N_6130);
or U10718 (N_10718,N_5302,N_9510);
nor U10719 (N_10719,N_5076,N_7070);
nor U10720 (N_10720,N_6211,N_6191);
nor U10721 (N_10721,N_9562,N_5797);
nand U10722 (N_10722,N_9881,N_7535);
nand U10723 (N_10723,N_8349,N_8060);
or U10724 (N_10724,N_7726,N_8924);
and U10725 (N_10725,N_5229,N_7852);
nand U10726 (N_10726,N_9313,N_8293);
and U10727 (N_10727,N_8224,N_9606);
or U10728 (N_10728,N_5558,N_8466);
or U10729 (N_10729,N_7178,N_9714);
or U10730 (N_10730,N_9279,N_9431);
or U10731 (N_10731,N_5538,N_6892);
nand U10732 (N_10732,N_6474,N_8998);
and U10733 (N_10733,N_6013,N_6678);
and U10734 (N_10734,N_8754,N_9789);
or U10735 (N_10735,N_5685,N_5602);
xor U10736 (N_10736,N_7966,N_7793);
xor U10737 (N_10737,N_8424,N_7108);
nand U10738 (N_10738,N_9318,N_8640);
nand U10739 (N_10739,N_6538,N_7404);
xor U10740 (N_10740,N_8058,N_8205);
nor U10741 (N_10741,N_9162,N_6178);
nor U10742 (N_10742,N_9619,N_7173);
or U10743 (N_10743,N_5533,N_9759);
nand U10744 (N_10744,N_8589,N_6104);
nand U10745 (N_10745,N_6877,N_5385);
xnor U10746 (N_10746,N_5395,N_7548);
nor U10747 (N_10747,N_8630,N_8629);
nor U10748 (N_10748,N_5733,N_8874);
nand U10749 (N_10749,N_6469,N_8281);
nand U10750 (N_10750,N_9467,N_7819);
nor U10751 (N_10751,N_6014,N_7489);
or U10752 (N_10752,N_5757,N_7458);
nand U10753 (N_10753,N_6092,N_6138);
and U10754 (N_10754,N_8760,N_8498);
and U10755 (N_10755,N_6607,N_8445);
nor U10756 (N_10756,N_6985,N_5273);
nand U10757 (N_10757,N_6478,N_5147);
and U10758 (N_10758,N_8179,N_5600);
or U10759 (N_10759,N_8696,N_7076);
nand U10760 (N_10760,N_5163,N_5669);
nor U10761 (N_10761,N_5514,N_7481);
xor U10762 (N_10762,N_7926,N_9183);
nand U10763 (N_10763,N_7363,N_8598);
nand U10764 (N_10764,N_5077,N_9419);
xnor U10765 (N_10765,N_5148,N_8348);
or U10766 (N_10766,N_5063,N_9488);
or U10767 (N_10767,N_7824,N_6815);
nand U10768 (N_10768,N_6953,N_6340);
nor U10769 (N_10769,N_6322,N_5210);
nor U10770 (N_10770,N_8800,N_5409);
or U10771 (N_10771,N_9607,N_9339);
xnor U10772 (N_10772,N_5078,N_6654);
nor U10773 (N_10773,N_5748,N_6930);
or U10774 (N_10774,N_8273,N_8002);
or U10775 (N_10775,N_5657,N_7992);
or U10776 (N_10776,N_6190,N_9154);
and U10777 (N_10777,N_6660,N_6088);
nand U10778 (N_10778,N_9852,N_8426);
nor U10779 (N_10779,N_9076,N_9613);
nor U10780 (N_10780,N_9550,N_6000);
nor U10781 (N_10781,N_8717,N_8425);
nor U10782 (N_10782,N_9885,N_8789);
nand U10783 (N_10783,N_9961,N_8242);
nand U10784 (N_10784,N_7919,N_5784);
nor U10785 (N_10785,N_9970,N_9080);
nand U10786 (N_10786,N_6979,N_9225);
or U10787 (N_10787,N_8576,N_9202);
nand U10788 (N_10788,N_9114,N_7955);
or U10789 (N_10789,N_9747,N_7860);
nand U10790 (N_10790,N_5755,N_6163);
and U10791 (N_10791,N_7001,N_5114);
nor U10792 (N_10792,N_5336,N_9040);
nor U10793 (N_10793,N_8862,N_6443);
or U10794 (N_10794,N_6732,N_8126);
or U10795 (N_10795,N_5213,N_6545);
or U10796 (N_10796,N_8039,N_6411);
xor U10797 (N_10797,N_6571,N_5979);
nand U10798 (N_10798,N_8892,N_5905);
nor U10799 (N_10799,N_5295,N_7823);
and U10800 (N_10800,N_8218,N_8770);
and U10801 (N_10801,N_9719,N_7485);
nor U10802 (N_10802,N_9898,N_5298);
nor U10803 (N_10803,N_8236,N_9455);
xnor U10804 (N_10804,N_6125,N_5001);
nor U10805 (N_10805,N_9591,N_9722);
xnor U10806 (N_10806,N_5242,N_9669);
and U10807 (N_10807,N_8907,N_5420);
nand U10808 (N_10808,N_9828,N_8121);
or U10809 (N_10809,N_8291,N_5759);
or U10810 (N_10810,N_8713,N_8950);
nand U10811 (N_10811,N_6203,N_8516);
or U10812 (N_10812,N_7171,N_9068);
xor U10813 (N_10813,N_9509,N_5581);
or U10814 (N_10814,N_6102,N_6889);
or U10815 (N_10815,N_6318,N_5625);
and U10816 (N_10816,N_5536,N_8297);
nand U10817 (N_10817,N_6754,N_7880);
nand U10818 (N_10818,N_9756,N_7952);
and U10819 (N_10819,N_9060,N_7284);
nand U10820 (N_10820,N_8608,N_7593);
nand U10821 (N_10821,N_5016,N_5895);
or U10822 (N_10822,N_5389,N_8914);
xnor U10823 (N_10823,N_7835,N_9827);
or U10824 (N_10824,N_9350,N_8787);
and U10825 (N_10825,N_9501,N_8030);
xor U10826 (N_10826,N_6989,N_9710);
or U10827 (N_10827,N_8738,N_6458);
nand U10828 (N_10828,N_9457,N_5331);
or U10829 (N_10829,N_9182,N_5972);
and U10830 (N_10830,N_5580,N_5739);
nand U10831 (N_10831,N_8517,N_9723);
xor U10832 (N_10832,N_6356,N_5056);
xor U10833 (N_10833,N_8220,N_6295);
nor U10834 (N_10834,N_6615,N_6231);
nand U10835 (N_10835,N_7811,N_6639);
nor U10836 (N_10836,N_8481,N_5086);
xor U10837 (N_10837,N_8618,N_9809);
nand U10838 (N_10838,N_5999,N_6071);
nor U10839 (N_10839,N_8727,N_6870);
and U10840 (N_10840,N_6038,N_7152);
nor U10841 (N_10841,N_7889,N_7541);
nand U10842 (N_10842,N_7621,N_9832);
nand U10843 (N_10843,N_8035,N_9297);
and U10844 (N_10844,N_7425,N_6964);
nand U10845 (N_10845,N_9805,N_8407);
nor U10846 (N_10846,N_9099,N_9396);
nand U10847 (N_10847,N_8723,N_6164);
or U10848 (N_10848,N_5456,N_8837);
nor U10849 (N_10849,N_7922,N_7733);
and U10850 (N_10850,N_9748,N_5688);
and U10851 (N_10851,N_5612,N_5629);
nor U10852 (N_10852,N_9919,N_8098);
and U10853 (N_10853,N_8878,N_5938);
nand U10854 (N_10854,N_9415,N_6131);
nand U10855 (N_10855,N_6796,N_8125);
nand U10856 (N_10856,N_8370,N_7609);
and U10857 (N_10857,N_9764,N_7812);
and U10858 (N_10858,N_9609,N_5749);
or U10859 (N_10859,N_7981,N_7866);
nand U10860 (N_10860,N_6664,N_9094);
nand U10861 (N_10861,N_9625,N_9141);
and U10862 (N_10862,N_7775,N_8099);
or U10863 (N_10863,N_6377,N_5427);
or U10864 (N_10864,N_5703,N_6832);
nor U10865 (N_10865,N_7349,N_9532);
nor U10866 (N_10866,N_6762,N_5415);
or U10867 (N_10867,N_5777,N_7545);
and U10868 (N_10868,N_9325,N_6245);
or U10869 (N_10869,N_7222,N_7137);
or U10870 (N_10870,N_8418,N_6810);
and U10871 (N_10871,N_7361,N_5458);
nand U10872 (N_10872,N_6249,N_8356);
xnor U10873 (N_10873,N_7958,N_7858);
nand U10874 (N_10874,N_7920,N_8553);
nand U10875 (N_10875,N_9763,N_8267);
or U10876 (N_10876,N_6848,N_9494);
nor U10877 (N_10877,N_7473,N_6908);
nand U10878 (N_10878,N_8755,N_9688);
nand U10879 (N_10879,N_5054,N_8470);
or U10880 (N_10880,N_7753,N_5579);
or U10881 (N_10881,N_5645,N_5238);
nand U10882 (N_10882,N_8665,N_9880);
nor U10883 (N_10883,N_7507,N_9192);
and U10884 (N_10884,N_6412,N_6725);
nand U10885 (N_10885,N_8353,N_8097);
nand U10886 (N_10886,N_7028,N_8288);
or U10887 (N_10887,N_9287,N_6004);
nor U10888 (N_10888,N_5734,N_9946);
xnor U10889 (N_10889,N_9681,N_5928);
or U10890 (N_10890,N_6099,N_5027);
nor U10891 (N_10891,N_8328,N_6776);
or U10892 (N_10892,N_6799,N_8521);
nor U10893 (N_10893,N_5542,N_9716);
and U10894 (N_10894,N_5554,N_8469);
nand U10895 (N_10895,N_5351,N_8040);
xnor U10896 (N_10896,N_8554,N_6220);
nor U10897 (N_10897,N_6526,N_8479);
nor U10898 (N_10898,N_9024,N_6805);
nor U10899 (N_10899,N_8901,N_9521);
xnor U10900 (N_10900,N_5386,N_6548);
nor U10901 (N_10901,N_8559,N_8626);
or U10902 (N_10902,N_8776,N_6927);
and U10903 (N_10903,N_8556,N_8542);
or U10904 (N_10904,N_7213,N_7737);
nand U10905 (N_10905,N_5058,N_5358);
nor U10906 (N_10906,N_6008,N_5008);
nor U10907 (N_10907,N_6064,N_8580);
or U10908 (N_10908,N_6086,N_5997);
or U10909 (N_10909,N_6680,N_6233);
or U10910 (N_10910,N_8246,N_9132);
nand U10911 (N_10911,N_7064,N_6380);
or U10912 (N_10912,N_9376,N_7089);
or U10913 (N_10913,N_5803,N_8460);
or U10914 (N_10914,N_8652,N_5987);
nand U10915 (N_10915,N_6352,N_6861);
nand U10916 (N_10916,N_6108,N_9718);
nor U10917 (N_10917,N_7884,N_9427);
and U10918 (N_10918,N_9818,N_7462);
and U10919 (N_10919,N_9301,N_8557);
nor U10920 (N_10920,N_5102,N_6449);
nand U10921 (N_10921,N_9357,N_5790);
or U10922 (N_10922,N_7146,N_5670);
or U10923 (N_10923,N_9814,N_9634);
or U10924 (N_10924,N_5157,N_5808);
and U10925 (N_10925,N_7680,N_9096);
nor U10926 (N_10926,N_8594,N_8913);
or U10927 (N_10927,N_5112,N_7526);
or U10928 (N_10928,N_5467,N_7296);
nor U10929 (N_10929,N_5193,N_5472);
or U10930 (N_10930,N_9030,N_8255);
or U10931 (N_10931,N_9702,N_5714);
nor U10932 (N_10932,N_7707,N_6994);
nor U10933 (N_10933,N_5974,N_7887);
nor U10934 (N_10934,N_5800,N_8784);
nand U10935 (N_10935,N_9360,N_8315);
xnor U10936 (N_10936,N_9198,N_9563);
or U10937 (N_10937,N_8587,N_8747);
nand U10938 (N_10938,N_9704,N_8806);
or U10939 (N_10939,N_6788,N_8586);
and U10940 (N_10940,N_8722,N_8773);
and U10941 (N_10941,N_9354,N_7106);
or U10942 (N_10942,N_9017,N_8585);
nor U10943 (N_10943,N_5713,N_8966);
xnor U10944 (N_10944,N_5452,N_9560);
and U10945 (N_10945,N_8122,N_7232);
nand U10946 (N_10946,N_8724,N_9237);
nor U10947 (N_10947,N_6143,N_7094);
nand U10948 (N_10948,N_5642,N_9594);
nand U10949 (N_10949,N_9940,N_6853);
nand U10950 (N_10950,N_6780,N_9343);
xnor U10951 (N_10951,N_8452,N_7979);
and U10952 (N_10952,N_7385,N_5244);
or U10953 (N_10953,N_9819,N_8639);
nand U10954 (N_10954,N_8728,N_7639);
nand U10955 (N_10955,N_5187,N_6733);
or U10956 (N_10956,N_7755,N_9700);
xnor U10957 (N_10957,N_6259,N_6437);
nand U10958 (N_10958,N_7888,N_9971);
nand U10959 (N_10959,N_8474,N_9196);
nor U10960 (N_10960,N_8658,N_5668);
nand U10961 (N_10961,N_8938,N_6613);
and U10962 (N_10962,N_6005,N_7854);
and U10963 (N_10963,N_8663,N_5862);
nor U10964 (N_10964,N_7465,N_5178);
or U10965 (N_10965,N_6427,N_5543);
or U10966 (N_10966,N_6970,N_9288);
or U10967 (N_10967,N_6743,N_7459);
nand U10968 (N_10968,N_6618,N_6127);
nor U10969 (N_10969,N_5357,N_6201);
or U10970 (N_10970,N_5827,N_5694);
xnor U10971 (N_10971,N_6579,N_8935);
or U10972 (N_10972,N_8614,N_6828);
nand U10973 (N_10973,N_9321,N_8214);
xnor U10974 (N_10974,N_9272,N_5199);
and U10975 (N_10975,N_9250,N_8084);
nand U10976 (N_10976,N_6291,N_7120);
or U10977 (N_10977,N_9643,N_9048);
and U10978 (N_10978,N_8053,N_5949);
xnor U10979 (N_10979,N_9660,N_7026);
or U10980 (N_10980,N_9187,N_8141);
nor U10981 (N_10981,N_8169,N_6386);
nor U10982 (N_10982,N_9020,N_8822);
or U10983 (N_10983,N_6124,N_9004);
xnor U10984 (N_10984,N_8633,N_9945);
and U10985 (N_10985,N_8270,N_6656);
nand U10986 (N_10986,N_5447,N_7257);
nor U10987 (N_10987,N_8310,N_8561);
xnor U10988 (N_10988,N_7575,N_6708);
and U10989 (N_10989,N_5263,N_8720);
and U10990 (N_10990,N_8583,N_8790);
and U10991 (N_10991,N_7873,N_5234);
or U10992 (N_10992,N_7062,N_5424);
nor U10993 (N_10993,N_5735,N_5141);
nor U10994 (N_10994,N_5416,N_8961);
or U10995 (N_10995,N_9934,N_6268);
nor U10996 (N_10996,N_8379,N_7713);
nand U10997 (N_10997,N_8385,N_9559);
nand U10998 (N_10998,N_6928,N_9884);
nor U10999 (N_10999,N_6710,N_9456);
or U11000 (N_11000,N_5744,N_6120);
or U11001 (N_11001,N_6087,N_8795);
or U11002 (N_11002,N_7233,N_6763);
xor U11003 (N_11003,N_6556,N_6090);
nand U11004 (N_11004,N_5531,N_9189);
and U11005 (N_11005,N_5101,N_5317);
nor U11006 (N_11006,N_7374,N_7405);
and U11007 (N_11007,N_7295,N_6076);
or U11008 (N_11008,N_6765,N_7907);
and U11009 (N_11009,N_5050,N_6272);
nor U11010 (N_11010,N_7790,N_7795);
or U11011 (N_11011,N_9938,N_8296);
and U11012 (N_11012,N_6026,N_7551);
xnor U11013 (N_11013,N_5555,N_8893);
and U11014 (N_11014,N_5515,N_5470);
or U11015 (N_11015,N_5320,N_5173);
nand U11016 (N_11016,N_8688,N_9974);
xnor U11017 (N_11017,N_6842,N_9033);
nand U11018 (N_11018,N_6914,N_6974);
nand U11019 (N_11019,N_7219,N_6931);
nand U11020 (N_11020,N_7021,N_5397);
or U11021 (N_11021,N_5523,N_5540);
or U11022 (N_11022,N_9912,N_9735);
nor U11023 (N_11023,N_6806,N_8320);
or U11024 (N_11024,N_6369,N_8451);
or U11025 (N_11025,N_7338,N_6224);
nor U11026 (N_11026,N_8880,N_5497);
nor U11027 (N_11027,N_9403,N_7806);
or U11028 (N_11028,N_8846,N_7235);
xnor U11029 (N_11029,N_7643,N_9166);
or U11030 (N_11030,N_5552,N_8312);
nor U11031 (N_11031,N_6497,N_7126);
and U11032 (N_11032,N_8532,N_8563);
nor U11033 (N_11033,N_7878,N_8490);
or U11034 (N_11034,N_5136,N_6757);
nor U11035 (N_11035,N_6081,N_5232);
nor U11036 (N_11036,N_9101,N_7751);
or U11037 (N_11037,N_5209,N_9109);
and U11038 (N_11038,N_9720,N_5471);
nor U11039 (N_11039,N_5422,N_9191);
or U11040 (N_11040,N_7181,N_7894);
or U11041 (N_11041,N_6053,N_5304);
or U11042 (N_11042,N_6292,N_7647);
nor U11043 (N_11043,N_6894,N_8086);
nor U11044 (N_11044,N_5893,N_8551);
nand U11045 (N_11045,N_8753,N_5153);
xor U11046 (N_11046,N_6915,N_7718);
or U11047 (N_11047,N_6444,N_5066);
nand U11048 (N_11048,N_5407,N_8891);
and U11049 (N_11049,N_8196,N_6898);
nor U11050 (N_11050,N_8087,N_7638);
nand U11051 (N_11051,N_5116,N_7653);
nand U11052 (N_11052,N_5200,N_9600);
nand U11053 (N_11053,N_9676,N_9602);
xor U11054 (N_11054,N_6457,N_8958);
and U11055 (N_11055,N_9491,N_6991);
and U11056 (N_11056,N_8780,N_7587);
and U11057 (N_11057,N_7475,N_8061);
or U11058 (N_11058,N_5942,N_9116);
or U11059 (N_11059,N_5046,N_5207);
and U11060 (N_11060,N_5594,N_5894);
or U11061 (N_11061,N_9911,N_7466);
and U11062 (N_11062,N_6887,N_7248);
or U11063 (N_11063,N_9776,N_6311);
xor U11064 (N_11064,N_5484,N_6112);
nor U11065 (N_11065,N_5751,N_8307);
nand U11066 (N_11066,N_6117,N_6273);
and U11067 (N_11067,N_9348,N_6531);
nor U11068 (N_11068,N_8887,N_5836);
or U11069 (N_11069,N_9699,N_8750);
nand U11070 (N_11070,N_6401,N_6864);
or U11071 (N_11071,N_8990,N_6749);
xnor U11072 (N_11072,N_6911,N_8301);
and U11073 (N_11073,N_5583,N_9471);
nand U11074 (N_11074,N_5237,N_5044);
nand U11075 (N_11075,N_8994,N_6730);
nand U11076 (N_11076,N_8101,N_9793);
nand U11077 (N_11077,N_5760,N_9893);
nor U11078 (N_11078,N_9942,N_9465);
and U11079 (N_11079,N_7163,N_9428);
nand U11080 (N_11080,N_6909,N_5087);
and U11081 (N_11081,N_7836,N_8109);
or U11082 (N_11082,N_6646,N_8852);
nand U11083 (N_11083,N_8657,N_9205);
and U11084 (N_11084,N_7455,N_8858);
nand U11085 (N_11085,N_5075,N_7035);
or U11086 (N_11086,N_7198,N_7759);
nand U11087 (N_11087,N_9355,N_6069);
and U11088 (N_11088,N_6872,N_8290);
nor U11089 (N_11089,N_9601,N_8079);
xnor U11090 (N_11090,N_5125,N_5194);
or U11091 (N_11091,N_9243,N_5296);
or U11092 (N_11092,N_8791,N_7924);
nor U11093 (N_11093,N_9558,N_9863);
or U11094 (N_11094,N_6782,N_5553);
nor U11095 (N_11095,N_7616,N_6530);
and U11096 (N_11096,N_7496,N_9973);
nor U11097 (N_11097,N_7596,N_5560);
nand U11098 (N_11098,N_7869,N_8974);
and U11099 (N_11099,N_8573,N_8751);
nor U11100 (N_11100,N_8417,N_7074);
and U11101 (N_11101,N_6051,N_9965);
or U11102 (N_11102,N_5885,N_6206);
or U11103 (N_11103,N_8212,N_6016);
nand U11104 (N_11104,N_8772,N_5239);
nand U11105 (N_11105,N_7603,N_5278);
or U11106 (N_11106,N_6591,N_8671);
or U11107 (N_11107,N_9380,N_5728);
nor U11108 (N_11108,N_6826,N_7103);
nor U11109 (N_11109,N_6758,N_7696);
and U11110 (N_11110,N_9705,N_8413);
nand U11111 (N_11111,N_5493,N_5911);
and U11112 (N_11112,N_7515,N_5822);
or U11113 (N_11113,N_8019,N_6286);
and U11114 (N_11114,N_5923,N_9812);
nor U11115 (N_11115,N_7993,N_5994);
nor U11116 (N_11116,N_8515,N_7560);
or U11117 (N_11117,N_7084,N_5444);
and U11118 (N_11118,N_7969,N_6459);
or U11119 (N_11119,N_6929,N_5010);
and U11120 (N_11120,N_8799,N_9975);
and U11121 (N_11121,N_5705,N_6057);
nor U11122 (N_11122,N_6650,N_7841);
nand U11123 (N_11123,N_5253,N_5897);
and U11124 (N_11124,N_9157,N_6675);
xor U11125 (N_11125,N_6303,N_7681);
or U11126 (N_11126,N_9623,N_7683);
or U11127 (N_11127,N_5665,N_9869);
nor U11128 (N_11128,N_5335,N_6936);
or U11129 (N_11129,N_7710,N_5146);
nand U11130 (N_11130,N_5494,N_5812);
and U11131 (N_11131,N_5823,N_6651);
and U11132 (N_11132,N_8178,N_5940);
or U11133 (N_11133,N_8689,N_6939);
nor U11134 (N_11134,N_7169,N_6263);
and U11135 (N_11135,N_7829,N_9356);
nor U11136 (N_11136,N_5469,N_9954);
nor U11137 (N_11137,N_7788,N_8287);
xor U11138 (N_11138,N_5562,N_8016);
nor U11139 (N_11139,N_7464,N_9171);
nand U11140 (N_11140,N_7636,N_5610);
nor U11141 (N_11141,N_7960,N_5220);
nor U11142 (N_11142,N_7532,N_8934);
and U11143 (N_11143,N_8361,N_8465);
xor U11144 (N_11144,N_6455,N_6649);
nor U11145 (N_11145,N_6154,N_6494);
nand U11146 (N_11146,N_7167,N_8812);
nor U11147 (N_11147,N_5111,N_5650);
nand U11148 (N_11148,N_6355,N_7063);
nor U11149 (N_11149,N_6399,N_8237);
nand U11150 (N_11150,N_7127,N_9316);
nor U11151 (N_11151,N_7769,N_7416);
nor U11152 (N_11152,N_6232,N_5216);
and U11153 (N_11153,N_7487,N_8505);
nor U11154 (N_11154,N_8455,N_5325);
or U11155 (N_11155,N_6772,N_5850);
nand U11156 (N_11156,N_9131,N_7523);
and U11157 (N_11157,N_8719,N_8835);
nor U11158 (N_11158,N_8072,N_7959);
nand U11159 (N_11159,N_7215,N_6415);
and U11160 (N_11160,N_5479,N_7728);
nor U11161 (N_11161,N_9309,N_8368);
or U11162 (N_11162,N_5231,N_8051);
nand U11163 (N_11163,N_8697,N_9835);
or U11164 (N_11164,N_6933,N_8289);
and U11165 (N_11165,N_8037,N_6236);
and U11166 (N_11166,N_6841,N_5563);
nor U11167 (N_11167,N_9762,N_5864);
nand U11168 (N_11168,N_8162,N_5039);
or U11169 (N_11169,N_9939,N_5955);
and U11170 (N_11170,N_7659,N_7119);
and U11171 (N_11171,N_7482,N_6653);
or U11172 (N_11172,N_7516,N_6720);
and U11173 (N_11173,N_7657,N_9583);
nor U11174 (N_11174,N_9382,N_7577);
nand U11175 (N_11175,N_8952,N_5384);
nand U11176 (N_11176,N_7399,N_8898);
and U11177 (N_11177,N_7088,N_8518);
xor U11178 (N_11178,N_6152,N_9599);
or U11179 (N_11179,N_5953,N_8180);
and U11180 (N_11180,N_5785,N_9866);
nand U11181 (N_11181,N_7027,N_5095);
and U11182 (N_11182,N_6851,N_8213);
and U11183 (N_11183,N_7149,N_8050);
nand U11184 (N_11184,N_5380,N_9349);
nand U11185 (N_11185,N_6098,N_5350);
or U11186 (N_11186,N_8473,N_5962);
or U11187 (N_11187,N_8017,N_7386);
nor U11188 (N_11188,N_9542,N_9561);
or U11189 (N_11189,N_8670,N_6450);
and U11190 (N_11190,N_5985,N_5852);
or U11191 (N_11191,N_7319,N_9984);
nand U11192 (N_11192,N_9682,N_7005);
xor U11193 (N_11193,N_9654,N_6945);
nand U11194 (N_11194,N_5503,N_6535);
or U11195 (N_11195,N_8376,N_9074);
xnor U11196 (N_11196,N_7382,N_8280);
or U11197 (N_11197,N_6375,N_8807);
nand U11198 (N_11198,N_9994,N_6199);
nor U11199 (N_11199,N_9646,N_8906);
xor U11200 (N_11200,N_7559,N_8369);
nand U11201 (N_11201,N_5909,N_6666);
nor U11202 (N_11202,N_7267,N_7573);
xnor U11203 (N_11203,N_6717,N_7043);
or U11204 (N_11204,N_8329,N_8263);
nand U11205 (N_11205,N_9618,N_5402);
nor U11206 (N_11206,N_7986,N_5000);
or U11207 (N_11207,N_7561,N_9761);
nand U11208 (N_11208,N_8954,N_8358);
or U11209 (N_11209,N_5952,N_8052);
nand U11210 (N_11210,N_6333,N_9139);
and U11211 (N_11211,N_8384,N_8979);
and U11212 (N_11212,N_6153,N_6490);
and U11213 (N_11213,N_8783,N_6838);
xor U11214 (N_11214,N_7265,N_9833);
and U11215 (N_11215,N_7114,N_8764);
nand U11216 (N_11216,N_6062,N_5720);
nor U11217 (N_11217,N_5123,N_5372);
or U11218 (N_11218,N_5104,N_7446);
nand U11219 (N_11219,N_9312,N_7618);
and U11220 (N_11220,N_6023,N_9441);
or U11221 (N_11221,N_9540,N_9072);
or U11222 (N_11222,N_9696,N_6922);
xor U11223 (N_11223,N_5828,N_8829);
nand U11224 (N_11224,N_5585,N_9913);
and U11225 (N_11225,N_9595,N_5608);
nand U11226 (N_11226,N_6198,N_7128);
or U11227 (N_11227,N_5341,N_9340);
and U11228 (N_11228,N_6800,N_9556);
xnor U11229 (N_11229,N_6783,N_6073);
nor U11230 (N_11230,N_9090,N_5332);
xnor U11231 (N_11231,N_9421,N_6818);
and U11232 (N_11232,N_9555,N_9344);
nand U11233 (N_11233,N_5613,N_7347);
or U11234 (N_11234,N_6850,N_7699);
nand U11235 (N_11235,N_5906,N_8539);
nor U11236 (N_11236,N_8450,N_6669);
xnor U11237 (N_11237,N_6821,N_7393);
and U11238 (N_11238,N_5567,N_6445);
nor U11239 (N_11239,N_8201,N_5883);
nand U11240 (N_11240,N_8552,N_9407);
nand U11241 (N_11241,N_6903,N_5519);
nor U11242 (N_11242,N_9215,N_7805);
or U11243 (N_11243,N_6501,N_6349);
and U11244 (N_11244,N_8931,N_8217);
or U11245 (N_11245,N_7183,N_9001);
xnor U11246 (N_11246,N_9679,N_9506);
nor U11247 (N_11247,N_5014,N_8046);
and U11248 (N_11248,N_6134,N_7654);
nor U11249 (N_11249,N_9173,N_9174);
or U11250 (N_11250,N_7153,N_7082);
or U11251 (N_11251,N_6969,N_8555);
and U11252 (N_11252,N_8282,N_8698);
or U11253 (N_11253,N_9061,N_8311);
nor U11254 (N_11254,N_5423,N_9334);
and U11255 (N_11255,N_5226,N_5106);
nand U11256 (N_11256,N_9468,N_7061);
nor U11257 (N_11257,N_9960,N_5099);
and U11258 (N_11258,N_9890,N_8989);
or U11259 (N_11259,N_8117,N_9148);
or U11260 (N_11260,N_5653,N_9514);
nand U11261 (N_11261,N_9572,N_9200);
nor U11262 (N_11262,N_8195,N_5513);
or U11263 (N_11263,N_6992,N_8433);
nand U11264 (N_11264,N_8323,N_9906);
nor U11265 (N_11265,N_5903,N_8223);
and U11266 (N_11266,N_6376,N_9300);
and U11267 (N_11267,N_7037,N_7228);
and U11268 (N_11268,N_7073,N_6358);
and U11269 (N_11269,N_9102,N_7943);
and U11270 (N_11270,N_9768,N_6812);
nor U11271 (N_11271,N_7421,N_8423);
and U11272 (N_11272,N_9760,N_5313);
nor U11273 (N_11273,N_9539,N_8792);
nor U11274 (N_11274,N_8443,N_6797);
nor U11275 (N_11275,N_8226,N_5995);
nand U11276 (N_11276,N_6496,N_5743);
nor U11277 (N_11277,N_9876,N_8940);
nand U11278 (N_11278,N_8674,N_5958);
and U11279 (N_11279,N_5221,N_5574);
nand U11280 (N_11280,N_5191,N_6031);
or U11281 (N_11281,N_9861,N_8546);
and U11282 (N_11282,N_5487,N_8983);
or U11283 (N_11283,N_5391,N_5804);
and U11284 (N_11284,N_5333,N_9274);
or U11285 (N_11285,N_5920,N_8992);
or U11286 (N_11286,N_5990,N_8972);
or U11287 (N_11287,N_8192,N_8883);
and U11288 (N_11288,N_9227,N_8360);
nand U11289 (N_11289,N_6508,N_5224);
nor U11290 (N_11290,N_6343,N_6852);
xor U11291 (N_11291,N_9990,N_6320);
or U11292 (N_11292,N_9851,N_5085);
nand U11293 (N_11293,N_8656,N_9743);
and U11294 (N_11294,N_6095,N_8047);
xnor U11295 (N_11295,N_7809,N_5666);
and U11296 (N_11296,N_7735,N_6218);
xor U11297 (N_11297,N_7565,N_8005);
nor U11298 (N_11298,N_5120,N_7134);
nand U11299 (N_11299,N_8285,N_6260);
nor U11300 (N_11300,N_5068,N_9372);
nor U11301 (N_11301,N_9329,N_6997);
and U11302 (N_11302,N_7440,N_5449);
and U11303 (N_11303,N_9774,N_6440);
and U11304 (N_11304,N_7527,N_8003);
or U11305 (N_11305,N_9637,N_9119);
nand U11306 (N_11306,N_7083,N_9821);
or U11307 (N_11307,N_8786,N_9765);
and U11308 (N_11308,N_9498,N_5110);
or U11309 (N_11309,N_6294,N_5442);
nand U11310 (N_11310,N_6588,N_7367);
and U11311 (N_11311,N_8809,N_8411);
or U11312 (N_11312,N_7049,N_9152);
nor U11313 (N_11313,N_6434,N_6219);
or U11314 (N_11314,N_6803,N_8529);
nand U11315 (N_11315,N_8911,N_6682);
nor U11316 (N_11316,N_7427,N_6638);
nor U11317 (N_11317,N_8298,N_9149);
or U11318 (N_11318,N_8390,N_5107);
or U11319 (N_11319,N_5766,N_6723);
and U11320 (N_11320,N_7433,N_6559);
xor U11321 (N_11321,N_6961,N_6467);
or U11322 (N_11322,N_5556,N_8181);
nand U11323 (N_11323,N_8080,N_9414);
nand U11324 (N_11324,N_7214,N_8245);
nor U11325 (N_11325,N_8923,N_9840);
and U11326 (N_11326,N_5400,N_9397);
xnor U11327 (N_11327,N_7397,N_6916);
nor U11328 (N_11328,N_5877,N_6256);
and U11329 (N_11329,N_7143,N_7375);
or U11330 (N_11330,N_8678,N_8895);
nor U11331 (N_11331,N_8193,N_6247);
and U11332 (N_11332,N_8113,N_8104);
nor U11333 (N_11333,N_6901,N_7580);
and U11334 (N_11334,N_7717,N_8654);
xnor U11335 (N_11335,N_6512,N_7444);
or U11336 (N_11336,N_8682,N_9689);
and U11337 (N_11337,N_9206,N_5868);
nand U11338 (N_11338,N_6600,N_7493);
or U11339 (N_11339,N_9892,N_9395);
or U11340 (N_11340,N_8206,N_6306);
and U11341 (N_11341,N_5809,N_7848);
and U11342 (N_11342,N_7372,N_7086);
nand U11343 (N_11343,N_9430,N_8152);
nand U11344 (N_11344,N_6481,N_5217);
and U11345 (N_11345,N_6149,N_9864);
or U11346 (N_11346,N_8993,N_5584);
nand U11347 (N_11347,N_5206,N_7766);
xor U11348 (N_11348,N_7140,N_5434);
nand U11349 (N_11349,N_5963,N_8164);
xnor U11350 (N_11350,N_9740,N_6580);
and U11351 (N_11351,N_9063,N_6718);
nor U11352 (N_11352,N_8197,N_8959);
xor U11353 (N_11353,N_6040,N_9734);
nor U11354 (N_11354,N_7175,N_9423);
nor U11355 (N_11355,N_7289,N_8059);
xnor U11356 (N_11356,N_5290,N_8980);
nand U11357 (N_11357,N_5222,N_8769);
or U11358 (N_11358,N_9234,N_6599);
nand U11359 (N_11359,N_7916,N_5108);
nor U11360 (N_11360,N_6432,N_7716);
nand U11361 (N_11361,N_9390,N_9474);
nor U11362 (N_11362,N_5024,N_6867);
xnor U11363 (N_11363,N_5816,N_5012);
nor U11364 (N_11364,N_8114,N_5649);
or U11365 (N_11365,N_6363,N_9104);
nor U11366 (N_11366,N_5887,N_9044);
nand U11367 (N_11367,N_5931,N_8830);
nand U11368 (N_11368,N_7343,N_9697);
nand U11369 (N_11369,N_7644,N_8137);
xor U11370 (N_11370,N_7970,N_7392);
nor U11371 (N_11371,N_6644,N_9551);
nor U11372 (N_11372,N_7221,N_7413);
nand U11373 (N_11373,N_9437,N_9841);
and U11374 (N_11374,N_6461,N_8190);
nand U11375 (N_11375,N_9622,N_5867);
and U11376 (N_11376,N_8591,N_9608);
and U11377 (N_11377,N_6871,N_7160);
and U11378 (N_11378,N_5437,N_8215);
nand U11379 (N_11379,N_8584,N_5914);
or U11380 (N_11380,N_7471,N_7668);
or U11381 (N_11381,N_6876,N_7217);
nand U11382 (N_11382,N_8886,N_8824);
nor U11383 (N_11383,N_7488,N_7156);
nand U11384 (N_11384,N_6802,N_9087);
nor U11385 (N_11385,N_6539,N_7709);
or U11386 (N_11386,N_7281,N_5029);
nor U11387 (N_11387,N_5227,N_7885);
and U11388 (N_11388,N_6093,N_7139);
or U11389 (N_11389,N_7815,N_6402);
or U11390 (N_11390,N_9472,N_7895);
and U11391 (N_11391,N_6910,N_9655);
nor U11392 (N_11392,N_5377,N_9981);
xor U11393 (N_11393,N_5266,N_7057);
nor U11394 (N_11394,N_5064,N_5183);
or U11395 (N_11395,N_7158,N_7932);
nand U11396 (N_11396,N_7945,N_8023);
or U11397 (N_11397,N_7827,N_9281);
nand U11398 (N_11398,N_9665,N_7906);
nand U11399 (N_11399,N_7451,N_6417);
or U11400 (N_11400,N_7905,N_6557);
and U11401 (N_11401,N_7510,N_8625);
nand U11402 (N_11402,N_7513,N_6920);
and U11403 (N_11403,N_8441,N_9400);
nand U11404 (N_11404,N_6959,N_5142);
nand U11405 (N_11405,N_7941,N_6751);
nand U11406 (N_11406,N_8074,N_8144);
or U11407 (N_11407,N_9278,N_9117);
nor U11408 (N_11408,N_7632,N_5898);
and U11409 (N_11409,N_6612,N_6185);
or U11410 (N_11410,N_9185,N_9255);
nor U11411 (N_11411,N_8313,N_6170);
or U11412 (N_11412,N_5300,N_9553);
nor U11413 (N_11413,N_5892,N_6699);
nand U11414 (N_11414,N_5432,N_6324);
nand U11415 (N_11415,N_6351,N_5838);
or U11416 (N_11416,N_7452,N_9290);
or U11417 (N_11417,N_7400,N_7937);
xnor U11418 (N_11418,N_9327,N_6276);
xor U11419 (N_11419,N_9304,N_8386);
and U11420 (N_11420,N_9846,N_6338);
or U11421 (N_11421,N_5932,N_9633);
and U11422 (N_11422,N_8611,N_9388);
and U11423 (N_11423,N_5499,N_5446);
and U11424 (N_11424,N_8000,N_5524);
or U11425 (N_11425,N_9692,N_8480);
and U11426 (N_11426,N_7754,N_9617);
xnor U11427 (N_11427,N_9879,N_9728);
xnor U11428 (N_11428,N_9582,N_6523);
and U11429 (N_11429,N_6900,N_9347);
nand U11430 (N_11430,N_8429,N_9257);
or U11431 (N_11431,N_6534,N_5279);
nand U11432 (N_11432,N_7525,N_6906);
or U11433 (N_11433,N_6084,N_8127);
nor U11434 (N_11434,N_7401,N_7929);
xnor U11435 (N_11435,N_6735,N_9635);
or U11436 (N_11436,N_5884,N_6724);
and U11437 (N_11437,N_5530,N_5363);
or U11438 (N_11438,N_6407,N_5712);
nor U11439 (N_11439,N_9322,N_7009);
xor U11440 (N_11440,N_5726,N_6817);
or U11441 (N_11441,N_7196,N_7739);
nand U11442 (N_11442,N_9589,N_7534);
nand U11443 (N_11443,N_6468,N_8506);
xor U11444 (N_11444,N_6942,N_8012);
nand U11445 (N_11445,N_6202,N_7069);
or U11446 (N_11446,N_9811,N_6657);
or U11447 (N_11447,N_9218,N_9978);
and U11448 (N_11448,N_7412,N_5924);
nor U11449 (N_11449,N_5366,N_9586);
nor U11450 (N_11450,N_9712,N_8978);
or U11451 (N_11451,N_9557,N_6315);
or U11452 (N_11452,N_5052,N_7395);
and U11453 (N_11453,N_8899,N_5282);
nor U11454 (N_11454,N_8391,N_9997);
nand U11455 (N_11455,N_7456,N_9476);
or U11456 (N_11456,N_9212,N_7402);
or U11457 (N_11457,N_9446,N_8139);
or U11458 (N_11458,N_6119,N_9259);
nor U11459 (N_11459,N_7467,N_7317);
nor U11460 (N_11460,N_7501,N_9611);
nand U11461 (N_11461,N_5090,N_6510);
or U11462 (N_11462,N_5820,N_9078);
nand U11463 (N_11463,N_9224,N_5088);
or U11464 (N_11464,N_7821,N_5618);
or U11465 (N_11465,N_6243,N_8233);
nand U11466 (N_11466,N_5756,N_6347);
and U11467 (N_11467,N_8419,N_7944);
xor U11468 (N_11468,N_8272,N_5262);
nor U11469 (N_11469,N_7570,N_8286);
xor U11470 (N_11470,N_5872,N_9052);
or U11471 (N_11471,N_9026,N_8653);
nor U11472 (N_11472,N_5988,N_8322);
and U11473 (N_11473,N_9877,N_6570);
nand U11474 (N_11474,N_7697,N_9566);
nand U11475 (N_11475,N_5324,N_5084);
and U11476 (N_11476,N_5750,N_9022);
and U11477 (N_11477,N_5754,N_6068);
xnor U11478 (N_11478,N_8741,N_8200);
xnor U11479 (N_11479,N_7498,N_9482);
and U11480 (N_11480,N_9433,N_8945);
nor U11481 (N_11481,N_7436,N_8011);
or U11482 (N_11482,N_8303,N_7115);
nor U11483 (N_11483,N_7211,N_8844);
xor U11484 (N_11484,N_6673,N_7369);
or U11485 (N_11485,N_7355,N_5083);
nand U11486 (N_11486,N_7886,N_8774);
xnor U11487 (N_11487,N_8672,N_5082);
or U11488 (N_11488,N_7975,N_8679);
xnor U11489 (N_11489,N_7964,N_8252);
nand U11490 (N_11490,N_8477,N_5976);
nor U11491 (N_11491,N_6691,N_9404);
nand U11492 (N_11492,N_6205,N_8211);
and U11493 (N_11493,N_7965,N_7761);
nand U11494 (N_11494,N_6687,N_5203);
and U11495 (N_11495,N_5092,N_9439);
nand U11496 (N_11496,N_6560,N_9909);
and U11497 (N_11497,N_9980,N_9517);
nor U11498 (N_11498,N_6966,N_6890);
nand U11499 (N_11499,N_5788,N_5621);
nand U11500 (N_11500,N_5250,N_6151);
nor U11501 (N_11501,N_5667,N_7315);
and U11502 (N_11502,N_5170,N_7672);
and U11503 (N_11503,N_8565,N_7306);
and U11504 (N_11504,N_7448,N_9194);
nand U11505 (N_11505,N_8155,N_9252);
xnor U11506 (N_11506,N_9178,N_5539);
nand U11507 (N_11507,N_6787,N_9989);
or U11508 (N_11508,N_7220,N_9616);
xor U11509 (N_11509,N_8746,N_8504);
and U11510 (N_11510,N_8756,N_6849);
xor U11511 (N_11511,N_8928,N_5171);
and U11512 (N_11512,N_8937,N_9330);
nand U11513 (N_11513,N_5376,N_6882);
xnor U11514 (N_11514,N_7044,N_6674);
and U11515 (N_11515,N_6176,N_9204);
nor U11516 (N_11516,N_8859,N_6003);
and U11517 (N_11517,N_9389,N_5260);
nand U11518 (N_11518,N_9785,N_9803);
or U11519 (N_11519,N_6778,N_7253);
xor U11520 (N_11520,N_6171,N_7917);
or U11521 (N_11521,N_6150,N_6121);
nand U11522 (N_11522,N_8947,N_7582);
nand U11523 (N_11523,N_7862,N_8645);
nor U11524 (N_11524,N_5719,N_9508);
and U11525 (N_11525,N_5811,N_7748);
nand U11526 (N_11526,N_9604,N_7415);
xnor U11527 (N_11527,N_7241,N_6298);
or U11528 (N_11528,N_8363,N_8335);
or U11529 (N_11529,N_7524,N_9417);
or U11530 (N_11530,N_5950,N_9947);
xor U11531 (N_11531,N_8903,N_9543);
nand U11532 (N_11532,N_8593,N_8921);
nand U11533 (N_11533,N_9708,N_7112);
nor U11534 (N_11534,N_9129,N_7388);
nand U11535 (N_11535,N_9570,N_5164);
and U11536 (N_11536,N_8699,N_5701);
nand U11537 (N_11537,N_5902,N_5873);
or U11538 (N_11538,N_7195,N_7780);
xor U11539 (N_11539,N_6148,N_6307);
xnor U11540 (N_11540,N_7568,N_6204);
or U11541 (N_11541,N_7556,N_8615);
xor U11542 (N_11542,N_7705,N_5119);
xnor U11543 (N_11543,N_6493,N_9056);
nor U11544 (N_11544,N_7828,N_8703);
and U11545 (N_11545,N_7337,N_8612);
xnor U11546 (N_11546,N_5405,N_8621);
xor U11547 (N_11547,N_7637,N_8856);
xnor U11548 (N_11548,N_8278,N_5655);
xor U11549 (N_11549,N_9727,N_6551);
and U11550 (N_11550,N_7692,N_5165);
nor U11551 (N_11551,N_6626,N_9338);
nor U11552 (N_11552,N_5501,N_8683);
nor U11553 (N_11553,N_8138,N_8684);
xor U11554 (N_11554,N_5306,N_8771);
and U11555 (N_11555,N_6950,N_9817);
nand U11556 (N_11556,N_8752,N_7660);
or U11557 (N_11557,N_9053,N_8710);
and U11558 (N_11558,N_8294,N_7238);
or U11559 (N_11559,N_9657,N_6819);
nor U11560 (N_11560,N_9918,N_8814);
or U11561 (N_11561,N_8675,N_7387);
and U11562 (N_11562,N_7453,N_8110);
nand U11563 (N_11563,N_8577,N_8032);
and U11564 (N_11564,N_9088,N_7165);
or U11565 (N_11565,N_9955,N_7264);
nand U11566 (N_11566,N_9641,N_9266);
and U11567 (N_11567,N_7817,N_9358);
nor U11568 (N_11568,N_6353,N_6874);
and U11569 (N_11569,N_6285,N_7628);
xnor U11570 (N_11570,N_8650,N_8366);
or U11571 (N_11571,N_6129,N_5781);
nor U11572 (N_11572,N_9936,N_5861);
xor U11573 (N_11573,N_5387,N_9000);
nor U11574 (N_11574,N_5817,N_7007);
and U11575 (N_11575,N_6971,N_8582);
nor U11576 (N_11576,N_6594,N_9379);
or U11577 (N_11577,N_7236,N_5343);
xor U11578 (N_11578,N_8985,N_9435);
or U11579 (N_11579,N_7991,N_8140);
or U11580 (N_11580,N_6010,N_6740);
or U11581 (N_11581,N_7159,N_6955);
nor U11582 (N_11582,N_8130,N_6899);
xnor U11583 (N_11583,N_8841,N_9425);
xor U11584 (N_11584,N_6891,N_6770);
nor U11585 (N_11585,N_9548,N_5658);
nand U11586 (N_11586,N_7938,N_5247);
and U11587 (N_11587,N_6262,N_6196);
nor U11588 (N_11588,N_9751,N_9959);
and U11589 (N_11589,N_6297,N_9409);
and U11590 (N_11590,N_6350,N_5742);
and U11591 (N_11591,N_5097,N_6035);
or U11592 (N_11592,N_7234,N_8116);
xor U11593 (N_11593,N_5677,N_6502);
nor U11594 (N_11594,N_6863,N_7113);
nand U11595 (N_11595,N_7714,N_6825);
or U11596 (N_11596,N_5845,N_5031);
or U11597 (N_11597,N_9093,N_9651);
nand U11598 (N_11598,N_6631,N_9426);
nor U11599 (N_11599,N_6648,N_5435);
and U11600 (N_11600,N_7802,N_5839);
nor U11601 (N_11601,N_6610,N_8642);
nor U11602 (N_11602,N_8120,N_6917);
nor U11603 (N_11603,N_6167,N_8560);
nor U11604 (N_11604,N_5019,N_7206);
xnor U11605 (N_11605,N_7934,N_9069);
or U11606 (N_11606,N_8308,N_5578);
and U11607 (N_11607,N_6329,N_8171);
nand U11608 (N_11608,N_8873,N_7607);
nand U11609 (N_11609,N_6265,N_6500);
nand U11610 (N_11610,N_6606,N_5059);
or U11611 (N_11611,N_8049,N_5457);
or U11612 (N_11612,N_9715,N_8033);
nand U11613 (N_11613,N_8038,N_6033);
or U11614 (N_11614,N_8953,N_6868);
and U11615 (N_11615,N_7209,N_7913);
nor U11616 (N_11616,N_8882,N_5604);
nand U11617 (N_11617,N_7771,N_7947);
or U11618 (N_11618,N_5305,N_9750);
or U11619 (N_11619,N_5225,N_6034);
or U11620 (N_11620,N_9276,N_7876);
nand U11621 (N_11621,N_7879,N_9703);
and U11622 (N_11622,N_6925,N_7188);
nand U11623 (N_11623,N_5876,N_9449);
nand U11624 (N_11624,N_6499,N_8908);
nand U11625 (N_11625,N_7391,N_8700);
or U11626 (N_11626,N_6144,N_8948);
nand U11627 (N_11627,N_6252,N_5365);
nor U11628 (N_11628,N_6904,N_6836);
or U11629 (N_11629,N_8271,N_7095);
xor U11630 (N_11630,N_8777,N_8971);
and U11631 (N_11631,N_5986,N_5274);
xnor U11632 (N_11632,N_9336,N_9135);
or U11633 (N_11633,N_5502,N_5854);
and U11634 (N_11634,N_8364,N_7746);
nor U11635 (N_11635,N_7351,N_9235);
nand U11636 (N_11636,N_6630,N_9693);
and U11637 (N_11637,N_7131,N_5271);
nor U11638 (N_11638,N_5258,N_5967);
or U11639 (N_11639,N_8715,N_5259);
and U11640 (N_11640,N_8396,N_6423);
and U11641 (N_11641,N_9487,N_5532);
nand U11642 (N_11642,N_8510,N_6587);
nor U11643 (N_11643,N_7976,N_8706);
nand U11644 (N_11644,N_5628,N_5401);
nor U11645 (N_11645,N_5767,N_8471);
nor U11646 (N_11646,N_8669,N_8128);
and U11647 (N_11647,N_6348,N_7334);
or U11648 (N_11648,N_5167,N_5155);
nand U11649 (N_11649,N_5028,N_6416);
and U11650 (N_11650,N_7227,N_7623);
or U11651 (N_11651,N_7294,N_9434);
nor U11652 (N_11652,N_7439,N_7147);
or U11653 (N_11653,N_5198,N_8823);
and U11654 (N_11654,N_9905,N_8627);
nand U11655 (N_11655,N_7032,N_7989);
and U11656 (N_11656,N_7606,N_7138);
or U11657 (N_11657,N_6515,N_9406);
or U11658 (N_11658,N_9392,N_7252);
xor U11659 (N_11659,N_5591,N_5347);
or U11660 (N_11660,N_8231,N_5037);
and U11661 (N_11661,N_9512,N_8499);
nor U11662 (N_11662,N_8172,N_7890);
nor U11663 (N_11663,N_8745,N_8008);
and U11664 (N_11664,N_7077,N_5393);
and U11665 (N_11665,N_9834,N_6420);
nand U11666 (N_11666,N_7724,N_8721);
and U11667 (N_11667,N_5172,N_8991);
nor U11668 (N_11668,N_9659,N_8649);
nand U11669 (N_11669,N_8705,N_7060);
nor U11670 (N_11670,N_6700,N_5007);
or U11671 (N_11671,N_5355,N_7087);
nand U11672 (N_11672,N_5072,N_9282);
or U11673 (N_11673,N_7608,N_8251);
or U11674 (N_11674,N_9245,N_5643);
nand U11675 (N_11675,N_7631,N_7231);
and U11676 (N_11676,N_6790,N_9479);
xnor U11677 (N_11677,N_9644,N_7908);
xnor U11678 (N_11678,N_8602,N_9284);
xor U11679 (N_11679,N_9648,N_8955);
and U11680 (N_11680,N_6592,N_9100);
or U11681 (N_11681,N_8832,N_9883);
or U11682 (N_11682,N_5853,N_6015);
and U11683 (N_11683,N_6085,N_6296);
nand U11684 (N_11684,N_9326,N_5053);
or U11685 (N_11685,N_6981,N_5412);
or U11686 (N_11686,N_7576,N_7279);
or U11687 (N_11687,N_7942,N_6603);
nand U11688 (N_11688,N_9084,N_6246);
nor U11689 (N_11689,N_5572,N_7822);
and U11690 (N_11690,N_9238,N_8187);
nor U11691 (N_11691,N_6174,N_5841);
and U11692 (N_11692,N_8641,N_6784);
nor U11693 (N_11693,N_5143,N_6689);
nand U11694 (N_11694,N_9787,N_7013);
and U11695 (N_11695,N_8326,N_7679);
nand U11696 (N_11696,N_5890,N_8817);
nand U11697 (N_11697,N_5036,N_7567);
and U11698 (N_11698,N_5937,N_6907);
nor U11699 (N_11699,N_5089,N_5801);
xor U11700 (N_11700,N_8651,N_9098);
and U11701 (N_11701,N_7776,N_9066);
and U11702 (N_11702,N_7333,N_9070);
and U11703 (N_11703,N_9370,N_6546);
nor U11704 (N_11704,N_7101,N_9213);
xnor U11705 (N_11705,N_6677,N_5832);
nand U11706 (N_11706,N_6028,N_6536);
nor U11707 (N_11707,N_6561,N_6484);
or U11708 (N_11708,N_7406,N_9573);
nand U11709 (N_11709,N_5204,N_9788);
or U11710 (N_11710,N_5152,N_9771);
xor U11711 (N_11711,N_5799,N_7855);
nor U11712 (N_11712,N_5736,N_8221);
and U11713 (N_11713,N_7359,N_7336);
nor U11714 (N_11714,N_7261,N_6895);
and U11715 (N_11715,N_6395,N_7111);
or U11716 (N_11716,N_6564,N_9062);
nand U11717 (N_11717,N_7204,N_6403);
nor U11718 (N_11718,N_9826,N_8119);
nand U11719 (N_11719,N_6083,N_9675);
nand U11720 (N_11720,N_8015,N_8463);
and U11721 (N_11721,N_6079,N_7071);
and U11722 (N_11722,N_5323,N_9577);
or U11723 (N_11723,N_7528,N_5517);
xor U11724 (N_11724,N_8375,N_5002);
or U11725 (N_11725,N_8274,N_7474);
or U11726 (N_11726,N_5096,N_6862);
nor U11727 (N_11727,N_7058,N_7490);
nor U11728 (N_11728,N_5354,N_5697);
or U11729 (N_11729,N_7383,N_6632);
or U11730 (N_11730,N_9124,N_7538);
nand U11731 (N_11731,N_5436,N_5219);
and U11732 (N_11732,N_7899,N_5474);
xnor U11733 (N_11733,N_6058,N_8840);
nand U11734 (N_11734,N_7002,N_7461);
nand U11735 (N_11735,N_9079,N_6498);
and U11736 (N_11736,N_8043,N_7918);
and U11737 (N_11737,N_7669,N_9496);
and U11738 (N_11738,N_7518,N_8637);
xnor U11739 (N_11739,N_5829,N_7850);
and U11740 (N_11740,N_9216,N_7166);
nor U11741 (N_11741,N_8147,N_6756);
nor U11742 (N_11742,N_7605,N_7423);
and U11743 (N_11743,N_8975,N_5071);
nand U11744 (N_11744,N_6789,N_5848);
and U11745 (N_11745,N_6250,N_9673);
nand U11746 (N_11746,N_6346,N_5280);
or U11747 (N_11747,N_6425,N_8102);
and U11748 (N_11748,N_9163,N_5732);
or U11749 (N_11749,N_9738,N_6767);
nor U11750 (N_11750,N_5855,N_9949);
or U11751 (N_11751,N_9420,N_7954);
xnor U11752 (N_11752,N_7666,N_9729);
nand U11753 (N_11753,N_9310,N_6077);
nand U11754 (N_11754,N_7831,N_9645);
and U11755 (N_11755,N_5061,N_7307);
or U11756 (N_11756,N_7449,N_5664);
nor U11757 (N_11757,N_7998,N_7030);
or U11758 (N_11758,N_9059,N_5489);
nor U11759 (N_11759,N_8737,N_8592);
nand U11760 (N_11760,N_7882,N_5671);
nand U11761 (N_11761,N_6951,N_5127);
and U11762 (N_11762,N_6960,N_7029);
and U11763 (N_11763,N_9769,N_5181);
nor U11764 (N_11764,N_7450,N_7266);
or U11765 (N_11765,N_8739,N_5557);
and U11766 (N_11766,N_8545,N_8894);
and U11767 (N_11767,N_9042,N_7796);
nand U11768 (N_11768,N_7164,N_8374);
or U11769 (N_11769,N_9569,N_8444);
or U11770 (N_11770,N_6487,N_8159);
nor U11771 (N_11771,N_5721,N_7770);
and U11772 (N_11772,N_8458,N_9337);
and U11773 (N_11773,N_6912,N_9118);
or U11774 (N_11774,N_5135,N_7339);
nor U11775 (N_11775,N_8496,N_6601);
and U11776 (N_11776,N_7721,N_9907);
nand U11777 (N_11777,N_6886,N_8820);
and U11778 (N_11778,N_6801,N_7651);
and U11779 (N_11779,N_7320,N_9473);
and U11780 (N_11780,N_6172,N_7648);
nand U11781 (N_11781,N_9170,N_6814);
nor U11782 (N_11782,N_7706,N_8967);
and U11783 (N_11783,N_7348,N_6921);
nand U11784 (N_11784,N_8601,N_5771);
nand U11785 (N_11785,N_9081,N_6200);
and U11786 (N_11786,N_7097,N_5741);
xnor U11787 (N_11787,N_9242,N_9485);
or U11788 (N_11788,N_7614,N_9598);
or U11789 (N_11789,N_5003,N_5647);
and U11790 (N_11790,N_9534,N_9089);
nand U11791 (N_11791,N_7529,N_6614);
or U11792 (N_11792,N_9167,N_5948);
and U11793 (N_11793,N_9315,N_7237);
and U11794 (N_11794,N_7602,N_8926);
nor U11795 (N_11795,N_9620,N_5005);
or U11796 (N_11796,N_8234,N_5527);
and U11797 (N_11797,N_5074,N_9972);
or U11798 (N_11798,N_5055,N_8410);
and U11799 (N_11799,N_5115,N_5404);
nand U11800 (N_11800,N_6393,N_8595);
and U11801 (N_11801,N_7589,N_8377);
nor U11802 (N_11802,N_9962,N_5875);
nor U11803 (N_11803,N_8412,N_6993);
or U11804 (N_11804,N_6602,N_8083);
and U11805 (N_11805,N_7734,N_5738);
and U11806 (N_11806,N_9450,N_6661);
nand U11807 (N_11807,N_5783,N_6366);
nand U11808 (N_11808,N_7673,N_9085);
nand U11809 (N_11809,N_7983,N_5476);
and U11810 (N_11810,N_5455,N_8744);
nand U11811 (N_11811,N_9520,N_7604);
xnor U11812 (N_11812,N_8530,N_8327);
nand U11813 (N_11813,N_6574,N_9302);
nand U11814 (N_11814,N_5569,N_8646);
nor U11815 (N_11815,N_9813,N_6958);
nor U11816 (N_11816,N_7655,N_5626);
nor U11817 (N_11817,N_6540,N_7135);
nand U11818 (N_11818,N_9484,N_8568);
xor U11819 (N_11819,N_6194,N_5430);
nand U11820 (N_11820,N_9891,N_6257);
or U11821 (N_11821,N_7326,N_7422);
and U11822 (N_11822,N_6009,N_8393);
and U11823 (N_11823,N_6785,N_7280);
and U11824 (N_11824,N_5426,N_9527);
nor U11825 (N_11825,N_7939,N_8351);
nand U11826 (N_11826,N_5233,N_8095);
or U11827 (N_11827,N_5098,N_8798);
and U11828 (N_11828,N_8090,N_5133);
nor U11829 (N_11829,N_8870,N_9848);
nand U11830 (N_11830,N_5410,N_6946);
and U11831 (N_11831,N_6771,N_7794);
xor U11832 (N_11832,N_7125,N_5128);
nand U11833 (N_11833,N_8183,N_7340);
nor U11834 (N_11834,N_5711,N_6759);
xor U11835 (N_11835,N_7210,N_7897);
nor U11836 (N_11836,N_5881,N_5535);
or U11837 (N_11837,N_5094,N_7867);
or U11838 (N_11838,N_7016,N_8647);
nand U11839 (N_11839,N_6983,N_9755);
nand U11840 (N_11840,N_9956,N_8123);
and U11841 (N_11841,N_7840,N_5627);
or U11842 (N_11842,N_5866,N_9039);
nor U11843 (N_11843,N_5568,N_6816);
or U11844 (N_11844,N_9220,N_8456);
or U11845 (N_11845,N_6491,N_6304);
or U11846 (N_11846,N_9671,N_5352);
or U11847 (N_11847,N_7711,N_6517);
or U11848 (N_11848,N_8485,N_9966);
or U11849 (N_11849,N_9706,N_8634);
nand U11850 (N_11850,N_7936,N_8869);
and U11851 (N_11851,N_8677,N_9535);
and U11852 (N_11852,N_7701,N_6020);
or U11853 (N_11853,N_8543,N_6132);
and U11854 (N_11854,N_5945,N_5025);
or U11855 (N_11855,N_7760,N_5882);
nor U11856 (N_11856,N_5683,N_9590);
xnor U11857 (N_11857,N_9684,N_8987);
xor U11858 (N_11858,N_9528,N_6938);
and U11859 (N_11859,N_5322,N_7107);
or U11860 (N_11860,N_5718,N_6007);
nor U11861 (N_11861,N_6503,N_6645);
or U11862 (N_11862,N_5849,N_7332);
nand U11863 (N_11863,N_8318,N_7297);
nand U11864 (N_11864,N_7476,N_5283);
nand U11865 (N_11865,N_9988,N_6693);
or U11866 (N_11866,N_5314,N_7784);
and U11867 (N_11867,N_7497,N_5687);
or U11868 (N_11868,N_7537,N_8063);
nand U11869 (N_11869,N_5593,N_9612);
or U11870 (N_11870,N_7849,N_5286);
xor U11871 (N_11871,N_5646,N_5461);
nand U11872 (N_11872,N_7931,N_7373);
nor U11873 (N_11873,N_7262,N_6002);
nor U11874 (N_11874,N_9968,N_5137);
xnor U11875 (N_11875,N_7109,N_9385);
xnor U11876 (N_11876,N_6714,N_7861);
and U11877 (N_11877,N_6722,N_5623);
or U11878 (N_11878,N_5835,N_8863);
xnor U11879 (N_11879,N_6240,N_8334);
or U11880 (N_11880,N_7781,N_9453);
nor U11881 (N_11881,N_7075,N_8399);
or U11882 (N_11882,N_5182,N_8673);
nor U11883 (N_11883,N_9503,N_8842);
and U11884 (N_11884,N_7055,N_6046);
nor U11885 (N_11885,N_5408,N_7352);
xnor U11886 (N_11886,N_9901,N_7047);
and U11887 (N_11887,N_6180,N_5505);
nand U11888 (N_11888,N_5326,N_9412);
or U11889 (N_11889,N_6982,N_8761);
and U11890 (N_11890,N_9571,N_5270);
nor U11891 (N_11891,N_7845,N_7786);
and U11892 (N_11892,N_8112,N_8567);
and U11893 (N_11893,N_6843,N_5731);
nand U11894 (N_11894,N_7470,N_5208);
or U11895 (N_11895,N_8861,N_5631);
nand U11896 (N_11896,N_7259,N_9749);
nand U11897 (N_11897,N_9144,N_5464);
xor U11898 (N_11898,N_9596,N_5761);
nor U11899 (N_11899,N_8537,N_6495);
nor U11900 (N_11900,N_7662,N_8013);
nand U11901 (N_11901,N_7665,N_7624);
and U11902 (N_11902,N_8600,N_5765);
and U11903 (N_11903,N_9855,N_5992);
or U11904 (N_11904,N_5980,N_9038);
nand U11905 (N_11905,N_5796,N_8951);
or U11906 (N_11906,N_6943,N_6846);
or U11907 (N_11907,N_8572,N_6547);
or U11908 (N_11908,N_5912,N_7611);
or U11909 (N_11909,N_8249,N_6406);
nand U11910 (N_11910,N_9777,N_7687);
and U11911 (N_11911,N_6181,N_9181);
nand U11912 (N_11912,N_5425,N_6439);
or U11913 (N_11913,N_7912,N_7677);
nor U11914 (N_11914,N_5465,N_8166);
nand U11915 (N_11915,N_6334,N_9362);
and U11916 (N_11916,N_5510,N_8279);
and U11917 (N_11917,N_8093,N_5947);
nor U11918 (N_11918,N_5185,N_7053);
or U11919 (N_11919,N_5596,N_8482);
nand U11920 (N_11920,N_8597,N_6394);
nor U11921 (N_11921,N_9798,N_7951);
nand U11922 (N_11922,N_6623,N_9377);
or U11923 (N_11923,N_6663,N_7927);
and U11924 (N_11924,N_6934,N_8383);
or U11925 (N_11925,N_5004,N_7881);
xnor U11926 (N_11926,N_6302,N_6786);
or U11927 (N_11927,N_7100,N_8707);
nor U11928 (N_11928,N_8797,N_9443);
and U11929 (N_11929,N_5321,N_9695);
xor U11930 (N_11930,N_5858,N_8227);
nand U11931 (N_11931,N_7300,N_5248);
or U11932 (N_11932,N_5545,N_8716);
xnor U11933 (N_11933,N_6505,N_8775);
xnor U11934 (N_11934,N_8062,N_9333);
nor U11935 (N_11935,N_5813,N_5724);
and U11936 (N_11936,N_9862,N_5547);
and U11937 (N_11937,N_7594,N_5100);
or U11938 (N_11938,N_6210,N_8478);
nand U11939 (N_11939,N_5805,N_7154);
and U11940 (N_11940,N_9391,N_6729);
xor U11941 (N_11941,N_9296,N_7844);
or U11942 (N_11942,N_7557,N_7645);
nor U11943 (N_11943,N_5481,N_9314);
and U11944 (N_11944,N_6339,N_7896);
or U11945 (N_11945,N_9307,N_8575);
nand U11946 (N_11946,N_9991,N_8262);
or U11947 (N_11947,N_6629,N_9576);
nor U11948 (N_11948,N_7006,N_9806);
nand U11949 (N_11949,N_7212,N_9405);
or U11950 (N_11950,N_7004,N_7443);
or U11951 (N_11951,N_9145,N_6300);
nand U11952 (N_11952,N_6238,N_9267);
nand U11953 (N_11953,N_5151,N_9095);
and U11954 (N_11954,N_7615,N_9887);
or U11955 (N_11955,N_6589,N_5485);
and U11956 (N_11956,N_7270,N_8803);
and U11957 (N_11957,N_8057,N_7990);
nor U11958 (N_11958,N_9353,N_5609);
nand U11959 (N_11959,N_9854,N_7997);
xor U11960 (N_11960,N_8488,N_6229);
nor U11961 (N_11961,N_6775,N_6021);
or U11962 (N_11962,N_8643,N_6616);
and U11963 (N_11963,N_9724,N_7948);
nor U11964 (N_11964,N_5779,N_5899);
xor U11965 (N_11965,N_5399,N_8522);
nor U11966 (N_11966,N_6627,N_8438);
xnor U11967 (N_11967,N_5145,N_6694);
or U11968 (N_11968,N_5211,N_5696);
or U11969 (N_11969,N_9367,N_6954);
or U11970 (N_11970,N_7271,N_9822);
nor U11971 (N_11971,N_9459,N_6998);
nor U11972 (N_11972,N_6223,N_7994);
and U11973 (N_11973,N_9364,N_9115);
and U11974 (N_11974,N_6137,N_7245);
and U11975 (N_11975,N_5889,N_8890);
or U11976 (N_11976,N_8838,N_6044);
and U11977 (N_11977,N_7162,N_9902);
or U11978 (N_11978,N_7597,N_8659);
or U11979 (N_11979,N_8367,N_9345);
nor U11980 (N_11980,N_9663,N_9260);
and U11981 (N_11981,N_5792,N_5392);
nor U11982 (N_11982,N_7743,N_5869);
or U11983 (N_11983,N_6410,N_5564);
or U11984 (N_11984,N_5205,N_9670);
and U11985 (N_11985,N_6896,N_5630);
nor U11986 (N_11986,N_6595,N_6372);
nand U11987 (N_11987,N_7670,N_8610);
nand U11988 (N_11988,N_8495,N_9368);
or U11989 (N_11989,N_6279,N_5512);
and U11990 (N_11990,N_5011,N_5396);
or U11991 (N_11991,N_8403,N_7254);
nand U11992 (N_11992,N_9371,N_8247);
nor U11993 (N_11993,N_5023,N_6373);
nor U11994 (N_11994,N_7224,N_9943);
or U11995 (N_11995,N_9951,N_6641);
and U11996 (N_11996,N_9140,N_7968);
nor U11997 (N_11997,N_7757,N_8230);
xnor U11998 (N_11998,N_6902,N_9359);
xor U11999 (N_11999,N_7398,N_5969);
nor U12000 (N_12000,N_9630,N_9547);
or U12001 (N_12001,N_7834,N_5778);
xnor U12002 (N_12002,N_9308,N_6408);
nor U12003 (N_12003,N_7354,N_7122);
nor U12004 (N_12004,N_8305,N_7066);
nor U12005 (N_12005,N_5319,N_5026);
or U12006 (N_12006,N_8889,N_8283);
xor U12007 (N_12007,N_7208,N_8153);
nand U12008 (N_12008,N_5202,N_6507);
nand U12009 (N_12009,N_6968,N_5762);
and U12010 (N_12010,N_5034,N_9674);
and U12011 (N_12011,N_5041,N_5660);
nor U12012 (N_12012,N_6055,N_7194);
nand U12013 (N_12013,N_7546,N_9270);
and U12014 (N_12014,N_6101,N_6973);
or U12015 (N_12015,N_5069,N_6822);
nand U12016 (N_12016,N_8813,N_8667);
nor U12017 (N_12017,N_8588,N_7871);
nand U12018 (N_12018,N_7472,N_5230);
nand U12019 (N_12019,N_9847,N_9150);
nand U12020 (N_12020,N_8468,N_7949);
or U12021 (N_12021,N_7303,N_8006);
xnor U12022 (N_12022,N_6793,N_7973);
nor U12023 (N_12023,N_6577,N_8526);
nor U12024 (N_12024,N_7875,N_9442);
nand U12025 (N_12025,N_8523,N_5956);
nand U12026 (N_12026,N_7729,N_7996);
nand U12027 (N_12027,N_9615,N_8622);
or U12028 (N_12028,N_9525,N_8704);
nand U12029 (N_12029,N_9567,N_8718);
nor U12030 (N_12030,N_5070,N_8381);
nand U12031 (N_12031,N_8571,N_5913);
and U12032 (N_12032,N_9565,N_9016);
nor U12033 (N_12033,N_5390,N_8802);
nand U12034 (N_12034,N_9745,N_9025);
nor U12035 (N_12035,N_5605,N_7313);
nand U12036 (N_12036,N_5169,N_9164);
nand U12037 (N_12037,N_5926,N_6049);
or U12038 (N_12038,N_5518,N_5918);
nand U12039 (N_12039,N_6575,N_5520);
or U12040 (N_12040,N_6869,N_8142);
nand U12041 (N_12041,N_6391,N_8373);
or U12042 (N_12042,N_6774,N_9979);
nand U12043 (N_12043,N_7688,N_9839);
or U12044 (N_12044,N_5706,N_7048);
xor U12045 (N_12045,N_9605,N_9009);
nand U12046 (N_12046,N_5281,N_5715);
nand U12047 (N_12047,N_5597,N_7034);
and U12048 (N_12048,N_7184,N_9195);
nand U12049 (N_12049,N_7902,N_6734);
xnor U12050 (N_12050,N_7054,N_8511);
nand U12051 (N_12051,N_9908,N_5373);
nand U12052 (N_12052,N_9895,N_7052);
nand U12053 (N_12053,N_8544,N_8209);
or U12054 (N_12054,N_7741,N_7747);
and U12055 (N_12055,N_5632,N_6447);
nor U12056 (N_12056,N_8920,N_6652);
xnor U12057 (N_12057,N_9824,N_9424);
xor U12058 (N_12058,N_7085,N_8352);
or U12059 (N_12059,N_8208,N_6962);
and U12060 (N_12060,N_5648,N_5951);
nand U12061 (N_12061,N_5981,N_9536);
or U12062 (N_12062,N_6984,N_9875);
or U12063 (N_12063,N_7192,N_5186);
or U12064 (N_12064,N_5498,N_7763);
or U12065 (N_12065,N_6690,N_5901);
or U12066 (N_12066,N_6305,N_7758);
nor U12067 (N_12067,N_9143,N_7193);
or U12068 (N_12068,N_6935,N_5908);
and U12069 (N_12069,N_8081,N_8881);
or U12070 (N_12070,N_5060,N_9843);
nand U12071 (N_12071,N_6436,N_7649);
and U12072 (N_12072,N_9754,N_5847);
xor U12073 (N_12073,N_6847,N_7820);
and U12074 (N_12074,N_5440,N_5795);
and U12075 (N_12075,N_9773,N_5576);
or U12076 (N_12076,N_9996,N_7275);
nor U12077 (N_12077,N_9031,N_5603);
nand U12078 (N_12078,N_8860,N_8550);
xnor U12079 (N_12079,N_9447,N_9791);
nand U12080 (N_12080,N_5699,N_9381);
and U12081 (N_12081,N_9265,N_5723);
nor U12082 (N_12082,N_8486,N_6883);
nand U12083 (N_12083,N_5309,N_7712);
and U12084 (N_12084,N_5904,N_9523);
nor U12085 (N_12085,N_5118,N_9823);
nand U12086 (N_12086,N_6309,N_8316);
and U12087 (N_12087,N_7892,N_8619);
and U12088 (N_12088,N_8202,N_9197);
nand U12089 (N_12089,N_5177,N_6314);
or U12090 (N_12090,N_5546,N_5922);
nor U12091 (N_12091,N_7684,N_6701);
and U12092 (N_12092,N_5370,N_8888);
and U12093 (N_12093,N_9002,N_5431);
or U12094 (N_12094,N_6473,N_9023);
nand U12095 (N_12095,N_6746,N_7704);
nor U12096 (N_12096,N_8321,N_7335);
or U12097 (N_12097,N_9236,N_6948);
or U12098 (N_12098,N_5360,N_6239);
or U12099 (N_12099,N_8885,N_6792);
nor U12100 (N_12100,N_5729,N_7364);
xor U12101 (N_12101,N_5140,N_9780);
and U12102 (N_12102,N_5768,N_5429);
xnor U12103 (N_12103,N_7864,N_9299);
and U12104 (N_12104,N_6075,N_5192);
and U12105 (N_12105,N_8439,N_9394);
xnor U12106 (N_12106,N_8900,N_9128);
or U12107 (N_12107,N_5158,N_6216);
nor U12108 (N_12108,N_5473,N_7229);
and U12109 (N_12109,N_7634,N_6374);
nor U12110 (N_12110,N_6511,N_5356);
nand U12111 (N_12111,N_9365,N_9678);
xnor U12112 (N_12112,N_5846,N_5067);
xor U12113 (N_12113,N_7182,N_9289);
and U12114 (N_12114,N_5989,N_5195);
nand U12115 (N_12115,N_5496,N_6537);
nor U12116 (N_12116,N_9742,N_9055);
or U12117 (N_12117,N_5327,N_9507);
nor U12118 (N_12118,N_9219,N_9857);
nand U12119 (N_12119,N_9910,N_5121);
or U12120 (N_12120,N_9208,N_5983);
nor U12121 (N_12121,N_8825,N_8569);
nand U12122 (N_12122,N_9463,N_9151);
and U12123 (N_12123,N_6918,N_6466);
or U12124 (N_12124,N_7251,N_5361);
or U12125 (N_12125,N_6128,N_9516);
and U12126 (N_12126,N_8435,N_5654);
nand U12127 (N_12127,N_8828,N_9928);
and U12128 (N_12128,N_8520,N_9306);
nor U12129 (N_12129,N_8875,N_6905);
xnor U12130 (N_12130,N_6080,N_7024);
and U12131 (N_12131,N_6858,N_7946);
and U12132 (N_12132,N_5537,N_8124);
nor U12133 (N_12133,N_5672,N_8936);
and U12134 (N_12134,N_5463,N_8238);
and U12135 (N_12135,N_7093,N_9210);
xor U12136 (N_12136,N_7810,N_7318);
and U12137 (N_12137,N_9649,N_5477);
nor U12138 (N_12138,N_8535,N_8031);
nor U12139 (N_12139,N_6957,N_9277);
or U12140 (N_12140,N_6254,N_5091);
nor U12141 (N_12141,N_5810,N_6827);
and U12142 (N_12142,N_6237,N_8711);
nor U12143 (N_12143,N_6839,N_6859);
or U12144 (N_12144,N_5752,N_5960);
or U12145 (N_12145,N_6913,N_7903);
nand U12146 (N_12146,N_8028,N_7909);
nand U12147 (N_12147,N_6956,N_6312);
nand U12148 (N_12148,N_5381,N_8988);
xor U12149 (N_12149,N_7911,N_9926);
xnor U12150 (N_12150,N_6001,N_8805);
nor U12151 (N_12151,N_5015,N_6293);
nor U12152 (N_12152,N_8158,N_9147);
xor U12153 (N_12153,N_5681,N_6284);
and U12154 (N_12154,N_6157,N_6713);
or U12155 (N_12155,N_8416,N_5105);
nand U12156 (N_12156,N_7454,N_6024);
nor U12157 (N_12157,N_9398,N_9522);
nor U12158 (N_12158,N_7187,N_8816);
or U12159 (N_12159,N_8562,N_5837);
xnor U12160 (N_12160,N_5659,N_7725);
xnor U12161 (N_12161,N_9184,N_9454);
or U12162 (N_12162,N_6683,N_5316);
and U12163 (N_12163,N_9838,N_6888);
and U12164 (N_12164,N_7250,N_6845);
and U12165 (N_12165,N_6022,N_9529);
nor U12166 (N_12166,N_5062,N_6214);
xnor U12167 (N_12167,N_9008,N_6065);
nand U12168 (N_12168,N_6404,N_5977);
and U12169 (N_12169,N_5299,N_9860);
or U12170 (N_12170,N_6967,N_5710);
and U12171 (N_12171,N_6747,N_8922);
nand U12172 (N_12172,N_7950,N_8655);
and U12173 (N_12173,N_5124,N_5921);
and U12174 (N_12174,N_8203,N_5577);
or U12175 (N_12175,N_8134,N_8538);
or U12176 (N_12176,N_9346,N_5793);
and U12177 (N_12177,N_6054,N_6529);
nand U12178 (N_12178,N_6676,N_7564);
nor U12179 (N_12179,N_8759,N_7833);
or U12180 (N_12180,N_5065,N_6706);
nand U12181 (N_12181,N_5197,N_8194);
nor U12182 (N_12182,N_5725,N_9568);
nand U12183 (N_12183,N_6113,N_8317);
nor U12184 (N_12184,N_9578,N_6671);
and U12185 (N_12185,N_8818,N_7563);
or U12186 (N_12186,N_6221,N_9136);
or U12187 (N_12187,N_6253,N_5398);
nand U12188 (N_12188,N_9878,N_8624);
and U12189 (N_12189,N_8422,N_8044);
and U12190 (N_12190,N_5126,N_5443);
nor U12191 (N_12191,N_8793,N_7291);
nand U12192 (N_12192,N_6593,N_7772);
or U12193 (N_12193,N_9092,N_6813);
nor U12194 (N_12194,N_9986,N_9386);
nor U12195 (N_12195,N_7080,N_9105);
or U12196 (N_12196,N_7301,N_5915);
xnor U12197 (N_12197,N_9458,N_9180);
xnor U12198 (N_12198,N_6118,N_8045);
nand U12199 (N_12199,N_6367,N_7121);
and U12200 (N_12200,N_5824,N_5747);
nor U12201 (N_12201,N_8406,N_6705);
nor U12202 (N_12202,N_5454,N_8916);
and U12203 (N_12203,N_6987,N_8188);
or U12204 (N_12204,N_8884,N_7956);
nand U12205 (N_12205,N_6453,N_9466);
xor U12206 (N_12206,N_6752,N_7017);
or U12207 (N_12207,N_9490,N_5548);
and U12208 (N_12208,N_9253,N_9677);
or U12209 (N_12209,N_9752,N_7286);
and U12210 (N_12210,N_8487,N_5831);
nand U12211 (N_12211,N_9480,N_9295);
nor U12212 (N_12212,N_6808,N_8508);
nor U12213 (N_12213,N_8076,N_6658);
and U12214 (N_12214,N_9293,N_6636);
nor U12215 (N_12215,N_5009,N_9146);
and U12216 (N_12216,N_7921,N_7018);
or U12217 (N_12217,N_9065,N_6396);
or U12218 (N_12218,N_6647,N_6418);
nor U12219 (N_12219,N_5774,N_7868);
nor U12220 (N_12220,N_7096,N_6844);
nor U12221 (N_12221,N_7272,N_7180);
or U12222 (N_12222,N_6504,N_7533);
nand U12223 (N_12223,N_6189,N_8927);
and U12224 (N_12224,N_7092,N_7914);
or U12225 (N_12225,N_9944,N_8493);
or U12226 (N_12226,N_7928,N_9373);
or U12227 (N_12227,N_7814,N_9291);
or U12228 (N_12228,N_6078,N_6520);
and U12229 (N_12229,N_7191,N_6543);
nand U12230 (N_12230,N_5678,N_7463);
nand U12231 (N_12231,N_7511,N_6271);
and U12232 (N_12232,N_9438,N_6359);
and U12233 (N_12233,N_6006,N_6413);
nor U12234 (N_12234,N_7601,N_7676);
and U12235 (N_12235,N_9029,N_7341);
and U12236 (N_12236,N_7731,N_8067);
or U12237 (N_12237,N_6442,N_7857);
nor U12238 (N_12238,N_7619,N_6472);
nor U12239 (N_12239,N_7247,N_5131);
nor U12240 (N_12240,N_7730,N_9653);
or U12241 (N_12241,N_6622,N_9481);
nand U12242 (N_12242,N_8163,N_7389);
and U12243 (N_12243,N_7105,N_9709);
nand U12244 (N_12244,N_5240,N_7693);
nand U12245 (N_12245,N_8946,N_8865);
nand U12246 (N_12246,N_6986,N_9113);
xnor U12247 (N_12247,N_7090,N_5218);
nor U12248 (N_12248,N_6248,N_8778);
or U12249 (N_12249,N_8331,N_8464);
xor U12250 (N_12250,N_7328,N_9418);
or U12251 (N_12251,N_9801,N_9859);
nand U12252 (N_12252,N_5264,N_9574);
nand U12253 (N_12253,N_8240,N_8574);
nand U12254 (N_12254,N_9500,N_6317);
or U12255 (N_12255,N_7329,N_8548);
and U12256 (N_12256,N_9012,N_6370);
and U12257 (N_12257,N_5525,N_9086);
nor U12258 (N_12258,N_6326,N_8105);
nor U12259 (N_12259,N_8932,N_6860);
nor U12260 (N_12260,N_7832,N_6990);
or U12261 (N_12261,N_6365,N_9440);
xnor U12262 (N_12262,N_7242,N_7893);
xor U12263 (N_12263,N_7274,N_6542);
nand U12264 (N_12264,N_5433,N_5149);
or U12265 (N_12265,N_9158,N_9800);
nand U12266 (N_12266,N_6048,N_6924);
or U12267 (N_12267,N_9448,N_6766);
and U12268 (N_12268,N_6146,N_7640);
or U12269 (N_12269,N_8064,N_6807);
nor U12270 (N_12270,N_8204,N_6976);
nor U12271 (N_12271,N_8709,N_5040);
or U12272 (N_12272,N_7974,N_9661);
xor U12273 (N_12273,N_9830,N_7205);
and U12274 (N_12274,N_7273,N_9904);
nor U12275 (N_12275,N_5722,N_7783);
and U12276 (N_12276,N_9753,N_6140);
nor U12277 (N_12277,N_5276,N_9707);
nor U12278 (N_12278,N_8136,N_7110);
nor U12279 (N_12279,N_6655,N_6562);
and U12280 (N_12280,N_7613,N_8065);
xnor U12281 (N_12281,N_7749,N_8877);
xnor U12282 (N_12282,N_5620,N_6779);
nor U12283 (N_12283,N_6703,N_8631);
and U12284 (N_12284,N_7630,N_5946);
nand U12285 (N_12285,N_6999,N_6662);
or U12286 (N_12286,N_7019,N_8708);
nand U12287 (N_12287,N_9744,N_7357);
or U12288 (N_12288,N_7664,N_6063);
and U12289 (N_12289,N_5168,N_6768);
or U12290 (N_12290,N_5261,N_6398);
nor U12291 (N_12291,N_5374,N_5294);
or U12292 (N_12292,N_8872,N_8748);
and U12293 (N_12293,N_8827,N_7915);
nor U12294 (N_12294,N_6572,N_6183);
or U12295 (N_12295,N_9091,N_9153);
or U12296 (N_12296,N_8336,N_5684);
nor U12297 (N_12297,N_8635,N_6155);
xor U12298 (N_12298,N_8026,N_5117);
nor U12299 (N_12299,N_8145,N_6544);
nor U12300 (N_12300,N_6241,N_8919);
and U12301 (N_12301,N_7174,N_5780);
nand U12302 (N_12302,N_9108,N_9958);
and U12303 (N_12303,N_8191,N_7199);
or U12304 (N_12304,N_7324,N_7025);
or U12305 (N_12305,N_6748,N_9112);
xor U12306 (N_12306,N_6106,N_9190);
nor U12307 (N_12307,N_7437,N_6288);
or U12308 (N_12308,N_5450,N_9844);
and U12309 (N_12309,N_7145,N_5379);
nand U12310 (N_12310,N_7434,N_8330);
or U12311 (N_12311,N_6875,N_6387);
and U12312 (N_12312,N_9977,N_9445);
nand U12313 (N_12313,N_5624,N_9207);
nor U12314 (N_12314,N_7322,N_9320);
or U12315 (N_12315,N_6126,N_8089);
nand U12316 (N_12316,N_7750,N_5344);
nand U12317 (N_12317,N_6230,N_8489);
nor U12318 (N_12318,N_8449,N_6621);
nand U12319 (N_12319,N_5636,N_5698);
or U12320 (N_12320,N_5709,N_8849);
nand U12321 (N_12321,N_6452,N_7691);
xnor U12322 (N_12322,N_9579,N_7046);
and U12323 (N_12323,N_7118,N_6668);
xor U12324 (N_12324,N_9921,N_5122);
nor U12325 (N_12325,N_6193,N_8115);
or U12326 (N_12326,N_7719,N_8389);
nand U12327 (N_12327,N_8029,N_5189);
or U12328 (N_12328,N_6269,N_8007);
or U12329 (N_12329,N_6061,N_8997);
or U12330 (N_12330,N_9931,N_9179);
or U12331 (N_12331,N_5249,N_9903);
nand U12332 (N_12332,N_5675,N_9460);
nand U12333 (N_12333,N_8765,N_6212);
or U12334 (N_12334,N_6215,N_7039);
and U12335 (N_12335,N_8362,N_6435);
xnor U12336 (N_12336,N_9808,N_8603);
nor U12337 (N_12337,N_8781,N_9168);
or U12338 (N_12338,N_6025,N_9603);
or U12339 (N_12339,N_5150,N_8836);
and U12340 (N_12340,N_7626,N_7522);
xnor U12341 (N_12341,N_7045,N_9324);
and U12342 (N_12342,N_5236,N_6135);
nand U12343 (N_12343,N_5348,N_6441);
and U12344 (N_12344,N_5900,N_5134);
nand U12345 (N_12345,N_9672,N_9082);
nor U12346 (N_12346,N_7558,N_9047);
and U12347 (N_12347,N_7041,N_9010);
nor U12348 (N_12348,N_9160,N_8819);
nor U12349 (N_12349,N_8131,N_8309);
and U12350 (N_12350,N_6831,N_7407);
nor U12351 (N_12351,N_6341,N_8266);
or U12352 (N_12352,N_9701,N_8077);
nand U12353 (N_12353,N_7492,N_8380);
or U12354 (N_12354,N_8091,N_8692);
or U12355 (N_12355,N_7331,N_8986);
nor U12356 (N_12356,N_8457,N_9868);
or U12357 (N_12357,N_7136,N_8170);
and U12358 (N_12358,N_7036,N_8225);
nand U12359 (N_12359,N_6397,N_7067);
nand U12360 (N_12360,N_8299,N_6764);
xnor U12361 (N_12361,N_9998,N_9248);
xnor U12362 (N_12362,N_7663,N_8942);
nand U12363 (N_12363,N_5475,N_8623);
and U12364 (N_12364,N_6475,N_5787);
or U12365 (N_12365,N_7091,N_9626);
or U12366 (N_12366,N_8378,N_9223);
and U12367 (N_12367,N_9767,N_5896);
or U12368 (N_12368,N_5362,N_9621);
xnor U12369 (N_12369,N_5371,N_9375);
or U12370 (N_12370,N_5815,N_8292);
and U12371 (N_12371,N_5441,N_5917);
and U12372 (N_12372,N_5297,N_8175);
or U12373 (N_12373,N_6361,N_8333);
and U12374 (N_12374,N_7698,N_7429);
or U12375 (N_12375,N_7269,N_8342);
nor U12376 (N_12376,N_8453,N_9784);
nand U12377 (N_12377,N_8714,N_7260);
nor U12378 (N_12378,N_6136,N_9037);
or U12379 (N_12379,N_5311,N_7255);
xor U12380 (N_12380,N_5541,N_8491);
and U12381 (N_12381,N_8354,N_7767);
and U12382 (N_12382,N_5018,N_8904);
or U12383 (N_12383,N_9656,N_9873);
or U12384 (N_12384,N_9351,N_9950);
and U12385 (N_12385,N_7428,N_6972);
and U12386 (N_12386,N_6182,N_6731);
and U12387 (N_12387,N_6533,N_8300);
xnor U12388 (N_12388,N_5772,N_9211);
nand U12389 (N_12389,N_8277,N_9804);
or U12390 (N_12390,N_6941,N_7499);
or U12391 (N_12391,N_8210,N_9201);
and U12392 (N_12392,N_6188,N_8616);
nor U12393 (N_12393,N_7170,N_8371);
xor U12394 (N_12394,N_7877,N_8833);
or U12395 (N_12395,N_7368,N_9175);
and U12396 (N_12396,N_8388,N_5534);
and U12397 (N_12397,N_5693,N_6045);
nand U12398 (N_12398,N_7256,N_5611);
nor U12399 (N_12399,N_5991,N_6368);
or U12400 (N_12400,N_7685,N_5057);
or U12401 (N_12401,N_5277,N_7299);
nor U12402 (N_12402,N_5851,N_8960);
nor U12403 (N_12403,N_9698,N_9021);
xnor U12404 (N_12404,N_8691,N_7883);
and U12405 (N_12405,N_8071,N_7599);
or U12406 (N_12406,N_8845,N_6739);
or U12407 (N_12407,N_8638,N_5966);
or U12408 (N_12408,N_8306,N_5859);
or U12409 (N_12409,N_9730,N_7148);
nor U12410 (N_12410,N_8636,N_9013);
nor U12411 (N_12411,N_7768,N_7543);
xor U12412 (N_12412,N_9393,N_8025);
nor U12413 (N_12413,N_9733,N_6096);
or U12414 (N_12414,N_8401,N_5607);
xnor U12415 (N_12415,N_6566,N_6830);
xor U12416 (N_12416,N_6866,N_8868);
xnor U12417 (N_12417,N_6737,N_7962);
nand U12418 (N_12418,N_5561,N_7514);
nand U12419 (N_12419,N_5633,N_7314);
xor U12420 (N_12420,N_9588,N_5910);
and U12421 (N_12421,N_7176,N_6428);
and U12422 (N_12422,N_8041,N_8108);
xor U12423 (N_12423,N_8314,N_5445);
nand U12424 (N_12424,N_5448,N_8628);
nor U12425 (N_12425,N_9050,N_7305);
or U12426 (N_12426,N_7000,N_9680);
nor U12427 (N_12427,N_9584,N_8915);
nand U12428 (N_12428,N_7325,N_7674);
xnor U12429 (N_12429,N_6509,N_9794);
and U12430 (N_12430,N_8632,N_5212);
nand U12431 (N_12431,N_6255,N_9103);
or U12432 (N_12432,N_6573,N_5954);
or U12433 (N_12433,N_6596,N_5930);
and U12434 (N_12434,N_7756,N_9011);
and U12435 (N_12435,N_6438,N_7745);
nor U12436 (N_12436,N_7612,N_8604);
and U12437 (N_12437,N_9193,N_7671);
or U12438 (N_12438,N_7292,N_9363);
and U12439 (N_12439,N_6598,N_5491);
and U12440 (N_12440,N_6114,N_6066);
nor U12441 (N_12441,N_5338,N_6670);
nand U12442 (N_12442,N_7342,N_5413);
and U12443 (N_12443,N_8729,N_9366);
nand U12444 (N_12444,N_7478,N_8500);
nand U12445 (N_12445,N_6581,N_6354);
or U12446 (N_12446,N_8405,N_6017);
nand U12447 (N_12447,N_7552,N_8344);
or U12448 (N_12448,N_7185,N_7445);
and U12449 (N_12449,N_9261,N_6672);
or U12450 (N_12450,N_6965,N_5843);
nor U12451 (N_12451,N_5919,N_7040);
nor U12452 (N_12452,N_5704,N_6829);
nand U12453 (N_12453,N_6692,N_7506);
or U12454 (N_12454,N_5691,N_6837);
xnor U12455 (N_12455,N_7846,N_7732);
nor U12456 (N_12456,N_5616,N_7980);
and U12457 (N_12457,N_6142,N_7484);
nor U12458 (N_12458,N_6060,N_5865);
nor U12459 (N_12459,N_6162,N_9126);
and U12460 (N_12460,N_6695,N_5745);
nor U12461 (N_12461,N_8512,N_5791);
and U12462 (N_12462,N_9983,N_7495);
and U12463 (N_12463,N_9953,N_8157);
nand U12464 (N_12464,N_9792,N_5737);
and U12465 (N_12465,N_7394,N_8103);
or U12466 (N_12466,N_6105,N_5907);
and U12467 (N_12467,N_7736,N_9992);
nand U12468 (N_12468,N_6261,N_5223);
nor U12469 (N_12469,N_6184,N_9331);
nand U12470 (N_12470,N_9592,N_8668);
nor U12471 (N_12471,N_8447,N_9628);
nand U12472 (N_12472,N_6158,N_9585);
or U12473 (N_12473,N_6234,N_8135);
nor U12474 (N_12474,N_7595,N_7197);
nor U12475 (N_12475,N_5129,N_7099);
nand U12476 (N_12476,N_8467,N_6308);
and U12477 (N_12477,N_8302,N_7773);
or U12478 (N_12478,N_7977,N_7141);
or U12479 (N_12479,N_6266,N_9610);
nor U12480 (N_12480,N_7411,N_5179);
xnor U12481 (N_12481,N_9067,N_7978);
and U12482 (N_12482,N_5673,N_9580);
nor U12483 (N_12483,N_5727,N_5159);
xnor U12484 (N_12484,N_6274,N_7851);
nor U12485 (N_12485,N_6978,N_6833);
nor U12486 (N_12486,N_6103,N_7371);
nor U12487 (N_12487,N_5550,N_5334);
or U12488 (N_12488,N_6337,N_9632);
nor U12489 (N_12489,N_9046,N_9006);
nand U12490 (N_12490,N_5516,N_7967);
and U12491 (N_12491,N_6605,N_6186);
or U12492 (N_12492,N_6919,N_9352);
and U12493 (N_12493,N_7468,N_7277);
nor U12494 (N_12494,N_6624,N_7553);
or U12495 (N_12495,N_5582,N_6056);
nand U12496 (N_12496,N_7161,N_7033);
nor U12497 (N_12497,N_8933,N_9294);
nor U12498 (N_12498,N_7321,N_5740);
or U12499 (N_12499,N_8018,N_5421);
and U12500 (N_12500,N_6512,N_5748);
nand U12501 (N_12501,N_6617,N_6240);
and U12502 (N_12502,N_7749,N_7094);
xor U12503 (N_12503,N_5840,N_5072);
nand U12504 (N_12504,N_9859,N_6934);
nor U12505 (N_12505,N_7743,N_9186);
and U12506 (N_12506,N_6386,N_9986);
nor U12507 (N_12507,N_9819,N_5741);
and U12508 (N_12508,N_9102,N_7689);
nor U12509 (N_12509,N_7022,N_5557);
and U12510 (N_12510,N_7108,N_9290);
nand U12511 (N_12511,N_5365,N_9055);
and U12512 (N_12512,N_7605,N_5406);
nor U12513 (N_12513,N_6956,N_5433);
nor U12514 (N_12514,N_6564,N_6629);
nor U12515 (N_12515,N_8212,N_6241);
nor U12516 (N_12516,N_8515,N_5584);
nor U12517 (N_12517,N_7390,N_9493);
nand U12518 (N_12518,N_5331,N_6523);
or U12519 (N_12519,N_5117,N_8762);
nor U12520 (N_12520,N_9413,N_8786);
or U12521 (N_12521,N_8072,N_5499);
nor U12522 (N_12522,N_6156,N_9972);
xor U12523 (N_12523,N_8525,N_9818);
nand U12524 (N_12524,N_6084,N_9978);
nor U12525 (N_12525,N_7945,N_8055);
nand U12526 (N_12526,N_9022,N_9878);
or U12527 (N_12527,N_7357,N_8486);
nand U12528 (N_12528,N_8635,N_8852);
and U12529 (N_12529,N_6820,N_7160);
nor U12530 (N_12530,N_9639,N_8831);
nand U12531 (N_12531,N_8142,N_5543);
nand U12532 (N_12532,N_5049,N_9075);
or U12533 (N_12533,N_7235,N_5376);
and U12534 (N_12534,N_5430,N_6796);
or U12535 (N_12535,N_6761,N_6312);
or U12536 (N_12536,N_5100,N_7527);
nand U12537 (N_12537,N_5961,N_8184);
and U12538 (N_12538,N_5141,N_5815);
and U12539 (N_12539,N_9680,N_5624);
nand U12540 (N_12540,N_6239,N_5307);
and U12541 (N_12541,N_7123,N_6002);
or U12542 (N_12542,N_7710,N_7927);
nor U12543 (N_12543,N_8862,N_7816);
and U12544 (N_12544,N_9727,N_9968);
nand U12545 (N_12545,N_8184,N_9027);
nor U12546 (N_12546,N_7172,N_9621);
xor U12547 (N_12547,N_5760,N_7657);
nand U12548 (N_12548,N_9721,N_6839);
xor U12549 (N_12549,N_8503,N_7365);
nor U12550 (N_12550,N_9041,N_7716);
nor U12551 (N_12551,N_5008,N_7622);
or U12552 (N_12552,N_5226,N_9063);
and U12553 (N_12553,N_5914,N_9185);
and U12554 (N_12554,N_7803,N_7332);
nand U12555 (N_12555,N_7637,N_9203);
and U12556 (N_12556,N_6563,N_6328);
nor U12557 (N_12557,N_6621,N_5862);
or U12558 (N_12558,N_7427,N_5532);
xnor U12559 (N_12559,N_7148,N_5202);
or U12560 (N_12560,N_5079,N_6142);
and U12561 (N_12561,N_8646,N_8779);
or U12562 (N_12562,N_9658,N_9809);
nand U12563 (N_12563,N_9436,N_7342);
xor U12564 (N_12564,N_5025,N_6104);
nand U12565 (N_12565,N_8357,N_8230);
or U12566 (N_12566,N_9002,N_8244);
or U12567 (N_12567,N_8254,N_8617);
and U12568 (N_12568,N_9711,N_5404);
and U12569 (N_12569,N_8917,N_9039);
nand U12570 (N_12570,N_6295,N_8251);
nand U12571 (N_12571,N_8623,N_6274);
nor U12572 (N_12572,N_5975,N_5317);
nor U12573 (N_12573,N_5309,N_7170);
and U12574 (N_12574,N_7483,N_9197);
nor U12575 (N_12575,N_5241,N_6554);
or U12576 (N_12576,N_5698,N_7034);
or U12577 (N_12577,N_5569,N_8865);
nor U12578 (N_12578,N_7090,N_8050);
nand U12579 (N_12579,N_9210,N_9314);
nand U12580 (N_12580,N_5136,N_9787);
or U12581 (N_12581,N_6309,N_5975);
and U12582 (N_12582,N_5324,N_7099);
nor U12583 (N_12583,N_9500,N_5461);
xor U12584 (N_12584,N_9763,N_8814);
nor U12585 (N_12585,N_6307,N_7273);
nor U12586 (N_12586,N_7143,N_6384);
nor U12587 (N_12587,N_6798,N_9686);
xor U12588 (N_12588,N_7583,N_5560);
nand U12589 (N_12589,N_7944,N_9498);
or U12590 (N_12590,N_9918,N_5796);
xor U12591 (N_12591,N_8070,N_9423);
or U12592 (N_12592,N_6131,N_9483);
xnor U12593 (N_12593,N_9975,N_6206);
nand U12594 (N_12594,N_6232,N_6531);
or U12595 (N_12595,N_8202,N_8816);
or U12596 (N_12596,N_9533,N_7016);
and U12597 (N_12597,N_7536,N_6176);
and U12598 (N_12598,N_5667,N_7638);
nand U12599 (N_12599,N_6159,N_9657);
nand U12600 (N_12600,N_8905,N_7838);
nand U12601 (N_12601,N_8277,N_8271);
or U12602 (N_12602,N_5043,N_9497);
or U12603 (N_12603,N_8307,N_9483);
nand U12604 (N_12604,N_9652,N_6041);
and U12605 (N_12605,N_6143,N_6346);
or U12606 (N_12606,N_9042,N_6143);
or U12607 (N_12607,N_6477,N_7389);
nor U12608 (N_12608,N_6140,N_5991);
nor U12609 (N_12609,N_5231,N_5459);
xor U12610 (N_12610,N_9238,N_8379);
or U12611 (N_12611,N_7114,N_8420);
and U12612 (N_12612,N_8200,N_7616);
or U12613 (N_12613,N_7063,N_5852);
or U12614 (N_12614,N_6206,N_6039);
and U12615 (N_12615,N_6578,N_6950);
nand U12616 (N_12616,N_6482,N_6598);
xnor U12617 (N_12617,N_7638,N_5290);
or U12618 (N_12618,N_7159,N_8948);
or U12619 (N_12619,N_8818,N_9161);
nand U12620 (N_12620,N_8199,N_8599);
xor U12621 (N_12621,N_8257,N_6735);
and U12622 (N_12622,N_7499,N_6617);
xnor U12623 (N_12623,N_8000,N_5335);
xor U12624 (N_12624,N_6502,N_9336);
or U12625 (N_12625,N_6193,N_8767);
and U12626 (N_12626,N_9217,N_7730);
nand U12627 (N_12627,N_9030,N_5751);
and U12628 (N_12628,N_5421,N_6809);
nor U12629 (N_12629,N_5600,N_7386);
and U12630 (N_12630,N_8906,N_6420);
xnor U12631 (N_12631,N_5417,N_8604);
nand U12632 (N_12632,N_8207,N_6048);
or U12633 (N_12633,N_7796,N_9919);
and U12634 (N_12634,N_8329,N_8064);
and U12635 (N_12635,N_7454,N_8569);
nor U12636 (N_12636,N_7893,N_5981);
nor U12637 (N_12637,N_9618,N_7924);
and U12638 (N_12638,N_9312,N_9418);
nor U12639 (N_12639,N_5675,N_7454);
nand U12640 (N_12640,N_8547,N_6068);
nor U12641 (N_12641,N_9293,N_8281);
or U12642 (N_12642,N_5230,N_7327);
nand U12643 (N_12643,N_8228,N_5010);
nor U12644 (N_12644,N_9809,N_8695);
nand U12645 (N_12645,N_7617,N_7660);
nor U12646 (N_12646,N_8975,N_6880);
nand U12647 (N_12647,N_9791,N_7435);
nand U12648 (N_12648,N_9117,N_7111);
nand U12649 (N_12649,N_8302,N_5592);
nand U12650 (N_12650,N_8735,N_8990);
and U12651 (N_12651,N_6164,N_7565);
xor U12652 (N_12652,N_5012,N_6720);
nor U12653 (N_12653,N_7233,N_9057);
xnor U12654 (N_12654,N_8946,N_8856);
nand U12655 (N_12655,N_6161,N_9935);
nand U12656 (N_12656,N_6755,N_9239);
or U12657 (N_12657,N_8514,N_7758);
or U12658 (N_12658,N_6709,N_6331);
and U12659 (N_12659,N_6046,N_7032);
nor U12660 (N_12660,N_6496,N_5951);
or U12661 (N_12661,N_6673,N_8528);
and U12662 (N_12662,N_8866,N_5186);
nand U12663 (N_12663,N_8388,N_5472);
nand U12664 (N_12664,N_6733,N_8898);
nor U12665 (N_12665,N_7196,N_8428);
and U12666 (N_12666,N_6756,N_5705);
and U12667 (N_12667,N_6366,N_7323);
nand U12668 (N_12668,N_8516,N_6853);
and U12669 (N_12669,N_6705,N_7048);
and U12670 (N_12670,N_7066,N_6218);
and U12671 (N_12671,N_9879,N_8757);
nor U12672 (N_12672,N_7937,N_7496);
or U12673 (N_12673,N_9317,N_6034);
nor U12674 (N_12674,N_8699,N_9681);
or U12675 (N_12675,N_5872,N_5049);
or U12676 (N_12676,N_6704,N_9767);
or U12677 (N_12677,N_8605,N_9667);
xnor U12678 (N_12678,N_7035,N_5852);
and U12679 (N_12679,N_5377,N_5992);
and U12680 (N_12680,N_8288,N_5379);
nor U12681 (N_12681,N_5783,N_8887);
and U12682 (N_12682,N_6250,N_7232);
xor U12683 (N_12683,N_8253,N_8970);
nand U12684 (N_12684,N_5774,N_7258);
nor U12685 (N_12685,N_9179,N_6861);
or U12686 (N_12686,N_7728,N_8994);
nand U12687 (N_12687,N_7844,N_9159);
nand U12688 (N_12688,N_5258,N_5637);
nand U12689 (N_12689,N_9719,N_5308);
nand U12690 (N_12690,N_8899,N_5872);
or U12691 (N_12691,N_9492,N_6233);
nand U12692 (N_12692,N_9367,N_5626);
or U12693 (N_12693,N_5045,N_7741);
nand U12694 (N_12694,N_6043,N_5185);
nand U12695 (N_12695,N_8293,N_9073);
nor U12696 (N_12696,N_7011,N_7648);
nand U12697 (N_12697,N_9392,N_9653);
and U12698 (N_12698,N_8965,N_7939);
nand U12699 (N_12699,N_5299,N_5979);
nand U12700 (N_12700,N_5994,N_7353);
nor U12701 (N_12701,N_9697,N_6260);
nor U12702 (N_12702,N_6838,N_7122);
nand U12703 (N_12703,N_8999,N_9522);
nand U12704 (N_12704,N_7049,N_9759);
or U12705 (N_12705,N_9638,N_6455);
nand U12706 (N_12706,N_7640,N_9041);
nand U12707 (N_12707,N_9011,N_8666);
nor U12708 (N_12708,N_8159,N_7108);
or U12709 (N_12709,N_9783,N_8170);
xnor U12710 (N_12710,N_7123,N_7056);
xnor U12711 (N_12711,N_5725,N_8314);
and U12712 (N_12712,N_7695,N_8305);
or U12713 (N_12713,N_9820,N_5025);
or U12714 (N_12714,N_7945,N_8959);
and U12715 (N_12715,N_9088,N_9440);
or U12716 (N_12716,N_7075,N_7091);
and U12717 (N_12717,N_9744,N_5321);
or U12718 (N_12718,N_9597,N_6121);
nor U12719 (N_12719,N_5441,N_5345);
nand U12720 (N_12720,N_6614,N_6004);
xnor U12721 (N_12721,N_5534,N_6450);
or U12722 (N_12722,N_9567,N_7947);
nor U12723 (N_12723,N_9139,N_8995);
and U12724 (N_12724,N_7256,N_7695);
and U12725 (N_12725,N_8757,N_7860);
nand U12726 (N_12726,N_7659,N_9284);
or U12727 (N_12727,N_7403,N_6929);
and U12728 (N_12728,N_9336,N_8040);
or U12729 (N_12729,N_8139,N_9784);
and U12730 (N_12730,N_6278,N_6457);
nor U12731 (N_12731,N_9008,N_9348);
nand U12732 (N_12732,N_7902,N_6121);
nand U12733 (N_12733,N_6797,N_5703);
or U12734 (N_12734,N_7169,N_9128);
or U12735 (N_12735,N_5048,N_6590);
nand U12736 (N_12736,N_5700,N_9971);
nor U12737 (N_12737,N_5804,N_8840);
nor U12738 (N_12738,N_5831,N_7750);
nand U12739 (N_12739,N_8546,N_8520);
nor U12740 (N_12740,N_5569,N_7104);
xor U12741 (N_12741,N_9263,N_5342);
and U12742 (N_12742,N_9449,N_5968);
nor U12743 (N_12743,N_9792,N_6187);
and U12744 (N_12744,N_7651,N_7917);
or U12745 (N_12745,N_8035,N_8020);
and U12746 (N_12746,N_8427,N_7251);
or U12747 (N_12747,N_9129,N_7750);
nor U12748 (N_12748,N_6175,N_9279);
or U12749 (N_12749,N_5498,N_8188);
xnor U12750 (N_12750,N_9809,N_5403);
nor U12751 (N_12751,N_8866,N_8807);
nand U12752 (N_12752,N_7687,N_5230);
and U12753 (N_12753,N_8765,N_6530);
nor U12754 (N_12754,N_8139,N_5062);
or U12755 (N_12755,N_6265,N_7012);
nand U12756 (N_12756,N_7158,N_8985);
and U12757 (N_12757,N_8981,N_6510);
nor U12758 (N_12758,N_6685,N_7760);
and U12759 (N_12759,N_6511,N_5558);
or U12760 (N_12760,N_5357,N_6862);
nand U12761 (N_12761,N_7766,N_7774);
nor U12762 (N_12762,N_8021,N_9863);
and U12763 (N_12763,N_9167,N_7949);
or U12764 (N_12764,N_6605,N_8591);
xor U12765 (N_12765,N_8030,N_9940);
and U12766 (N_12766,N_7471,N_7290);
or U12767 (N_12767,N_5060,N_6655);
xor U12768 (N_12768,N_8083,N_7801);
nand U12769 (N_12769,N_5742,N_6952);
and U12770 (N_12770,N_9627,N_9321);
or U12771 (N_12771,N_7026,N_7548);
or U12772 (N_12772,N_9761,N_7374);
and U12773 (N_12773,N_9859,N_7225);
and U12774 (N_12774,N_5028,N_9539);
and U12775 (N_12775,N_6386,N_7784);
xor U12776 (N_12776,N_8330,N_6244);
nand U12777 (N_12777,N_6644,N_8886);
xor U12778 (N_12778,N_8385,N_9744);
nand U12779 (N_12779,N_8587,N_6509);
and U12780 (N_12780,N_5141,N_7700);
nand U12781 (N_12781,N_9434,N_6208);
nor U12782 (N_12782,N_9522,N_8471);
nand U12783 (N_12783,N_8141,N_9219);
nand U12784 (N_12784,N_6214,N_5132);
xnor U12785 (N_12785,N_6557,N_9724);
or U12786 (N_12786,N_9482,N_7722);
nor U12787 (N_12787,N_7775,N_5343);
and U12788 (N_12788,N_9941,N_6318);
xnor U12789 (N_12789,N_7021,N_6652);
nor U12790 (N_12790,N_5035,N_9687);
xnor U12791 (N_12791,N_9108,N_6135);
or U12792 (N_12792,N_5928,N_7561);
and U12793 (N_12793,N_9915,N_8047);
nand U12794 (N_12794,N_6240,N_5799);
nor U12795 (N_12795,N_7675,N_7490);
nand U12796 (N_12796,N_8976,N_6918);
or U12797 (N_12797,N_5913,N_5735);
xor U12798 (N_12798,N_8040,N_7589);
nand U12799 (N_12799,N_9396,N_5018);
nor U12800 (N_12800,N_5915,N_7518);
nor U12801 (N_12801,N_7477,N_8528);
nand U12802 (N_12802,N_8376,N_6932);
and U12803 (N_12803,N_5474,N_9919);
or U12804 (N_12804,N_5669,N_9610);
xnor U12805 (N_12805,N_7644,N_9635);
nand U12806 (N_12806,N_7385,N_8836);
nor U12807 (N_12807,N_9650,N_7588);
nand U12808 (N_12808,N_8239,N_9832);
and U12809 (N_12809,N_8451,N_8741);
or U12810 (N_12810,N_9335,N_8091);
nor U12811 (N_12811,N_7148,N_6010);
nor U12812 (N_12812,N_5483,N_5044);
and U12813 (N_12813,N_6738,N_9804);
nor U12814 (N_12814,N_8105,N_9053);
nand U12815 (N_12815,N_6810,N_6419);
xnor U12816 (N_12816,N_8043,N_6467);
or U12817 (N_12817,N_7313,N_7270);
nor U12818 (N_12818,N_5146,N_5914);
and U12819 (N_12819,N_7123,N_5746);
nand U12820 (N_12820,N_6349,N_6386);
or U12821 (N_12821,N_8184,N_6494);
nor U12822 (N_12822,N_7499,N_7060);
and U12823 (N_12823,N_6731,N_9877);
and U12824 (N_12824,N_7662,N_5186);
xnor U12825 (N_12825,N_8658,N_8132);
and U12826 (N_12826,N_5174,N_5572);
nand U12827 (N_12827,N_8323,N_5439);
and U12828 (N_12828,N_8557,N_7662);
or U12829 (N_12829,N_5771,N_6772);
nor U12830 (N_12830,N_7780,N_8206);
nor U12831 (N_12831,N_7330,N_5790);
or U12832 (N_12832,N_9863,N_7034);
or U12833 (N_12833,N_6116,N_8340);
nand U12834 (N_12834,N_5560,N_9445);
and U12835 (N_12835,N_6136,N_6247);
nor U12836 (N_12836,N_8830,N_9025);
nor U12837 (N_12837,N_6778,N_6606);
nor U12838 (N_12838,N_7061,N_9921);
and U12839 (N_12839,N_7111,N_8438);
nand U12840 (N_12840,N_5044,N_7603);
and U12841 (N_12841,N_6442,N_6550);
nor U12842 (N_12842,N_6678,N_7971);
xnor U12843 (N_12843,N_7129,N_7577);
and U12844 (N_12844,N_5856,N_6090);
or U12845 (N_12845,N_8168,N_7405);
or U12846 (N_12846,N_8800,N_6269);
nor U12847 (N_12847,N_6934,N_7700);
and U12848 (N_12848,N_8009,N_8322);
nand U12849 (N_12849,N_9495,N_7961);
or U12850 (N_12850,N_5945,N_8473);
or U12851 (N_12851,N_6706,N_6087);
nand U12852 (N_12852,N_6318,N_8803);
nand U12853 (N_12853,N_6488,N_6143);
nor U12854 (N_12854,N_6844,N_5641);
and U12855 (N_12855,N_8204,N_7753);
and U12856 (N_12856,N_8560,N_5468);
nor U12857 (N_12857,N_8986,N_9596);
nor U12858 (N_12858,N_6958,N_6556);
and U12859 (N_12859,N_9708,N_5133);
nand U12860 (N_12860,N_6605,N_9769);
nor U12861 (N_12861,N_6347,N_8066);
nor U12862 (N_12862,N_7820,N_5480);
and U12863 (N_12863,N_8341,N_6306);
or U12864 (N_12864,N_5997,N_9703);
and U12865 (N_12865,N_6363,N_9561);
or U12866 (N_12866,N_9390,N_8539);
xnor U12867 (N_12867,N_7342,N_8855);
or U12868 (N_12868,N_6965,N_6761);
nor U12869 (N_12869,N_9295,N_7380);
or U12870 (N_12870,N_7099,N_5373);
nand U12871 (N_12871,N_6526,N_5824);
nand U12872 (N_12872,N_8393,N_9551);
xnor U12873 (N_12873,N_8733,N_6296);
nor U12874 (N_12874,N_6988,N_9860);
nand U12875 (N_12875,N_9775,N_9430);
or U12876 (N_12876,N_8196,N_9094);
nor U12877 (N_12877,N_7018,N_6539);
and U12878 (N_12878,N_7309,N_9512);
and U12879 (N_12879,N_7670,N_7594);
nand U12880 (N_12880,N_5274,N_6753);
nor U12881 (N_12881,N_6036,N_8382);
nor U12882 (N_12882,N_6054,N_8548);
nor U12883 (N_12883,N_8345,N_9230);
nor U12884 (N_12884,N_6653,N_8439);
nor U12885 (N_12885,N_5162,N_6098);
nand U12886 (N_12886,N_5869,N_7900);
or U12887 (N_12887,N_5965,N_8211);
xnor U12888 (N_12888,N_9397,N_8051);
or U12889 (N_12889,N_5694,N_7802);
nor U12890 (N_12890,N_6546,N_9666);
nand U12891 (N_12891,N_8901,N_9160);
nor U12892 (N_12892,N_7332,N_9163);
nor U12893 (N_12893,N_6373,N_5665);
or U12894 (N_12894,N_8418,N_6785);
nand U12895 (N_12895,N_8805,N_8995);
nand U12896 (N_12896,N_5379,N_5711);
nand U12897 (N_12897,N_9052,N_7878);
nand U12898 (N_12898,N_8927,N_6656);
or U12899 (N_12899,N_9725,N_8892);
nand U12900 (N_12900,N_8751,N_8671);
and U12901 (N_12901,N_7352,N_9855);
nor U12902 (N_12902,N_9507,N_8521);
and U12903 (N_12903,N_5176,N_6723);
nor U12904 (N_12904,N_8302,N_7665);
nand U12905 (N_12905,N_7760,N_7864);
nand U12906 (N_12906,N_8115,N_9306);
xor U12907 (N_12907,N_9465,N_8527);
and U12908 (N_12908,N_7032,N_6523);
nor U12909 (N_12909,N_9498,N_6447);
nand U12910 (N_12910,N_7440,N_9343);
or U12911 (N_12911,N_5102,N_8582);
nand U12912 (N_12912,N_9687,N_7938);
or U12913 (N_12913,N_5199,N_6402);
nor U12914 (N_12914,N_7066,N_7113);
nand U12915 (N_12915,N_5536,N_9822);
nand U12916 (N_12916,N_5519,N_7150);
or U12917 (N_12917,N_8741,N_6384);
xnor U12918 (N_12918,N_9595,N_8996);
and U12919 (N_12919,N_8388,N_9537);
nand U12920 (N_12920,N_5644,N_5744);
nor U12921 (N_12921,N_9142,N_5466);
nor U12922 (N_12922,N_5101,N_7671);
nand U12923 (N_12923,N_9108,N_8374);
nand U12924 (N_12924,N_5010,N_9771);
nor U12925 (N_12925,N_5872,N_7280);
nor U12926 (N_12926,N_5931,N_8711);
and U12927 (N_12927,N_9523,N_6580);
nor U12928 (N_12928,N_8800,N_8798);
and U12929 (N_12929,N_5831,N_9485);
nor U12930 (N_12930,N_8368,N_9611);
xnor U12931 (N_12931,N_6021,N_8820);
nor U12932 (N_12932,N_5653,N_6294);
or U12933 (N_12933,N_5521,N_8252);
and U12934 (N_12934,N_9791,N_7232);
nand U12935 (N_12935,N_9824,N_6796);
nor U12936 (N_12936,N_6963,N_5055);
or U12937 (N_12937,N_9968,N_6679);
xnor U12938 (N_12938,N_9464,N_7117);
nor U12939 (N_12939,N_8103,N_5788);
or U12940 (N_12940,N_9860,N_6306);
nand U12941 (N_12941,N_9492,N_6730);
and U12942 (N_12942,N_8809,N_5778);
or U12943 (N_12943,N_6458,N_5026);
nor U12944 (N_12944,N_6996,N_5470);
or U12945 (N_12945,N_5931,N_7980);
nand U12946 (N_12946,N_9007,N_6938);
nand U12947 (N_12947,N_7684,N_6853);
nand U12948 (N_12948,N_9120,N_8996);
and U12949 (N_12949,N_7641,N_7924);
or U12950 (N_12950,N_6978,N_9943);
nor U12951 (N_12951,N_8470,N_7644);
nor U12952 (N_12952,N_9866,N_9749);
xnor U12953 (N_12953,N_8621,N_7450);
and U12954 (N_12954,N_5260,N_5354);
nor U12955 (N_12955,N_7162,N_9897);
nand U12956 (N_12956,N_6688,N_6316);
nand U12957 (N_12957,N_8087,N_9879);
nand U12958 (N_12958,N_8768,N_6199);
nor U12959 (N_12959,N_9424,N_6811);
or U12960 (N_12960,N_5046,N_6570);
or U12961 (N_12961,N_6525,N_8357);
nor U12962 (N_12962,N_8653,N_7064);
nor U12963 (N_12963,N_5038,N_9801);
nor U12964 (N_12964,N_6742,N_9607);
or U12965 (N_12965,N_5469,N_6114);
or U12966 (N_12966,N_7736,N_6852);
xnor U12967 (N_12967,N_6962,N_8223);
and U12968 (N_12968,N_7835,N_9662);
xnor U12969 (N_12969,N_7538,N_5549);
nand U12970 (N_12970,N_7865,N_8692);
nor U12971 (N_12971,N_5528,N_8212);
nand U12972 (N_12972,N_9785,N_7799);
nor U12973 (N_12973,N_5880,N_9688);
xnor U12974 (N_12974,N_8888,N_9422);
and U12975 (N_12975,N_9794,N_5641);
or U12976 (N_12976,N_8478,N_9104);
or U12977 (N_12977,N_7233,N_6533);
xnor U12978 (N_12978,N_6642,N_9422);
nor U12979 (N_12979,N_8230,N_8542);
nor U12980 (N_12980,N_7118,N_8958);
nand U12981 (N_12981,N_6470,N_9825);
or U12982 (N_12982,N_7492,N_7154);
xnor U12983 (N_12983,N_7437,N_8358);
nor U12984 (N_12984,N_8556,N_9462);
or U12985 (N_12985,N_6233,N_8524);
xnor U12986 (N_12986,N_9715,N_6357);
and U12987 (N_12987,N_8916,N_9170);
nand U12988 (N_12988,N_8169,N_9853);
nand U12989 (N_12989,N_8793,N_8602);
and U12990 (N_12990,N_7103,N_6618);
xor U12991 (N_12991,N_7995,N_5773);
nor U12992 (N_12992,N_7674,N_6827);
nand U12993 (N_12993,N_7173,N_6404);
or U12994 (N_12994,N_5612,N_5391);
or U12995 (N_12995,N_5449,N_5910);
nor U12996 (N_12996,N_7794,N_7756);
or U12997 (N_12997,N_6913,N_7600);
or U12998 (N_12998,N_8358,N_8407);
and U12999 (N_12999,N_7908,N_5832);
or U13000 (N_13000,N_6432,N_7639);
xor U13001 (N_13001,N_5339,N_9572);
nor U13002 (N_13002,N_7747,N_6442);
or U13003 (N_13003,N_6646,N_7837);
and U13004 (N_13004,N_8375,N_6743);
nand U13005 (N_13005,N_5506,N_6780);
nor U13006 (N_13006,N_8598,N_8329);
nor U13007 (N_13007,N_9679,N_8712);
and U13008 (N_13008,N_6411,N_7745);
or U13009 (N_13009,N_7936,N_8994);
nor U13010 (N_13010,N_7336,N_6436);
nand U13011 (N_13011,N_8703,N_5126);
nand U13012 (N_13012,N_7498,N_8115);
nand U13013 (N_13013,N_8485,N_7499);
nand U13014 (N_13014,N_6947,N_6022);
nand U13015 (N_13015,N_6444,N_5305);
nand U13016 (N_13016,N_6516,N_5017);
nor U13017 (N_13017,N_8367,N_6606);
or U13018 (N_13018,N_5135,N_5962);
or U13019 (N_13019,N_6558,N_9196);
or U13020 (N_13020,N_9429,N_6425);
nor U13021 (N_13021,N_8729,N_8238);
or U13022 (N_13022,N_7693,N_8671);
nand U13023 (N_13023,N_6686,N_7355);
or U13024 (N_13024,N_6055,N_5755);
xor U13025 (N_13025,N_5472,N_5319);
nand U13026 (N_13026,N_7091,N_8642);
nand U13027 (N_13027,N_8289,N_7209);
and U13028 (N_13028,N_8298,N_9867);
and U13029 (N_13029,N_9532,N_6775);
nand U13030 (N_13030,N_9715,N_8355);
and U13031 (N_13031,N_6163,N_9563);
nor U13032 (N_13032,N_6535,N_7694);
xor U13033 (N_13033,N_7438,N_7804);
nor U13034 (N_13034,N_8351,N_8655);
nor U13035 (N_13035,N_8430,N_6248);
nand U13036 (N_13036,N_5257,N_9835);
nor U13037 (N_13037,N_6317,N_9970);
nor U13038 (N_13038,N_8278,N_6308);
xnor U13039 (N_13039,N_9429,N_6147);
nand U13040 (N_13040,N_6183,N_9334);
or U13041 (N_13041,N_5842,N_9895);
and U13042 (N_13042,N_6674,N_9712);
nand U13043 (N_13043,N_5833,N_5904);
or U13044 (N_13044,N_5666,N_8033);
nand U13045 (N_13045,N_9562,N_7188);
xnor U13046 (N_13046,N_5379,N_9677);
and U13047 (N_13047,N_9014,N_9207);
or U13048 (N_13048,N_6407,N_8296);
and U13049 (N_13049,N_7900,N_7722);
xor U13050 (N_13050,N_5508,N_9178);
nor U13051 (N_13051,N_7749,N_6764);
nand U13052 (N_13052,N_5377,N_9533);
or U13053 (N_13053,N_8733,N_8639);
nand U13054 (N_13054,N_6169,N_9505);
or U13055 (N_13055,N_5434,N_5627);
nand U13056 (N_13056,N_8579,N_5296);
xor U13057 (N_13057,N_7847,N_7925);
or U13058 (N_13058,N_8177,N_5669);
nand U13059 (N_13059,N_7996,N_7430);
nor U13060 (N_13060,N_5869,N_9578);
or U13061 (N_13061,N_8301,N_8072);
or U13062 (N_13062,N_9556,N_5208);
and U13063 (N_13063,N_9783,N_9160);
nand U13064 (N_13064,N_6196,N_8653);
nand U13065 (N_13065,N_9501,N_9431);
or U13066 (N_13066,N_8967,N_7370);
or U13067 (N_13067,N_8391,N_9802);
nand U13068 (N_13068,N_9556,N_9703);
or U13069 (N_13069,N_8392,N_8724);
or U13070 (N_13070,N_8651,N_5640);
and U13071 (N_13071,N_9215,N_7988);
nand U13072 (N_13072,N_8806,N_8203);
nand U13073 (N_13073,N_6518,N_5391);
and U13074 (N_13074,N_7707,N_5673);
xnor U13075 (N_13075,N_5179,N_5701);
nand U13076 (N_13076,N_9325,N_7785);
or U13077 (N_13077,N_7948,N_6843);
or U13078 (N_13078,N_8751,N_9685);
nand U13079 (N_13079,N_7928,N_5908);
nand U13080 (N_13080,N_7126,N_6900);
or U13081 (N_13081,N_9438,N_9150);
or U13082 (N_13082,N_6457,N_6377);
nor U13083 (N_13083,N_9459,N_6345);
or U13084 (N_13084,N_9400,N_8206);
xor U13085 (N_13085,N_7903,N_6942);
and U13086 (N_13086,N_8618,N_8967);
and U13087 (N_13087,N_9852,N_5068);
and U13088 (N_13088,N_5595,N_6277);
nor U13089 (N_13089,N_6021,N_9671);
nor U13090 (N_13090,N_9205,N_9754);
or U13091 (N_13091,N_5182,N_9450);
nor U13092 (N_13092,N_7692,N_6977);
nand U13093 (N_13093,N_8649,N_7685);
xor U13094 (N_13094,N_9524,N_9377);
and U13095 (N_13095,N_9023,N_5857);
nand U13096 (N_13096,N_8896,N_8146);
or U13097 (N_13097,N_7630,N_7404);
and U13098 (N_13098,N_7684,N_8359);
nand U13099 (N_13099,N_5544,N_6637);
and U13100 (N_13100,N_5589,N_5259);
or U13101 (N_13101,N_5734,N_7391);
or U13102 (N_13102,N_8109,N_8382);
nand U13103 (N_13103,N_8816,N_5903);
xor U13104 (N_13104,N_8539,N_7910);
nand U13105 (N_13105,N_7424,N_6147);
or U13106 (N_13106,N_6979,N_7487);
nor U13107 (N_13107,N_7727,N_8465);
nor U13108 (N_13108,N_9558,N_7296);
nor U13109 (N_13109,N_6892,N_9290);
or U13110 (N_13110,N_8198,N_9067);
and U13111 (N_13111,N_7754,N_8709);
nand U13112 (N_13112,N_9318,N_8425);
nor U13113 (N_13113,N_5798,N_8263);
nor U13114 (N_13114,N_8317,N_8468);
nor U13115 (N_13115,N_6261,N_8319);
nor U13116 (N_13116,N_7999,N_6519);
xor U13117 (N_13117,N_7418,N_5588);
nand U13118 (N_13118,N_8351,N_7106);
xor U13119 (N_13119,N_5698,N_7663);
nand U13120 (N_13120,N_7423,N_7986);
nand U13121 (N_13121,N_8574,N_8141);
and U13122 (N_13122,N_9855,N_7995);
and U13123 (N_13123,N_9235,N_6655);
and U13124 (N_13124,N_7353,N_6892);
and U13125 (N_13125,N_5434,N_6189);
nor U13126 (N_13126,N_7835,N_7022);
nor U13127 (N_13127,N_6566,N_9659);
nand U13128 (N_13128,N_6439,N_5011);
or U13129 (N_13129,N_5410,N_5949);
and U13130 (N_13130,N_6023,N_6281);
nand U13131 (N_13131,N_9876,N_9527);
and U13132 (N_13132,N_9101,N_8176);
or U13133 (N_13133,N_7346,N_5013);
or U13134 (N_13134,N_6556,N_6468);
and U13135 (N_13135,N_7995,N_6976);
nor U13136 (N_13136,N_5517,N_9521);
xnor U13137 (N_13137,N_7130,N_8962);
nand U13138 (N_13138,N_5499,N_6003);
xor U13139 (N_13139,N_6647,N_9244);
nor U13140 (N_13140,N_7845,N_5997);
nand U13141 (N_13141,N_6599,N_9065);
and U13142 (N_13142,N_6253,N_9418);
and U13143 (N_13143,N_8060,N_7840);
or U13144 (N_13144,N_8678,N_6933);
nor U13145 (N_13145,N_7352,N_8386);
xnor U13146 (N_13146,N_5490,N_6316);
and U13147 (N_13147,N_9626,N_5841);
and U13148 (N_13148,N_6109,N_7825);
and U13149 (N_13149,N_6226,N_5009);
or U13150 (N_13150,N_5036,N_6078);
and U13151 (N_13151,N_9398,N_7530);
or U13152 (N_13152,N_7217,N_8163);
and U13153 (N_13153,N_8178,N_6566);
xnor U13154 (N_13154,N_8404,N_8138);
xnor U13155 (N_13155,N_5536,N_7828);
nand U13156 (N_13156,N_5127,N_9654);
xor U13157 (N_13157,N_5634,N_9816);
xnor U13158 (N_13158,N_9660,N_6861);
and U13159 (N_13159,N_7375,N_5708);
or U13160 (N_13160,N_5353,N_5659);
nor U13161 (N_13161,N_5236,N_6168);
nor U13162 (N_13162,N_6138,N_5812);
and U13163 (N_13163,N_9999,N_9721);
and U13164 (N_13164,N_6789,N_6803);
nand U13165 (N_13165,N_5398,N_9776);
nand U13166 (N_13166,N_8289,N_5959);
nor U13167 (N_13167,N_7836,N_7890);
nand U13168 (N_13168,N_6415,N_8845);
nor U13169 (N_13169,N_8260,N_8026);
xor U13170 (N_13170,N_6974,N_8317);
nor U13171 (N_13171,N_6060,N_5081);
xnor U13172 (N_13172,N_6397,N_5611);
or U13173 (N_13173,N_7518,N_9909);
nor U13174 (N_13174,N_8426,N_7740);
nor U13175 (N_13175,N_8831,N_9224);
xor U13176 (N_13176,N_8782,N_5310);
nand U13177 (N_13177,N_6756,N_7943);
nand U13178 (N_13178,N_8359,N_7263);
and U13179 (N_13179,N_5704,N_9482);
and U13180 (N_13180,N_6285,N_6273);
or U13181 (N_13181,N_9207,N_7393);
or U13182 (N_13182,N_6722,N_9120);
nor U13183 (N_13183,N_9238,N_7189);
nand U13184 (N_13184,N_6343,N_7416);
or U13185 (N_13185,N_9285,N_7773);
and U13186 (N_13186,N_7540,N_9831);
nand U13187 (N_13187,N_8280,N_6288);
nor U13188 (N_13188,N_8997,N_8193);
nand U13189 (N_13189,N_9777,N_8632);
nand U13190 (N_13190,N_5061,N_9755);
nor U13191 (N_13191,N_7213,N_8562);
nor U13192 (N_13192,N_8259,N_7276);
and U13193 (N_13193,N_8608,N_9151);
nor U13194 (N_13194,N_7205,N_9473);
nor U13195 (N_13195,N_9401,N_8705);
and U13196 (N_13196,N_6901,N_7210);
and U13197 (N_13197,N_5891,N_8253);
nand U13198 (N_13198,N_5048,N_8411);
nand U13199 (N_13199,N_7031,N_9628);
or U13200 (N_13200,N_8704,N_6561);
or U13201 (N_13201,N_9279,N_6274);
and U13202 (N_13202,N_7460,N_5184);
or U13203 (N_13203,N_6676,N_8928);
nand U13204 (N_13204,N_6269,N_5574);
nand U13205 (N_13205,N_7732,N_9822);
or U13206 (N_13206,N_5106,N_9864);
nand U13207 (N_13207,N_6305,N_5464);
nor U13208 (N_13208,N_9958,N_6792);
nand U13209 (N_13209,N_6359,N_7474);
xor U13210 (N_13210,N_7887,N_6646);
nand U13211 (N_13211,N_7422,N_8647);
nand U13212 (N_13212,N_5338,N_5630);
and U13213 (N_13213,N_7852,N_7738);
xnor U13214 (N_13214,N_5310,N_7817);
nor U13215 (N_13215,N_5404,N_7037);
nand U13216 (N_13216,N_5243,N_7553);
xnor U13217 (N_13217,N_7739,N_7017);
and U13218 (N_13218,N_7449,N_6638);
or U13219 (N_13219,N_6203,N_9382);
or U13220 (N_13220,N_5976,N_6250);
and U13221 (N_13221,N_5614,N_6168);
nand U13222 (N_13222,N_9788,N_9803);
and U13223 (N_13223,N_9466,N_9962);
nand U13224 (N_13224,N_6970,N_5614);
nand U13225 (N_13225,N_7132,N_8359);
xnor U13226 (N_13226,N_9239,N_8288);
nor U13227 (N_13227,N_7758,N_8842);
nor U13228 (N_13228,N_8035,N_5398);
nor U13229 (N_13229,N_7869,N_9376);
nand U13230 (N_13230,N_7918,N_5135);
or U13231 (N_13231,N_7004,N_6634);
nor U13232 (N_13232,N_5209,N_9935);
nor U13233 (N_13233,N_9292,N_6065);
or U13234 (N_13234,N_5924,N_9746);
nor U13235 (N_13235,N_6149,N_6438);
and U13236 (N_13236,N_7682,N_6165);
nand U13237 (N_13237,N_8251,N_7536);
and U13238 (N_13238,N_9626,N_5302);
nor U13239 (N_13239,N_5727,N_8994);
and U13240 (N_13240,N_7397,N_8690);
nand U13241 (N_13241,N_8700,N_7161);
nor U13242 (N_13242,N_7751,N_9536);
and U13243 (N_13243,N_9485,N_9165);
nand U13244 (N_13244,N_6938,N_7334);
and U13245 (N_13245,N_8347,N_5356);
and U13246 (N_13246,N_6390,N_7316);
nor U13247 (N_13247,N_8946,N_9118);
or U13248 (N_13248,N_7070,N_6148);
nand U13249 (N_13249,N_7162,N_7452);
or U13250 (N_13250,N_7746,N_9046);
nand U13251 (N_13251,N_6409,N_9408);
or U13252 (N_13252,N_8934,N_5629);
or U13253 (N_13253,N_7538,N_8478);
and U13254 (N_13254,N_5100,N_6724);
or U13255 (N_13255,N_7357,N_7844);
xnor U13256 (N_13256,N_7277,N_5667);
and U13257 (N_13257,N_6769,N_6014);
or U13258 (N_13258,N_9629,N_5842);
and U13259 (N_13259,N_9389,N_8157);
or U13260 (N_13260,N_8312,N_6126);
nor U13261 (N_13261,N_5737,N_8905);
or U13262 (N_13262,N_9158,N_5365);
nand U13263 (N_13263,N_9202,N_8361);
and U13264 (N_13264,N_5848,N_7086);
or U13265 (N_13265,N_9055,N_6601);
xor U13266 (N_13266,N_9451,N_5257);
nor U13267 (N_13267,N_5905,N_7527);
xnor U13268 (N_13268,N_7853,N_9965);
nor U13269 (N_13269,N_6472,N_6388);
nor U13270 (N_13270,N_8671,N_5486);
xnor U13271 (N_13271,N_5300,N_9632);
nand U13272 (N_13272,N_7182,N_8809);
nor U13273 (N_13273,N_9449,N_8713);
nand U13274 (N_13274,N_9305,N_7432);
or U13275 (N_13275,N_9745,N_5985);
nor U13276 (N_13276,N_7371,N_7148);
or U13277 (N_13277,N_8023,N_7577);
or U13278 (N_13278,N_8864,N_7530);
or U13279 (N_13279,N_9330,N_7478);
xnor U13280 (N_13280,N_6381,N_9317);
and U13281 (N_13281,N_7675,N_9390);
or U13282 (N_13282,N_6977,N_7536);
and U13283 (N_13283,N_6668,N_8370);
nor U13284 (N_13284,N_5387,N_8106);
xor U13285 (N_13285,N_9093,N_7287);
nand U13286 (N_13286,N_8143,N_6277);
nand U13287 (N_13287,N_7367,N_6408);
nor U13288 (N_13288,N_7297,N_9851);
nor U13289 (N_13289,N_6001,N_7562);
and U13290 (N_13290,N_6052,N_5575);
xnor U13291 (N_13291,N_5426,N_9856);
nand U13292 (N_13292,N_7488,N_7441);
nor U13293 (N_13293,N_7952,N_6023);
nand U13294 (N_13294,N_6631,N_9312);
or U13295 (N_13295,N_8713,N_6271);
nand U13296 (N_13296,N_8245,N_7067);
and U13297 (N_13297,N_5502,N_9531);
or U13298 (N_13298,N_8619,N_9376);
nand U13299 (N_13299,N_7496,N_8450);
nand U13300 (N_13300,N_6008,N_9364);
nor U13301 (N_13301,N_5970,N_7813);
nor U13302 (N_13302,N_7099,N_8906);
or U13303 (N_13303,N_8229,N_7813);
nand U13304 (N_13304,N_8367,N_9359);
and U13305 (N_13305,N_6473,N_6117);
nor U13306 (N_13306,N_7537,N_9692);
nor U13307 (N_13307,N_9465,N_8382);
and U13308 (N_13308,N_7881,N_8252);
nor U13309 (N_13309,N_6547,N_7307);
nor U13310 (N_13310,N_9615,N_9086);
or U13311 (N_13311,N_6178,N_7361);
or U13312 (N_13312,N_5375,N_8868);
and U13313 (N_13313,N_5916,N_9634);
nor U13314 (N_13314,N_7081,N_7018);
xor U13315 (N_13315,N_8164,N_6962);
nand U13316 (N_13316,N_8909,N_5724);
or U13317 (N_13317,N_9986,N_9981);
or U13318 (N_13318,N_7219,N_6983);
nand U13319 (N_13319,N_6344,N_8406);
and U13320 (N_13320,N_6328,N_8490);
nor U13321 (N_13321,N_9144,N_9780);
nand U13322 (N_13322,N_9088,N_8554);
nor U13323 (N_13323,N_6192,N_8283);
or U13324 (N_13324,N_8872,N_6244);
or U13325 (N_13325,N_5569,N_7644);
nor U13326 (N_13326,N_8444,N_5482);
and U13327 (N_13327,N_9611,N_7988);
nor U13328 (N_13328,N_9414,N_6169);
and U13329 (N_13329,N_7972,N_9592);
xnor U13330 (N_13330,N_5104,N_5891);
nor U13331 (N_13331,N_7120,N_6774);
or U13332 (N_13332,N_5730,N_5572);
or U13333 (N_13333,N_9115,N_6077);
nor U13334 (N_13334,N_5041,N_7315);
or U13335 (N_13335,N_8557,N_7065);
nand U13336 (N_13336,N_9709,N_8076);
and U13337 (N_13337,N_6227,N_8738);
nand U13338 (N_13338,N_9501,N_8815);
and U13339 (N_13339,N_6594,N_9953);
and U13340 (N_13340,N_8169,N_5033);
or U13341 (N_13341,N_8126,N_6828);
or U13342 (N_13342,N_6560,N_9534);
nor U13343 (N_13343,N_8671,N_8106);
xor U13344 (N_13344,N_5360,N_8028);
and U13345 (N_13345,N_6992,N_9577);
and U13346 (N_13346,N_9267,N_6883);
or U13347 (N_13347,N_8601,N_9645);
or U13348 (N_13348,N_6030,N_6154);
xnor U13349 (N_13349,N_7101,N_8272);
nand U13350 (N_13350,N_8219,N_5706);
nor U13351 (N_13351,N_5060,N_7056);
or U13352 (N_13352,N_7011,N_6611);
nor U13353 (N_13353,N_6461,N_6060);
xor U13354 (N_13354,N_6482,N_5608);
or U13355 (N_13355,N_5052,N_8531);
or U13356 (N_13356,N_5750,N_9530);
nor U13357 (N_13357,N_6974,N_9570);
nor U13358 (N_13358,N_7371,N_6160);
nor U13359 (N_13359,N_6936,N_7904);
or U13360 (N_13360,N_6168,N_6914);
nand U13361 (N_13361,N_7701,N_9612);
and U13362 (N_13362,N_6203,N_9826);
xor U13363 (N_13363,N_9028,N_8061);
nor U13364 (N_13364,N_5843,N_5373);
nor U13365 (N_13365,N_5898,N_9902);
and U13366 (N_13366,N_5706,N_6066);
nor U13367 (N_13367,N_9522,N_5396);
and U13368 (N_13368,N_7715,N_7925);
or U13369 (N_13369,N_9712,N_7347);
and U13370 (N_13370,N_7697,N_6936);
and U13371 (N_13371,N_8268,N_8954);
nand U13372 (N_13372,N_7594,N_8694);
xnor U13373 (N_13373,N_7768,N_5462);
nand U13374 (N_13374,N_5603,N_8532);
or U13375 (N_13375,N_8320,N_6448);
nor U13376 (N_13376,N_8508,N_9253);
nor U13377 (N_13377,N_9563,N_7758);
nor U13378 (N_13378,N_8393,N_7191);
nand U13379 (N_13379,N_6725,N_5608);
and U13380 (N_13380,N_7559,N_6232);
nand U13381 (N_13381,N_9288,N_8880);
or U13382 (N_13382,N_9691,N_5485);
xnor U13383 (N_13383,N_6162,N_8615);
and U13384 (N_13384,N_8865,N_6096);
nand U13385 (N_13385,N_7883,N_5451);
nand U13386 (N_13386,N_6925,N_5688);
nand U13387 (N_13387,N_7982,N_7043);
or U13388 (N_13388,N_9985,N_6913);
nor U13389 (N_13389,N_6221,N_6664);
nor U13390 (N_13390,N_7314,N_6814);
nor U13391 (N_13391,N_6885,N_5619);
nor U13392 (N_13392,N_6543,N_6583);
or U13393 (N_13393,N_6452,N_7636);
nand U13394 (N_13394,N_9341,N_6818);
and U13395 (N_13395,N_6195,N_9385);
nand U13396 (N_13396,N_5787,N_7735);
or U13397 (N_13397,N_8426,N_8535);
or U13398 (N_13398,N_5214,N_5191);
nor U13399 (N_13399,N_9406,N_9676);
and U13400 (N_13400,N_5261,N_5594);
nor U13401 (N_13401,N_6186,N_5495);
xnor U13402 (N_13402,N_9170,N_9885);
or U13403 (N_13403,N_5580,N_8941);
nor U13404 (N_13404,N_9021,N_7294);
xor U13405 (N_13405,N_8618,N_8605);
nand U13406 (N_13406,N_8380,N_9426);
or U13407 (N_13407,N_7841,N_8247);
or U13408 (N_13408,N_8220,N_8752);
or U13409 (N_13409,N_9245,N_9330);
nand U13410 (N_13410,N_8293,N_5408);
or U13411 (N_13411,N_8947,N_7804);
nand U13412 (N_13412,N_8111,N_8189);
nand U13413 (N_13413,N_5397,N_8574);
xnor U13414 (N_13414,N_7575,N_7765);
nand U13415 (N_13415,N_8665,N_7582);
or U13416 (N_13416,N_6667,N_7840);
nor U13417 (N_13417,N_7243,N_8934);
and U13418 (N_13418,N_8698,N_9890);
xnor U13419 (N_13419,N_6366,N_6199);
nor U13420 (N_13420,N_9579,N_5095);
nand U13421 (N_13421,N_6243,N_6411);
xnor U13422 (N_13422,N_8646,N_8264);
or U13423 (N_13423,N_8812,N_9705);
and U13424 (N_13424,N_7605,N_7183);
or U13425 (N_13425,N_6522,N_8494);
and U13426 (N_13426,N_8622,N_8116);
or U13427 (N_13427,N_5530,N_7201);
and U13428 (N_13428,N_6254,N_7980);
and U13429 (N_13429,N_8222,N_8576);
and U13430 (N_13430,N_8760,N_8515);
and U13431 (N_13431,N_7709,N_5219);
or U13432 (N_13432,N_9473,N_7429);
and U13433 (N_13433,N_9602,N_8085);
or U13434 (N_13434,N_7987,N_7290);
or U13435 (N_13435,N_8674,N_9934);
nand U13436 (N_13436,N_8624,N_9040);
nand U13437 (N_13437,N_9086,N_8202);
nand U13438 (N_13438,N_6504,N_8180);
or U13439 (N_13439,N_5345,N_8201);
or U13440 (N_13440,N_8981,N_6502);
nor U13441 (N_13441,N_7964,N_5384);
and U13442 (N_13442,N_8982,N_8413);
nand U13443 (N_13443,N_8952,N_6818);
nand U13444 (N_13444,N_5226,N_5017);
nand U13445 (N_13445,N_7144,N_9179);
nand U13446 (N_13446,N_8618,N_8473);
nand U13447 (N_13447,N_7304,N_8278);
nand U13448 (N_13448,N_7904,N_7441);
nor U13449 (N_13449,N_9780,N_6685);
or U13450 (N_13450,N_8480,N_9221);
and U13451 (N_13451,N_9097,N_7438);
and U13452 (N_13452,N_6268,N_6313);
nand U13453 (N_13453,N_8383,N_6770);
nor U13454 (N_13454,N_6299,N_9012);
and U13455 (N_13455,N_7609,N_9295);
or U13456 (N_13456,N_8038,N_5224);
and U13457 (N_13457,N_6909,N_9740);
nor U13458 (N_13458,N_8195,N_6232);
or U13459 (N_13459,N_8774,N_6319);
nor U13460 (N_13460,N_6147,N_5483);
nor U13461 (N_13461,N_7415,N_9009);
and U13462 (N_13462,N_7003,N_8729);
xor U13463 (N_13463,N_8081,N_5738);
nor U13464 (N_13464,N_6114,N_6689);
and U13465 (N_13465,N_9135,N_7987);
xor U13466 (N_13466,N_7673,N_7156);
nor U13467 (N_13467,N_6207,N_6620);
or U13468 (N_13468,N_5314,N_5873);
and U13469 (N_13469,N_5552,N_7528);
xor U13470 (N_13470,N_5137,N_6550);
or U13471 (N_13471,N_5374,N_8538);
nand U13472 (N_13472,N_7913,N_6327);
and U13473 (N_13473,N_8217,N_8677);
nor U13474 (N_13474,N_7259,N_5874);
nor U13475 (N_13475,N_8961,N_7657);
nor U13476 (N_13476,N_9458,N_5928);
or U13477 (N_13477,N_8941,N_9834);
nand U13478 (N_13478,N_8415,N_7595);
or U13479 (N_13479,N_8480,N_5985);
xnor U13480 (N_13480,N_7970,N_5688);
and U13481 (N_13481,N_5557,N_7835);
nand U13482 (N_13482,N_9842,N_8217);
and U13483 (N_13483,N_7901,N_5148);
xnor U13484 (N_13484,N_6964,N_7398);
or U13485 (N_13485,N_5051,N_8545);
or U13486 (N_13486,N_9799,N_8015);
and U13487 (N_13487,N_7724,N_9932);
nand U13488 (N_13488,N_9125,N_6346);
nor U13489 (N_13489,N_6450,N_8695);
nor U13490 (N_13490,N_6893,N_7482);
or U13491 (N_13491,N_6360,N_7441);
and U13492 (N_13492,N_7446,N_8036);
nand U13493 (N_13493,N_6916,N_5811);
nand U13494 (N_13494,N_9876,N_7943);
nor U13495 (N_13495,N_6910,N_9754);
nor U13496 (N_13496,N_8232,N_8746);
nor U13497 (N_13497,N_5450,N_6705);
nor U13498 (N_13498,N_5113,N_9416);
nor U13499 (N_13499,N_6439,N_5045);
and U13500 (N_13500,N_5139,N_6678);
xnor U13501 (N_13501,N_5903,N_9239);
nor U13502 (N_13502,N_6709,N_9088);
nand U13503 (N_13503,N_7437,N_9536);
or U13504 (N_13504,N_8608,N_9579);
and U13505 (N_13505,N_5778,N_8709);
or U13506 (N_13506,N_6323,N_9065);
nor U13507 (N_13507,N_5737,N_7417);
nand U13508 (N_13508,N_7595,N_9207);
nand U13509 (N_13509,N_9670,N_9535);
nor U13510 (N_13510,N_7464,N_9879);
nand U13511 (N_13511,N_8979,N_8660);
and U13512 (N_13512,N_5812,N_8534);
nor U13513 (N_13513,N_9110,N_9420);
nor U13514 (N_13514,N_5666,N_8742);
or U13515 (N_13515,N_9687,N_9694);
nand U13516 (N_13516,N_5755,N_6733);
nand U13517 (N_13517,N_7001,N_7939);
xor U13518 (N_13518,N_5144,N_7821);
nor U13519 (N_13519,N_8912,N_5463);
nand U13520 (N_13520,N_7488,N_6847);
nor U13521 (N_13521,N_6752,N_7170);
or U13522 (N_13522,N_8485,N_6099);
nand U13523 (N_13523,N_7390,N_6978);
and U13524 (N_13524,N_9212,N_9324);
nor U13525 (N_13525,N_5002,N_9275);
xor U13526 (N_13526,N_7998,N_7688);
or U13527 (N_13527,N_8915,N_9844);
nand U13528 (N_13528,N_6351,N_8264);
nand U13529 (N_13529,N_9824,N_9936);
and U13530 (N_13530,N_6273,N_9891);
and U13531 (N_13531,N_8614,N_9578);
nand U13532 (N_13532,N_9510,N_8856);
nand U13533 (N_13533,N_6068,N_5124);
and U13534 (N_13534,N_5124,N_8419);
nor U13535 (N_13535,N_7265,N_9967);
and U13536 (N_13536,N_5309,N_5494);
nand U13537 (N_13537,N_8193,N_8152);
nand U13538 (N_13538,N_5088,N_6827);
xor U13539 (N_13539,N_7956,N_9488);
or U13540 (N_13540,N_7507,N_7981);
nor U13541 (N_13541,N_8122,N_9950);
or U13542 (N_13542,N_8208,N_5905);
nor U13543 (N_13543,N_7503,N_8276);
xor U13544 (N_13544,N_8526,N_7092);
nor U13545 (N_13545,N_7407,N_5201);
xor U13546 (N_13546,N_8876,N_6674);
nor U13547 (N_13547,N_6466,N_9966);
and U13548 (N_13548,N_6260,N_6688);
xor U13549 (N_13549,N_8990,N_7615);
nor U13550 (N_13550,N_8114,N_6230);
or U13551 (N_13551,N_9874,N_5277);
and U13552 (N_13552,N_6146,N_8935);
xnor U13553 (N_13553,N_5736,N_8379);
and U13554 (N_13554,N_8011,N_7361);
nor U13555 (N_13555,N_6711,N_6036);
nand U13556 (N_13556,N_9289,N_8092);
or U13557 (N_13557,N_9345,N_8968);
or U13558 (N_13558,N_6631,N_5187);
and U13559 (N_13559,N_5289,N_9865);
and U13560 (N_13560,N_6071,N_6713);
xor U13561 (N_13561,N_6116,N_8011);
and U13562 (N_13562,N_7446,N_8722);
or U13563 (N_13563,N_7243,N_9236);
nand U13564 (N_13564,N_7775,N_7689);
nor U13565 (N_13565,N_8940,N_5540);
or U13566 (N_13566,N_7935,N_7058);
or U13567 (N_13567,N_6515,N_5394);
and U13568 (N_13568,N_9799,N_5441);
or U13569 (N_13569,N_6929,N_7131);
and U13570 (N_13570,N_9867,N_6716);
nand U13571 (N_13571,N_5180,N_5496);
nand U13572 (N_13572,N_9225,N_8560);
nand U13573 (N_13573,N_6036,N_9637);
nor U13574 (N_13574,N_5283,N_5359);
and U13575 (N_13575,N_9552,N_7531);
or U13576 (N_13576,N_6384,N_6777);
or U13577 (N_13577,N_6234,N_6265);
and U13578 (N_13578,N_8266,N_6056);
or U13579 (N_13579,N_6411,N_5363);
nand U13580 (N_13580,N_6999,N_7979);
nand U13581 (N_13581,N_7151,N_8008);
xnor U13582 (N_13582,N_6671,N_5162);
and U13583 (N_13583,N_8321,N_6328);
and U13584 (N_13584,N_9213,N_7624);
nand U13585 (N_13585,N_7351,N_7993);
nor U13586 (N_13586,N_6280,N_8159);
or U13587 (N_13587,N_5804,N_8681);
nor U13588 (N_13588,N_9409,N_8976);
nand U13589 (N_13589,N_7088,N_6274);
nor U13590 (N_13590,N_9628,N_8042);
and U13591 (N_13591,N_8752,N_6110);
nand U13592 (N_13592,N_6954,N_6115);
nor U13593 (N_13593,N_6921,N_9465);
nand U13594 (N_13594,N_6883,N_6090);
or U13595 (N_13595,N_5750,N_5391);
xor U13596 (N_13596,N_7613,N_6060);
xor U13597 (N_13597,N_7720,N_7350);
or U13598 (N_13598,N_7227,N_6629);
or U13599 (N_13599,N_6002,N_6895);
or U13600 (N_13600,N_7122,N_7448);
nand U13601 (N_13601,N_6953,N_6918);
nand U13602 (N_13602,N_6931,N_6334);
nand U13603 (N_13603,N_5498,N_8917);
and U13604 (N_13604,N_8141,N_5826);
xnor U13605 (N_13605,N_5662,N_6835);
nor U13606 (N_13606,N_9204,N_6138);
or U13607 (N_13607,N_5487,N_5744);
and U13608 (N_13608,N_8763,N_5871);
and U13609 (N_13609,N_9402,N_6169);
and U13610 (N_13610,N_5350,N_5225);
and U13611 (N_13611,N_8958,N_7321);
nand U13612 (N_13612,N_8411,N_7206);
nand U13613 (N_13613,N_7373,N_5502);
and U13614 (N_13614,N_5415,N_7626);
nand U13615 (N_13615,N_9737,N_5998);
nand U13616 (N_13616,N_7410,N_8355);
xor U13617 (N_13617,N_5231,N_8635);
nand U13618 (N_13618,N_6683,N_9821);
or U13619 (N_13619,N_9826,N_5549);
nand U13620 (N_13620,N_9044,N_8808);
or U13621 (N_13621,N_5215,N_6777);
nand U13622 (N_13622,N_8694,N_8340);
or U13623 (N_13623,N_7898,N_8617);
or U13624 (N_13624,N_6197,N_8207);
and U13625 (N_13625,N_9623,N_6819);
nor U13626 (N_13626,N_5182,N_6814);
or U13627 (N_13627,N_8822,N_8308);
and U13628 (N_13628,N_9957,N_9077);
xor U13629 (N_13629,N_5065,N_8754);
nor U13630 (N_13630,N_7320,N_6002);
nor U13631 (N_13631,N_7374,N_5619);
or U13632 (N_13632,N_7205,N_5029);
and U13633 (N_13633,N_8843,N_9422);
nor U13634 (N_13634,N_7412,N_7475);
or U13635 (N_13635,N_5364,N_5072);
nor U13636 (N_13636,N_9784,N_5337);
or U13637 (N_13637,N_6878,N_9452);
xnor U13638 (N_13638,N_5668,N_7752);
and U13639 (N_13639,N_5374,N_9750);
nand U13640 (N_13640,N_5637,N_5816);
and U13641 (N_13641,N_8102,N_8464);
or U13642 (N_13642,N_8437,N_6162);
nor U13643 (N_13643,N_9645,N_9634);
and U13644 (N_13644,N_7938,N_5493);
xnor U13645 (N_13645,N_5007,N_9462);
nand U13646 (N_13646,N_7077,N_9680);
and U13647 (N_13647,N_9734,N_7183);
xnor U13648 (N_13648,N_9249,N_9472);
nand U13649 (N_13649,N_6815,N_5599);
nor U13650 (N_13650,N_5087,N_8701);
nor U13651 (N_13651,N_9666,N_5400);
nand U13652 (N_13652,N_8962,N_6558);
nand U13653 (N_13653,N_8815,N_7121);
nor U13654 (N_13654,N_6671,N_8502);
nand U13655 (N_13655,N_8776,N_7846);
xnor U13656 (N_13656,N_6615,N_9299);
nand U13657 (N_13657,N_7194,N_7679);
and U13658 (N_13658,N_9500,N_6600);
nor U13659 (N_13659,N_9824,N_5095);
and U13660 (N_13660,N_6422,N_9537);
xor U13661 (N_13661,N_6348,N_8133);
or U13662 (N_13662,N_5219,N_6146);
and U13663 (N_13663,N_6629,N_9344);
and U13664 (N_13664,N_7058,N_5987);
nor U13665 (N_13665,N_9566,N_8894);
and U13666 (N_13666,N_5257,N_8407);
nand U13667 (N_13667,N_5633,N_7598);
and U13668 (N_13668,N_7539,N_6983);
or U13669 (N_13669,N_5753,N_8523);
nor U13670 (N_13670,N_7498,N_6954);
nand U13671 (N_13671,N_7759,N_8651);
and U13672 (N_13672,N_9304,N_6663);
nor U13673 (N_13673,N_5203,N_7668);
nand U13674 (N_13674,N_5288,N_9111);
nor U13675 (N_13675,N_6662,N_5387);
nor U13676 (N_13676,N_7652,N_6515);
nor U13677 (N_13677,N_8453,N_8291);
nand U13678 (N_13678,N_5858,N_7502);
nor U13679 (N_13679,N_5334,N_6995);
and U13680 (N_13680,N_9245,N_7077);
nor U13681 (N_13681,N_5026,N_7586);
nor U13682 (N_13682,N_8035,N_8450);
xnor U13683 (N_13683,N_6718,N_6129);
nand U13684 (N_13684,N_7079,N_6867);
nand U13685 (N_13685,N_5742,N_6655);
and U13686 (N_13686,N_6312,N_9691);
xor U13687 (N_13687,N_8572,N_7904);
nand U13688 (N_13688,N_6551,N_6674);
nor U13689 (N_13689,N_7997,N_9245);
nor U13690 (N_13690,N_7108,N_8474);
or U13691 (N_13691,N_8454,N_8630);
or U13692 (N_13692,N_8183,N_8125);
nand U13693 (N_13693,N_8089,N_9550);
nand U13694 (N_13694,N_7789,N_9671);
nand U13695 (N_13695,N_9209,N_7759);
nor U13696 (N_13696,N_7654,N_6642);
or U13697 (N_13697,N_9478,N_8814);
or U13698 (N_13698,N_5704,N_6844);
nor U13699 (N_13699,N_5838,N_9907);
nand U13700 (N_13700,N_9344,N_5166);
nand U13701 (N_13701,N_7440,N_6579);
nand U13702 (N_13702,N_9627,N_9453);
xnor U13703 (N_13703,N_7586,N_8605);
nand U13704 (N_13704,N_5377,N_8725);
or U13705 (N_13705,N_5325,N_6149);
nand U13706 (N_13706,N_6933,N_9107);
or U13707 (N_13707,N_7247,N_5180);
nor U13708 (N_13708,N_8228,N_7107);
xor U13709 (N_13709,N_6972,N_7036);
nor U13710 (N_13710,N_6735,N_9993);
or U13711 (N_13711,N_9082,N_6736);
or U13712 (N_13712,N_5874,N_7097);
nand U13713 (N_13713,N_6843,N_6775);
xor U13714 (N_13714,N_8198,N_7437);
or U13715 (N_13715,N_9328,N_8743);
nor U13716 (N_13716,N_5318,N_9114);
nand U13717 (N_13717,N_8343,N_7793);
nor U13718 (N_13718,N_8229,N_9531);
nand U13719 (N_13719,N_8234,N_9059);
nor U13720 (N_13720,N_9188,N_9401);
nand U13721 (N_13721,N_7441,N_9107);
xnor U13722 (N_13722,N_6692,N_5372);
or U13723 (N_13723,N_7809,N_8106);
and U13724 (N_13724,N_9347,N_9600);
and U13725 (N_13725,N_8323,N_7540);
nor U13726 (N_13726,N_5163,N_6581);
or U13727 (N_13727,N_7613,N_9329);
nand U13728 (N_13728,N_5626,N_9004);
and U13729 (N_13729,N_8168,N_5064);
nand U13730 (N_13730,N_5598,N_5290);
and U13731 (N_13731,N_9741,N_9945);
or U13732 (N_13732,N_7510,N_6360);
nand U13733 (N_13733,N_8010,N_9493);
and U13734 (N_13734,N_6786,N_9189);
nor U13735 (N_13735,N_6854,N_7789);
nor U13736 (N_13736,N_8523,N_5930);
or U13737 (N_13737,N_9252,N_5854);
nand U13738 (N_13738,N_7209,N_5647);
xor U13739 (N_13739,N_9859,N_6527);
xor U13740 (N_13740,N_5419,N_9130);
nand U13741 (N_13741,N_7961,N_7439);
and U13742 (N_13742,N_7790,N_8413);
and U13743 (N_13743,N_8260,N_7459);
and U13744 (N_13744,N_7384,N_8798);
nor U13745 (N_13745,N_7491,N_5265);
and U13746 (N_13746,N_9691,N_6113);
nor U13747 (N_13747,N_5559,N_8750);
or U13748 (N_13748,N_8564,N_5325);
xnor U13749 (N_13749,N_5400,N_8096);
nand U13750 (N_13750,N_7764,N_7538);
and U13751 (N_13751,N_8840,N_9435);
or U13752 (N_13752,N_9866,N_5007);
nor U13753 (N_13753,N_8406,N_7258);
nand U13754 (N_13754,N_5331,N_6342);
nor U13755 (N_13755,N_8282,N_6953);
or U13756 (N_13756,N_7928,N_7048);
and U13757 (N_13757,N_5104,N_9812);
nor U13758 (N_13758,N_5719,N_7511);
or U13759 (N_13759,N_8963,N_5590);
and U13760 (N_13760,N_7928,N_7257);
and U13761 (N_13761,N_5850,N_6870);
and U13762 (N_13762,N_8946,N_9465);
nor U13763 (N_13763,N_5618,N_9457);
and U13764 (N_13764,N_5176,N_5722);
or U13765 (N_13765,N_7858,N_6309);
or U13766 (N_13766,N_9614,N_9966);
or U13767 (N_13767,N_7680,N_5092);
nor U13768 (N_13768,N_7507,N_9028);
nor U13769 (N_13769,N_6076,N_5689);
nand U13770 (N_13770,N_5450,N_7202);
nand U13771 (N_13771,N_5601,N_7693);
or U13772 (N_13772,N_8276,N_6354);
nand U13773 (N_13773,N_8286,N_5195);
and U13774 (N_13774,N_9358,N_5076);
or U13775 (N_13775,N_8301,N_6931);
nand U13776 (N_13776,N_5447,N_5036);
and U13777 (N_13777,N_9768,N_9648);
nand U13778 (N_13778,N_9779,N_7914);
or U13779 (N_13779,N_6275,N_9280);
and U13780 (N_13780,N_6812,N_6786);
or U13781 (N_13781,N_7704,N_8772);
and U13782 (N_13782,N_5511,N_5776);
nor U13783 (N_13783,N_5776,N_9293);
nand U13784 (N_13784,N_6908,N_8328);
nor U13785 (N_13785,N_8103,N_5137);
and U13786 (N_13786,N_7447,N_8399);
nand U13787 (N_13787,N_8450,N_5607);
and U13788 (N_13788,N_9316,N_9038);
xnor U13789 (N_13789,N_9020,N_9845);
nor U13790 (N_13790,N_9631,N_8319);
nor U13791 (N_13791,N_6004,N_5328);
nor U13792 (N_13792,N_7896,N_8967);
nor U13793 (N_13793,N_5751,N_9762);
nand U13794 (N_13794,N_6903,N_5087);
or U13795 (N_13795,N_6464,N_9288);
nor U13796 (N_13796,N_9788,N_6022);
nand U13797 (N_13797,N_5186,N_7267);
and U13798 (N_13798,N_8828,N_6527);
or U13799 (N_13799,N_7294,N_8188);
or U13800 (N_13800,N_8330,N_6607);
nand U13801 (N_13801,N_7590,N_5156);
and U13802 (N_13802,N_6856,N_7426);
nand U13803 (N_13803,N_8573,N_8449);
nand U13804 (N_13804,N_9347,N_9327);
nand U13805 (N_13805,N_9851,N_8447);
nand U13806 (N_13806,N_9738,N_8624);
nand U13807 (N_13807,N_5520,N_7747);
nand U13808 (N_13808,N_9134,N_8954);
nor U13809 (N_13809,N_9166,N_5149);
and U13810 (N_13810,N_9080,N_9283);
nand U13811 (N_13811,N_6316,N_5714);
nor U13812 (N_13812,N_5895,N_9978);
nor U13813 (N_13813,N_7851,N_5762);
nor U13814 (N_13814,N_5845,N_6908);
nand U13815 (N_13815,N_8829,N_9741);
nor U13816 (N_13816,N_9844,N_7420);
or U13817 (N_13817,N_9095,N_7148);
nor U13818 (N_13818,N_9522,N_7715);
nand U13819 (N_13819,N_7442,N_8459);
or U13820 (N_13820,N_7578,N_7750);
nor U13821 (N_13821,N_9760,N_7700);
nor U13822 (N_13822,N_6030,N_8044);
xor U13823 (N_13823,N_9564,N_6758);
and U13824 (N_13824,N_9364,N_7975);
or U13825 (N_13825,N_8109,N_9654);
nand U13826 (N_13826,N_8546,N_6990);
and U13827 (N_13827,N_9304,N_5897);
nor U13828 (N_13828,N_8534,N_9956);
nand U13829 (N_13829,N_7164,N_7453);
xor U13830 (N_13830,N_9453,N_9771);
nor U13831 (N_13831,N_7976,N_9229);
and U13832 (N_13832,N_6259,N_6381);
or U13833 (N_13833,N_8565,N_7817);
or U13834 (N_13834,N_8011,N_6712);
nand U13835 (N_13835,N_8502,N_7812);
nor U13836 (N_13836,N_6529,N_5611);
xnor U13837 (N_13837,N_9523,N_8505);
nor U13838 (N_13838,N_9847,N_6925);
and U13839 (N_13839,N_6233,N_7560);
nand U13840 (N_13840,N_5999,N_6139);
xor U13841 (N_13841,N_6214,N_6118);
and U13842 (N_13842,N_6347,N_8956);
nand U13843 (N_13843,N_7685,N_6899);
and U13844 (N_13844,N_7109,N_5379);
xnor U13845 (N_13845,N_5643,N_5628);
nand U13846 (N_13846,N_5319,N_8722);
or U13847 (N_13847,N_9027,N_7790);
nor U13848 (N_13848,N_8466,N_7094);
nand U13849 (N_13849,N_9747,N_6611);
and U13850 (N_13850,N_6783,N_8124);
and U13851 (N_13851,N_7556,N_5023);
nand U13852 (N_13852,N_6782,N_7649);
nor U13853 (N_13853,N_6770,N_5229);
or U13854 (N_13854,N_7789,N_6660);
nor U13855 (N_13855,N_6929,N_5283);
nand U13856 (N_13856,N_7514,N_7314);
nand U13857 (N_13857,N_7173,N_5219);
nor U13858 (N_13858,N_7330,N_6677);
or U13859 (N_13859,N_7296,N_5914);
nand U13860 (N_13860,N_5143,N_9428);
nor U13861 (N_13861,N_8584,N_5679);
or U13862 (N_13862,N_6221,N_6586);
and U13863 (N_13863,N_6994,N_8097);
or U13864 (N_13864,N_5384,N_6177);
nor U13865 (N_13865,N_9166,N_5176);
xnor U13866 (N_13866,N_5650,N_6204);
or U13867 (N_13867,N_6744,N_6650);
nor U13868 (N_13868,N_7830,N_7691);
or U13869 (N_13869,N_7581,N_7526);
and U13870 (N_13870,N_6797,N_5754);
nand U13871 (N_13871,N_8202,N_5122);
nand U13872 (N_13872,N_5840,N_8613);
and U13873 (N_13873,N_8137,N_8492);
nor U13874 (N_13874,N_7071,N_6751);
and U13875 (N_13875,N_5438,N_5926);
nor U13876 (N_13876,N_7554,N_7075);
and U13877 (N_13877,N_9614,N_9835);
nor U13878 (N_13878,N_7330,N_6718);
nor U13879 (N_13879,N_7016,N_9039);
nor U13880 (N_13880,N_9693,N_7049);
xor U13881 (N_13881,N_8567,N_7426);
nor U13882 (N_13882,N_9559,N_9325);
xor U13883 (N_13883,N_9148,N_6544);
xor U13884 (N_13884,N_5273,N_8863);
nor U13885 (N_13885,N_6653,N_7179);
and U13886 (N_13886,N_9914,N_5063);
and U13887 (N_13887,N_6991,N_9487);
and U13888 (N_13888,N_6550,N_5357);
nor U13889 (N_13889,N_8426,N_7619);
nand U13890 (N_13890,N_6927,N_5292);
or U13891 (N_13891,N_9573,N_6180);
nand U13892 (N_13892,N_8623,N_6409);
nand U13893 (N_13893,N_9386,N_8095);
nor U13894 (N_13894,N_8816,N_5356);
nor U13895 (N_13895,N_9622,N_8074);
and U13896 (N_13896,N_7609,N_6215);
nor U13897 (N_13897,N_7370,N_7441);
and U13898 (N_13898,N_9442,N_7884);
xor U13899 (N_13899,N_5232,N_8258);
or U13900 (N_13900,N_5507,N_8532);
nor U13901 (N_13901,N_6502,N_8036);
nand U13902 (N_13902,N_8444,N_9359);
nor U13903 (N_13903,N_6952,N_5438);
and U13904 (N_13904,N_9867,N_6583);
or U13905 (N_13905,N_7640,N_5101);
or U13906 (N_13906,N_9945,N_8818);
and U13907 (N_13907,N_7075,N_6546);
nand U13908 (N_13908,N_9539,N_8035);
and U13909 (N_13909,N_6793,N_8656);
nor U13910 (N_13910,N_8118,N_6320);
nand U13911 (N_13911,N_7462,N_7703);
xnor U13912 (N_13912,N_6930,N_5616);
nand U13913 (N_13913,N_7816,N_5437);
and U13914 (N_13914,N_5731,N_6876);
nor U13915 (N_13915,N_7597,N_6039);
or U13916 (N_13916,N_5035,N_9858);
nor U13917 (N_13917,N_9496,N_5313);
xor U13918 (N_13918,N_9496,N_7892);
or U13919 (N_13919,N_8465,N_9989);
nand U13920 (N_13920,N_7473,N_8299);
nor U13921 (N_13921,N_7497,N_9674);
and U13922 (N_13922,N_9996,N_6349);
nor U13923 (N_13923,N_9919,N_6886);
nor U13924 (N_13924,N_7131,N_6157);
and U13925 (N_13925,N_9998,N_7770);
or U13926 (N_13926,N_7016,N_7099);
or U13927 (N_13927,N_6073,N_6270);
or U13928 (N_13928,N_9070,N_8074);
nor U13929 (N_13929,N_7817,N_7340);
xor U13930 (N_13930,N_5149,N_7811);
or U13931 (N_13931,N_5091,N_5819);
xor U13932 (N_13932,N_8573,N_7769);
nand U13933 (N_13933,N_7555,N_5412);
and U13934 (N_13934,N_5708,N_6288);
nand U13935 (N_13935,N_8257,N_7156);
nand U13936 (N_13936,N_9600,N_8273);
or U13937 (N_13937,N_6467,N_7990);
xor U13938 (N_13938,N_7135,N_5191);
nor U13939 (N_13939,N_7219,N_7285);
or U13940 (N_13940,N_5824,N_6612);
and U13941 (N_13941,N_8106,N_8773);
nor U13942 (N_13942,N_6786,N_8680);
or U13943 (N_13943,N_7944,N_7965);
xnor U13944 (N_13944,N_6009,N_8318);
xor U13945 (N_13945,N_6974,N_6089);
nor U13946 (N_13946,N_8053,N_6580);
nor U13947 (N_13947,N_7583,N_8298);
xnor U13948 (N_13948,N_7207,N_5167);
or U13949 (N_13949,N_9533,N_9852);
or U13950 (N_13950,N_7862,N_8000);
nor U13951 (N_13951,N_7899,N_6250);
and U13952 (N_13952,N_7266,N_8746);
and U13953 (N_13953,N_8477,N_7115);
nor U13954 (N_13954,N_7364,N_5467);
and U13955 (N_13955,N_8577,N_5032);
and U13956 (N_13956,N_9599,N_7312);
nand U13957 (N_13957,N_9478,N_8084);
or U13958 (N_13958,N_5310,N_9309);
and U13959 (N_13959,N_6024,N_5416);
nand U13960 (N_13960,N_8527,N_7295);
nand U13961 (N_13961,N_5012,N_7056);
or U13962 (N_13962,N_6005,N_7526);
nor U13963 (N_13963,N_7464,N_6069);
and U13964 (N_13964,N_7387,N_6468);
and U13965 (N_13965,N_6584,N_8036);
xnor U13966 (N_13966,N_9698,N_6366);
or U13967 (N_13967,N_8651,N_7000);
or U13968 (N_13968,N_5142,N_6155);
or U13969 (N_13969,N_9561,N_6851);
or U13970 (N_13970,N_5735,N_6002);
or U13971 (N_13971,N_9628,N_8837);
nor U13972 (N_13972,N_9902,N_9267);
nor U13973 (N_13973,N_6899,N_8578);
nand U13974 (N_13974,N_5652,N_8552);
xnor U13975 (N_13975,N_6796,N_7622);
nand U13976 (N_13976,N_6857,N_5462);
nand U13977 (N_13977,N_7545,N_5155);
nor U13978 (N_13978,N_5196,N_6795);
and U13979 (N_13979,N_8384,N_6884);
or U13980 (N_13980,N_5041,N_8695);
and U13981 (N_13981,N_6533,N_5091);
nand U13982 (N_13982,N_6650,N_6159);
or U13983 (N_13983,N_9837,N_9396);
or U13984 (N_13984,N_5709,N_9914);
and U13985 (N_13985,N_7818,N_9039);
nand U13986 (N_13986,N_6967,N_5838);
and U13987 (N_13987,N_6294,N_7809);
or U13988 (N_13988,N_5987,N_9131);
or U13989 (N_13989,N_9195,N_7284);
and U13990 (N_13990,N_5191,N_5706);
nand U13991 (N_13991,N_7500,N_5494);
or U13992 (N_13992,N_7303,N_5184);
and U13993 (N_13993,N_8171,N_8992);
or U13994 (N_13994,N_7542,N_7601);
nand U13995 (N_13995,N_8487,N_5660);
and U13996 (N_13996,N_6208,N_6913);
nand U13997 (N_13997,N_7832,N_6619);
and U13998 (N_13998,N_8496,N_8504);
nand U13999 (N_13999,N_5262,N_5297);
and U14000 (N_14000,N_9819,N_7172);
nor U14001 (N_14001,N_6341,N_5143);
or U14002 (N_14002,N_7459,N_9384);
and U14003 (N_14003,N_5013,N_9934);
nor U14004 (N_14004,N_8363,N_6141);
or U14005 (N_14005,N_6180,N_6407);
nand U14006 (N_14006,N_7740,N_8672);
nor U14007 (N_14007,N_7288,N_7566);
nor U14008 (N_14008,N_5848,N_6776);
nor U14009 (N_14009,N_7454,N_7396);
nand U14010 (N_14010,N_9136,N_5377);
nor U14011 (N_14011,N_6690,N_7048);
nor U14012 (N_14012,N_5526,N_8535);
and U14013 (N_14013,N_9174,N_6657);
nor U14014 (N_14014,N_6035,N_6806);
xnor U14015 (N_14015,N_9014,N_5803);
nor U14016 (N_14016,N_5966,N_8081);
and U14017 (N_14017,N_8865,N_8453);
nand U14018 (N_14018,N_9808,N_6945);
xor U14019 (N_14019,N_8576,N_7375);
nand U14020 (N_14020,N_6827,N_9834);
and U14021 (N_14021,N_7777,N_7179);
nor U14022 (N_14022,N_8318,N_8891);
and U14023 (N_14023,N_7827,N_8567);
and U14024 (N_14024,N_9302,N_6234);
nand U14025 (N_14025,N_9053,N_7278);
nor U14026 (N_14026,N_9940,N_7575);
nand U14027 (N_14027,N_7767,N_9633);
and U14028 (N_14028,N_5074,N_9003);
and U14029 (N_14029,N_7196,N_5737);
or U14030 (N_14030,N_7107,N_8581);
nand U14031 (N_14031,N_8459,N_5680);
nor U14032 (N_14032,N_7658,N_7116);
nand U14033 (N_14033,N_9291,N_5598);
nor U14034 (N_14034,N_5826,N_8925);
nor U14035 (N_14035,N_9274,N_6319);
nand U14036 (N_14036,N_6977,N_5297);
and U14037 (N_14037,N_5930,N_6617);
and U14038 (N_14038,N_6954,N_5417);
nand U14039 (N_14039,N_8743,N_6973);
nor U14040 (N_14040,N_6244,N_8656);
or U14041 (N_14041,N_6970,N_8343);
and U14042 (N_14042,N_6362,N_9002);
nor U14043 (N_14043,N_6282,N_8261);
and U14044 (N_14044,N_9547,N_7935);
nor U14045 (N_14045,N_9389,N_9532);
and U14046 (N_14046,N_9765,N_8561);
and U14047 (N_14047,N_5407,N_6130);
nand U14048 (N_14048,N_7222,N_7443);
nand U14049 (N_14049,N_8542,N_9572);
nand U14050 (N_14050,N_6059,N_5002);
or U14051 (N_14051,N_6021,N_8201);
or U14052 (N_14052,N_8855,N_8264);
nor U14053 (N_14053,N_9986,N_8929);
nor U14054 (N_14054,N_5911,N_6905);
or U14055 (N_14055,N_7378,N_7166);
nor U14056 (N_14056,N_6813,N_6721);
nor U14057 (N_14057,N_6347,N_9580);
nor U14058 (N_14058,N_6920,N_9354);
or U14059 (N_14059,N_7765,N_6039);
nor U14060 (N_14060,N_9339,N_6466);
or U14061 (N_14061,N_5419,N_5679);
and U14062 (N_14062,N_8542,N_5572);
or U14063 (N_14063,N_9911,N_5446);
or U14064 (N_14064,N_5092,N_7847);
xor U14065 (N_14065,N_9587,N_8809);
xnor U14066 (N_14066,N_5586,N_5843);
nor U14067 (N_14067,N_5212,N_6305);
or U14068 (N_14068,N_9328,N_6687);
nor U14069 (N_14069,N_6662,N_6918);
nand U14070 (N_14070,N_8292,N_5741);
nor U14071 (N_14071,N_7150,N_5207);
nand U14072 (N_14072,N_7231,N_5936);
and U14073 (N_14073,N_7490,N_6322);
nor U14074 (N_14074,N_8222,N_6375);
nand U14075 (N_14075,N_5164,N_6809);
nor U14076 (N_14076,N_5480,N_7249);
or U14077 (N_14077,N_8149,N_6676);
or U14078 (N_14078,N_6500,N_6491);
nor U14079 (N_14079,N_9920,N_5518);
nand U14080 (N_14080,N_6904,N_7565);
nor U14081 (N_14081,N_9927,N_7393);
nand U14082 (N_14082,N_9249,N_6305);
or U14083 (N_14083,N_8673,N_9491);
or U14084 (N_14084,N_8983,N_7718);
xor U14085 (N_14085,N_5712,N_7941);
nand U14086 (N_14086,N_5229,N_8586);
nand U14087 (N_14087,N_5647,N_8536);
xor U14088 (N_14088,N_8496,N_8253);
and U14089 (N_14089,N_7371,N_7924);
xnor U14090 (N_14090,N_6728,N_5127);
or U14091 (N_14091,N_6289,N_6031);
or U14092 (N_14092,N_5488,N_8919);
or U14093 (N_14093,N_9262,N_6125);
nand U14094 (N_14094,N_9386,N_6201);
nor U14095 (N_14095,N_8369,N_5719);
or U14096 (N_14096,N_8721,N_8457);
nor U14097 (N_14097,N_6766,N_7477);
and U14098 (N_14098,N_9870,N_6837);
nand U14099 (N_14099,N_5060,N_6612);
nor U14100 (N_14100,N_7045,N_9409);
nand U14101 (N_14101,N_5678,N_8241);
or U14102 (N_14102,N_5114,N_5256);
xor U14103 (N_14103,N_7921,N_6416);
nor U14104 (N_14104,N_5350,N_6538);
and U14105 (N_14105,N_9685,N_5699);
nand U14106 (N_14106,N_7649,N_9960);
nor U14107 (N_14107,N_5323,N_9563);
nor U14108 (N_14108,N_8982,N_7301);
or U14109 (N_14109,N_7383,N_9192);
nor U14110 (N_14110,N_5301,N_9966);
and U14111 (N_14111,N_9638,N_6173);
or U14112 (N_14112,N_7509,N_9119);
or U14113 (N_14113,N_7188,N_7391);
or U14114 (N_14114,N_8932,N_5417);
and U14115 (N_14115,N_6626,N_9141);
nand U14116 (N_14116,N_7953,N_8221);
and U14117 (N_14117,N_9805,N_5920);
nand U14118 (N_14118,N_8292,N_5023);
and U14119 (N_14119,N_6600,N_6363);
nand U14120 (N_14120,N_6740,N_6329);
and U14121 (N_14121,N_7120,N_8554);
nand U14122 (N_14122,N_6746,N_5780);
nor U14123 (N_14123,N_8398,N_5254);
and U14124 (N_14124,N_8617,N_9500);
and U14125 (N_14125,N_5850,N_9299);
nand U14126 (N_14126,N_5862,N_8185);
nand U14127 (N_14127,N_9939,N_5176);
or U14128 (N_14128,N_5670,N_9026);
or U14129 (N_14129,N_5578,N_5903);
or U14130 (N_14130,N_6715,N_8675);
or U14131 (N_14131,N_6212,N_7798);
or U14132 (N_14132,N_5202,N_7848);
and U14133 (N_14133,N_8999,N_6579);
nor U14134 (N_14134,N_9448,N_9885);
nor U14135 (N_14135,N_6447,N_9120);
nor U14136 (N_14136,N_5220,N_8254);
nor U14137 (N_14137,N_5830,N_9549);
nor U14138 (N_14138,N_7196,N_5595);
and U14139 (N_14139,N_9241,N_8522);
and U14140 (N_14140,N_8504,N_8097);
nor U14141 (N_14141,N_9314,N_7616);
or U14142 (N_14142,N_5271,N_9391);
nand U14143 (N_14143,N_6769,N_6673);
nand U14144 (N_14144,N_6958,N_7481);
and U14145 (N_14145,N_9029,N_8029);
nor U14146 (N_14146,N_8046,N_5918);
nor U14147 (N_14147,N_9081,N_6264);
nand U14148 (N_14148,N_5519,N_6944);
or U14149 (N_14149,N_5323,N_8536);
and U14150 (N_14150,N_6903,N_5418);
nor U14151 (N_14151,N_7931,N_5713);
nor U14152 (N_14152,N_9274,N_5973);
or U14153 (N_14153,N_8963,N_9729);
nand U14154 (N_14154,N_5078,N_8066);
nand U14155 (N_14155,N_9358,N_6382);
or U14156 (N_14156,N_5995,N_7049);
nand U14157 (N_14157,N_7038,N_5937);
nor U14158 (N_14158,N_8033,N_7282);
and U14159 (N_14159,N_5392,N_7564);
nor U14160 (N_14160,N_5722,N_6503);
and U14161 (N_14161,N_8159,N_6440);
or U14162 (N_14162,N_8019,N_6954);
nand U14163 (N_14163,N_9936,N_8440);
nor U14164 (N_14164,N_8627,N_7896);
and U14165 (N_14165,N_6417,N_7304);
xnor U14166 (N_14166,N_8272,N_6270);
nand U14167 (N_14167,N_5495,N_7034);
nand U14168 (N_14168,N_9833,N_6439);
nand U14169 (N_14169,N_7658,N_9224);
or U14170 (N_14170,N_9637,N_9008);
nand U14171 (N_14171,N_8363,N_6168);
nand U14172 (N_14172,N_9332,N_7563);
and U14173 (N_14173,N_7480,N_7520);
and U14174 (N_14174,N_8004,N_8813);
xnor U14175 (N_14175,N_9000,N_7977);
nor U14176 (N_14176,N_5555,N_7399);
or U14177 (N_14177,N_7727,N_7746);
and U14178 (N_14178,N_5224,N_9055);
and U14179 (N_14179,N_9497,N_5427);
or U14180 (N_14180,N_6975,N_5650);
and U14181 (N_14181,N_7931,N_7064);
and U14182 (N_14182,N_9045,N_9977);
nor U14183 (N_14183,N_9151,N_9713);
or U14184 (N_14184,N_7035,N_5207);
or U14185 (N_14185,N_6592,N_6484);
or U14186 (N_14186,N_8636,N_8158);
nand U14187 (N_14187,N_8980,N_7936);
nand U14188 (N_14188,N_9925,N_7388);
or U14189 (N_14189,N_6447,N_5469);
nor U14190 (N_14190,N_6318,N_7312);
xor U14191 (N_14191,N_9801,N_8950);
nand U14192 (N_14192,N_9215,N_9413);
nor U14193 (N_14193,N_8586,N_8862);
and U14194 (N_14194,N_8620,N_9396);
and U14195 (N_14195,N_5799,N_9524);
nand U14196 (N_14196,N_9934,N_8648);
nor U14197 (N_14197,N_6314,N_7885);
nand U14198 (N_14198,N_9735,N_5885);
or U14199 (N_14199,N_7264,N_6379);
nand U14200 (N_14200,N_5259,N_7247);
or U14201 (N_14201,N_9409,N_6930);
xor U14202 (N_14202,N_5256,N_8051);
nor U14203 (N_14203,N_8666,N_9671);
nor U14204 (N_14204,N_5399,N_8414);
nor U14205 (N_14205,N_8315,N_5888);
nor U14206 (N_14206,N_9253,N_5531);
nand U14207 (N_14207,N_7487,N_7565);
nor U14208 (N_14208,N_6556,N_9395);
nand U14209 (N_14209,N_7352,N_5260);
nand U14210 (N_14210,N_7389,N_8228);
or U14211 (N_14211,N_5493,N_6880);
nand U14212 (N_14212,N_6408,N_8881);
and U14213 (N_14213,N_5702,N_9408);
nand U14214 (N_14214,N_5637,N_8840);
and U14215 (N_14215,N_6007,N_8361);
and U14216 (N_14216,N_8987,N_9713);
nor U14217 (N_14217,N_8139,N_7167);
or U14218 (N_14218,N_8982,N_8252);
and U14219 (N_14219,N_9445,N_9191);
nand U14220 (N_14220,N_9960,N_8936);
nand U14221 (N_14221,N_8651,N_6126);
or U14222 (N_14222,N_6337,N_6941);
and U14223 (N_14223,N_7226,N_9911);
xnor U14224 (N_14224,N_8761,N_6484);
and U14225 (N_14225,N_8080,N_7159);
nor U14226 (N_14226,N_6231,N_8253);
nand U14227 (N_14227,N_8286,N_5696);
and U14228 (N_14228,N_9108,N_6253);
nor U14229 (N_14229,N_5414,N_9820);
nor U14230 (N_14230,N_7967,N_9674);
nand U14231 (N_14231,N_7134,N_6411);
nor U14232 (N_14232,N_5083,N_7486);
nor U14233 (N_14233,N_5394,N_7133);
and U14234 (N_14234,N_6015,N_7814);
or U14235 (N_14235,N_9400,N_8626);
and U14236 (N_14236,N_5910,N_6103);
or U14237 (N_14237,N_5611,N_8064);
or U14238 (N_14238,N_8500,N_6705);
or U14239 (N_14239,N_5051,N_5881);
nor U14240 (N_14240,N_7729,N_7516);
nor U14241 (N_14241,N_7421,N_8087);
nand U14242 (N_14242,N_6991,N_7827);
nand U14243 (N_14243,N_6386,N_9686);
xnor U14244 (N_14244,N_9086,N_8719);
xor U14245 (N_14245,N_9469,N_5643);
nor U14246 (N_14246,N_8372,N_9729);
and U14247 (N_14247,N_7338,N_7950);
nor U14248 (N_14248,N_5110,N_5991);
nand U14249 (N_14249,N_8316,N_5824);
or U14250 (N_14250,N_9052,N_5315);
nor U14251 (N_14251,N_9158,N_6142);
and U14252 (N_14252,N_9629,N_7130);
and U14253 (N_14253,N_7587,N_9390);
or U14254 (N_14254,N_8994,N_9631);
and U14255 (N_14255,N_5295,N_5044);
and U14256 (N_14256,N_5278,N_9236);
or U14257 (N_14257,N_6845,N_7392);
xor U14258 (N_14258,N_6254,N_9155);
xnor U14259 (N_14259,N_5606,N_6959);
or U14260 (N_14260,N_7985,N_8244);
xor U14261 (N_14261,N_8118,N_7057);
xor U14262 (N_14262,N_7562,N_9823);
nor U14263 (N_14263,N_7461,N_8496);
nand U14264 (N_14264,N_6766,N_6631);
nand U14265 (N_14265,N_8490,N_5377);
nor U14266 (N_14266,N_6937,N_9537);
nand U14267 (N_14267,N_6520,N_7857);
and U14268 (N_14268,N_7831,N_8097);
nand U14269 (N_14269,N_6672,N_8192);
nor U14270 (N_14270,N_9447,N_6235);
or U14271 (N_14271,N_8395,N_7533);
xnor U14272 (N_14272,N_9369,N_7104);
xor U14273 (N_14273,N_5241,N_8451);
nor U14274 (N_14274,N_8654,N_5173);
xnor U14275 (N_14275,N_6296,N_5641);
nor U14276 (N_14276,N_8371,N_8487);
and U14277 (N_14277,N_6129,N_6351);
nor U14278 (N_14278,N_9561,N_8514);
nand U14279 (N_14279,N_6304,N_5088);
and U14280 (N_14280,N_9688,N_6010);
or U14281 (N_14281,N_9336,N_6985);
nand U14282 (N_14282,N_7759,N_8250);
nand U14283 (N_14283,N_5372,N_5701);
nand U14284 (N_14284,N_8811,N_8473);
or U14285 (N_14285,N_6219,N_9856);
nand U14286 (N_14286,N_6208,N_9820);
nand U14287 (N_14287,N_7847,N_9380);
xnor U14288 (N_14288,N_5315,N_7553);
nand U14289 (N_14289,N_6323,N_7561);
and U14290 (N_14290,N_8533,N_8897);
nor U14291 (N_14291,N_7258,N_8737);
and U14292 (N_14292,N_5555,N_7667);
nand U14293 (N_14293,N_9980,N_8001);
nor U14294 (N_14294,N_9646,N_9134);
and U14295 (N_14295,N_6279,N_7486);
nand U14296 (N_14296,N_7404,N_5159);
and U14297 (N_14297,N_8599,N_7464);
or U14298 (N_14298,N_9583,N_7503);
and U14299 (N_14299,N_6247,N_9559);
xor U14300 (N_14300,N_8296,N_7384);
nor U14301 (N_14301,N_9830,N_8532);
and U14302 (N_14302,N_8782,N_5548);
nand U14303 (N_14303,N_6271,N_9777);
nor U14304 (N_14304,N_7667,N_6006);
nand U14305 (N_14305,N_7085,N_6831);
xnor U14306 (N_14306,N_5490,N_6508);
nor U14307 (N_14307,N_7628,N_7320);
nand U14308 (N_14308,N_5283,N_9294);
nand U14309 (N_14309,N_8930,N_6069);
and U14310 (N_14310,N_7839,N_9751);
or U14311 (N_14311,N_7015,N_7662);
nand U14312 (N_14312,N_6392,N_9414);
nand U14313 (N_14313,N_7679,N_5461);
xnor U14314 (N_14314,N_7174,N_5783);
and U14315 (N_14315,N_9800,N_9355);
nor U14316 (N_14316,N_5932,N_7328);
nor U14317 (N_14317,N_8852,N_5302);
nand U14318 (N_14318,N_8768,N_9847);
nand U14319 (N_14319,N_5748,N_5960);
and U14320 (N_14320,N_7685,N_6627);
or U14321 (N_14321,N_7169,N_6813);
xor U14322 (N_14322,N_9671,N_6355);
nand U14323 (N_14323,N_7274,N_7747);
and U14324 (N_14324,N_6308,N_7763);
and U14325 (N_14325,N_6716,N_9930);
nand U14326 (N_14326,N_6794,N_8609);
or U14327 (N_14327,N_7649,N_5161);
nand U14328 (N_14328,N_5290,N_8183);
nor U14329 (N_14329,N_5564,N_7375);
nand U14330 (N_14330,N_7416,N_9777);
nor U14331 (N_14331,N_6295,N_5264);
nor U14332 (N_14332,N_9826,N_7132);
and U14333 (N_14333,N_8910,N_7916);
or U14334 (N_14334,N_5545,N_5960);
nor U14335 (N_14335,N_7881,N_5009);
or U14336 (N_14336,N_8517,N_9487);
or U14337 (N_14337,N_6490,N_6737);
nand U14338 (N_14338,N_8367,N_5393);
xor U14339 (N_14339,N_6146,N_6041);
xnor U14340 (N_14340,N_6344,N_5009);
nor U14341 (N_14341,N_6639,N_9326);
or U14342 (N_14342,N_8502,N_8935);
xor U14343 (N_14343,N_5796,N_5867);
xor U14344 (N_14344,N_9913,N_8466);
and U14345 (N_14345,N_8963,N_5201);
nor U14346 (N_14346,N_7460,N_8507);
nor U14347 (N_14347,N_7896,N_7841);
nor U14348 (N_14348,N_8812,N_6851);
nor U14349 (N_14349,N_9327,N_6962);
and U14350 (N_14350,N_8550,N_5582);
or U14351 (N_14351,N_7667,N_7472);
xnor U14352 (N_14352,N_7494,N_6350);
nor U14353 (N_14353,N_6954,N_9993);
nor U14354 (N_14354,N_7161,N_8145);
nand U14355 (N_14355,N_8235,N_9254);
nor U14356 (N_14356,N_6418,N_5406);
or U14357 (N_14357,N_6245,N_6195);
and U14358 (N_14358,N_7208,N_5796);
or U14359 (N_14359,N_5631,N_9069);
nand U14360 (N_14360,N_6938,N_5139);
xnor U14361 (N_14361,N_7837,N_5329);
and U14362 (N_14362,N_6309,N_7296);
and U14363 (N_14363,N_9646,N_9933);
or U14364 (N_14364,N_7314,N_8395);
nand U14365 (N_14365,N_7642,N_9350);
or U14366 (N_14366,N_8523,N_9276);
nand U14367 (N_14367,N_9752,N_5680);
xor U14368 (N_14368,N_5055,N_7208);
nand U14369 (N_14369,N_5215,N_8715);
or U14370 (N_14370,N_5761,N_8949);
or U14371 (N_14371,N_5247,N_5801);
or U14372 (N_14372,N_9784,N_7749);
and U14373 (N_14373,N_8043,N_8602);
nand U14374 (N_14374,N_5068,N_5922);
nor U14375 (N_14375,N_6045,N_9915);
nor U14376 (N_14376,N_8069,N_9623);
nor U14377 (N_14377,N_5546,N_6373);
or U14378 (N_14378,N_8640,N_5935);
or U14379 (N_14379,N_7473,N_9585);
nand U14380 (N_14380,N_7197,N_9190);
nor U14381 (N_14381,N_6946,N_6072);
and U14382 (N_14382,N_8101,N_7904);
nor U14383 (N_14383,N_6738,N_9070);
and U14384 (N_14384,N_7645,N_7076);
xor U14385 (N_14385,N_9917,N_7642);
nor U14386 (N_14386,N_8138,N_8267);
and U14387 (N_14387,N_8706,N_7559);
nor U14388 (N_14388,N_5579,N_6241);
or U14389 (N_14389,N_5702,N_8954);
and U14390 (N_14390,N_9389,N_9912);
nand U14391 (N_14391,N_8938,N_8248);
xor U14392 (N_14392,N_7498,N_7021);
and U14393 (N_14393,N_9652,N_7440);
nand U14394 (N_14394,N_7427,N_9681);
nand U14395 (N_14395,N_6782,N_7536);
nand U14396 (N_14396,N_8607,N_5915);
and U14397 (N_14397,N_6709,N_7236);
nand U14398 (N_14398,N_8639,N_6877);
or U14399 (N_14399,N_6347,N_7097);
nor U14400 (N_14400,N_7535,N_8938);
and U14401 (N_14401,N_5216,N_5053);
nor U14402 (N_14402,N_8754,N_8477);
nand U14403 (N_14403,N_8348,N_7196);
or U14404 (N_14404,N_7170,N_9518);
nand U14405 (N_14405,N_6063,N_9590);
nand U14406 (N_14406,N_6662,N_8484);
and U14407 (N_14407,N_9187,N_7679);
or U14408 (N_14408,N_6453,N_8197);
or U14409 (N_14409,N_5862,N_7170);
nor U14410 (N_14410,N_8082,N_5310);
or U14411 (N_14411,N_7218,N_5486);
nand U14412 (N_14412,N_7894,N_6166);
or U14413 (N_14413,N_5820,N_9733);
nand U14414 (N_14414,N_5533,N_5086);
xnor U14415 (N_14415,N_6418,N_9703);
nor U14416 (N_14416,N_6490,N_9650);
and U14417 (N_14417,N_9982,N_7755);
nor U14418 (N_14418,N_9416,N_7746);
or U14419 (N_14419,N_5684,N_9779);
nor U14420 (N_14420,N_8818,N_6030);
and U14421 (N_14421,N_5969,N_6619);
nor U14422 (N_14422,N_6991,N_7466);
nand U14423 (N_14423,N_5488,N_8951);
nand U14424 (N_14424,N_8636,N_8193);
nand U14425 (N_14425,N_7001,N_6224);
nor U14426 (N_14426,N_7464,N_9956);
or U14427 (N_14427,N_5523,N_6483);
nand U14428 (N_14428,N_8318,N_7270);
nand U14429 (N_14429,N_5279,N_8974);
or U14430 (N_14430,N_6475,N_6220);
nor U14431 (N_14431,N_5139,N_5070);
nand U14432 (N_14432,N_5933,N_6607);
and U14433 (N_14433,N_6179,N_6161);
and U14434 (N_14434,N_6595,N_7882);
nor U14435 (N_14435,N_5905,N_8748);
and U14436 (N_14436,N_5579,N_8194);
or U14437 (N_14437,N_8930,N_9676);
or U14438 (N_14438,N_9192,N_9913);
and U14439 (N_14439,N_5959,N_8748);
or U14440 (N_14440,N_6197,N_9882);
or U14441 (N_14441,N_9957,N_9361);
and U14442 (N_14442,N_9689,N_6250);
nand U14443 (N_14443,N_6414,N_6391);
or U14444 (N_14444,N_8179,N_6145);
nor U14445 (N_14445,N_5610,N_5408);
or U14446 (N_14446,N_6129,N_9187);
nor U14447 (N_14447,N_7070,N_7764);
and U14448 (N_14448,N_5474,N_5551);
and U14449 (N_14449,N_7515,N_8506);
xor U14450 (N_14450,N_8145,N_5360);
or U14451 (N_14451,N_9439,N_8464);
nor U14452 (N_14452,N_5774,N_8411);
nor U14453 (N_14453,N_5469,N_6932);
or U14454 (N_14454,N_6291,N_9710);
and U14455 (N_14455,N_8060,N_7431);
and U14456 (N_14456,N_7185,N_6436);
nand U14457 (N_14457,N_5791,N_9639);
nor U14458 (N_14458,N_6811,N_6765);
and U14459 (N_14459,N_8607,N_9303);
and U14460 (N_14460,N_7922,N_5344);
or U14461 (N_14461,N_9462,N_6953);
or U14462 (N_14462,N_7110,N_9500);
nor U14463 (N_14463,N_9352,N_7348);
nor U14464 (N_14464,N_8781,N_8111);
nand U14465 (N_14465,N_6886,N_9387);
nor U14466 (N_14466,N_7392,N_9458);
nand U14467 (N_14467,N_5956,N_9492);
nor U14468 (N_14468,N_7073,N_9713);
nor U14469 (N_14469,N_6236,N_8959);
nor U14470 (N_14470,N_5677,N_5615);
nand U14471 (N_14471,N_6139,N_5846);
nand U14472 (N_14472,N_9120,N_5053);
xor U14473 (N_14473,N_5694,N_5096);
and U14474 (N_14474,N_5879,N_9929);
and U14475 (N_14475,N_7536,N_9292);
or U14476 (N_14476,N_9049,N_5724);
or U14477 (N_14477,N_8333,N_7809);
and U14478 (N_14478,N_8274,N_7152);
nand U14479 (N_14479,N_6715,N_6516);
nor U14480 (N_14480,N_7725,N_9931);
and U14481 (N_14481,N_7570,N_9274);
or U14482 (N_14482,N_6513,N_5081);
and U14483 (N_14483,N_5894,N_6817);
and U14484 (N_14484,N_7348,N_6226);
nand U14485 (N_14485,N_5004,N_5119);
nor U14486 (N_14486,N_7408,N_5217);
and U14487 (N_14487,N_9842,N_6874);
or U14488 (N_14488,N_9307,N_8739);
nand U14489 (N_14489,N_5065,N_6130);
or U14490 (N_14490,N_8894,N_9474);
or U14491 (N_14491,N_8638,N_8283);
or U14492 (N_14492,N_8071,N_5670);
and U14493 (N_14493,N_8232,N_7613);
and U14494 (N_14494,N_8628,N_8002);
or U14495 (N_14495,N_6320,N_5740);
or U14496 (N_14496,N_6305,N_6642);
nand U14497 (N_14497,N_5502,N_5349);
or U14498 (N_14498,N_7362,N_8769);
nand U14499 (N_14499,N_7060,N_5470);
nand U14500 (N_14500,N_9077,N_8521);
or U14501 (N_14501,N_5228,N_9147);
or U14502 (N_14502,N_7870,N_8145);
or U14503 (N_14503,N_7972,N_9675);
and U14504 (N_14504,N_5329,N_9577);
nor U14505 (N_14505,N_9002,N_6262);
xnor U14506 (N_14506,N_8310,N_9770);
xor U14507 (N_14507,N_8682,N_8321);
nor U14508 (N_14508,N_7033,N_8219);
nor U14509 (N_14509,N_9671,N_6947);
nor U14510 (N_14510,N_5151,N_6603);
and U14511 (N_14511,N_6532,N_5301);
and U14512 (N_14512,N_9127,N_5951);
nor U14513 (N_14513,N_5320,N_7516);
xnor U14514 (N_14514,N_5323,N_7155);
nand U14515 (N_14515,N_9720,N_8959);
and U14516 (N_14516,N_9925,N_9257);
or U14517 (N_14517,N_7647,N_7832);
and U14518 (N_14518,N_7092,N_6191);
nand U14519 (N_14519,N_6937,N_9331);
xnor U14520 (N_14520,N_9280,N_8613);
nand U14521 (N_14521,N_7752,N_9950);
or U14522 (N_14522,N_5917,N_7248);
nand U14523 (N_14523,N_7902,N_5572);
nor U14524 (N_14524,N_7069,N_7341);
nor U14525 (N_14525,N_9614,N_7132);
nand U14526 (N_14526,N_5971,N_7831);
and U14527 (N_14527,N_7127,N_7169);
or U14528 (N_14528,N_5123,N_8157);
and U14529 (N_14529,N_7110,N_5312);
nand U14530 (N_14530,N_6310,N_8691);
nand U14531 (N_14531,N_7374,N_6005);
nand U14532 (N_14532,N_9461,N_7473);
nand U14533 (N_14533,N_9763,N_6878);
or U14534 (N_14534,N_6327,N_6007);
nor U14535 (N_14535,N_6431,N_8731);
or U14536 (N_14536,N_8146,N_6008);
and U14537 (N_14537,N_6516,N_7199);
or U14538 (N_14538,N_9208,N_7062);
nor U14539 (N_14539,N_5870,N_8346);
or U14540 (N_14540,N_5426,N_6481);
nand U14541 (N_14541,N_7208,N_6025);
nand U14542 (N_14542,N_7332,N_7625);
or U14543 (N_14543,N_9220,N_6790);
or U14544 (N_14544,N_9075,N_8299);
xnor U14545 (N_14545,N_7699,N_8528);
and U14546 (N_14546,N_7932,N_5039);
or U14547 (N_14547,N_6388,N_6755);
nand U14548 (N_14548,N_7200,N_9225);
nor U14549 (N_14549,N_7656,N_5824);
or U14550 (N_14550,N_6852,N_5619);
and U14551 (N_14551,N_8538,N_5745);
nor U14552 (N_14552,N_9496,N_8856);
nor U14553 (N_14553,N_8642,N_5243);
and U14554 (N_14554,N_7900,N_5437);
nand U14555 (N_14555,N_7178,N_6157);
nor U14556 (N_14556,N_5894,N_8914);
or U14557 (N_14557,N_7915,N_5232);
nand U14558 (N_14558,N_6362,N_9622);
or U14559 (N_14559,N_9903,N_6461);
and U14560 (N_14560,N_8136,N_7537);
nor U14561 (N_14561,N_6714,N_7191);
or U14562 (N_14562,N_8665,N_7047);
and U14563 (N_14563,N_8529,N_7023);
or U14564 (N_14564,N_5478,N_5550);
and U14565 (N_14565,N_8430,N_6910);
and U14566 (N_14566,N_7635,N_9287);
xnor U14567 (N_14567,N_5889,N_6582);
nor U14568 (N_14568,N_7821,N_6771);
xor U14569 (N_14569,N_6235,N_5913);
nor U14570 (N_14570,N_6225,N_7914);
or U14571 (N_14571,N_6799,N_7334);
xnor U14572 (N_14572,N_8361,N_5692);
nor U14573 (N_14573,N_7109,N_9190);
or U14574 (N_14574,N_6507,N_5958);
nand U14575 (N_14575,N_7708,N_7955);
nand U14576 (N_14576,N_6390,N_9909);
nor U14577 (N_14577,N_5466,N_6329);
xnor U14578 (N_14578,N_8896,N_8369);
xor U14579 (N_14579,N_6872,N_8710);
or U14580 (N_14580,N_9061,N_6126);
xor U14581 (N_14581,N_7010,N_8817);
or U14582 (N_14582,N_9453,N_6926);
and U14583 (N_14583,N_5974,N_7223);
xor U14584 (N_14584,N_5735,N_9273);
nand U14585 (N_14585,N_5869,N_5846);
nand U14586 (N_14586,N_6622,N_6525);
and U14587 (N_14587,N_6740,N_8088);
or U14588 (N_14588,N_6341,N_8032);
nor U14589 (N_14589,N_7845,N_7683);
xor U14590 (N_14590,N_7612,N_5350);
and U14591 (N_14591,N_5871,N_8160);
nor U14592 (N_14592,N_9258,N_6749);
nor U14593 (N_14593,N_6811,N_6941);
nand U14594 (N_14594,N_9577,N_6194);
nand U14595 (N_14595,N_9324,N_7555);
or U14596 (N_14596,N_8199,N_6019);
nand U14597 (N_14597,N_7059,N_8473);
or U14598 (N_14598,N_6327,N_9479);
and U14599 (N_14599,N_6006,N_9482);
xor U14600 (N_14600,N_9173,N_9051);
nor U14601 (N_14601,N_5600,N_8147);
nand U14602 (N_14602,N_9084,N_5572);
or U14603 (N_14603,N_9785,N_8154);
nand U14604 (N_14604,N_5953,N_7975);
xnor U14605 (N_14605,N_9841,N_5125);
and U14606 (N_14606,N_6910,N_9330);
or U14607 (N_14607,N_9318,N_7990);
xor U14608 (N_14608,N_9831,N_6585);
nor U14609 (N_14609,N_5380,N_5137);
nor U14610 (N_14610,N_8406,N_9167);
or U14611 (N_14611,N_5801,N_8837);
or U14612 (N_14612,N_9625,N_9830);
nand U14613 (N_14613,N_9651,N_9465);
and U14614 (N_14614,N_8987,N_9392);
and U14615 (N_14615,N_6282,N_6218);
and U14616 (N_14616,N_7130,N_6707);
nand U14617 (N_14617,N_8060,N_9521);
nor U14618 (N_14618,N_9145,N_5331);
nand U14619 (N_14619,N_7707,N_9305);
xor U14620 (N_14620,N_7617,N_8209);
and U14621 (N_14621,N_7109,N_7094);
or U14622 (N_14622,N_6975,N_5073);
or U14623 (N_14623,N_8830,N_7523);
and U14624 (N_14624,N_7314,N_9852);
or U14625 (N_14625,N_5159,N_6550);
nor U14626 (N_14626,N_7868,N_8658);
nand U14627 (N_14627,N_7107,N_9188);
xnor U14628 (N_14628,N_7074,N_5865);
and U14629 (N_14629,N_5240,N_5310);
and U14630 (N_14630,N_5106,N_6818);
or U14631 (N_14631,N_9024,N_6268);
and U14632 (N_14632,N_9290,N_8661);
xnor U14633 (N_14633,N_5964,N_9359);
xnor U14634 (N_14634,N_5367,N_6555);
nor U14635 (N_14635,N_8448,N_8378);
or U14636 (N_14636,N_5181,N_9449);
and U14637 (N_14637,N_8920,N_6480);
nand U14638 (N_14638,N_8634,N_8066);
nor U14639 (N_14639,N_6434,N_5383);
or U14640 (N_14640,N_8218,N_6367);
xor U14641 (N_14641,N_5385,N_9972);
or U14642 (N_14642,N_9770,N_5792);
or U14643 (N_14643,N_9228,N_7598);
nand U14644 (N_14644,N_5405,N_8702);
nand U14645 (N_14645,N_5538,N_5746);
or U14646 (N_14646,N_6958,N_6665);
nand U14647 (N_14647,N_9647,N_7105);
nand U14648 (N_14648,N_8587,N_6339);
nor U14649 (N_14649,N_6436,N_6867);
nand U14650 (N_14650,N_7811,N_8462);
xnor U14651 (N_14651,N_8523,N_8456);
nor U14652 (N_14652,N_6372,N_6650);
and U14653 (N_14653,N_5286,N_5767);
or U14654 (N_14654,N_8511,N_9298);
and U14655 (N_14655,N_9073,N_8398);
nand U14656 (N_14656,N_8741,N_7939);
xnor U14657 (N_14657,N_8182,N_7655);
nor U14658 (N_14658,N_7144,N_9502);
or U14659 (N_14659,N_5477,N_6699);
nor U14660 (N_14660,N_6849,N_5586);
or U14661 (N_14661,N_8833,N_5894);
and U14662 (N_14662,N_8054,N_5843);
nor U14663 (N_14663,N_9200,N_9342);
nor U14664 (N_14664,N_6902,N_6930);
nor U14665 (N_14665,N_5055,N_9569);
nand U14666 (N_14666,N_6384,N_8804);
or U14667 (N_14667,N_9802,N_5275);
xnor U14668 (N_14668,N_6244,N_8572);
and U14669 (N_14669,N_9147,N_9555);
nand U14670 (N_14670,N_8137,N_8920);
and U14671 (N_14671,N_9528,N_5338);
nor U14672 (N_14672,N_7554,N_9560);
or U14673 (N_14673,N_8705,N_9588);
nand U14674 (N_14674,N_9816,N_6453);
nand U14675 (N_14675,N_7933,N_9121);
xor U14676 (N_14676,N_5099,N_7611);
or U14677 (N_14677,N_5188,N_5990);
nor U14678 (N_14678,N_5385,N_6117);
and U14679 (N_14679,N_9661,N_5827);
and U14680 (N_14680,N_9920,N_7602);
nand U14681 (N_14681,N_9105,N_8562);
or U14682 (N_14682,N_8264,N_6822);
nor U14683 (N_14683,N_7380,N_9603);
nand U14684 (N_14684,N_9696,N_9719);
or U14685 (N_14685,N_5980,N_7195);
nand U14686 (N_14686,N_8924,N_9597);
nand U14687 (N_14687,N_7606,N_7006);
and U14688 (N_14688,N_7926,N_9357);
nand U14689 (N_14689,N_9384,N_6932);
or U14690 (N_14690,N_9027,N_5057);
nand U14691 (N_14691,N_9024,N_5356);
and U14692 (N_14692,N_7451,N_9067);
and U14693 (N_14693,N_6509,N_9268);
or U14694 (N_14694,N_9326,N_8398);
nor U14695 (N_14695,N_5595,N_7912);
nor U14696 (N_14696,N_6957,N_8514);
nand U14697 (N_14697,N_6099,N_7710);
and U14698 (N_14698,N_7343,N_6973);
nand U14699 (N_14699,N_7208,N_8643);
nor U14700 (N_14700,N_7344,N_6547);
xnor U14701 (N_14701,N_6399,N_6738);
or U14702 (N_14702,N_6385,N_6422);
and U14703 (N_14703,N_8378,N_8936);
nor U14704 (N_14704,N_6695,N_9949);
or U14705 (N_14705,N_7677,N_6563);
and U14706 (N_14706,N_5357,N_9742);
or U14707 (N_14707,N_7592,N_5605);
or U14708 (N_14708,N_8664,N_9560);
xor U14709 (N_14709,N_7503,N_8835);
or U14710 (N_14710,N_7811,N_9994);
nand U14711 (N_14711,N_7741,N_9598);
nor U14712 (N_14712,N_6666,N_6004);
nor U14713 (N_14713,N_5205,N_5100);
nand U14714 (N_14714,N_7085,N_6657);
nand U14715 (N_14715,N_8645,N_7439);
nand U14716 (N_14716,N_6344,N_9307);
nor U14717 (N_14717,N_6477,N_8923);
nor U14718 (N_14718,N_7392,N_6122);
and U14719 (N_14719,N_8093,N_5123);
or U14720 (N_14720,N_8110,N_7352);
nand U14721 (N_14721,N_5530,N_8089);
or U14722 (N_14722,N_6894,N_9817);
or U14723 (N_14723,N_8259,N_6073);
nor U14724 (N_14724,N_7350,N_7908);
nand U14725 (N_14725,N_8724,N_9217);
and U14726 (N_14726,N_6683,N_5845);
or U14727 (N_14727,N_7568,N_6870);
nor U14728 (N_14728,N_7705,N_9644);
and U14729 (N_14729,N_8740,N_7325);
nor U14730 (N_14730,N_5707,N_6189);
or U14731 (N_14731,N_5111,N_9542);
or U14732 (N_14732,N_5753,N_8634);
nor U14733 (N_14733,N_8403,N_7991);
xor U14734 (N_14734,N_7396,N_9125);
or U14735 (N_14735,N_8740,N_8345);
or U14736 (N_14736,N_6601,N_8666);
or U14737 (N_14737,N_8774,N_6133);
nand U14738 (N_14738,N_5451,N_6489);
nor U14739 (N_14739,N_8249,N_6240);
nor U14740 (N_14740,N_7503,N_6380);
nand U14741 (N_14741,N_9205,N_9800);
nand U14742 (N_14742,N_8305,N_9974);
nor U14743 (N_14743,N_7124,N_7839);
and U14744 (N_14744,N_9909,N_5730);
nor U14745 (N_14745,N_8858,N_9833);
or U14746 (N_14746,N_8976,N_6818);
and U14747 (N_14747,N_5382,N_5103);
nor U14748 (N_14748,N_5752,N_6803);
nor U14749 (N_14749,N_6782,N_5758);
and U14750 (N_14750,N_6434,N_6495);
nor U14751 (N_14751,N_8875,N_5907);
nand U14752 (N_14752,N_7507,N_7245);
and U14753 (N_14753,N_8746,N_7417);
nor U14754 (N_14754,N_5247,N_8613);
or U14755 (N_14755,N_5317,N_9553);
and U14756 (N_14756,N_8649,N_5701);
nand U14757 (N_14757,N_8079,N_9689);
nand U14758 (N_14758,N_9608,N_5377);
or U14759 (N_14759,N_8859,N_5986);
nor U14760 (N_14760,N_9223,N_5456);
or U14761 (N_14761,N_5778,N_9775);
nand U14762 (N_14762,N_8483,N_5507);
and U14763 (N_14763,N_5257,N_5931);
nand U14764 (N_14764,N_8928,N_9167);
and U14765 (N_14765,N_6798,N_9106);
or U14766 (N_14766,N_5825,N_9395);
nand U14767 (N_14767,N_9990,N_6821);
or U14768 (N_14768,N_8432,N_5476);
and U14769 (N_14769,N_8699,N_8108);
or U14770 (N_14770,N_5442,N_7932);
xor U14771 (N_14771,N_8880,N_8023);
or U14772 (N_14772,N_5828,N_8788);
xor U14773 (N_14773,N_5944,N_5862);
or U14774 (N_14774,N_6427,N_9579);
and U14775 (N_14775,N_6808,N_8290);
and U14776 (N_14776,N_8398,N_5085);
xnor U14777 (N_14777,N_6479,N_5626);
nor U14778 (N_14778,N_6580,N_7126);
nor U14779 (N_14779,N_6240,N_8088);
and U14780 (N_14780,N_9567,N_6967);
and U14781 (N_14781,N_9739,N_7313);
nand U14782 (N_14782,N_5190,N_9848);
xor U14783 (N_14783,N_9462,N_7352);
nor U14784 (N_14784,N_6249,N_8319);
and U14785 (N_14785,N_8326,N_5997);
or U14786 (N_14786,N_9418,N_8659);
xor U14787 (N_14787,N_9373,N_7976);
nor U14788 (N_14788,N_7215,N_7560);
nor U14789 (N_14789,N_6892,N_6942);
xnor U14790 (N_14790,N_5742,N_9622);
and U14791 (N_14791,N_8507,N_6650);
and U14792 (N_14792,N_9164,N_6654);
nand U14793 (N_14793,N_6754,N_8377);
or U14794 (N_14794,N_8072,N_5085);
or U14795 (N_14795,N_7765,N_8955);
and U14796 (N_14796,N_9971,N_7479);
nor U14797 (N_14797,N_9638,N_5788);
or U14798 (N_14798,N_6943,N_5277);
and U14799 (N_14799,N_7726,N_8947);
xnor U14800 (N_14800,N_8721,N_5441);
nor U14801 (N_14801,N_6655,N_8439);
nand U14802 (N_14802,N_7721,N_8899);
nor U14803 (N_14803,N_8000,N_8068);
nor U14804 (N_14804,N_9197,N_7779);
and U14805 (N_14805,N_5902,N_5681);
and U14806 (N_14806,N_9249,N_9318);
nand U14807 (N_14807,N_8146,N_8834);
xor U14808 (N_14808,N_7476,N_8815);
xnor U14809 (N_14809,N_5752,N_5536);
or U14810 (N_14810,N_8609,N_9303);
or U14811 (N_14811,N_6589,N_8598);
nand U14812 (N_14812,N_7509,N_9366);
and U14813 (N_14813,N_5402,N_6706);
nor U14814 (N_14814,N_9165,N_7217);
nor U14815 (N_14815,N_9923,N_8371);
nor U14816 (N_14816,N_6769,N_5580);
and U14817 (N_14817,N_7560,N_7129);
or U14818 (N_14818,N_5769,N_9849);
nor U14819 (N_14819,N_5503,N_7652);
nor U14820 (N_14820,N_6586,N_5067);
and U14821 (N_14821,N_6321,N_7225);
or U14822 (N_14822,N_5806,N_7214);
or U14823 (N_14823,N_9778,N_7624);
nor U14824 (N_14824,N_5491,N_8671);
nor U14825 (N_14825,N_5059,N_6037);
and U14826 (N_14826,N_6223,N_7392);
and U14827 (N_14827,N_9293,N_8549);
nor U14828 (N_14828,N_5033,N_6548);
xor U14829 (N_14829,N_6780,N_7670);
nor U14830 (N_14830,N_7364,N_8925);
nand U14831 (N_14831,N_6954,N_8054);
and U14832 (N_14832,N_6063,N_7434);
or U14833 (N_14833,N_6570,N_7527);
or U14834 (N_14834,N_8406,N_8399);
or U14835 (N_14835,N_8457,N_8936);
and U14836 (N_14836,N_9992,N_6859);
and U14837 (N_14837,N_5993,N_9310);
or U14838 (N_14838,N_8240,N_9880);
and U14839 (N_14839,N_9506,N_8845);
xnor U14840 (N_14840,N_5473,N_5926);
or U14841 (N_14841,N_7897,N_7676);
nand U14842 (N_14842,N_5064,N_8717);
or U14843 (N_14843,N_7294,N_8351);
or U14844 (N_14844,N_6641,N_9476);
nor U14845 (N_14845,N_5574,N_8096);
and U14846 (N_14846,N_7165,N_7994);
xnor U14847 (N_14847,N_6680,N_5944);
xnor U14848 (N_14848,N_5154,N_7616);
xnor U14849 (N_14849,N_6917,N_8987);
and U14850 (N_14850,N_8911,N_9457);
nand U14851 (N_14851,N_8725,N_8921);
and U14852 (N_14852,N_5162,N_7645);
or U14853 (N_14853,N_5248,N_6293);
and U14854 (N_14854,N_5798,N_5272);
nand U14855 (N_14855,N_8333,N_8336);
nor U14856 (N_14856,N_5481,N_5308);
nand U14857 (N_14857,N_5414,N_5648);
nand U14858 (N_14858,N_6602,N_9389);
and U14859 (N_14859,N_6533,N_9377);
or U14860 (N_14860,N_6958,N_5559);
or U14861 (N_14861,N_8459,N_6885);
and U14862 (N_14862,N_5114,N_5609);
and U14863 (N_14863,N_6850,N_7630);
nor U14864 (N_14864,N_9542,N_9391);
nor U14865 (N_14865,N_5339,N_5401);
nor U14866 (N_14866,N_7030,N_7860);
and U14867 (N_14867,N_7300,N_8679);
nor U14868 (N_14868,N_5847,N_5624);
nand U14869 (N_14869,N_5645,N_9742);
xnor U14870 (N_14870,N_7631,N_9339);
and U14871 (N_14871,N_8522,N_5973);
and U14872 (N_14872,N_9725,N_6608);
nor U14873 (N_14873,N_7657,N_5913);
and U14874 (N_14874,N_8379,N_5698);
nand U14875 (N_14875,N_5701,N_5941);
xor U14876 (N_14876,N_6600,N_7212);
and U14877 (N_14877,N_9588,N_8775);
nor U14878 (N_14878,N_8794,N_8883);
nand U14879 (N_14879,N_5418,N_5274);
and U14880 (N_14880,N_9001,N_5610);
or U14881 (N_14881,N_9727,N_7786);
or U14882 (N_14882,N_5963,N_8577);
and U14883 (N_14883,N_5415,N_7979);
xnor U14884 (N_14884,N_8256,N_8254);
or U14885 (N_14885,N_8158,N_5342);
xor U14886 (N_14886,N_7440,N_6851);
or U14887 (N_14887,N_7738,N_9864);
and U14888 (N_14888,N_6220,N_6418);
or U14889 (N_14889,N_9812,N_8745);
or U14890 (N_14890,N_6209,N_8579);
nand U14891 (N_14891,N_5261,N_9453);
and U14892 (N_14892,N_5133,N_9500);
and U14893 (N_14893,N_7352,N_9600);
xnor U14894 (N_14894,N_6304,N_9246);
or U14895 (N_14895,N_9537,N_8326);
nand U14896 (N_14896,N_6847,N_7399);
nor U14897 (N_14897,N_8854,N_7930);
or U14898 (N_14898,N_8853,N_9725);
nand U14899 (N_14899,N_5211,N_5555);
or U14900 (N_14900,N_8548,N_5138);
nand U14901 (N_14901,N_9888,N_7578);
nand U14902 (N_14902,N_6238,N_6361);
nor U14903 (N_14903,N_7211,N_6014);
nor U14904 (N_14904,N_8170,N_6976);
nor U14905 (N_14905,N_8498,N_7238);
nand U14906 (N_14906,N_5007,N_6218);
nor U14907 (N_14907,N_8262,N_7004);
nand U14908 (N_14908,N_7296,N_9376);
nor U14909 (N_14909,N_8850,N_9046);
nand U14910 (N_14910,N_6297,N_5626);
nand U14911 (N_14911,N_7909,N_9187);
nand U14912 (N_14912,N_5553,N_6762);
nor U14913 (N_14913,N_7892,N_9323);
and U14914 (N_14914,N_5847,N_6093);
or U14915 (N_14915,N_7873,N_6424);
nor U14916 (N_14916,N_9776,N_8820);
or U14917 (N_14917,N_9470,N_8389);
nor U14918 (N_14918,N_9520,N_6524);
or U14919 (N_14919,N_6432,N_7502);
nor U14920 (N_14920,N_9376,N_7182);
or U14921 (N_14921,N_5433,N_8613);
or U14922 (N_14922,N_7677,N_7899);
or U14923 (N_14923,N_6166,N_9086);
nand U14924 (N_14924,N_7203,N_6292);
nor U14925 (N_14925,N_5189,N_6263);
or U14926 (N_14926,N_5804,N_9531);
nor U14927 (N_14927,N_9621,N_8505);
nand U14928 (N_14928,N_7901,N_7920);
nor U14929 (N_14929,N_8423,N_8530);
nor U14930 (N_14930,N_5854,N_7403);
and U14931 (N_14931,N_9568,N_6847);
or U14932 (N_14932,N_8363,N_8526);
nor U14933 (N_14933,N_9111,N_8051);
or U14934 (N_14934,N_5223,N_5411);
or U14935 (N_14935,N_9434,N_8065);
nor U14936 (N_14936,N_5876,N_7135);
nand U14937 (N_14937,N_6597,N_8903);
nand U14938 (N_14938,N_7836,N_8668);
nor U14939 (N_14939,N_8980,N_8249);
or U14940 (N_14940,N_5230,N_5885);
nor U14941 (N_14941,N_9839,N_8911);
nand U14942 (N_14942,N_5256,N_9216);
and U14943 (N_14943,N_8853,N_7474);
xor U14944 (N_14944,N_7914,N_7854);
and U14945 (N_14945,N_7151,N_9297);
nor U14946 (N_14946,N_5542,N_5535);
or U14947 (N_14947,N_5274,N_7594);
nand U14948 (N_14948,N_6626,N_6481);
xnor U14949 (N_14949,N_5227,N_6988);
nor U14950 (N_14950,N_8522,N_9547);
or U14951 (N_14951,N_6925,N_5911);
and U14952 (N_14952,N_7545,N_7963);
xnor U14953 (N_14953,N_5372,N_7582);
or U14954 (N_14954,N_8010,N_6032);
xor U14955 (N_14955,N_6753,N_7987);
or U14956 (N_14956,N_7626,N_8958);
nor U14957 (N_14957,N_8738,N_9516);
xnor U14958 (N_14958,N_8274,N_5526);
and U14959 (N_14959,N_7038,N_5246);
or U14960 (N_14960,N_7087,N_8311);
or U14961 (N_14961,N_6463,N_9872);
nand U14962 (N_14962,N_8375,N_8762);
or U14963 (N_14963,N_6585,N_8073);
or U14964 (N_14964,N_8653,N_9042);
nor U14965 (N_14965,N_6224,N_9565);
and U14966 (N_14966,N_7376,N_9099);
nor U14967 (N_14967,N_5834,N_6092);
nand U14968 (N_14968,N_5529,N_5024);
and U14969 (N_14969,N_5010,N_7207);
nor U14970 (N_14970,N_5134,N_7427);
nor U14971 (N_14971,N_6512,N_5371);
and U14972 (N_14972,N_6200,N_5702);
and U14973 (N_14973,N_6124,N_8525);
nand U14974 (N_14974,N_8915,N_8294);
or U14975 (N_14975,N_6641,N_8416);
nand U14976 (N_14976,N_8712,N_9691);
nand U14977 (N_14977,N_8169,N_8077);
and U14978 (N_14978,N_9277,N_6172);
nand U14979 (N_14979,N_9181,N_6970);
and U14980 (N_14980,N_7177,N_6655);
xor U14981 (N_14981,N_8410,N_5218);
nor U14982 (N_14982,N_9567,N_9651);
nor U14983 (N_14983,N_9928,N_7729);
and U14984 (N_14984,N_7024,N_5667);
or U14985 (N_14985,N_7763,N_5871);
and U14986 (N_14986,N_6191,N_5262);
nand U14987 (N_14987,N_7216,N_9548);
and U14988 (N_14988,N_5349,N_9073);
and U14989 (N_14989,N_5700,N_7268);
or U14990 (N_14990,N_6811,N_7956);
nand U14991 (N_14991,N_5982,N_5961);
nor U14992 (N_14992,N_5717,N_9594);
nand U14993 (N_14993,N_9854,N_7621);
nand U14994 (N_14994,N_5490,N_9343);
and U14995 (N_14995,N_6432,N_8085);
nor U14996 (N_14996,N_9464,N_7868);
nor U14997 (N_14997,N_6134,N_8578);
nor U14998 (N_14998,N_9711,N_6115);
xor U14999 (N_14999,N_6588,N_7221);
nor U15000 (N_15000,N_11184,N_12411);
or U15001 (N_15001,N_11254,N_13279);
nand U15002 (N_15002,N_14120,N_12933);
nand U15003 (N_15003,N_14263,N_12452);
nor U15004 (N_15004,N_12986,N_11050);
nand U15005 (N_15005,N_10050,N_13084);
and U15006 (N_15006,N_14232,N_12430);
or U15007 (N_15007,N_10492,N_14694);
and U15008 (N_15008,N_14016,N_11152);
xnor U15009 (N_15009,N_13792,N_13385);
nand U15010 (N_15010,N_11740,N_14824);
or U15011 (N_15011,N_10458,N_13290);
and U15012 (N_15012,N_12977,N_12290);
nand U15013 (N_15013,N_13992,N_11348);
or U15014 (N_15014,N_11373,N_13317);
nand U15015 (N_15015,N_10933,N_13821);
or U15016 (N_15016,N_13304,N_12711);
and U15017 (N_15017,N_13810,N_13728);
nor U15018 (N_15018,N_13946,N_12293);
nand U15019 (N_15019,N_14836,N_11252);
xor U15020 (N_15020,N_10829,N_13022);
nor U15021 (N_15021,N_12283,N_14779);
nand U15022 (N_15022,N_11418,N_12767);
or U15023 (N_15023,N_14280,N_14076);
and U15024 (N_15024,N_13358,N_14791);
nor U15025 (N_15025,N_12410,N_13007);
and U15026 (N_15026,N_14431,N_11166);
or U15027 (N_15027,N_10183,N_14670);
or U15028 (N_15028,N_10021,N_13028);
nor U15029 (N_15029,N_14816,N_10557);
nor U15030 (N_15030,N_11539,N_12172);
or U15031 (N_15031,N_13510,N_12110);
or U15032 (N_15032,N_13701,N_10227);
and U15033 (N_15033,N_11022,N_14702);
nand U15034 (N_15034,N_11405,N_12478);
nand U15035 (N_15035,N_11753,N_10257);
nand U15036 (N_15036,N_13360,N_11726);
or U15037 (N_15037,N_14274,N_10284);
nor U15038 (N_15038,N_14672,N_11327);
nand U15039 (N_15039,N_12790,N_13220);
and U15040 (N_15040,N_11519,N_10983);
and U15041 (N_15041,N_14339,N_10433);
nand U15042 (N_15042,N_11182,N_11498);
or U15043 (N_15043,N_14030,N_12896);
or U15044 (N_15044,N_13911,N_12702);
nor U15045 (N_15045,N_10503,N_14290);
xor U15046 (N_15046,N_11932,N_11058);
nand U15047 (N_15047,N_14380,N_14495);
nand U15048 (N_15048,N_11385,N_10594);
and U15049 (N_15049,N_12085,N_13086);
or U15050 (N_15050,N_13345,N_11195);
nor U15051 (N_15051,N_13608,N_10036);
nor U15052 (N_15052,N_13841,N_14114);
and U15053 (N_15053,N_10443,N_10088);
xor U15054 (N_15054,N_13953,N_10316);
or U15055 (N_15055,N_11198,N_14344);
or U15056 (N_15056,N_14907,N_11009);
nor U15057 (N_15057,N_12610,N_11822);
or U15058 (N_15058,N_13104,N_12414);
nand U15059 (N_15059,N_14808,N_12061);
nor U15060 (N_15060,N_14342,N_10522);
nor U15061 (N_15061,N_12940,N_12277);
nand U15062 (N_15062,N_14399,N_12054);
or U15063 (N_15063,N_12901,N_12114);
xor U15064 (N_15064,N_10152,N_11424);
or U15065 (N_15065,N_11615,N_11447);
and U15066 (N_15066,N_10395,N_10236);
and U15067 (N_15067,N_12695,N_13714);
nand U15068 (N_15068,N_14612,N_12040);
nand U15069 (N_15069,N_10744,N_12162);
nor U15070 (N_15070,N_12882,N_13124);
and U15071 (N_15071,N_10352,N_11607);
and U15072 (N_15072,N_11588,N_10411);
or U15073 (N_15073,N_10926,N_14853);
nand U15074 (N_15074,N_11998,N_14767);
nor U15075 (N_15075,N_11005,N_14490);
nor U15076 (N_15076,N_11450,N_11041);
and U15077 (N_15077,N_14002,N_11493);
nand U15078 (N_15078,N_13499,N_12450);
nand U15079 (N_15079,N_14143,N_14148);
and U15080 (N_15080,N_10338,N_14810);
xor U15081 (N_15081,N_10978,N_12663);
or U15082 (N_15082,N_13447,N_14610);
and U15083 (N_15083,N_12871,N_10981);
nand U15084 (N_15084,N_10430,N_11426);
or U15085 (N_15085,N_11849,N_10684);
nor U15086 (N_15086,N_10051,N_14959);
and U15087 (N_15087,N_14046,N_14464);
and U15088 (N_15088,N_14243,N_11256);
and U15089 (N_15089,N_11392,N_10578);
or U15090 (N_15090,N_10565,N_11960);
or U15091 (N_15091,N_10157,N_11513);
and U15092 (N_15092,N_12113,N_11391);
and U15093 (N_15093,N_12617,N_12221);
xor U15094 (N_15094,N_14341,N_11043);
or U15095 (N_15095,N_14036,N_11913);
nor U15096 (N_15096,N_14206,N_13059);
xnor U15097 (N_15097,N_14322,N_14593);
nor U15098 (N_15098,N_13865,N_13416);
and U15099 (N_15099,N_10104,N_11582);
and U15100 (N_15100,N_10181,N_13078);
nand U15101 (N_15101,N_14604,N_10239);
or U15102 (N_15102,N_13346,N_10416);
xor U15103 (N_15103,N_13657,N_13577);
and U15104 (N_15104,N_12191,N_13139);
or U15105 (N_15105,N_10339,N_10555);
and U15106 (N_15106,N_13932,N_14879);
and U15107 (N_15107,N_14241,N_11407);
nand U15108 (N_15108,N_12751,N_14703);
or U15109 (N_15109,N_12125,N_13995);
nand U15110 (N_15110,N_11338,N_10817);
nand U15111 (N_15111,N_12703,N_14644);
nand U15112 (N_15112,N_13585,N_14864);
or U15113 (N_15113,N_13005,N_12334);
and U15114 (N_15114,N_11950,N_12868);
nand U15115 (N_15115,N_12320,N_14963);
xor U15116 (N_15116,N_11812,N_12893);
nor U15117 (N_15117,N_14218,N_13636);
or U15118 (N_15118,N_13235,N_14834);
and U15119 (N_15119,N_11130,N_11957);
nor U15120 (N_15120,N_10394,N_10679);
nor U15121 (N_15121,N_14771,N_10688);
nand U15122 (N_15122,N_10043,N_14924);
nor U15123 (N_15123,N_12417,N_11427);
or U15124 (N_15124,N_14656,N_14543);
xor U15125 (N_15125,N_12676,N_12988);
xor U15126 (N_15126,N_11160,N_10622);
nand U15127 (N_15127,N_11342,N_12499);
nand U15128 (N_15128,N_13341,N_11278);
nand U15129 (N_15129,N_12570,N_12200);
and U15130 (N_15130,N_14031,N_12649);
and U15131 (N_15131,N_10702,N_13214);
nand U15132 (N_15132,N_11180,N_13493);
nor U15133 (N_15133,N_11835,N_11949);
nand U15134 (N_15134,N_10590,N_13830);
nand U15135 (N_15135,N_11821,N_12029);
and U15136 (N_15136,N_10514,N_11484);
and U15137 (N_15137,N_13320,N_12843);
nand U15138 (N_15138,N_12673,N_13379);
nand U15139 (N_15139,N_10807,N_13102);
and U15140 (N_15140,N_10837,N_12508);
and U15141 (N_15141,N_11042,N_10536);
or U15142 (N_15142,N_11111,N_12133);
xor U15143 (N_15143,N_14580,N_10432);
xor U15144 (N_15144,N_13959,N_13227);
nand U15145 (N_15145,N_14067,N_10950);
or U15146 (N_15146,N_12388,N_10165);
and U15147 (N_15147,N_12352,N_10228);
and U15148 (N_15148,N_13938,N_12745);
nor U15149 (N_15149,N_14505,N_11717);
xor U15150 (N_15150,N_12108,N_12152);
nor U15151 (N_15151,N_14253,N_13167);
nand U15152 (N_15152,N_14208,N_12303);
nand U15153 (N_15153,N_13426,N_14449);
or U15154 (N_15154,N_12174,N_11367);
or U15155 (N_15155,N_13970,N_11759);
nand U15156 (N_15156,N_14482,N_10224);
and U15157 (N_15157,N_14625,N_13108);
or U15158 (N_15158,N_11301,N_10582);
nor U15159 (N_15159,N_12075,N_11078);
or U15160 (N_15160,N_10917,N_11732);
nand U15161 (N_15161,N_13515,N_13363);
nand U15162 (N_15162,N_10469,N_14020);
and U15163 (N_15163,N_11903,N_11203);
nand U15164 (N_15164,N_13618,N_10887);
nand U15165 (N_15165,N_12366,N_14546);
nor U15166 (N_15166,N_12158,N_11750);
or U15167 (N_15167,N_11564,N_11300);
or U15168 (N_15168,N_14088,N_10718);
nor U15169 (N_15169,N_11406,N_11125);
and U15170 (N_15170,N_13025,N_13757);
or U15171 (N_15171,N_14012,N_14429);
nor U15172 (N_15172,N_12138,N_10958);
nand U15173 (N_15173,N_10075,N_14397);
xnor U15174 (N_15174,N_12444,N_12719);
or U15175 (N_15175,N_10304,N_14157);
nand U15176 (N_15176,N_12203,N_14049);
xor U15177 (N_15177,N_13812,N_14154);
or U15178 (N_15178,N_12992,N_14083);
nand U15179 (N_15179,N_11270,N_11704);
or U15180 (N_15180,N_13692,N_11323);
and U15181 (N_15181,N_10741,N_10139);
and U15182 (N_15182,N_14686,N_10288);
or U15183 (N_15183,N_14726,N_12803);
nand U15184 (N_15184,N_10653,N_10844);
nand U15185 (N_15185,N_10577,N_14675);
nor U15186 (N_15186,N_13335,N_11233);
or U15187 (N_15187,N_10520,N_13113);
nor U15188 (N_15188,N_14704,N_12607);
or U15189 (N_15189,N_12015,N_13607);
nor U15190 (N_15190,N_11369,N_10879);
xnor U15191 (N_15191,N_13635,N_14210);
or U15192 (N_15192,N_10614,N_12214);
nand U15193 (N_15193,N_13737,N_14516);
and U15194 (N_15194,N_14296,N_11433);
or U15195 (N_15195,N_10621,N_14440);
or U15196 (N_15196,N_11928,N_13831);
xnor U15197 (N_15197,N_10572,N_14299);
or U15198 (N_15198,N_10846,N_14751);
nor U15199 (N_15199,N_10544,N_12681);
nor U15200 (N_15200,N_12361,N_12183);
nor U15201 (N_15201,N_10056,N_12735);
xnor U15202 (N_15202,N_10965,N_11400);
and U15203 (N_15203,N_12348,N_13572);
xor U15204 (N_15204,N_10992,N_10194);
and U15205 (N_15205,N_10897,N_12747);
nand U15206 (N_15206,N_14536,N_13408);
nor U15207 (N_15207,N_14842,N_13594);
or U15208 (N_15208,N_13818,N_11091);
nand U15209 (N_15209,N_12777,N_13748);
nand U15210 (N_15210,N_12837,N_13816);
and U15211 (N_15211,N_10550,N_11471);
nand U15212 (N_15212,N_14970,N_10721);
xor U15213 (N_15213,N_10039,N_13492);
nand U15214 (N_15214,N_10940,N_14601);
nor U15215 (N_15215,N_13226,N_11438);
and U15216 (N_15216,N_14504,N_10334);
nor U15217 (N_15217,N_10434,N_11538);
nand U15218 (N_15218,N_10853,N_11982);
nand U15219 (N_15219,N_10603,N_10843);
nand U15220 (N_15220,N_12278,N_13339);
and U15221 (N_15221,N_14971,N_12159);
and U15222 (N_15222,N_11275,N_12879);
nand U15223 (N_15223,N_10025,N_13438);
nor U15224 (N_15224,N_13565,N_13421);
nand U15225 (N_15225,N_11721,N_14502);
xnor U15226 (N_15226,N_10629,N_11977);
and U15227 (N_15227,N_10365,N_11016);
and U15228 (N_15228,N_14064,N_10264);
and U15229 (N_15229,N_10361,N_10064);
or U15230 (N_15230,N_10249,N_14596);
nor U15231 (N_15231,N_13172,N_14700);
nand U15232 (N_15232,N_12389,N_13160);
nor U15233 (N_15233,N_13234,N_12425);
or U15234 (N_15234,N_11993,N_12525);
and U15235 (N_15235,N_13982,N_10366);
or U15236 (N_15236,N_11806,N_10930);
nand U15237 (N_15237,N_10059,N_10420);
or U15238 (N_15238,N_13344,N_14822);
or U15239 (N_15239,N_13722,N_13811);
nor U15240 (N_15240,N_13276,N_10027);
nand U15241 (N_15241,N_11241,N_13130);
and U15242 (N_15242,N_13806,N_11886);
and U15243 (N_15243,N_13547,N_11332);
or U15244 (N_15244,N_14178,N_12161);
and U15245 (N_15245,N_12081,N_10901);
nand U15246 (N_15246,N_10727,N_11144);
and U15247 (N_15247,N_13870,N_11202);
or U15248 (N_15248,N_13163,N_14781);
nand U15249 (N_15249,N_14663,N_10802);
nor U15250 (N_15250,N_12260,N_14239);
nand U15251 (N_15251,N_14607,N_11777);
nand U15252 (N_15252,N_11206,N_12382);
nand U15253 (N_15253,N_11505,N_10066);
and U15254 (N_15254,N_14371,N_12249);
xnor U15255 (N_15255,N_10403,N_10600);
or U15256 (N_15256,N_13321,N_14620);
nand U15257 (N_15257,N_11908,N_10473);
xor U15258 (N_15258,N_11659,N_12635);
or U15259 (N_15259,N_13422,N_11414);
and U15260 (N_15260,N_11923,N_11371);
and U15261 (N_15261,N_10226,N_10273);
or U15262 (N_15262,N_14891,N_14425);
nand U15263 (N_15263,N_12684,N_14956);
nor U15264 (N_15264,N_13480,N_10117);
and U15265 (N_15265,N_11996,N_11896);
xnor U15266 (N_15266,N_14676,N_13719);
nor U15267 (N_15267,N_14542,N_10595);
and U15268 (N_15268,N_13239,N_14988);
or U15269 (N_15269,N_10882,N_10609);
or U15270 (N_15270,N_13936,N_10184);
or U15271 (N_15271,N_10715,N_12069);
nor U15272 (N_15272,N_11098,N_10467);
xor U15273 (N_15273,N_14950,N_10201);
or U15274 (N_15274,N_13117,N_13655);
xor U15275 (N_15275,N_10488,N_12936);
nand U15276 (N_15276,N_13926,N_12563);
and U15277 (N_15277,N_11987,N_14874);
xnor U15278 (N_15278,N_12937,N_14926);
and U15279 (N_15279,N_11212,N_10731);
or U15280 (N_15280,N_14749,N_10602);
and U15281 (N_15281,N_14573,N_11216);
or U15282 (N_15282,N_11366,N_10814);
and U15283 (N_15283,N_11116,N_10742);
or U15284 (N_15284,N_11349,N_11415);
xnor U15285 (N_15285,N_10709,N_10344);
or U15286 (N_15286,N_11359,N_14271);
nand U15287 (N_15287,N_11641,N_14320);
or U15288 (N_15288,N_12005,N_12853);
or U15289 (N_15289,N_11133,N_14129);
and U15290 (N_15290,N_14392,N_14739);
xnor U15291 (N_15291,N_13778,N_13538);
nand U15292 (N_15292,N_14105,N_10714);
nand U15293 (N_15293,N_14600,N_12854);
nand U15294 (N_15294,N_14078,N_11047);
xnor U15295 (N_15295,N_12543,N_10337);
and U15296 (N_15296,N_14940,N_11158);
nor U15297 (N_15297,N_10764,N_12722);
and U15298 (N_15298,N_13660,N_10728);
or U15299 (N_15299,N_14171,N_12641);
and U15300 (N_15300,N_11893,N_14494);
and U15301 (N_15301,N_14854,N_10658);
nor U15302 (N_15302,N_10539,N_12875);
nand U15303 (N_15303,N_11561,N_10235);
or U15304 (N_15304,N_10074,N_13285);
and U15305 (N_15305,N_11827,N_14861);
xnor U15306 (N_15306,N_13079,N_14230);
and U15307 (N_15307,N_10654,N_10285);
and U15308 (N_15308,N_14878,N_14977);
nor U15309 (N_15309,N_13218,N_14015);
and U15310 (N_15310,N_12304,N_12862);
nand U15311 (N_15311,N_14086,N_10055);
nand U15312 (N_15312,N_13735,N_11872);
or U15313 (N_15313,N_12620,N_14732);
nand U15314 (N_15314,N_12529,N_10706);
nand U15315 (N_15315,N_14382,N_14708);
and U15316 (N_15316,N_11985,N_11293);
nand U15317 (N_15317,N_14617,N_10296);
nand U15318 (N_15318,N_14586,N_13207);
or U15319 (N_15319,N_11796,N_13734);
nand U15320 (N_15320,N_13186,N_10008);
xnor U15321 (N_15321,N_14453,N_10724);
nor U15322 (N_15322,N_12236,N_12899);
and U15323 (N_15323,N_14205,N_11947);
nor U15324 (N_15324,N_11266,N_10608);
or U15325 (N_15325,N_11757,N_13798);
and U15326 (N_15326,N_12954,N_14817);
or U15327 (N_15327,N_10450,N_11689);
or U15328 (N_15328,N_10923,N_11313);
xnor U15329 (N_15329,N_12384,N_12874);
nand U15330 (N_15330,N_10125,N_10824);
nor U15331 (N_15331,N_13009,N_14850);
or U15332 (N_15332,N_13103,N_12393);
nor U15333 (N_15333,N_10905,N_14717);
nand U15334 (N_15334,N_12416,N_14754);
or U15335 (N_15335,N_10569,N_11019);
or U15336 (N_15336,N_11416,N_13015);
nor U15337 (N_15337,N_13824,N_12036);
and U15338 (N_15338,N_12042,N_11147);
nand U15339 (N_15339,N_14736,N_13498);
nor U15340 (N_15340,N_13138,N_11535);
or U15341 (N_15341,N_10092,N_12014);
nor U15342 (N_15342,N_12422,N_13500);
or U15343 (N_15343,N_14646,N_14925);
and U15344 (N_15344,N_13779,N_10561);
and U15345 (N_15345,N_11110,N_12698);
nand U15346 (N_15346,N_13347,N_13817);
xnor U15347 (N_15347,N_13296,N_13567);
nor U15348 (N_15348,N_10110,N_10348);
or U15349 (N_15349,N_13298,N_11673);
nand U15350 (N_15350,N_14485,N_11818);
nor U15351 (N_15351,N_11051,N_12934);
and U15352 (N_15352,N_13229,N_12506);
xnor U15353 (N_15353,N_11475,N_10279);
nor U15354 (N_15354,N_12800,N_10091);
or U15355 (N_15355,N_11077,N_11245);
xnor U15356 (N_15356,N_14975,N_14457);
nand U15357 (N_15357,N_14109,N_10346);
nand U15358 (N_15358,N_14848,N_14233);
or U15359 (N_15359,N_11653,N_12582);
nor U15360 (N_15360,N_10392,N_14969);
or U15361 (N_15361,N_10665,N_10875);
and U15362 (N_15362,N_12820,N_12622);
or U15363 (N_15363,N_10632,N_14099);
and U15364 (N_15364,N_12510,N_11397);
and U15365 (N_15365,N_11646,N_12978);
nand U15366 (N_15366,N_12064,N_12816);
or U15367 (N_15367,N_10476,N_12920);
or U15368 (N_15368,N_13908,N_14869);
xnor U15369 (N_15369,N_11946,N_12644);
or U15370 (N_15370,N_12754,N_10297);
nor U15371 (N_15371,N_12006,N_14643);
or U15372 (N_15372,N_14489,N_11999);
xnor U15373 (N_15373,N_12243,N_12420);
nor U15374 (N_15374,N_13013,N_11226);
and U15375 (N_15375,N_12058,N_10996);
and U15376 (N_15376,N_11488,N_14651);
and U15377 (N_15377,N_12718,N_11532);
nor U15378 (N_15378,N_14436,N_14730);
and U15379 (N_15379,N_10779,N_12048);
and U15380 (N_15380,N_10190,N_11457);
nand U15381 (N_15381,N_12938,N_13813);
or U15382 (N_15382,N_13836,N_13713);
and U15383 (N_15383,N_14500,N_10592);
and U15384 (N_15384,N_12629,N_12507);
nand U15385 (N_15385,N_10451,N_11106);
nor U15386 (N_15386,N_14943,N_10024);
and U15387 (N_15387,N_10705,N_12687);
nor U15388 (N_15388,N_12844,N_10694);
and U15389 (N_15389,N_13255,N_11071);
nand U15390 (N_15390,N_14325,N_14035);
nand U15391 (N_15391,N_14662,N_11594);
nand U15392 (N_15392,N_10740,N_14585);
nand U15393 (N_15393,N_11634,N_10359);
nor U15394 (N_15394,N_13943,N_12606);
and U15395 (N_15395,N_11527,N_14430);
nor U15396 (N_15396,N_10885,N_12415);
nand U15397 (N_15397,N_10294,N_12878);
xor U15398 (N_15398,N_11602,N_10221);
nand U15399 (N_15399,N_11725,N_14862);
nor U15400 (N_15400,N_13787,N_13769);
or U15401 (N_15401,N_11428,N_12924);
or U15402 (N_15402,N_10154,N_11976);
nand U15403 (N_15403,N_12599,N_10186);
or U15404 (N_15404,N_14551,N_10510);
and U15405 (N_15405,N_13266,N_14785);
xor U15406 (N_15406,N_11423,N_14289);
nor U15407 (N_15407,N_13136,N_10680);
nand U15408 (N_15408,N_11755,N_12608);
or U15409 (N_15409,N_10326,N_11517);
or U15410 (N_15410,N_11191,N_11250);
and U15411 (N_15411,N_13435,N_13294);
or U15412 (N_15412,N_14932,N_12489);
or U15413 (N_15413,N_10435,N_14760);
nand U15414 (N_15414,N_11183,N_10357);
nand U15415 (N_15415,N_13378,N_11108);
nand U15416 (N_15416,N_12400,N_10868);
nor U15417 (N_15417,N_12202,N_13740);
and U15418 (N_15418,N_11643,N_11134);
or U15419 (N_15419,N_10966,N_11525);
and U15420 (N_15420,N_14427,N_12928);
nor U15421 (N_15421,N_14252,N_12791);
nand U15422 (N_15422,N_10571,N_13731);
or U15423 (N_15423,N_12550,N_14630);
nor U15424 (N_15424,N_13308,N_12432);
nand U15425 (N_15425,N_11097,N_14138);
nand U15426 (N_15426,N_13661,N_14533);
nor U15427 (N_15427,N_12013,N_13945);
or U15428 (N_15428,N_11062,N_10149);
nand U15429 (N_15429,N_14367,N_14527);
nand U15430 (N_15430,N_13236,N_14042);
nor U15431 (N_15431,N_12030,N_13825);
or U15432 (N_15432,N_11853,N_13886);
and U15433 (N_15433,N_13502,N_11742);
and U15434 (N_15434,N_13128,N_13762);
and U15435 (N_15435,N_10260,N_10501);
and U15436 (N_15436,N_13931,N_12554);
or U15437 (N_15437,N_13061,N_12813);
or U15438 (N_15438,N_13224,N_14990);
and U15439 (N_15439,N_11870,N_11364);
nor U15440 (N_15440,N_13947,N_12638);
nor U15441 (N_15441,N_12194,N_12519);
nand U15442 (N_15442,N_12119,N_11638);
and U15443 (N_15443,N_12639,N_13329);
and U15444 (N_15444,N_12808,N_11865);
xor U15445 (N_15445,N_14889,N_10823);
nor U15446 (N_15446,N_10943,N_10922);
nand U15447 (N_15447,N_14329,N_14835);
and U15448 (N_15448,N_11374,N_13682);
and U15449 (N_15449,N_12276,N_13193);
nor U15450 (N_15450,N_10813,N_13131);
or U15451 (N_15451,N_14055,N_11489);
nand U15452 (N_15452,N_11687,N_14886);
or U15453 (N_15453,N_10095,N_11176);
and U15454 (N_15454,N_13794,N_10808);
or U15455 (N_15455,N_10170,N_14841);
nand U15456 (N_15456,N_13702,N_10401);
nor U15457 (N_15457,N_13809,N_14634);
and U15458 (N_15458,N_12011,N_10038);
nand U15459 (N_15459,N_11131,N_11410);
nor U15460 (N_15460,N_13887,N_14649);
nor U15461 (N_15461,N_13462,N_10325);
and U15462 (N_15462,N_12520,N_13683);
nor U15463 (N_15463,N_12238,N_10355);
and U15464 (N_15464,N_11377,N_14865);
and U15465 (N_15465,N_12877,N_12070);
or U15466 (N_15466,N_10144,N_13981);
or U15467 (N_15467,N_10234,N_13307);
and U15468 (N_15468,N_13249,N_12761);
nand U15469 (N_15469,N_13645,N_12780);
xnor U15470 (N_15470,N_11432,N_12841);
nor U15471 (N_15471,N_13230,N_12852);
nor U15472 (N_15472,N_14727,N_10131);
nor U15473 (N_15473,N_13373,N_13393);
or U15474 (N_15474,N_11070,N_12835);
and U15475 (N_15475,N_12109,N_13629);
xnor U15476 (N_15476,N_14819,N_12679);
and U15477 (N_15477,N_11117,N_10858);
nor U15478 (N_15478,N_14776,N_14085);
xnor U15479 (N_15479,N_12713,N_12332);
nand U15480 (N_15480,N_11580,N_14687);
and U15481 (N_15481,N_11151,N_11684);
nor U15482 (N_15482,N_14098,N_11860);
nand U15483 (N_15483,N_14911,N_11626);
and U15484 (N_15484,N_10013,N_14000);
nor U15485 (N_15485,N_12322,N_13840);
nand U15486 (N_15486,N_12471,N_14522);
or U15487 (N_15487,N_10692,N_13600);
nand U15488 (N_15488,N_14893,N_14103);
nor U15489 (N_15489,N_12760,N_13553);
nand U15490 (N_15490,N_13788,N_14372);
and U15491 (N_15491,N_12749,N_14731);
and U15492 (N_15492,N_10368,N_11807);
xnor U15493 (N_15493,N_13286,N_14111);
xnor U15494 (N_15494,N_10552,N_10069);
nor U15495 (N_15495,N_10205,N_12618);
and U15496 (N_15496,N_10369,N_13647);
nor U15497 (N_15497,N_13240,N_13529);
nand U15498 (N_15498,N_14664,N_11897);
nand U15499 (N_15499,N_13900,N_12763);
xor U15500 (N_15500,N_14053,N_12714);
and U15501 (N_15501,N_13114,N_11696);
or U15502 (N_15502,N_14052,N_10697);
nor U15503 (N_15503,N_12337,N_12118);
and U15504 (N_15504,N_12908,N_12910);
xor U15505 (N_15505,N_13472,N_12675);
nor U15506 (N_15506,N_11174,N_10271);
and U15507 (N_15507,N_13057,N_12463);
and U15508 (N_15508,N_12205,N_13796);
nor U15509 (N_15509,N_13175,N_12245);
and U15510 (N_15510,N_14317,N_10020);
nand U15511 (N_15511,N_11675,N_10143);
and U15512 (N_15512,N_14096,N_13711);
or U15513 (N_15513,N_10016,N_14706);
nand U15514 (N_15514,N_13076,N_12019);
or U15515 (N_15515,N_10011,N_10438);
and U15516 (N_15516,N_12930,N_13602);
and U15517 (N_15517,N_14570,N_14302);
or U15518 (N_15518,N_11002,N_11558);
xor U15519 (N_15519,N_14837,N_13099);
nand U15520 (N_15520,N_14336,N_13143);
nor U15521 (N_15521,N_14383,N_11697);
nand U15522 (N_15522,N_13881,N_10517);
xor U15523 (N_15523,N_11255,N_10804);
nor U15524 (N_15524,N_10547,N_10895);
or U15525 (N_15525,N_12107,N_11497);
or U15526 (N_15526,N_13725,N_14282);
or U15527 (N_15527,N_13054,N_14711);
nor U15528 (N_15528,N_10525,N_14518);
or U15529 (N_15529,N_13374,N_13141);
or U15530 (N_15530,N_12996,N_13039);
or U15531 (N_15531,N_14199,N_13974);
nor U15532 (N_15532,N_13659,N_10738);
nand U15533 (N_15533,N_10907,N_11591);
or U15534 (N_15534,N_12010,N_12092);
nand U15535 (N_15535,N_10388,N_12516);
xnor U15536 (N_15536,N_11633,N_12786);
xnor U15537 (N_15537,N_13384,N_13859);
or U15538 (N_15538,N_13723,N_13431);
nand U15539 (N_15539,N_11503,N_13715);
xnor U15540 (N_15540,N_13720,N_13309);
or U15541 (N_15541,N_10002,N_12812);
xor U15542 (N_15542,N_13450,N_10980);
and U15543 (N_15543,N_14650,N_13724);
nor U15544 (N_15544,N_13544,N_12209);
and U15545 (N_15545,N_11231,N_14618);
nand U15546 (N_15546,N_10437,N_11540);
nand U15547 (N_15547,N_14821,N_11705);
nand U15548 (N_15548,N_12783,N_10431);
or U15549 (N_15549,N_10830,N_10040);
or U15550 (N_15550,N_11587,N_12350);
or U15551 (N_15551,N_10867,N_13717);
xor U15552 (N_15552,N_10398,N_11983);
and U15553 (N_15553,N_11666,N_14270);
nor U15554 (N_15554,N_11844,N_14194);
and U15555 (N_15555,N_10619,N_10891);
or U15556 (N_15556,N_10763,N_11730);
or U15557 (N_15557,N_12459,N_11798);
nand U15558 (N_15558,N_13222,N_10105);
nand U15559 (N_15559,N_13634,N_11287);
or U15560 (N_15560,N_12482,N_13872);
and U15561 (N_15561,N_12915,N_14398);
and U15562 (N_15562,N_10613,N_11001);
nand U15563 (N_15563,N_12424,N_13561);
nor U15564 (N_15564,N_12285,N_14520);
nand U15565 (N_15565,N_12625,N_14758);
or U15566 (N_15566,N_12307,N_13611);
nand U15567 (N_15567,N_10321,N_11399);
xnor U15568 (N_15568,N_14778,N_11441);
and U15569 (N_15569,N_12686,N_13156);
or U15570 (N_15570,N_12299,N_12511);
or U15571 (N_15571,N_14584,N_10022);
or U15572 (N_15572,N_10031,N_13972);
nand U15573 (N_15573,N_10761,N_14247);
or U15574 (N_15574,N_12849,N_12251);
nand U15575 (N_15575,N_13852,N_13834);
nand U15576 (N_15576,N_11335,N_11140);
nor U15577 (N_15577,N_14168,N_10307);
nor U15578 (N_15578,N_14404,N_10159);
and U15579 (N_15579,N_14059,N_13261);
and U15580 (N_15580,N_14236,N_14069);
and U15581 (N_15581,N_14187,N_10806);
nand U15582 (N_15582,N_10893,N_10311);
nor U15583 (N_15583,N_10350,N_14359);
and U15584 (N_15584,N_14742,N_11531);
nor U15585 (N_15585,N_13210,N_13353);
nor U15586 (N_15586,N_13165,N_11227);
and U15587 (N_15587,N_12441,N_14568);
or U15588 (N_15588,N_14623,N_10356);
nand U15589 (N_15589,N_10623,N_12768);
and U15590 (N_15590,N_11453,N_11326);
nor U15591 (N_15591,N_12890,N_10380);
and U15592 (N_15592,N_13473,N_12811);
nand U15593 (N_15593,N_13018,N_12568);
or U15594 (N_15594,N_13756,N_12726);
or U15595 (N_15595,N_14305,N_11900);
xor U15596 (N_15596,N_14659,N_12733);
nand U15597 (N_15597,N_10545,N_13771);
nand U15598 (N_15598,N_14021,N_14897);
and U15599 (N_15599,N_10751,N_13080);
and U15600 (N_15600,N_14539,N_13050);
and U15601 (N_15601,N_11839,N_14598);
nand U15602 (N_15602,N_11273,N_12975);
and U15603 (N_15603,N_13270,N_12440);
and U15604 (N_15604,N_11627,N_10734);
and U15605 (N_15605,N_11123,N_12032);
or U15606 (N_15606,N_10861,N_11351);
xor U15607 (N_15607,N_13376,N_14567);
nand U15608 (N_15608,N_12445,N_11846);
or U15609 (N_15609,N_12403,N_11018);
nor U15610 (N_15610,N_11063,N_10507);
or U15611 (N_15611,N_10601,N_10852);
nor U15612 (N_15612,N_13892,N_13404);
or U15613 (N_15613,N_14162,N_10865);
nor U15614 (N_15614,N_13698,N_14572);
or U15615 (N_15615,N_11857,N_14633);
and U15616 (N_15616,N_14803,N_12116);
nand U15617 (N_15617,N_10314,N_12434);
nor U15618 (N_15618,N_14638,N_10335);
and U15619 (N_15619,N_13732,N_11829);
nor U15620 (N_15620,N_14345,N_14066);
and U15621 (N_15621,N_13781,N_10128);
nor U15622 (N_15622,N_10642,N_11027);
nor U15623 (N_15623,N_12822,N_12208);
nand U15624 (N_15624,N_14616,N_14235);
or U15625 (N_15625,N_13467,N_14478);
and U15626 (N_15626,N_11989,N_10585);
xnor U15627 (N_15627,N_11772,N_14082);
or U15628 (N_15628,N_12990,N_10477);
nor U15629 (N_15629,N_14309,N_14514);
or U15630 (N_15630,N_14904,N_12926);
nand U15631 (N_15631,N_14992,N_11378);
nand U15632 (N_15632,N_13666,N_10902);
nand U15633 (N_15633,N_14418,N_11127);
nand U15634 (N_15634,N_14037,N_10323);
xnor U15635 (N_15635,N_14407,N_12836);
xor U15636 (N_15636,N_14639,N_13451);
and U15637 (N_15637,N_14097,N_10872);
and U15638 (N_15638,N_12916,N_12549);
nor U15639 (N_15639,N_14456,N_10795);
nand U15640 (N_15640,N_11775,N_10854);
nor U15641 (N_15641,N_14818,N_11925);
xnor U15642 (N_15642,N_10072,N_10597);
xnor U15643 (N_15643,N_13518,N_14335);
or U15644 (N_15644,N_12518,N_13070);
and U15645 (N_15645,N_11248,N_14581);
and U15646 (N_15646,N_10256,N_12451);
nand U15647 (N_15647,N_12677,N_14370);
or U15648 (N_15648,N_13632,N_11592);
or U15649 (N_15649,N_12475,N_10928);
xnor U15650 (N_15650,N_10672,N_10485);
xnor U15651 (N_15651,N_13775,N_14314);
or U15652 (N_15652,N_11389,N_14851);
or U15653 (N_15653,N_12333,N_14029);
nand U15654 (N_15654,N_10424,N_14652);
and U15655 (N_15655,N_13687,N_10809);
xnor U15656 (N_15656,N_10230,N_11863);
nand U15657 (N_15657,N_13545,N_13284);
xor U15658 (N_15658,N_13004,N_13033);
or U15659 (N_15659,N_12188,N_14843);
xnor U15660 (N_15660,N_11345,N_10566);
nor U15661 (N_15661,N_13688,N_10635);
nor U15662 (N_15662,N_13760,N_12356);
xor U15663 (N_15663,N_12865,N_13513);
or U15664 (N_15664,N_10029,N_11482);
nand U15665 (N_15665,N_10405,N_13343);
xor U15666 (N_15666,N_14019,N_12317);
nand U15667 (N_15667,N_14094,N_11911);
nor U15668 (N_15668,N_10674,N_14039);
and U15669 (N_15669,N_12242,N_14081);
nand U15670 (N_15670,N_11355,N_14166);
nand U15671 (N_15671,N_10341,N_14292);
and U15672 (N_15672,N_11825,N_13073);
xor U15673 (N_15673,N_10755,N_10417);
nor U15674 (N_15674,N_13153,N_13331);
nor U15675 (N_15675,N_11205,N_13988);
nor U15676 (N_15676,N_10426,N_11636);
and U15677 (N_15677,N_12613,N_14722);
or U15678 (N_15678,N_14006,N_14051);
nor U15679 (N_15679,N_10987,N_13223);
or U15680 (N_15680,N_14691,N_12740);
nor U15681 (N_15681,N_11711,N_13199);
nor U15682 (N_15682,N_13790,N_11648);
and U15683 (N_15683,N_12364,N_12645);
nor U15684 (N_15684,N_13237,N_13400);
nand U15685 (N_15685,N_10776,N_13232);
nor U15686 (N_15686,N_13453,N_12115);
nor U15687 (N_15687,N_11836,N_12222);
nor U15688 (N_15688,N_12594,N_14259);
nor U15689 (N_15689,N_10204,N_11404);
nor U15690 (N_15690,N_11253,N_11990);
or U15691 (N_15691,N_12087,N_12009);
xor U15692 (N_15692,N_14466,N_11746);
xor U15693 (N_15693,N_10233,N_11429);
nor U15694 (N_15694,N_11708,N_11126);
xnor U15695 (N_15695,N_10797,N_13644);
or U15696 (N_15696,N_13318,N_12166);
and U15697 (N_15697,N_10440,N_12694);
or U15698 (N_15698,N_14566,N_14434);
nand U15699 (N_15699,N_10938,N_10062);
xnor U15700 (N_15700,N_14743,N_11437);
and U15701 (N_15701,N_14802,N_13192);
or U15702 (N_15702,N_10548,N_11902);
nand U15703 (N_15703,N_14279,N_13989);
or U15704 (N_15704,N_10287,N_13263);
nor U15705 (N_15705,N_10777,N_10449);
or U15706 (N_15706,N_13332,N_11560);
xor U15707 (N_15707,N_13568,N_10496);
xnor U15708 (N_15708,N_14564,N_13396);
nor U15709 (N_15709,N_11884,N_14857);
or U15710 (N_15710,N_12288,N_11008);
nor U15711 (N_15711,N_12171,N_11670);
xnor U15712 (N_15712,N_14858,N_12891);
and U15713 (N_15713,N_11628,N_14991);
xnor U15714 (N_15714,N_12369,N_13388);
xor U15715 (N_15715,N_10457,N_11820);
nand U15716 (N_15716,N_11213,N_14144);
nor U15717 (N_15717,N_10362,N_10012);
or U15718 (N_15718,N_11652,N_14882);
nor U15719 (N_15719,N_10726,N_13804);
and U15720 (N_15720,N_13587,N_10540);
nor U15721 (N_15721,N_12330,N_10899);
nor U15722 (N_15722,N_12439,N_13764);
nor U15723 (N_15723,N_13036,N_12785);
nand U15724 (N_15724,N_13686,N_14010);
and U15725 (N_15725,N_12286,N_10372);
nor U15726 (N_15726,N_11676,N_11828);
and U15727 (N_15727,N_10267,N_13802);
and U15728 (N_15728,N_10818,N_12026);
nand U15729 (N_15729,N_11284,N_12746);
nor U15730 (N_15730,N_11290,N_10533);
nor U15731 (N_15731,N_10820,N_14193);
xor U15732 (N_15732,N_10275,N_12797);
nand U15733 (N_15733,N_10584,N_10598);
and U15734 (N_15734,N_11204,N_14683);
or U15735 (N_15735,N_11760,N_10720);
xor U15736 (N_15736,N_12246,N_13528);
and U15737 (N_15737,N_14531,N_11703);
or U15738 (N_15738,N_12267,N_12932);
nand U15739 (N_15739,N_13487,N_10769);
or U15740 (N_15740,N_12313,N_14435);
nand U15741 (N_15741,N_13503,N_11907);
and U15742 (N_15742,N_10666,N_10390);
or U15743 (N_15743,N_11966,N_14377);
and U15744 (N_15744,N_13217,N_12965);
nand U15745 (N_15745,N_13326,N_13843);
nor U15746 (N_15746,N_12576,N_11094);
nand U15747 (N_15747,N_12121,N_12633);
nand U15748 (N_15748,N_12864,N_13580);
nor U15749 (N_15749,N_13407,N_14357);
and U15750 (N_15750,N_13228,N_10789);
xor U15751 (N_15751,N_11099,N_13559);
nand U15752 (N_15752,N_10651,N_10689);
nor U15753 (N_15753,N_13672,N_11880);
or U15754 (N_15754,N_14931,N_10291);
nor U15755 (N_15755,N_14461,N_10864);
nor U15756 (N_15756,N_13405,N_14674);
xor U15757 (N_15757,N_13055,N_11197);
nor U15758 (N_15758,N_14738,N_13807);
and U15759 (N_15759,N_11232,N_11477);
or U15760 (N_15760,N_11137,N_11096);
nand U15761 (N_15761,N_13693,N_12235);
or U15762 (N_15762,N_10081,N_14679);
or U15763 (N_15763,N_14993,N_11655);
and U15764 (N_15764,N_12717,N_10161);
or U15765 (N_15765,N_11472,N_12468);
nor U15766 (N_15766,N_14805,N_13173);
nand U15767 (N_15767,N_14153,N_14792);
nor U15768 (N_15768,N_10174,N_13606);
nand U15769 (N_15769,N_13709,N_14590);
and U15770 (N_15770,N_10863,N_12589);
and U15771 (N_15771,N_10167,N_14146);
and U15772 (N_15772,N_11347,N_12187);
nand U15773 (N_15773,N_11593,N_10849);
and U15774 (N_15774,N_11115,N_12918);
nor U15775 (N_15775,N_13201,N_13615);
nand U15776 (N_15776,N_10148,N_10290);
or U15777 (N_15777,N_12074,N_10093);
nand U15778 (N_15778,N_12281,N_12524);
nand U15779 (N_15779,N_13853,N_12473);
nand U15780 (N_15780,N_13803,N_13386);
nor U15781 (N_15781,N_11714,N_12976);
xor U15782 (N_15782,N_14388,N_13844);
nor U15783 (N_15783,N_10508,N_11199);
or U15784 (N_15784,N_10707,N_13017);
or U15785 (N_15785,N_14734,N_14393);
and U15786 (N_15786,N_14748,N_14951);
nand U15787 (N_15787,N_12234,N_11021);
and U15788 (N_15788,N_11052,N_10107);
nor U15789 (N_15789,N_12741,N_10445);
or U15790 (N_15790,N_12083,N_12637);
xnor U15791 (N_15791,N_11782,N_12145);
nor U15792 (N_15792,N_10649,N_14790);
nor U15793 (N_15793,N_14277,N_11056);
nor U15794 (N_15794,N_14909,N_10172);
nand U15795 (N_15795,N_10003,N_13777);
nor U15796 (N_15796,N_11305,N_14460);
nand U15797 (N_15797,N_12998,N_13468);
or U15798 (N_15798,N_10904,N_12049);
or U15799 (N_15799,N_11065,N_11167);
and U15800 (N_15800,N_14765,N_10472);
nor U15801 (N_15801,N_13670,N_13375);
and U15802 (N_15802,N_10399,N_12900);
nor U15803 (N_15803,N_13680,N_14626);
xnor U15804 (N_15804,N_14063,N_13913);
nand U15805 (N_15805,N_12156,N_10900);
nand U15806 (N_15806,N_10209,N_12082);
nand U15807 (N_15807,N_11909,N_11238);
xor U15808 (N_15808,N_10444,N_13758);
nor U15809 (N_15809,N_11919,N_14333);
and U15810 (N_15810,N_13440,N_13442);
nor U15811 (N_15811,N_13785,N_12247);
or U15812 (N_15812,N_11080,N_11067);
nand U15813 (N_15813,N_10716,N_12970);
or U15814 (N_15814,N_14890,N_12354);
xnor U15815 (N_15815,N_11735,N_12257);
and U15816 (N_15816,N_10644,N_14198);
nand U15817 (N_15817,N_14395,N_14151);
or U15818 (N_15818,N_13948,N_14327);
or U15819 (N_15819,N_13008,N_12056);
or U15820 (N_15820,N_12093,N_11328);
or U15821 (N_15821,N_10617,N_13191);
nor U15822 (N_15822,N_13389,N_14040);
nand U15823 (N_15823,N_12265,N_14696);
nor U15824 (N_15824,N_10018,N_10766);
or U15825 (N_15825,N_13525,N_10301);
and U15826 (N_15826,N_11937,N_14641);
nor U15827 (N_15827,N_13597,N_12948);
or U15828 (N_15828,N_10466,N_13805);
and U15829 (N_15829,N_13557,N_10164);
or U15830 (N_15830,N_10760,N_13361);
and U15831 (N_15831,N_12540,N_11930);
or U15832 (N_15832,N_14467,N_14443);
nor U15833 (N_15833,N_13797,N_11644);
and U15834 (N_15834,N_13311,N_12496);
and U15835 (N_15835,N_13414,N_14025);
nand U15836 (N_15836,N_13282,N_14477);
xor U15837 (N_15837,N_11635,N_14286);
or U15838 (N_15838,N_14352,N_11445);
and U15839 (N_15839,N_12963,N_14881);
nand U15840 (N_15840,N_11921,N_10252);
or U15841 (N_15841,N_11964,N_10960);
and U15842 (N_15842,N_12493,N_14655);
and U15843 (N_15843,N_10101,N_11136);
nand U15844 (N_15844,N_13292,N_13850);
and U15845 (N_15845,N_13786,N_11639);
nand U15846 (N_15846,N_14047,N_12614);
and U15847 (N_15847,N_13906,N_10415);
nor U15848 (N_15848,N_11320,N_10176);
nand U15849 (N_15849,N_11915,N_11630);
nand U15850 (N_15850,N_12071,N_12521);
and U15851 (N_15851,N_10178,N_10237);
or U15852 (N_15852,N_10903,N_11286);
or U15853 (N_15853,N_13044,N_13949);
nor U15854 (N_15854,N_13514,N_13252);
and U15855 (N_15855,N_14454,N_12945);
and U15856 (N_15856,N_11953,N_12817);
and U15857 (N_15857,N_12057,N_13355);
nor U15858 (N_15858,N_11295,N_14387);
and U15859 (N_15859,N_12488,N_10752);
nor U15860 (N_15860,N_14310,N_12262);
and U15861 (N_15861,N_14125,N_11751);
nor U15862 (N_15862,N_13766,N_11442);
nand U15863 (N_15863,N_11795,N_13264);
nand U15864 (N_15864,N_12178,N_14276);
nand U15865 (N_15865,N_13774,N_10639);
nand U15866 (N_15866,N_14228,N_14552);
xnor U15867 (N_15867,N_11688,N_14953);
and U15868 (N_15868,N_13512,N_11752);
nand U15869 (N_15869,N_13507,N_10511);
nand U15870 (N_15870,N_10479,N_12419);
and U15871 (N_15871,N_13536,N_14648);
and U15872 (N_15872,N_13656,N_11575);
nand U15873 (N_15873,N_10210,N_13162);
nor U15874 (N_15874,N_11745,N_14422);
nor U15875 (N_15875,N_10199,N_12149);
nand U15876 (N_15876,N_14677,N_14588);
and U15877 (N_15877,N_14303,N_14017);
and U15878 (N_15878,N_12241,N_11451);
or U15879 (N_15879,N_11733,N_12887);
nand U15880 (N_15880,N_11912,N_12651);
or U15881 (N_15881,N_10634,N_11261);
nand U15882 (N_15882,N_12395,N_10876);
or U15883 (N_15883,N_11657,N_11105);
nand U15884 (N_15884,N_11211,N_10032);
nor U15885 (N_15885,N_10109,N_13526);
nand U15886 (N_15886,N_11340,N_12066);
nand U15887 (N_15887,N_14997,N_13876);
and U15888 (N_15888,N_12421,N_13914);
and U15889 (N_15889,N_12602,N_10646);
or U15890 (N_15890,N_11691,N_13000);
nand U15891 (N_15891,N_12532,N_11970);
and U15892 (N_15892,N_11769,N_11955);
xnor U15893 (N_15893,N_11368,N_13369);
nor U15894 (N_15894,N_12968,N_14343);
nor U15895 (N_15895,N_10324,N_11218);
and U15896 (N_15896,N_12699,N_10197);
or U15897 (N_15897,N_11573,N_11783);
nand U15898 (N_15898,N_12662,N_11514);
nor U15899 (N_15899,N_11201,N_12409);
or U15900 (N_15900,N_12548,N_11502);
and U15901 (N_15901,N_13768,N_11901);
nand U15902 (N_15902,N_11786,N_14603);
and U15903 (N_15903,N_10217,N_13863);
nand U15904 (N_15904,N_13340,N_12601);
and U15905 (N_15905,N_13157,N_13364);
and U15906 (N_15906,N_12593,N_14784);
nand U15907 (N_15907,N_13736,N_12690);
or U15908 (N_15908,N_12856,N_11663);
nor U15909 (N_15909,N_12557,N_11698);
or U15910 (N_15910,N_12362,N_12765);
nand U15911 (N_15911,N_10103,N_11390);
nand U15912 (N_15912,N_12960,N_12512);
nor U15913 (N_15913,N_13755,N_13694);
nor U15914 (N_15914,N_11858,N_12117);
nand U15915 (N_15915,N_10890,N_10839);
or U15916 (N_15916,N_13928,N_13047);
nor U15917 (N_15917,N_13368,N_11148);
nand U15918 (N_15918,N_10448,N_14428);
xnor U15919 (N_15919,N_12997,N_14538);
or U15920 (N_15920,N_13110,N_14949);
and U15921 (N_15921,N_13610,N_10811);
and U15922 (N_15922,N_12423,N_14245);
xor U15923 (N_15923,N_13069,N_10397);
nand U15924 (N_15924,N_10353,N_11794);
or U15925 (N_15925,N_12653,N_11465);
nor U15926 (N_15926,N_13744,N_12873);
or U15927 (N_15927,N_12600,N_11868);
nor U15928 (N_15928,N_14952,N_12476);
nor U15929 (N_15929,N_10054,N_11692);
xor U15930 (N_15930,N_11220,N_13704);
nand U15931 (N_15931,N_13791,N_14657);
nand U15932 (N_15932,N_14709,N_11685);
and U15933 (N_15933,N_11102,N_11931);
nor U15934 (N_15934,N_11504,N_10327);
and U15935 (N_15935,N_11879,N_12953);
or U15936 (N_15936,N_12305,N_12311);
xor U15937 (N_15937,N_13269,N_12958);
or U15938 (N_15938,N_11141,N_10211);
or U15939 (N_15939,N_12815,N_14622);
xnor U15940 (N_15940,N_11544,N_14695);
and U15941 (N_15941,N_11764,N_10272);
nor U15942 (N_15942,N_11524,N_12268);
nand U15943 (N_15943,N_11495,N_13918);
or U15944 (N_15944,N_11483,N_12043);
or U15945 (N_15945,N_14315,N_10048);
nor U15946 (N_15946,N_11375,N_11461);
nor U15947 (N_15947,N_12407,N_12588);
or U15948 (N_15948,N_12683,N_10583);
or U15949 (N_15949,N_12213,N_14713);
or U15950 (N_15950,N_13342,N_10219);
nor U15951 (N_15951,N_12007,N_12595);
nand U15952 (N_15952,N_12226,N_11601);
and U15953 (N_15953,N_11263,N_11942);
nand U15954 (N_15954,N_10785,N_14575);
or U15955 (N_15955,N_10691,N_12884);
or U15956 (N_15956,N_14262,N_11804);
nand U15957 (N_15957,N_13048,N_12142);
nor U15958 (N_15958,N_11551,N_11612);
nor U15959 (N_15959,N_13323,N_14346);
or U15960 (N_15960,N_13272,N_12623);
nand U15961 (N_15961,N_10888,N_10026);
nand U15962 (N_15962,N_12656,N_13277);
or U15963 (N_15963,N_14745,N_10626);
and U15964 (N_15964,N_12143,N_10413);
and U15965 (N_15965,N_14983,N_10722);
and U15966 (N_15966,N_13019,N_14014);
nor U15967 (N_15967,N_11848,N_13106);
nand U15968 (N_15968,N_10962,N_11329);
and U15969 (N_15969,N_12555,N_14179);
or U15970 (N_15970,N_12528,N_13489);
xnor U15971 (N_15971,N_12779,N_14621);
xnor U15972 (N_15972,N_11621,N_12798);
and U15973 (N_15973,N_10749,N_14008);
nor U15974 (N_15974,N_11500,N_11910);
and U15975 (N_15975,N_13997,N_12647);
xnor U15976 (N_15976,N_11613,N_12207);
and U15977 (N_15977,N_10778,N_10908);
or U15978 (N_15978,N_12310,N_12077);
nor U15979 (N_15979,N_10419,N_11843);
and U15980 (N_15980,N_11311,N_14326);
and U15981 (N_15981,N_13275,N_12094);
or U15982 (N_15982,N_10225,N_14962);
nand U15983 (N_15983,N_13205,N_10354);
nand U15984 (N_15984,N_11570,N_10340);
xor U15985 (N_15985,N_14401,N_11622);
and U15986 (N_15986,N_11173,N_10493);
nor U15987 (N_15987,N_12212,N_13842);
and U15988 (N_15988,N_11124,N_12168);
and U15989 (N_15989,N_10974,N_10652);
and U15990 (N_15990,N_12436,N_12024);
or U15991 (N_15991,N_11595,N_12217);
nor U15992 (N_15992,N_13648,N_10007);
nor U15993 (N_15993,N_10096,N_14576);
nand U15994 (N_15994,N_10358,N_12845);
nand U15995 (N_15995,N_14374,N_14050);
nand U15996 (N_15996,N_12185,N_14795);
and U15997 (N_15997,N_14979,N_10733);
xnor U15998 (N_15998,N_12139,N_11647);
or U15999 (N_15999,N_13837,N_11143);
nand U16000 (N_16000,N_14297,N_12671);
nand U16001 (N_16001,N_13466,N_12840);
or U16002 (N_16002,N_10067,N_13459);
and U16003 (N_16003,N_13155,N_12544);
nand U16004 (N_16004,N_11439,N_14658);
xnor U16005 (N_16005,N_14065,N_11869);
and U16006 (N_16006,N_10342,N_13251);
nor U16007 (N_16007,N_12558,N_13087);
nand U16008 (N_16008,N_13903,N_14071);
or U16009 (N_16009,N_14996,N_11623);
or U16010 (N_16010,N_12335,N_10136);
nand U16011 (N_16011,N_12263,N_10627);
and U16012 (N_16012,N_12380,N_14448);
nor U16013 (N_16013,N_12824,N_13604);
nor U16014 (N_16014,N_14506,N_14534);
and U16015 (N_16015,N_11464,N_14589);
nand U16016 (N_16016,N_11487,N_12255);
nor U16017 (N_16017,N_12244,N_13371);
xnor U16018 (N_16018,N_14764,N_14072);
nor U16019 (N_16019,N_14255,N_13952);
and U16020 (N_16020,N_13894,N_12626);
nor U16021 (N_16021,N_13316,N_10484);
or U16022 (N_16022,N_10113,N_10669);
and U16023 (N_16023,N_11006,N_10768);
and U16024 (N_16024,N_11061,N_11536);
or U16025 (N_16025,N_11952,N_13140);
nor U16026 (N_16026,N_14386,N_13016);
nand U16027 (N_16027,N_10506,N_10915);
nand U16028 (N_16028,N_12134,N_13665);
and U16029 (N_16029,N_12336,N_14127);
xor U16030 (N_16030,N_14507,N_12438);
nor U16031 (N_16031,N_12160,N_10574);
xnor U16032 (N_16032,N_14033,N_14761);
and U16033 (N_16033,N_10077,N_14635);
and U16034 (N_16034,N_13471,N_13213);
nand U16035 (N_16035,N_14678,N_13448);
nor U16036 (N_16036,N_12192,N_12474);
nor U16037 (N_16037,N_12669,N_12378);
and U16038 (N_16038,N_12292,N_13381);
nor U16039 (N_16039,N_12597,N_14707);
nand U16040 (N_16040,N_12892,N_10169);
and U16041 (N_16041,N_14186,N_13519);
nor U16042 (N_16042,N_13741,N_13146);
xor U16043 (N_16043,N_11149,N_10006);
nand U16044 (N_16044,N_14321,N_10650);
nor U16045 (N_16045,N_14414,N_14998);
or U16046 (N_16046,N_12559,N_11559);
nor U16047 (N_16047,N_12039,N_11064);
and U16048 (N_16048,N_12562,N_10292);
nor U16049 (N_16049,N_14579,N_10202);
and U16050 (N_16050,N_14275,N_12225);
nand U16051 (N_16051,N_13267,N_11230);
nand U16052 (N_16052,N_12955,N_14965);
nor U16053 (N_16053,N_13034,N_12697);
nand U16054 (N_16054,N_10929,N_11089);
nor U16055 (N_16055,N_14595,N_12923);
or U16056 (N_16056,N_13293,N_13883);
or U16057 (N_16057,N_13560,N_14933);
nand U16058 (N_16058,N_10166,N_13433);
nor U16059 (N_16059,N_12553,N_11334);
nand U16060 (N_16060,N_11474,N_13773);
nand U16061 (N_16061,N_11618,N_14712);
nand U16062 (N_16062,N_13819,N_14095);
and U16063 (N_16063,N_11092,N_11553);
and U16064 (N_16064,N_12712,N_11165);
or U16065 (N_16065,N_11935,N_11032);
nor U16066 (N_16066,N_13188,N_13366);
nor U16067 (N_16067,N_11851,N_11306);
and U16068 (N_16068,N_11282,N_12250);
and U16069 (N_16069,N_13395,N_14757);
or U16070 (N_16070,N_10835,N_11258);
and U16071 (N_16071,N_14946,N_11674);
and U16072 (N_16072,N_14432,N_14608);
nor U16073 (N_16073,N_12781,N_12230);
and U16074 (N_16074,N_10119,N_11882);
or U16075 (N_16075,N_10317,N_13268);
or U16076 (N_16076,N_12254,N_12787);
nor U16077 (N_16077,N_14966,N_13658);
or U16078 (N_16078,N_10195,N_13474);
or U16079 (N_16079,N_13823,N_12033);
nor U16080 (N_16080,N_10993,N_13463);
xnor U16081 (N_16081,N_12398,N_13753);
or U16082 (N_16082,N_11680,N_13481);
nand U16083 (N_16083,N_10300,N_10874);
nor U16084 (N_16084,N_12731,N_10274);
and U16085 (N_16085,N_11787,N_14459);
and U16086 (N_16086,N_10017,N_11875);
xnor U16087 (N_16087,N_12941,N_11396);
nand U16088 (N_16088,N_11159,N_11826);
nand U16089 (N_16089,N_14746,N_14209);
nand U16090 (N_16090,N_10035,N_10985);
and U16091 (N_16091,N_13351,N_13410);
nand U16092 (N_16092,N_12035,N_12052);
or U16093 (N_16093,N_13105,N_14486);
and U16094 (N_16094,N_12386,N_13653);
and U16095 (N_16095,N_10678,N_11280);
and U16096 (N_16096,N_14423,N_13579);
nor U16097 (N_16097,N_14793,N_12583);
nand U16098 (N_16098,N_12358,N_14562);
or U16099 (N_16099,N_13993,N_10360);
or U16100 (N_16100,N_14034,N_14496);
nand U16101 (N_16101,N_10333,N_12522);
nand U16102 (N_16102,N_10783,N_14470);
nor U16103 (N_16103,N_11381,N_14442);
nor U16104 (N_16104,N_10942,N_12433);
xnor U16105 (N_16105,N_11577,N_10343);
or U16106 (N_16106,N_10842,N_12556);
or U16107 (N_16107,N_10061,N_12981);
or U16108 (N_16108,N_10765,N_10312);
nand U16109 (N_16109,N_10964,N_11837);
nor U16110 (N_16110,N_10347,N_11112);
nand U16111 (N_16111,N_12737,N_10254);
and U16112 (N_16112,N_14445,N_10126);
or U16113 (N_16113,N_10871,N_14499);
xnor U16114 (N_16114,N_10192,N_11671);
nand U16115 (N_16115,N_11303,N_12757);
or U16116 (N_16116,N_11599,N_10563);
and U16117 (N_16117,N_13623,N_13977);
or U16118 (N_16118,N_14462,N_10638);
and U16119 (N_16119,N_13961,N_13027);
nor U16120 (N_16120,N_12821,N_14013);
nor U16121 (N_16121,N_11631,N_12391);
xnor U16122 (N_16122,N_11645,N_11283);
and U16123 (N_16123,N_14131,N_10042);
or U16124 (N_16124,N_14846,N_14092);
or U16125 (N_16125,N_13578,N_14116);
or U16126 (N_16126,N_14605,N_11974);
nand U16127 (N_16127,N_11963,N_11044);
nor U16128 (N_16128,N_13062,N_13563);
and U16129 (N_16129,N_14142,N_11516);
nor U16130 (N_16130,N_10800,N_13679);
nor U16131 (N_16131,N_12796,N_14512);
or U16132 (N_16132,N_13328,N_12264);
nand U16133 (N_16133,N_10833,N_10499);
or U16134 (N_16134,N_10976,N_13710);
or U16135 (N_16135,N_12338,N_10984);
xnor U16136 (N_16136,N_10238,N_11781);
nor U16137 (N_16137,N_13570,N_14766);
nand U16138 (N_16138,N_13258,N_12571);
or U16139 (N_16139,N_11864,N_14108);
nand U16140 (N_16140,N_11308,N_11454);
xor U16141 (N_16141,N_12502,N_10282);
nor U16142 (N_16142,N_14073,N_11132);
or U16143 (N_16143,N_12551,N_13743);
or U16144 (N_16144,N_14472,N_10979);
and U16145 (N_16145,N_12771,N_10001);
nor U16146 (N_16146,N_13633,N_10546);
and U16147 (N_16147,N_10560,N_14409);
or U16148 (N_16148,N_10746,N_13979);
or U16149 (N_16149,N_10685,N_13383);
xor U16150 (N_16150,N_12282,N_13430);
and U16151 (N_16151,N_11861,N_13910);
nor U16152 (N_16152,N_11574,N_14849);
xnor U16153 (N_16153,N_10305,N_13424);
or U16154 (N_16154,N_12561,N_14080);
or U16155 (N_16155,N_11425,N_10391);
and U16156 (N_16156,N_13185,N_13795);
or U16157 (N_16157,N_11866,N_12925);
xor U16158 (N_16158,N_11003,N_12274);
and U16159 (N_16159,N_11372,N_11060);
nand U16160 (N_16160,N_14602,N_14272);
or U16161 (N_16161,N_14197,N_14723);
and U16162 (N_16162,N_11572,N_13475);
and U16163 (N_16163,N_13783,N_14720);
or U16164 (N_16164,N_12615,N_10223);
nor U16165 (N_16165,N_10847,N_12592);
nand U16166 (N_16166,N_14528,N_11279);
nand U16167 (N_16167,N_12654,N_10421);
or U16168 (N_16168,N_12271,N_11754);
nor U16169 (N_16169,N_10610,N_10660);
xor U16170 (N_16170,N_10732,N_10123);
and U16171 (N_16171,N_12272,N_10468);
and U16172 (N_16172,N_10869,N_11129);
nand U16173 (N_16173,N_10182,N_11358);
and U16174 (N_16174,N_13046,N_13178);
nor U16175 (N_16175,N_13152,N_14967);
or U16176 (N_16176,N_12315,N_11948);
or U16177 (N_16177,N_12652,N_12266);
nand U16178 (N_16178,N_14140,N_13312);
nor U16179 (N_16179,N_11084,N_11718);
nor U16180 (N_16180,N_12706,N_11075);
or U16181 (N_16181,N_13884,N_13352);
xnor U16182 (N_16182,N_12709,N_14264);
and U16183 (N_16183,N_12944,N_11830);
and U16184 (N_16184,N_10079,N_14124);
or U16185 (N_16185,N_14213,N_13060);
and U16186 (N_16186,N_13180,N_13413);
and U16187 (N_16187,N_13415,N_10147);
nand U16188 (N_16188,N_14801,N_12098);
or U16189 (N_16189,N_13727,N_12483);
nand U16190 (N_16190,N_12269,N_14645);
and U16191 (N_16191,N_12572,N_12163);
or U16192 (N_16192,N_14724,N_13021);
nor U16193 (N_16193,N_11873,N_10471);
xnor U16194 (N_16194,N_11121,N_14668);
and U16195 (N_16195,N_14908,N_11229);
nand U16196 (N_16196,N_13933,N_14188);
nor U16197 (N_16197,N_13772,N_12885);
and U16198 (N_16198,N_13491,N_13002);
and U16199 (N_16199,N_12612,N_14163);
nor U16200 (N_16200,N_11243,N_11421);
nor U16201 (N_16201,N_11277,N_13799);
or U16202 (N_16202,N_10482,N_13135);
or U16203 (N_16203,N_13082,N_12501);
or U16204 (N_16204,N_11020,N_13089);
nor U16205 (N_16205,N_11920,N_11768);
or U16206 (N_16206,N_13278,N_14365);
or U16207 (N_16207,N_13902,N_12140);
and U16208 (N_16208,N_12983,N_13195);
xor U16209 (N_16209,N_13595,N_14458);
and U16210 (N_16210,N_13609,N_14060);
nand U16211 (N_16211,N_12406,N_13700);
and U16212 (N_16212,N_10155,N_12090);
or U16213 (N_16213,N_13780,N_13556);
nand U16214 (N_16214,N_12631,N_13123);
nor U16215 (N_16215,N_13980,N_14559);
nand U16216 (N_16216,N_10389,N_10094);
and U16217 (N_16217,N_13449,N_11701);
or U16218 (N_16218,N_14421,N_11747);
nor U16219 (N_16219,N_10947,N_14939);
nor U16220 (N_16220,N_11597,N_10266);
or U16221 (N_16221,N_14164,N_11520);
nor U16222 (N_16222,N_13297,N_14930);
nand U16223 (N_16223,N_10670,N_14719);
and U16224 (N_16224,N_13965,N_11546);
nor U16225 (N_16225,N_10351,N_13259);
and U16226 (N_16226,N_13198,N_12072);
and U16227 (N_16227,N_13209,N_14682);
nor U16228 (N_16228,N_14101,N_11417);
nor U16229 (N_16229,N_10812,N_12905);
nand U16230 (N_16230,N_13695,N_12220);
and U16231 (N_16231,N_10483,N_10782);
and U16232 (N_16232,N_11892,N_11352);
or U16233 (N_16233,N_10995,N_10952);
or U16234 (N_16234,N_14170,N_14948);
and U16235 (N_16235,N_10661,N_14937);
nor U16236 (N_16236,N_12405,N_12870);
nor U16237 (N_16237,N_13912,N_13745);
nor U16238 (N_16238,N_10112,N_12708);
or U16239 (N_16239,N_14741,N_10188);
nand U16240 (N_16240,N_11926,N_13274);
or U16241 (N_16241,N_13202,N_14330);
xnor U16242 (N_16242,N_14439,N_10723);
nor U16243 (N_16243,N_10474,N_11387);
or U16244 (N_16244,N_14782,N_14844);
xor U16245 (N_16245,N_11679,N_13183);
nor U16246 (N_16246,N_12584,N_13516);
or U16247 (N_16247,N_14405,N_14755);
xnor U16248 (N_16248,N_10259,N_11773);
or U16249 (N_16249,N_14872,N_14560);
nand U16250 (N_16250,N_11491,N_10786);
and U16251 (N_16251,N_13651,N_10489);
xor U16252 (N_16252,N_14375,N_14599);
or U16253 (N_16253,N_13616,N_10229);
xor U16254 (N_16254,N_11219,N_11984);
and U16255 (N_16255,N_12931,N_13049);
xnor U16256 (N_16256,N_14597,N_10162);
or U16257 (N_16257,N_14820,N_11380);
or U16258 (N_16258,N_12240,N_13591);
or U16259 (N_16259,N_13377,N_10429);
nor U16260 (N_16260,N_10177,N_13429);
nand U16261 (N_16261,N_12342,N_13968);
nand U16262 (N_16262,N_11840,N_14556);
nand U16263 (N_16263,N_12345,N_11049);
or U16264 (N_16264,N_11420,N_11542);
nor U16265 (N_16265,N_10452,N_11678);
and U16266 (N_16266,N_13861,N_14809);
nor U16267 (N_16267,N_12806,N_13301);
and U16268 (N_16268,N_11883,N_14158);
nor U16269 (N_16269,N_13244,N_11774);
nand U16270 (N_16270,N_12756,N_14902);
nor U16271 (N_16271,N_13676,N_12155);
and U16272 (N_16272,N_12316,N_10819);
nand U16273 (N_16273,N_14883,N_11260);
nor U16274 (N_16274,N_13924,N_10349);
or U16275 (N_16275,N_13041,N_11153);
and U16276 (N_16276,N_13987,N_12539);
and U16277 (N_16277,N_10328,N_13746);
or U16278 (N_16278,N_13576,N_10883);
nor U16279 (N_16279,N_12943,N_13864);
xor U16280 (N_16280,N_10402,N_13357);
or U16281 (N_16281,N_14896,N_10616);
or U16282 (N_16282,N_12022,N_12341);
nor U16283 (N_16283,N_14877,N_13501);
nor U16284 (N_16284,N_13038,N_13622);
and U16285 (N_16285,N_11683,N_11651);
or U16286 (N_16286,N_13037,N_13158);
or U16287 (N_16287,N_10831,N_12807);
and U16288 (N_16288,N_13524,N_12729);
or U16289 (N_16289,N_14887,N_12755);
nand U16290 (N_16290,N_14815,N_12628);
or U16291 (N_16291,N_11834,N_14744);
or U16292 (N_16292,N_14747,N_11515);
and U16293 (N_16293,N_12866,N_14169);
nand U16294 (N_16294,N_13334,N_12701);
nand U16295 (N_16295,N_14914,N_12515);
or U16296 (N_16296,N_12859,N_12102);
nand U16297 (N_16297,N_14406,N_13671);
or U16298 (N_16298,N_12867,N_14798);
or U16299 (N_16299,N_14961,N_11914);
and U16300 (N_16300,N_10099,N_10116);
nand U16301 (N_16301,N_14102,N_13302);
and U16302 (N_16302,N_14353,N_10240);
and U16303 (N_16303,N_12318,N_12769);
xnor U16304 (N_16304,N_14007,N_10704);
nand U16305 (N_16305,N_14800,N_10193);
and U16306 (N_16306,N_14609,N_12604);
and U16307 (N_16307,N_13043,N_11449);
nor U16308 (N_16308,N_10894,N_13832);
nand U16309 (N_16309,N_13125,N_10866);
nand U16310 (N_16310,N_12088,N_12759);
and U16311 (N_16311,N_11765,N_10537);
and U16312 (N_16312,N_13398,N_11994);
and U16313 (N_16313,N_11462,N_13273);
nor U16314 (N_16314,N_14928,N_14637);
or U16315 (N_16315,N_12732,N_14769);
or U16316 (N_16316,N_11036,N_11478);
nor U16317 (N_16317,N_12379,N_12567);
nor U16318 (N_16318,N_13441,N_12340);
or U16319 (N_16319,N_13485,N_11771);
and U16320 (N_16320,N_10770,N_11563);
nor U16321 (N_16321,N_13531,N_10299);
nand U16322 (N_16322,N_11068,N_11712);
nor U16323 (N_16323,N_13390,N_10270);
or U16324 (N_16324,N_10559,N_10198);
xnor U16325 (N_16325,N_10605,N_14814);
and U16326 (N_16326,N_11079,N_12762);
or U16327 (N_16327,N_11333,N_12181);
and U16328 (N_16328,N_10138,N_13833);
nor U16329 (N_16329,N_11271,N_13203);
and U16330 (N_16330,N_12858,N_11972);
and U16331 (N_16331,N_11031,N_11235);
nand U16332 (N_16332,N_14875,N_13626);
and U16333 (N_16333,N_12141,N_13243);
xnor U16334 (N_16334,N_14175,N_14117);
xnor U16335 (N_16335,N_12533,N_10203);
nand U16336 (N_16336,N_11299,N_11014);
nand U16337 (N_16337,N_12261,N_14811);
and U16338 (N_16338,N_14294,N_12370);
nand U16339 (N_16339,N_14901,N_10509);
nor U16340 (N_16340,N_10977,N_14184);
or U16341 (N_16341,N_12027,N_10322);
or U16342 (N_16342,N_12700,N_13930);
and U16343 (N_16343,N_14107,N_12984);
or U16344 (N_16344,N_12464,N_10504);
or U16345 (N_16345,N_10133,N_12101);
nor U16346 (N_16346,N_14337,N_13014);
and U16347 (N_16347,N_11486,N_10191);
nor U16348 (N_16348,N_12127,N_10562);
nor U16349 (N_16349,N_12086,N_12466);
and U16350 (N_16350,N_10664,N_13641);
and U16351 (N_16351,N_12177,N_14026);
nor U16352 (N_16352,N_12738,N_13505);
nand U16353 (N_16353,N_10232,N_13362);
nor U16354 (N_16354,N_12175,N_12734);
or U16355 (N_16355,N_14517,N_10515);
nand U16356 (N_16356,N_13064,N_14839);
nor U16357 (N_16357,N_14480,N_11510);
xnor U16358 (N_16358,N_12300,N_14389);
nor U16359 (N_16359,N_14541,N_14348);
and U16360 (N_16360,N_14260,N_11819);
nor U16361 (N_16361,N_13673,N_12164);
nor U16362 (N_16362,N_10277,N_11354);
and U16363 (N_16363,N_11991,N_10567);
nand U16364 (N_16364,N_14415,N_11181);
and U16365 (N_16365,N_14710,N_13983);
or U16366 (N_16366,N_14565,N_13617);
or U16367 (N_16367,N_14450,N_10180);
nor U16368 (N_16368,N_10682,N_11249);
nor U16369 (N_16369,N_10207,N_12838);
and U16370 (N_16370,N_12609,N_12547);
or U16371 (N_16371,N_14452,N_12860);
or U16372 (N_16372,N_10408,N_13939);
nor U16373 (N_16373,N_13074,N_14673);
xnor U16374 (N_16374,N_14545,N_13654);
nand U16375 (N_16375,N_10535,N_10998);
and U16376 (N_16376,N_12895,N_11379);
nor U16377 (N_16377,N_14826,N_13954);
and U16378 (N_16378,N_10142,N_13121);
and U16379 (N_16379,N_14273,N_14483);
nand U16380 (N_16380,N_12964,N_10920);
and U16381 (N_16381,N_13219,N_13149);
or U16382 (N_16382,N_14384,N_14133);
and U16383 (N_16383,N_13040,N_12720);
nor U16384 (N_16384,N_12392,N_14147);
and U16385 (N_16385,N_13151,N_13994);
and U16386 (N_16386,N_11494,N_10102);
nand U16387 (N_16387,N_12128,N_11605);
xnor U16388 (N_16388,N_13822,N_12294);
nor U16389 (N_16389,N_13596,N_14136);
nor U16390 (N_16390,N_13242,N_11723);
nand U16391 (N_16391,N_10877,N_12089);
nand U16392 (N_16392,N_12888,N_12215);
nand U16393 (N_16393,N_12517,N_11267);
or U16394 (N_16394,N_13685,N_10085);
nor U16395 (N_16395,N_12349,N_11485);
nand U16396 (N_16396,N_12668,N_13857);
nor U16397 (N_16397,N_13315,N_12917);
or U16398 (N_16398,N_14508,N_11695);
nand U16399 (N_16399,N_13482,N_11398);
and U16400 (N_16400,N_11004,N_10945);
nand U16401 (N_16401,N_12799,N_14215);
nand U16402 (N_16402,N_10939,N_11624);
and U16403 (N_16403,N_10568,N_10315);
or U16404 (N_16404,N_14139,N_12935);
xnor U16405 (N_16405,N_14689,N_12051);
or U16406 (N_16406,N_10331,N_12148);
and U16407 (N_16407,N_14661,N_11555);
nor U16408 (N_16408,N_10826,N_11175);
nor U16409 (N_16409,N_12750,N_11403);
nor U16410 (N_16410,N_11448,N_10378);
and U16411 (N_16411,N_12399,N_10185);
or U16412 (N_16412,N_14917,N_14789);
nor U16413 (N_16413,N_13548,N_12453);
nand U16414 (N_16414,N_14920,N_13470);
and U16415 (N_16415,N_13072,N_10208);
nand U16416 (N_16416,N_12402,N_11710);
nor U16417 (N_16417,N_14426,N_11331);
nand U16418 (N_16418,N_10857,N_14115);
and U16419 (N_16419,N_14408,N_10163);
nor U16420 (N_16420,N_10886,N_13024);
and U16421 (N_16421,N_14681,N_11867);
nand U16422 (N_16422,N_11793,N_10242);
nand U16423 (N_16423,N_13990,N_14028);
nand U16424 (N_16424,N_13543,N_13399);
nor U16425 (N_16425,N_12097,N_13030);
nand U16426 (N_16426,N_14829,N_11610);
nor U16427 (N_16427,N_11629,N_14832);
and U16428 (N_16428,N_14987,N_12055);
nand U16429 (N_16429,N_12724,N_14182);
nand U16430 (N_16430,N_10607,N_12376);
nor U16431 (N_16431,N_14807,N_12743);
nand U16432 (N_16432,N_14929,N_12872);
nand U16433 (N_16433,N_10640,N_13897);
or U16434 (N_16434,N_12739,N_10014);
nor U16435 (N_16435,N_10396,N_13534);
or U16436 (N_16436,N_11000,N_13920);
and U16437 (N_16437,N_11604,N_10459);
or U16438 (N_16438,N_12124,N_10948);
nor U16439 (N_16439,N_12346,N_12834);
and U16440 (N_16440,N_11824,N_14995);
or U16441 (N_16441,N_13179,N_13401);
nand U16442 (N_16442,N_10878,N_10780);
nor U16443 (N_16443,N_10972,N_11492);
or U16444 (N_16444,N_10556,N_11583);
nor U16445 (N_16445,N_12753,N_13337);
nor U16446 (N_16446,N_12643,N_13957);
or U16447 (N_16447,N_13742,N_13973);
xor U16448 (N_16448,N_14396,N_10747);
xnor U16449 (N_16449,N_10481,N_14242);
and U16450 (N_16450,N_14191,N_12180);
or U16451 (N_16451,N_10604,N_10371);
nor U16452 (N_16452,N_10087,N_13662);
nand U16453 (N_16453,N_14481,N_14141);
nor U16454 (N_16454,N_11413,N_10906);
or U16455 (N_16455,N_10851,N_10076);
xnor U16456 (N_16456,N_14363,N_13182);
nand U16457 (N_16457,N_13118,N_12062);
nand U16458 (N_16458,N_11066,N_14787);
or U16459 (N_16459,N_11939,N_14955);
and U16460 (N_16460,N_12104,N_12197);
xor U16461 (N_16461,N_12500,N_13299);
nand U16462 (N_16462,N_11362,N_11876);
and U16463 (N_16463,N_14304,N_10409);
nor U16464 (N_16464,N_10773,N_13090);
nand U16465 (N_16465,N_11817,N_11749);
nor U16466 (N_16466,N_14692,N_13882);
and U16467 (N_16467,N_10033,N_13571);
and U16468 (N_16468,N_10329,N_10668);
nor U16469 (N_16469,N_14797,N_11028);
nor U16470 (N_16470,N_11038,N_12545);
and U16471 (N_16471,N_12788,N_11693);
nor U16472 (N_16472,N_11356,N_10124);
nand U16473 (N_16473,N_10427,N_10628);
or U16474 (N_16474,N_10701,N_14413);
and U16475 (N_16475,N_13091,N_12252);
nand U16476 (N_16476,N_12297,N_13095);
nor U16477 (N_16477,N_14509,N_12792);
nor U16478 (N_16478,N_13246,N_12199);
nor U16479 (N_16479,N_10251,N_11076);
xnor U16480 (N_16480,N_10675,N_12661);
xnor U16481 (N_16481,N_11393,N_13150);
nand U16482 (N_16482,N_12301,N_11285);
or U16483 (N_16483,N_13349,N_13784);
nand U16484 (N_16484,N_13901,N_12223);
and U16485 (N_16485,N_14118,N_10407);
and U16486 (N_16486,N_12165,N_12095);
and U16487 (N_16487,N_14278,N_11600);
or U16488 (N_16488,N_10896,N_10470);
nor U16489 (N_16489,N_13100,N_10862);
nand U16490 (N_16490,N_12969,N_14510);
nand U16491 (N_16491,N_12239,N_13212);
nand U16492 (N_16492,N_14119,N_11187);
and U16493 (N_16493,N_12123,N_12897);
xor U16494 (N_16494,N_14923,N_12456);
xnor U16495 (N_16495,N_12831,N_11756);
nor U16496 (N_16496,N_12758,N_11236);
and U16497 (N_16497,N_10794,N_14043);
or U16498 (N_16498,N_13540,N_13669);
nand U16499 (N_16499,N_13851,N_12084);
nor U16500 (N_16500,N_10028,N_14627);
nor U16501 (N_16501,N_13455,N_13109);
nand U16502 (N_16502,N_14980,N_11480);
or U16503 (N_16503,N_11809,N_12782);
or U16504 (N_16504,N_14204,N_10796);
nor U16505 (N_16505,N_11346,N_10631);
nor U16506 (N_16506,N_12999,N_10134);
nor U16507 (N_16507,N_13306,N_14176);
xnor U16508 (N_16508,N_13068,N_10214);
or U16509 (N_16509,N_14266,N_11669);
or U16510 (N_16510,N_10713,N_12927);
and U16511 (N_16511,N_14227,N_12067);
or U16512 (N_16512,N_14403,N_10792);
and U16513 (N_16513,N_10542,N_12826);
xor U16514 (N_16514,N_11040,N_11728);
nor U16515 (N_16515,N_11603,N_10588);
or U16516 (N_16516,N_12819,N_13546);
nand U16517 (N_16517,N_11967,N_10986);
or U16518 (N_16518,N_11319,N_13281);
nor U16519 (N_16519,N_10832,N_11877);
xor U16520 (N_16520,N_10889,N_14361);
nand U16521 (N_16521,N_14770,N_10383);
nand U16522 (N_16522,N_12028,N_13550);
or U16523 (N_16523,N_14249,N_10141);
nand U16524 (N_16524,N_11881,N_12137);
or U16525 (N_16525,N_10975,N_12312);
or U16526 (N_16526,N_11981,N_10171);
or U16527 (N_16527,N_14752,N_12397);
and U16528 (N_16528,N_13348,N_12428);
xnor U16529 (N_16529,N_12372,N_12233);
xnor U16530 (N_16530,N_11797,N_11552);
or U16531 (N_16531,N_13937,N_10748);
nand U16532 (N_16532,N_12667,N_13668);
or U16533 (N_16533,N_14876,N_14503);
or U16534 (N_16534,N_11508,N_12921);
or U16535 (N_16535,N_11168,N_11720);
or U16536 (N_16536,N_14298,N_11916);
or U16537 (N_16537,N_14203,N_11737);
and U16538 (N_16538,N_12279,N_14226);
and U16539 (N_16539,N_10009,N_10636);
or U16540 (N_16540,N_10840,N_13896);
nand U16541 (N_16541,N_10516,N_10587);
nor U16542 (N_16542,N_10946,N_13478);
nor U16543 (N_16543,N_13161,N_11614);
nand U16544 (N_16544,N_13964,N_11459);
and U16545 (N_16545,N_14571,N_13184);
nand U16546 (N_16546,N_13934,N_13132);
or U16547 (N_16547,N_14159,N_11446);
nor U16548 (N_16548,N_13097,N_10319);
or U16549 (N_16549,N_13667,N_13530);
or U16550 (N_16550,N_10374,N_10573);
or U16551 (N_16551,N_13322,N_13564);
nor U16552 (N_16552,N_13631,N_14548);
or U16553 (N_16553,N_12193,N_11234);
xnor U16554 (N_16554,N_14319,N_10478);
and U16555 (N_16555,N_11534,N_11479);
and U16556 (N_16556,N_14786,N_10816);
and U16557 (N_16557,N_12846,N_12448);
or U16558 (N_16558,N_12616,N_10381);
xor U16559 (N_16559,N_10737,N_11072);
and U16560 (N_16560,N_14340,N_13601);
xor U16561 (N_16561,N_13452,N_13330);
nand U16562 (N_16562,N_11938,N_14806);
xnor U16563 (N_16563,N_10455,N_11541);
and U16564 (N_16564,N_11100,N_11309);
or U16565 (N_16565,N_13045,N_12534);
nor U16566 (N_16566,N_13488,N_14207);
or U16567 (N_16567,N_10253,N_14957);
nand U16568 (N_16568,N_12907,N_13250);
or U16569 (N_16569,N_10137,N_13115);
nand U16570 (N_16570,N_13283,N_10456);
nor U16571 (N_16571,N_14356,N_14910);
nor U16572 (N_16572,N_12390,N_14222);
nor U16573 (N_16573,N_13333,N_11138);
or U16574 (N_16574,N_13552,N_14606);
and U16575 (N_16575,N_12025,N_13508);
xnor U16576 (N_16576,N_14813,N_11189);
and U16577 (N_16577,N_13112,N_10803);
nand U16578 (N_16578,N_13523,N_13976);
nand U16579 (N_16579,N_13969,N_11321);
nand U16580 (N_16580,N_12721,N_10968);
nor U16581 (N_16581,N_13614,N_13751);
or U16582 (N_16582,N_13077,N_11221);
or U16583 (N_16583,N_11501,N_13581);
nand U16584 (N_16584,N_14265,N_11224);
and U16585 (N_16585,N_13216,N_10541);
nand U16586 (N_16586,N_10058,N_14256);
or U16587 (N_16587,N_11709,N_10410);
nor U16588 (N_16588,N_13174,N_11316);
nor U16589 (N_16589,N_11731,N_14328);
and U16590 (N_16590,N_13144,N_11035);
and U16591 (N_16591,N_11936,N_10787);
nor U16592 (N_16592,N_13484,N_12003);
or U16593 (N_16593,N_13893,N_11337);
nor U16594 (N_16594,N_13436,N_12861);
and U16595 (N_16595,N_14583,N_10412);
xnor U16596 (N_16596,N_11139,N_10084);
or U16597 (N_16597,N_11430,N_10097);
nor U16598 (N_16598,N_14553,N_12536);
nand U16599 (N_16599,N_11490,N_13582);
nand U16600 (N_16600,N_12443,N_12131);
or U16601 (N_16601,N_12326,N_13098);
and U16602 (N_16602,N_14161,N_10384);
nand U16603 (N_16603,N_14768,N_11026);
or U16604 (N_16604,N_13096,N_10918);
xor U16605 (N_16605,N_11496,N_12401);
and U16606 (N_16606,N_10114,N_11736);
and U16607 (N_16607,N_14737,N_11015);
or U16608 (N_16608,N_12122,N_10261);
or U16609 (N_16609,N_13854,N_13613);
nand U16610 (N_16610,N_12485,N_11109);
nor U16611 (N_16611,N_14027,N_14716);
and U16612 (N_16612,N_11686,N_13464);
nor U16613 (N_16613,N_14251,N_11713);
and U16614 (N_16614,N_12491,N_10439);
nand U16615 (N_16615,N_12224,N_13716);
nor U16616 (N_16616,N_13808,N_13916);
nand U16617 (N_16617,N_13354,N_14128);
nand U16618 (N_16618,N_10633,N_14056);
and U16619 (N_16619,N_14491,N_12995);
nand U16620 (N_16620,N_12189,N_10570);
xnor U16621 (N_16621,N_11707,N_14366);
and U16622 (N_16622,N_14497,N_10838);
or U16623 (N_16623,N_14899,N_12742);
or U16624 (N_16624,N_10931,N_14558);
nor U16625 (N_16625,N_11606,N_11365);
or U16626 (N_16626,N_13733,N_13944);
nor U16627 (N_16627,N_14827,N_14628);
or U16628 (N_16628,N_13300,N_10289);
or U16629 (N_16629,N_12314,N_12296);
nand U16630 (N_16630,N_11833,N_11383);
nor U16631 (N_16631,N_11292,N_11767);
or U16632 (N_16632,N_13747,N_10892);
and U16633 (N_16633,N_14550,N_10045);
nor U16634 (N_16634,N_14613,N_12728);
nand U16635 (N_16635,N_10736,N_13253);
nand U16636 (N_16636,N_13868,N_14200);
and U16637 (N_16637,N_13444,N_10586);
nand U16638 (N_16638,N_12446,N_10044);
nand U16639 (N_16639,N_14018,N_10529);
nand U16640 (N_16640,N_13391,N_12387);
and U16641 (N_16641,N_14311,N_11625);
nor U16642 (N_16642,N_14437,N_12966);
or U16643 (N_16643,N_14057,N_11724);
nor U16644 (N_16644,N_12693,N_14871);
xor U16645 (N_16645,N_11395,N_12530);
or U16646 (N_16646,N_13869,N_11434);
xnor U16647 (N_16647,N_14934,N_12195);
and U16648 (N_16648,N_11164,N_13003);
nor U16649 (N_16649,N_11589,N_11719);
xnor U16650 (N_16650,N_12021,N_10845);
nand U16651 (N_16651,N_14753,N_13147);
nand U16652 (N_16652,N_11894,N_14368);
nor U16653 (N_16653,N_11816,N_14024);
xnor U16654 (N_16654,N_10970,N_10010);
nor U16655 (N_16655,N_12880,N_10999);
xnor U16656 (N_16656,N_11556,N_11700);
xnor U16657 (N_16657,N_12621,N_11528);
and U16658 (N_16658,N_12480,N_11887);
or U16659 (N_16659,N_10379,N_12308);
and U16660 (N_16660,N_11083,N_13411);
nor U16661 (N_16661,N_13539,N_10156);
nand U16662 (N_16662,N_13051,N_10725);
and U16663 (N_16663,N_12355,N_12105);
or U16664 (N_16664,N_13603,N_10263);
or U16665 (N_16665,N_12396,N_14669);
nor U16666 (N_16666,N_11237,N_14563);
nand U16667 (N_16667,N_14838,N_11128);
nand U16668 (N_16668,N_13247,N_10531);
or U16669 (N_16669,N_10047,N_11336);
and U16670 (N_16670,N_11823,N_12091);
or U16671 (N_16671,N_10554,N_12065);
or U16672 (N_16672,N_10505,N_12579);
nor U16673 (N_16673,N_12736,N_11081);
and U16674 (N_16674,N_11339,N_11940);
xnor U16675 (N_16675,N_10060,N_14636);
or U16676 (N_16676,N_12648,N_10065);
or U16677 (N_16677,N_12598,N_10310);
nor U16678 (N_16678,N_14498,N_14022);
nor U16679 (N_16679,N_12479,N_12078);
nand U16680 (N_16680,N_10643,N_12232);
xnor U16681 (N_16681,N_11150,N_13885);
nand U16682 (N_16682,N_14927,N_11289);
and U16683 (N_16683,N_11832,N_14783);
nor U16684 (N_16684,N_13319,N_14149);
nor U16685 (N_16685,N_12259,N_14354);
or U16686 (N_16686,N_13365,N_12657);
nand U16687 (N_16687,N_14825,N_10268);
or U16688 (N_16688,N_11190,N_12766);
nor U16689 (N_16689,N_12495,N_13649);
and U16690 (N_16690,N_14680,N_10160);
and U16691 (N_16691,N_10558,N_12427);
nand U16692 (N_16692,N_11222,N_12537);
xnor U16693 (N_16693,N_11171,N_12573);
nor U16694 (N_16694,N_14799,N_10196);
or U16695 (N_16695,N_12962,N_14524);
nor U16696 (N_16696,N_14402,N_11871);
and U16697 (N_16697,N_12169,N_12206);
nor U16698 (N_16698,N_11511,N_13023);
nor U16699 (N_16699,N_12804,N_11037);
nor U16700 (N_16700,N_13215,N_11119);
nor U16701 (N_16701,N_14362,N_11370);
nor U16702 (N_16702,N_10519,N_11444);
or U16703 (N_16703,N_13166,N_12287);
nor U16704 (N_16704,N_11178,N_14391);
xnor U16705 (N_16705,N_10281,N_13170);
nand U16706 (N_16706,N_13295,N_12331);
nor U16707 (N_16707,N_10754,N_12689);
xor U16708 (N_16708,N_14373,N_11318);
and U16709 (N_16709,N_12135,N_12839);
or U16710 (N_16710,N_10370,N_10924);
nand U16711 (N_16711,N_10957,N_11155);
nor U16712 (N_16712,N_10969,N_10971);
nor U16713 (N_16713,N_11048,N_14160);
nor U16714 (N_16714,N_13955,N_12828);
nor U16715 (N_16715,N_11965,N_11246);
xor U16716 (N_16716,N_12538,N_14224);
or U16717 (N_16717,N_10959,N_14240);
nand U16718 (N_16718,N_11891,N_12343);
and U16719 (N_16719,N_12624,N_13042);
or U16720 (N_16720,N_10880,N_13782);
and U16721 (N_16721,N_10916,N_12412);
or U16722 (N_16722,N_12727,N_12776);
nand U16723 (N_16723,N_12949,N_14394);
nor U16724 (N_16724,N_12079,N_13573);
and U16725 (N_16725,N_13011,N_12902);
nor U16726 (N_16726,N_12642,N_13820);
or U16727 (N_16727,N_10298,N_13718);
or U16728 (N_16728,N_13001,N_13627);
nand U16729 (N_16729,N_11738,N_12939);
and U16730 (N_16730,N_11194,N_13638);
nor U16731 (N_16731,N_10656,N_11681);
nor U16732 (N_16732,N_11888,N_10283);
xor U16733 (N_16733,N_14004,N_14523);
or U16734 (N_16734,N_10673,N_11408);
nor U16735 (N_16735,N_10750,N_10127);
or U16736 (N_16736,N_10376,N_13231);
nand U16737 (N_16737,N_12980,N_11384);
nand U16738 (N_16738,N_14137,N_11473);
nand U16739 (N_16739,N_12157,N_10944);
nand U16740 (N_16740,N_13168,N_11163);
and U16741 (N_16741,N_12636,N_14733);
and U16742 (N_16742,N_11223,N_11609);
nor U16743 (N_16743,N_13815,N_11660);
or U16744 (N_16744,N_12045,N_13359);
or U16745 (N_16745,N_14177,N_13194);
nand U16746 (N_16746,N_12696,N_14267);
nor U16747 (N_16747,N_13697,N_14312);
and U16748 (N_16748,N_12605,N_10553);
and U16749 (N_16749,N_13029,N_10953);
or U16750 (N_16750,N_13310,N_11620);
or U16751 (N_16751,N_13063,N_13372);
nand U16752 (N_16752,N_11922,N_10618);
or U16753 (N_16753,N_12377,N_11467);
nand U16754 (N_16754,N_10318,N_11661);
nand U16755 (N_16755,N_13338,N_11192);
or U16756 (N_16756,N_13067,N_14986);
nand U16757 (N_16757,N_11007,N_13652);
xor U16758 (N_16758,N_13476,N_14295);
or U16759 (N_16759,N_12716,N_13922);
nand U16760 (N_16760,N_10135,N_14350);
nand U16761 (N_16761,N_14794,N_13527);
xnor U16762 (N_16762,N_12112,N_13065);
and U16763 (N_16763,N_10303,N_12967);
and U16764 (N_16764,N_14958,N_12634);
and U16765 (N_16765,N_10676,N_14756);
nand U16766 (N_16766,N_13752,N_10425);
or U16767 (N_16767,N_12147,N_10821);
and U16768 (N_16768,N_10551,N_14537);
and U16769 (N_16769,N_10367,N_11276);
and U16770 (N_16770,N_14729,N_11954);
nor U16771 (N_16771,N_13899,N_13877);
nand U16772 (N_16772,N_12132,N_11186);
nor U16773 (N_16773,N_14705,N_13460);
or U16774 (N_16774,N_14894,N_12574);
nor U16775 (N_16775,N_13012,N_13260);
and U16776 (N_16776,N_14614,N_13975);
nand U16777 (N_16777,N_14268,N_11968);
and U16778 (N_16778,N_14918,N_14697);
or U16779 (N_16779,N_11481,N_11642);
nand U16780 (N_16780,N_11010,N_13826);
or U16781 (N_16781,N_13446,N_13483);
or U16782 (N_16782,N_10801,N_12237);
nand U16783 (N_16783,N_11529,N_13923);
or U16784 (N_16784,N_10245,N_10465);
or U16785 (N_16785,N_11856,N_12630);
or U16786 (N_16786,N_11361,N_10647);
or U16787 (N_16787,N_11677,N_10881);
and U16788 (N_16788,N_12959,N_11784);
xnor U16789 (N_16789,N_10153,N_12784);
nor U16790 (N_16790,N_13871,N_11855);
or U16791 (N_16791,N_12008,N_13479);
xnor U16792 (N_16792,N_13122,N_10615);
nand U16793 (N_16793,N_12957,N_11715);
or U16794 (N_16794,N_12327,N_13962);
and U16795 (N_16795,N_13423,N_14866);
nand U16796 (N_16796,N_14631,N_10913);
or U16797 (N_16797,N_14529,N_11729);
or U16798 (N_16798,N_11980,N_14922);
nor U16799 (N_16799,N_12659,N_13708);
and U16800 (N_16800,N_13592,N_14411);
nand U16801 (N_16801,N_12365,N_11177);
and U16802 (N_16802,N_14351,N_10518);
nor U16803 (N_16803,N_12542,N_11522);
nand U16804 (N_16804,N_10189,N_11547);
nor U16805 (N_16805,N_10460,N_12196);
xnor U16806 (N_16806,N_12076,N_12770);
and U16807 (N_16807,N_14954,N_13569);
nand U16808 (N_16808,N_11422,N_10699);
or U16809 (N_16809,N_14530,N_10645);
nor U16810 (N_16810,N_12323,N_13402);
nor U16811 (N_16811,N_12004,N_14358);
or U16812 (N_16812,N_12457,N_13862);
nand U16813 (N_16813,N_13325,N_14855);
nor U16814 (N_16814,N_10083,N_13619);
nor U16815 (N_16815,N_12063,N_14438);
nand U16816 (N_16816,N_11095,N_14324);
or U16817 (N_16817,N_12477,N_10805);
nand U16818 (N_16818,N_14479,N_14699);
and U16819 (N_16819,N_12704,N_14211);
nor U16820 (N_16820,N_12481,N_12823);
nor U16821 (N_16821,N_11741,N_12658);
nor U16822 (N_16822,N_13991,N_13793);
or U16823 (N_16823,N_13575,N_10436);
and U16824 (N_16824,N_14823,N_12531);
and U16825 (N_16825,N_14237,N_13888);
and U16826 (N_16826,N_10122,N_13056);
nand U16827 (N_16827,N_12581,N_10659);
nand U16828 (N_16828,N_10850,N_11307);
and U16829 (N_16829,N_13674,N_12660);
nor U16830 (N_16830,N_12825,N_12569);
or U16831 (N_16831,N_14244,N_14968);
xnor U16832 (N_16832,N_10859,N_14526);
or U16833 (N_16833,N_10695,N_11706);
xor U16834 (N_16834,N_11904,N_12914);
and U16835 (N_16835,N_11665,N_14665);
xnor U16836 (N_16836,N_11811,N_11847);
nand U16837 (N_16837,N_14044,N_12566);
nor U16838 (N_16838,N_10967,N_12447);
or U16839 (N_16839,N_11046,N_12130);
nand U16840 (N_16840,N_12329,N_14611);
or U16841 (N_16841,N_10132,N_11012);
nor U16842 (N_16842,N_12947,N_12374);
xnor U16843 (N_16843,N_14898,N_14075);
and U16844 (N_16844,N_10935,N_14288);
and U16845 (N_16845,N_13075,N_12038);
nor U16846 (N_16846,N_13370,N_12184);
or U16847 (N_16847,N_12707,N_13966);
or U16848 (N_16848,N_11017,N_10700);
nor U16849 (N_16849,N_10841,N_10248);
and U16850 (N_16850,N_12503,N_12848);
xor U16851 (N_16851,N_14306,N_14513);
nor U16852 (N_16852,N_10078,N_14087);
nor U16853 (N_16853,N_14615,N_13624);
or U16854 (N_16854,N_13765,N_10954);
nor U16855 (N_16855,N_10662,N_13621);
nand U16856 (N_16856,N_10200,N_11265);
nor U16857 (N_16857,N_14519,N_10955);
and U16858 (N_16858,N_11157,N_10941);
nor U16859 (N_16859,N_12513,N_11854);
or U16860 (N_16860,N_13999,N_12275);
nand U16861 (N_16861,N_14400,N_13133);
and U16862 (N_16862,N_13406,N_10756);
nor U16863 (N_16863,N_11654,N_10241);
and U16864 (N_16864,N_14982,N_10810);
nor U16865 (N_16865,N_11550,N_14084);
or U16866 (N_16866,N_11571,N_11521);
and U16867 (N_16867,N_12951,N_11314);
and U16868 (N_16868,N_13598,N_14150);
xnor U16869 (N_16869,N_11086,N_14110);
or U16870 (N_16870,N_13403,N_11917);
nand U16871 (N_16871,N_13750,N_11030);
nand U16872 (N_16872,N_14985,N_14202);
or U16873 (N_16873,N_12041,N_11899);
and U16874 (N_16874,N_10453,N_11743);
nor U16875 (N_16875,N_12744,N_10428);
and U16876 (N_16876,N_12794,N_11789);
or U16877 (N_16877,N_11069,N_13006);
nand U16878 (N_16878,N_14145,N_11419);
nor U16879 (N_16879,N_10963,N_11862);
and U16880 (N_16880,N_10663,N_14135);
nand U16881 (N_16881,N_11842,N_12295);
nor U16882 (N_16882,N_11209,N_13845);
or U16883 (N_16883,N_13208,N_12805);
or U16884 (N_16884,N_11011,N_14671);
nor U16885 (N_16885,N_12216,N_14238);
xnor U16886 (N_16886,N_12881,N_12498);
and U16887 (N_16887,N_12906,N_10671);
and U16888 (N_16888,N_13313,N_14172);
nand U16889 (N_16889,N_10532,N_11554);
nor U16890 (N_16890,N_12670,N_11779);
or U16891 (N_16891,N_10175,N_14390);
and U16892 (N_16892,N_13148,N_10098);
nand U16893 (N_16893,N_11210,N_12552);
nor U16894 (N_16894,N_14313,N_13584);
and U16895 (N_16895,N_10951,N_13305);
xnor U16896 (N_16896,N_13940,N_10364);
nand U16897 (N_16897,N_14349,N_14921);
nor U16898 (N_16898,N_12942,N_12993);
and U16899 (N_16899,N_12284,N_12903);
or U16900 (N_16900,N_10624,N_14773);
nor U16901 (N_16901,N_11325,N_13190);
and U16902 (N_16902,N_11637,N_11156);
or U16903 (N_16903,N_10836,N_13838);
nor U16904 (N_16904,N_12682,N_13599);
nor U16905 (N_16905,N_14725,N_10994);
nand U16906 (N_16906,N_12886,N_11734);
or U16907 (N_16907,N_13895,N_12748);
or U16908 (N_16908,N_11402,N_11578);
nand U16909 (N_16909,N_11411,N_11053);
nor U16910 (N_16910,N_13336,N_11788);
nor U16911 (N_16911,N_11469,N_12404);
and U16912 (N_16912,N_14174,N_11274);
and U16913 (N_16913,N_14880,N_10870);
and U16914 (N_16914,N_12575,N_10708);
and U16915 (N_16915,N_11838,N_14577);
nor U16916 (N_16916,N_14667,N_14859);
nor U16917 (N_16917,N_10973,N_12818);
or U16918 (N_16918,N_14473,N_12590);
or U16919 (N_16919,N_11074,N_13904);
or U16920 (N_16920,N_11470,N_14167);
or U16921 (N_16921,N_14540,N_13169);
nand U16922 (N_16922,N_14180,N_11808);
nor U16923 (N_16923,N_14089,N_12596);
nand U16924 (N_16924,N_12367,N_14334);
or U16925 (N_16925,N_10579,N_14112);
and U16926 (N_16926,N_10255,N_14223);
and U16927 (N_16927,N_11850,N_11906);
xnor U16928 (N_16928,N_14331,N_12505);
and U16929 (N_16929,N_12211,N_13052);
nand U16930 (N_16930,N_10071,N_10686);
nor U16931 (N_16931,N_11088,N_12001);
or U16932 (N_16932,N_13625,N_12723);
or U16933 (N_16933,N_11055,N_10108);
or U16934 (N_16934,N_11353,N_12603);
and U16935 (N_16935,N_14061,N_11590);
xor U16936 (N_16936,N_12050,N_11169);
nand U16937 (N_16937,N_10222,N_11682);
nand U16938 (N_16938,N_14944,N_11085);
and U16939 (N_16939,N_10382,N_12182);
nand U16940 (N_16940,N_10265,N_11310);
nand U16941 (N_16941,N_12455,N_13504);
nor U16942 (N_16942,N_12991,N_12904);
nor U16943 (N_16943,N_10295,N_10696);
and U16944 (N_16944,N_10758,N_12179);
or U16945 (N_16945,N_11443,N_10989);
and U16946 (N_16946,N_12016,N_14947);
and U16947 (N_16947,N_13663,N_13458);
or U16948 (N_16948,N_11452,N_14714);
or U16949 (N_16949,N_13978,N_13248);
and U16950 (N_16950,N_11557,N_12431);
or U16951 (N_16951,N_12000,N_14189);
or U16952 (N_16952,N_12460,N_10464);
and U16953 (N_16953,N_10276,N_14077);
and U16954 (N_16954,N_14283,N_12150);
nor U16955 (N_16955,N_11969,N_13677);
and U16956 (N_16956,N_11034,N_12666);
nor U16957 (N_16957,N_14123,N_14557);
xnor U16958 (N_16958,N_14441,N_12685);
nor U16959 (N_16959,N_14892,N_10589);
and U16960 (N_16960,N_10015,N_14900);
and U16961 (N_16961,N_11188,N_11562);
nand U16962 (N_16962,N_10772,N_11135);
and U16963 (N_16963,N_10441,N_10280);
nand U16964 (N_16964,N_13929,N_10490);
and U16965 (N_16965,N_13549,N_10527);
or U16966 (N_16966,N_12023,N_10000);
and U16967 (N_16967,N_14715,N_10534);
nor U16968 (N_16968,N_14685,N_13554);
or U16969 (N_16969,N_13520,N_12321);
and U16970 (N_16970,N_10591,N_11566);
and U16971 (N_16971,N_14750,N_10512);
xor U16972 (N_16972,N_11929,N_14870);
and U16973 (N_16973,N_11294,N_13443);
and U16974 (N_16974,N_11699,N_10269);
and U16975 (N_16975,N_10454,N_12248);
nor U16976 (N_16976,N_10187,N_14156);
or U16977 (N_16977,N_11973,N_12302);
nand U16978 (N_16978,N_12173,N_13846);
nand U16979 (N_16979,N_13866,N_11344);
and U16980 (N_16980,N_10308,N_12710);
nand U16981 (N_16981,N_12044,N_10041);
and U16982 (N_16982,N_11523,N_13971);
and U16983 (N_16983,N_14501,N_14796);
nor U16984 (N_16984,N_12470,N_13490);
xor U16985 (N_16985,N_12664,N_12847);
xor U16986 (N_16986,N_13094,N_12231);
or U16987 (N_16987,N_11791,N_10735);
xor U16988 (N_16988,N_13562,N_10956);
and U16989 (N_16989,N_10168,N_11259);
and U16990 (N_16990,N_11207,N_13288);
and U16991 (N_16991,N_13583,N_14780);
xor U16992 (N_16992,N_11845,N_10667);
and U16993 (N_16993,N_13058,N_10363);
xor U16994 (N_16994,N_11889,N_11841);
and U16995 (N_16995,N_12979,N_10655);
and U16996 (N_16996,N_10934,N_12176);
nor U16997 (N_16997,N_11800,N_13889);
nand U16998 (N_16998,N_13107,N_11341);
or U16999 (N_16999,N_10997,N_12832);
nor U17000 (N_17000,N_10037,N_12985);
xnor U17001 (N_17001,N_13092,N_13703);
xnor U17002 (N_17002,N_13233,N_14285);
xnor U17003 (N_17003,N_13847,N_13800);
and U17004 (N_17004,N_13875,N_13566);
nor U17005 (N_17005,N_10345,N_14444);
or U17006 (N_17006,N_14554,N_10220);
nand U17007 (N_17007,N_13111,N_10937);
nor U17008 (N_17008,N_11330,N_11533);
nand U17009 (N_17009,N_10528,N_12486);
nand U17010 (N_17010,N_12484,N_13465);
nand U17011 (N_17011,N_10494,N_13691);
xor U17012 (N_17012,N_14847,N_11548);
or U17013 (N_17013,N_12876,N_14484);
nand U17014 (N_17014,N_11244,N_10791);
or U17015 (N_17015,N_11054,N_12253);
nand U17016 (N_17016,N_13590,N_11941);
nor U17017 (N_17017,N_12691,N_11059);
nor U17018 (N_17018,N_12688,N_14788);
and U17019 (N_17019,N_11831,N_12017);
or U17020 (N_17020,N_14845,N_10089);
nand U17021 (N_17021,N_14229,N_11934);
nor U17022 (N_17022,N_14451,N_14419);
xor U17023 (N_17023,N_10822,N_13409);
or U17024 (N_17024,N_10681,N_12344);
xnor U17025 (N_17025,N_13454,N_10884);
and U17026 (N_17026,N_14574,N_12280);
xnor U17027 (N_17027,N_11890,N_10486);
nand U17028 (N_17028,N_11118,N_11810);
nand U17029 (N_17029,N_10158,N_11933);
nand U17030 (N_17030,N_13289,N_13486);
nand U17031 (N_17031,N_11045,N_13271);
or U17032 (N_17032,N_12099,N_11304);
nor U17033 (N_17033,N_13860,N_13690);
and U17034 (N_17034,N_13088,N_10244);
or U17035 (N_17035,N_14759,N_12509);
and U17036 (N_17036,N_10599,N_14221);
nand U17037 (N_17037,N_12950,N_10611);
nor U17038 (N_17038,N_14001,N_14100);
nor U17039 (N_17039,N_11762,N_12426);
or U17040 (N_17040,N_11979,N_10825);
nand U17041 (N_17041,N_10145,N_12339);
and U17042 (N_17042,N_11154,N_10404);
and U17043 (N_17043,N_13425,N_14355);
nor U17044 (N_17044,N_12298,N_12375);
nor U17045 (N_17045,N_12919,N_11992);
or U17046 (N_17046,N_11196,N_14378);
nand U17047 (N_17047,N_10386,N_12850);
nand U17048 (N_17048,N_12363,N_10146);
nor U17049 (N_17049,N_11761,N_14698);
nor U17050 (N_17050,N_11770,N_10743);
or U17051 (N_17051,N_12273,N_14009);
nand U17052 (N_17052,N_14316,N_11951);
and U17053 (N_17053,N_12982,N_13588);
nor U17054 (N_17054,N_13905,N_14258);
and U17055 (N_17055,N_14192,N_12772);
and U17056 (N_17056,N_11537,N_14126);
nor U17057 (N_17057,N_11315,N_14544);
nor U17058 (N_17058,N_14974,N_14254);
nor U17059 (N_17059,N_11297,N_11179);
xnor U17060 (N_17060,N_11357,N_14777);
nor U17061 (N_17061,N_10910,N_11995);
nand U17062 (N_17062,N_14582,N_12514);
nand U17063 (N_17063,N_11943,N_10982);
and U17064 (N_17064,N_12580,N_14906);
and U17065 (N_17065,N_10781,N_10543);
nor U17066 (N_17066,N_12863,N_12802);
or U17067 (N_17067,N_11114,N_11616);
and U17068 (N_17068,N_12385,N_11023);
nor U17069 (N_17069,N_13996,N_14525);
xnor U17070 (N_17070,N_13681,N_14281);
nor U17071 (N_17071,N_13789,N_13324);
and U17072 (N_17072,N_12012,N_13593);
nor U17073 (N_17073,N_11617,N_12429);
xnor U17074 (N_17074,N_11217,N_10151);
nand U17075 (N_17075,N_12289,N_10990);
and U17076 (N_17076,N_11722,N_11961);
nand U17077 (N_17077,N_14293,N_10549);
xor U17078 (N_17078,N_11744,N_14134);
nor U17079 (N_17079,N_13586,N_12408);
or U17080 (N_17080,N_11611,N_10762);
xnor U17081 (N_17081,N_11269,N_12458);
or U17082 (N_17082,N_11988,N_11507);
or U17083 (N_17083,N_11298,N_13134);
nand U17084 (N_17084,N_13291,N_11962);
nand U17085 (N_17085,N_14469,N_12546);
xor U17086 (N_17086,N_14212,N_10513);
or U17087 (N_17087,N_12611,N_13511);
xnor U17088 (N_17088,N_13020,N_11388);
nor U17089 (N_17089,N_14666,N_11466);
and U17090 (N_17090,N_12994,N_13541);
nor U17091 (N_17091,N_13640,N_13848);
nor U17092 (N_17092,N_10400,N_11272);
and U17093 (N_17093,N_12778,N_13696);
and U17094 (N_17094,N_10745,N_12106);
nor U17095 (N_17095,N_13643,N_12911);
and U17096 (N_17096,N_11924,N_11813);
nand U17097 (N_17097,N_14291,N_11242);
or U17098 (N_17098,N_14936,N_11193);
and U17099 (N_17099,N_10111,N_13867);
or U17100 (N_17100,N_14981,N_12467);
or U17101 (N_17101,N_14976,N_10914);
nand U17102 (N_17102,N_12442,N_12198);
xnor U17103 (N_17103,N_14938,N_13763);
xnor U17104 (N_17104,N_11436,N_13828);
nor U17105 (N_17105,N_13496,N_12619);
or U17106 (N_17106,N_11748,N_12462);
nand U17107 (N_17107,N_12793,N_14217);
and U17108 (N_17108,N_12774,N_11945);
and U17109 (N_17109,N_14121,N_11025);
and U17110 (N_17110,N_14070,N_11376);
or U17111 (N_17111,N_12037,N_14775);
or U17112 (N_17112,N_10774,N_10082);
or U17113 (N_17113,N_14772,N_13835);
or U17114 (N_17114,N_10336,N_10173);
or U17115 (N_17115,N_10775,N_12678);
nand U17116 (N_17116,N_10790,N_13206);
or U17117 (N_17117,N_10004,N_13171);
nor U17118 (N_17118,N_11958,N_11024);
nand U17119 (N_17119,N_12096,N_13509);
and U17120 (N_17120,N_10302,N_11801);
nor U17121 (N_17121,N_14833,N_13941);
or U17122 (N_17122,N_10243,N_11512);
and U17123 (N_17123,N_12869,N_14515);
xor U17124 (N_17124,N_12291,N_10767);
or U17125 (N_17125,N_14521,N_12146);
nor U17126 (N_17126,N_10648,N_10212);
nand U17127 (N_17127,N_13726,N_10215);
nor U17128 (N_17128,N_10375,N_11455);
or U17129 (N_17129,N_10932,N_13739);
and U17130 (N_17130,N_10005,N_14165);
or U17131 (N_17131,N_10502,N_13730);
or U17132 (N_17132,N_12764,N_11885);
nor U17133 (N_17133,N_14888,N_13858);
xor U17134 (N_17134,N_10052,N_12465);
xnor U17135 (N_17135,N_10313,N_11350);
and U17136 (N_17136,N_14369,N_14003);
and U17137 (N_17137,N_11585,N_12144);
and U17138 (N_17138,N_10246,N_13427);
nand U17139 (N_17139,N_11815,N_14447);
xnor U17140 (N_17140,N_14475,N_11803);
and U17141 (N_17141,N_10447,N_11898);
and U17142 (N_17142,N_10385,N_13497);
and U17143 (N_17143,N_12535,N_12031);
nand U17144 (N_17144,N_13469,N_13265);
nor U17145 (N_17145,N_13032,N_11120);
nand U17146 (N_17146,N_11401,N_13196);
nor U17147 (N_17147,N_14220,N_13907);
and U17148 (N_17148,N_13558,N_13879);
nand U17149 (N_17149,N_12725,N_11506);
nor U17150 (N_17150,N_12730,N_14032);
and U17151 (N_17151,N_12306,N_10498);
and U17152 (N_17152,N_13699,N_11581);
nor U17153 (N_17153,N_13898,N_14465);
nand U17154 (N_17154,N_13646,N_13890);
nand U17155 (N_17155,N_10423,N_12674);
nor U17156 (N_17156,N_13035,N_10480);
and U17157 (N_17157,N_14721,N_11971);
and U17158 (N_17158,N_12973,N_12587);
xnor U17159 (N_17159,N_12564,N_14532);
or U17160 (N_17160,N_13126,N_13878);
and U17161 (N_17161,N_11090,N_14941);
or U17162 (N_17162,N_11567,N_11251);
xnor U17163 (N_17163,N_14640,N_13958);
or U17164 (N_17164,N_10827,N_14433);
nand U17165 (N_17165,N_10739,N_13856);
or U17166 (N_17166,N_14122,N_13495);
nor U17167 (N_17167,N_10759,N_10120);
nor U17168 (N_17168,N_13706,N_10049);
nand U17169 (N_17169,N_12018,N_13533);
and U17170 (N_17170,N_10919,N_10068);
nand U17171 (N_17171,N_11296,N_10140);
nor U17172 (N_17172,N_13241,N_10023);
or U17173 (N_17173,N_13684,N_12830);
and U17174 (N_17174,N_11778,N_13116);
or U17175 (N_17175,N_14994,N_11776);
and U17176 (N_17176,N_12154,N_14999);
nor U17177 (N_17177,N_14385,N_10179);
nor U17178 (N_17178,N_14804,N_10799);
nand U17179 (N_17179,N_12773,N_12136);
nand U17180 (N_17180,N_10575,N_11288);
xnor U17181 (N_17181,N_10576,N_12449);
nor U17182 (N_17182,N_13327,N_10856);
and U17183 (N_17183,N_14005,N_11146);
or U17184 (N_17184,N_13066,N_11458);
nand U17185 (N_17185,N_13238,N_12565);
or U17186 (N_17186,N_11247,N_12324);
nand U17187 (N_17187,N_10677,N_11363);
nor U17188 (N_17188,N_12229,N_13628);
xor U17189 (N_17189,N_14248,N_10730);
or U17190 (N_17190,N_13053,N_13280);
nor U17191 (N_17191,N_12795,N_14023);
or U17192 (N_17192,N_11568,N_10406);
nor U17193 (N_17193,N_11758,N_14104);
or U17194 (N_17194,N_12228,N_14660);
xnor U17195 (N_17195,N_12368,N_13419);
nand U17196 (N_17196,N_12111,N_14287);
nor U17197 (N_17197,N_12952,N_11170);
nor U17198 (N_17198,N_14511,N_13917);
or U17199 (N_17199,N_12060,N_11576);
and U17200 (N_17200,N_10393,N_13522);
nand U17201 (N_17201,N_13417,N_10703);
xor U17202 (N_17202,N_13738,N_11658);
and U17203 (N_17203,N_12974,N_10909);
nor U17204 (N_17204,N_11382,N_11878);
or U17205 (N_17205,N_12256,N_12585);
or U17206 (N_17206,N_14913,N_10693);
nor U17207 (N_17207,N_10828,N_10247);
and U17208 (N_17208,N_10712,N_12898);
or U17209 (N_17209,N_11598,N_14690);
xor U17210 (N_17210,N_12080,N_11814);
nor U17211 (N_17211,N_10216,N_14364);
xor U17212 (N_17212,N_13880,N_11596);
nand U17213 (N_17213,N_11852,N_11662);
nand U17214 (N_17214,N_11543,N_11632);
and U17215 (N_17215,N_10834,N_12627);
and U17216 (N_17216,N_14867,N_11859);
and U17217 (N_17217,N_10927,N_11145);
or U17218 (N_17218,N_14642,N_11087);
or U17219 (N_17219,N_14812,N_11107);
xnor U17220 (N_17220,N_12680,N_13382);
nor U17221 (N_17221,N_14038,N_11240);
xnor U17222 (N_17222,N_13612,N_12153);
nand U17223 (N_17223,N_14058,N_11104);
nand U17224 (N_17224,N_13984,N_12809);
nor U17225 (N_17225,N_14549,N_12167);
nand U17226 (N_17226,N_14152,N_11619);
nand U17227 (N_17227,N_14856,N_12526);
nor U17228 (N_17228,N_11584,N_14113);
and U17229 (N_17229,N_14903,N_11468);
nor U17230 (N_17230,N_11975,N_14225);
and U17231 (N_17231,N_10414,N_13387);
xor U17232 (N_17232,N_11456,N_12775);
nor U17233 (N_17233,N_14863,N_13154);
nand U17234 (N_17234,N_12454,N_13909);
and U17235 (N_17235,N_13461,N_10330);
or U17236 (N_17236,N_14250,N_10309);
nand U17237 (N_17237,N_11944,N_14487);
xnor U17238 (N_17238,N_12328,N_12829);
nor U17239 (N_17239,N_11268,N_12810);
or U17240 (N_17240,N_11918,N_11649);
nor U17241 (N_17241,N_11162,N_10855);
nand U17242 (N_17242,N_13712,N_10630);
nand U17243 (N_17243,N_10293,N_13456);
or U17244 (N_17244,N_10080,N_11281);
xor U17245 (N_17245,N_14195,N_14074);
nor U17246 (N_17246,N_13873,N_13749);
and U17247 (N_17247,N_11215,N_10523);
or U17248 (N_17248,N_10129,N_10538);
xor U17249 (N_17249,N_14688,N_12494);
nand U17250 (N_17250,N_14130,N_10463);
nand U17251 (N_17251,N_10698,N_10873);
or U17252 (N_17252,N_11927,N_13921);
and U17253 (N_17253,N_14915,N_14860);
or U17254 (N_17254,N_11785,N_14919);
xnor U17255 (N_17255,N_11608,N_10034);
and U17256 (N_17256,N_14830,N_13085);
xor U17257 (N_17257,N_14219,N_10564);
and U17258 (N_17258,N_14054,N_13521);
nand U17259 (N_17259,N_11142,N_13960);
nand U17260 (N_17260,N_13759,N_12527);
or U17261 (N_17261,N_12359,N_13925);
or U17262 (N_17262,N_14173,N_13729);
nand U17263 (N_17263,N_11694,N_13457);
nand U17264 (N_17264,N_13093,N_13254);
nand U17265 (N_17265,N_13891,N_13356);
and U17266 (N_17266,N_14740,N_13967);
nand U17267 (N_17267,N_10771,N_10320);
or U17268 (N_17268,N_13956,N_13031);
nor U17269 (N_17269,N_12461,N_11409);
or U17270 (N_17270,N_13350,N_14629);
nor U17271 (N_17271,N_12353,N_10286);
and U17272 (N_17272,N_11208,N_14569);
xor U17273 (N_17273,N_14960,N_11113);
xnor U17274 (N_17274,N_10690,N_14214);
or U17275 (N_17275,N_11509,N_14474);
or U17276 (N_17276,N_10100,N_14547);
nor U17277 (N_17277,N_12170,N_12394);
nor U17278 (N_17278,N_14488,N_14978);
nor U17279 (N_17279,N_14416,N_12715);
xor U17280 (N_17280,N_14594,N_11033);
and U17281 (N_17281,N_10278,N_13707);
and U17282 (N_17282,N_12351,N_10487);
nor U17283 (N_17283,N_10218,N_13380);
nand U17284 (N_17284,N_14183,N_10936);
and U17285 (N_17285,N_12922,N_12492);
nor U17286 (N_17286,N_14338,N_13101);
and U17287 (N_17287,N_12833,N_14106);
nor U17288 (N_17288,N_11161,N_14989);
and U17289 (N_17289,N_13394,N_11874);
nor U17290 (N_17290,N_10387,N_12046);
and U17291 (N_17291,N_14619,N_11702);
and U17292 (N_17292,N_14185,N_12586);
and U17293 (N_17293,N_13204,N_12913);
and U17294 (N_17294,N_12883,N_11302);
or U17295 (N_17295,N_10497,N_11225);
or U17296 (N_17296,N_11766,N_11545);
nand U17297 (N_17297,N_14561,N_11200);
nor U17298 (N_17298,N_13437,N_14376);
xor U17299 (N_17299,N_12020,N_10815);
nand U17300 (N_17300,N_14132,N_11672);
nor U17301 (N_17301,N_12752,N_14420);
nand U17302 (N_17302,N_12360,N_13827);
nor U17303 (N_17303,N_13142,N_14735);
xor U17304 (N_17304,N_14155,N_10070);
or U17305 (N_17305,N_13081,N_10446);
or U17306 (N_17306,N_14828,N_13950);
nand U17307 (N_17307,N_10086,N_11956);
xor U17308 (N_17308,N_12218,N_14424);
xor U17309 (N_17309,N_13767,N_13418);
or U17310 (N_17310,N_13986,N_14090);
nor U17311 (N_17311,N_11073,N_10530);
or U17312 (N_17312,N_13026,N_12357);
nor U17313 (N_17313,N_14693,N_13589);
nor U17314 (N_17314,N_13159,N_13637);
and U17315 (N_17315,N_10030,N_13814);
nand U17316 (N_17316,N_11780,N_10526);
nor U17317 (N_17317,N_14093,N_13574);
nor U17318 (N_17318,N_12270,N_14417);
or U17319 (N_17319,N_14935,N_10258);
nor U17320 (N_17320,N_12827,N_14840);
nor U17321 (N_17321,N_14774,N_14307);
or U17322 (N_17322,N_14446,N_14895);
nor U17323 (N_17323,N_13935,N_12210);
nand U17324 (N_17324,N_11093,N_14973);
nand U17325 (N_17325,N_14246,N_12151);
nand U17326 (N_17326,N_10500,N_10657);
xnor U17327 (N_17327,N_14379,N_14062);
and U17328 (N_17328,N_12646,N_10262);
nor U17329 (N_17329,N_12842,N_13829);
nand U17330 (N_17330,N_12650,N_13506);
and U17331 (N_17331,N_12961,N_10991);
nand U17332 (N_17332,N_14269,N_10625);
and U17333 (N_17333,N_12889,N_11640);
nand U17334 (N_17334,N_13985,N_12909);
nand U17335 (N_17335,N_11039,N_13177);
nand U17336 (N_17336,N_13770,N_11228);
nand U17337 (N_17337,N_13262,N_12490);
xnor U17338 (N_17338,N_14718,N_13517);
nor U17339 (N_17339,N_13664,N_10793);
nor U17340 (N_17340,N_13605,N_14624);
nand U17341 (N_17341,N_12435,N_11978);
and U17342 (N_17342,N_14984,N_10250);
or U17343 (N_17343,N_13951,N_11905);
nor U17344 (N_17344,N_12894,N_13200);
nor U17345 (N_17345,N_14942,N_10911);
or U17346 (N_17346,N_12309,N_14308);
nand U17347 (N_17347,N_13542,N_12855);
or U17348 (N_17348,N_14216,N_13083);
nor U17349 (N_17349,N_12034,N_11013);
or U17350 (N_17350,N_14535,N_12851);
and U17351 (N_17351,N_11029,N_11656);
nand U17352 (N_17352,N_11463,N_13221);
xnor U17353 (N_17353,N_13620,N_10115);
nand U17354 (N_17354,N_10925,N_13678);
nor U17355 (N_17355,N_11763,N_11122);
or U17356 (N_17356,N_10988,N_12789);
or U17357 (N_17357,N_12672,N_11959);
and U17358 (N_17358,N_11716,N_14591);
and U17359 (N_17359,N_13776,N_10090);
nor U17360 (N_17360,N_14763,N_13010);
nor U17361 (N_17361,N_11586,N_11499);
nand U17362 (N_17362,N_10418,N_14196);
xor U17363 (N_17363,N_13211,N_11386);
nand U17364 (N_17364,N_11101,N_13434);
or U17365 (N_17365,N_12469,N_11431);
or U17366 (N_17366,N_13432,N_13129);
nor U17367 (N_17367,N_12418,N_12705);
xor U17368 (N_17368,N_11518,N_11262);
or U17369 (N_17369,N_12325,N_11895);
xor U17370 (N_17370,N_13119,N_13998);
and U17371 (N_17371,N_12347,N_10596);
nand U17372 (N_17372,N_12381,N_12201);
or U17373 (N_17373,N_10580,N_11727);
or U17374 (N_17374,N_14455,N_14323);
or U17375 (N_17375,N_13942,N_14945);
and U17376 (N_17376,N_11435,N_13257);
or U17377 (N_17377,N_14592,N_12504);
xnor U17378 (N_17378,N_13551,N_11264);
or U17379 (N_17379,N_13420,N_11565);
nand U17380 (N_17380,N_10019,N_10848);
xor U17381 (N_17381,N_10206,N_14011);
or U17382 (N_17382,N_14728,N_10719);
nor U17383 (N_17383,N_11997,N_11185);
or U17384 (N_17384,N_14300,N_13367);
and U17385 (N_17385,N_13754,N_13650);
and U17386 (N_17386,N_13187,N_13477);
or U17387 (N_17387,N_14476,N_13397);
or U17388 (N_17388,N_11526,N_14045);
nand U17389 (N_17389,N_12972,N_11057);
nand U17390 (N_17390,N_14852,N_12190);
nand U17391 (N_17391,N_12002,N_13705);
nand U17392 (N_17392,N_12103,N_14347);
nor U17393 (N_17393,N_13532,N_12373);
or U17394 (N_17394,N_10332,N_13555);
nand U17395 (N_17395,N_14468,N_11792);
nand U17396 (N_17396,N_14410,N_13639);
and U17397 (N_17397,N_14884,N_11460);
or U17398 (N_17398,N_13874,N_12692);
and U17399 (N_17399,N_13145,N_14653);
and U17400 (N_17400,N_14181,N_11986);
and U17401 (N_17401,N_12946,N_10057);
nor U17402 (N_17402,N_13963,N_10641);
and U17403 (N_17403,N_12437,N_13630);
nor U17404 (N_17404,N_12100,N_14068);
and U17405 (N_17405,N_14868,N_10593);
nor U17406 (N_17406,N_14972,N_13181);
or U17407 (N_17407,N_10687,N_12129);
or U17408 (N_17408,N_13197,N_12665);
nand U17409 (N_17409,N_11739,N_14587);
nand U17410 (N_17410,N_13494,N_14647);
and U17411 (N_17411,N_12929,N_13761);
nand U17412 (N_17412,N_11172,N_12578);
nor U17413 (N_17413,N_14079,N_13801);
and U17414 (N_17414,N_10053,N_11239);
and U17415 (N_17415,N_11322,N_10798);
xnor U17416 (N_17416,N_11569,N_12073);
nand U17417 (N_17417,N_14257,N_13314);
nor U17418 (N_17418,N_14381,N_13919);
and U17419 (N_17419,N_12319,N_14041);
nor U17420 (N_17420,N_10118,N_10373);
or U17421 (N_17421,N_11324,N_13412);
nand U17422 (N_17422,N_12059,N_14701);
nand U17423 (N_17423,N_14048,N_12126);
nor U17424 (N_17424,N_12053,N_14471);
nand U17425 (N_17425,N_14762,N_10491);
nand U17426 (N_17426,N_10711,N_14332);
nor U17427 (N_17427,N_11291,N_10150);
or U17428 (N_17428,N_10788,N_14091);
nand U17429 (N_17429,N_10073,N_13127);
and U17430 (N_17430,N_11664,N_13445);
and U17431 (N_17431,N_12591,N_10495);
nor U17432 (N_17432,N_10753,N_11690);
and U17433 (N_17433,N_14201,N_13428);
nor U17434 (N_17434,N_12120,N_14632);
or U17435 (N_17435,N_14493,N_10757);
or U17436 (N_17436,N_10637,N_13915);
or U17437 (N_17437,N_13537,N_10521);
nor U17438 (N_17438,N_10612,N_13245);
and U17439 (N_17439,N_10683,N_11360);
nor U17440 (N_17440,N_12047,N_14831);
xor U17441 (N_17441,N_12987,N_13535);
nor U17442 (N_17442,N_12258,N_13287);
and U17443 (N_17443,N_14555,N_14284);
nand U17444 (N_17444,N_12472,N_12383);
and U17445 (N_17445,N_10461,N_10729);
nor U17446 (N_17446,N_12204,N_12989);
or U17447 (N_17447,N_12227,N_12219);
nand U17448 (N_17448,N_10912,N_12632);
xor U17449 (N_17449,N_11257,N_10784);
nor U17450 (N_17450,N_13927,N_14578);
nand U17451 (N_17451,N_13439,N_10475);
and U17452 (N_17452,N_11790,N_10581);
or U17453 (N_17453,N_12801,N_11394);
and U17454 (N_17454,N_10462,N_11802);
nand U17455 (N_17455,N_11412,N_10949);
or U17456 (N_17456,N_12971,N_14684);
and U17457 (N_17457,N_12814,N_10106);
or U17458 (N_17458,N_12912,N_14912);
and U17459 (N_17459,N_13137,N_11103);
or U17460 (N_17460,N_12956,N_10710);
and U17461 (N_17461,N_10524,N_10442);
and U17462 (N_17462,N_13849,N_11214);
and U17463 (N_17463,N_14234,N_12068);
nor U17464 (N_17464,N_10130,N_11343);
nor U17465 (N_17465,N_13642,N_10063);
or U17466 (N_17466,N_14916,N_14873);
and U17467 (N_17467,N_10860,N_11667);
and U17468 (N_17468,N_12413,N_14964);
nand U17469 (N_17469,N_14412,N_11799);
nor U17470 (N_17470,N_12186,N_11317);
or U17471 (N_17471,N_13303,N_14261);
or U17472 (N_17472,N_13675,N_10606);
nand U17473 (N_17473,N_14463,N_10306);
and U17474 (N_17474,N_14360,N_10121);
and U17475 (N_17475,N_11530,N_11312);
nor U17476 (N_17476,N_11579,N_11440);
nor U17477 (N_17477,N_11668,N_14231);
nand U17478 (N_17478,N_13392,N_12497);
nor U17479 (N_17479,N_11650,N_10620);
or U17480 (N_17480,N_11549,N_12523);
nand U17481 (N_17481,N_10961,N_14318);
or U17482 (N_17482,N_14885,N_10898);
and U17483 (N_17483,N_13120,N_12640);
nor U17484 (N_17484,N_12560,N_10046);
nand U17485 (N_17485,N_13256,N_12857);
nand U17486 (N_17486,N_11082,N_13176);
or U17487 (N_17487,N_11476,N_14492);
xor U17488 (N_17488,N_11805,N_13721);
and U17489 (N_17489,N_13689,N_10213);
or U17490 (N_17490,N_12541,N_12577);
or U17491 (N_17491,N_10717,N_10422);
and U17492 (N_17492,N_10231,N_12655);
or U17493 (N_17493,N_13839,N_12371);
or U17494 (N_17494,N_13855,N_14654);
or U17495 (N_17495,N_14301,N_13071);
nand U17496 (N_17496,N_10377,N_14905);
and U17497 (N_17497,N_13189,N_12487);
nor U17498 (N_17498,N_10921,N_13225);
nand U17499 (N_17499,N_13164,N_14190);
or U17500 (N_17500,N_10996,N_12133);
xnor U17501 (N_17501,N_10169,N_11946);
nand U17502 (N_17502,N_13822,N_12129);
nand U17503 (N_17503,N_14852,N_11664);
nor U17504 (N_17504,N_10869,N_11997);
nand U17505 (N_17505,N_13445,N_12602);
nand U17506 (N_17506,N_12177,N_13789);
and U17507 (N_17507,N_13015,N_11980);
and U17508 (N_17508,N_10375,N_10762);
and U17509 (N_17509,N_12506,N_12222);
nand U17510 (N_17510,N_14581,N_11468);
xor U17511 (N_17511,N_12091,N_13666);
and U17512 (N_17512,N_13774,N_13826);
nor U17513 (N_17513,N_10822,N_13030);
xnor U17514 (N_17514,N_12520,N_10082);
or U17515 (N_17515,N_14302,N_13319);
and U17516 (N_17516,N_13646,N_13231);
and U17517 (N_17517,N_11103,N_10781);
and U17518 (N_17518,N_11953,N_11949);
xor U17519 (N_17519,N_13025,N_14016);
nand U17520 (N_17520,N_10663,N_10844);
and U17521 (N_17521,N_13474,N_10498);
nand U17522 (N_17522,N_12177,N_12722);
or U17523 (N_17523,N_13592,N_14388);
and U17524 (N_17524,N_14813,N_11810);
and U17525 (N_17525,N_14049,N_12430);
or U17526 (N_17526,N_13915,N_12220);
or U17527 (N_17527,N_10138,N_11147);
or U17528 (N_17528,N_10627,N_10986);
and U17529 (N_17529,N_12174,N_10167);
nand U17530 (N_17530,N_13479,N_11963);
or U17531 (N_17531,N_14114,N_10099);
xor U17532 (N_17532,N_14517,N_14335);
and U17533 (N_17533,N_11441,N_14681);
xor U17534 (N_17534,N_10478,N_11374);
nand U17535 (N_17535,N_12841,N_10568);
or U17536 (N_17536,N_10935,N_14072);
or U17537 (N_17537,N_14785,N_12614);
nor U17538 (N_17538,N_12703,N_14594);
and U17539 (N_17539,N_14040,N_11760);
nand U17540 (N_17540,N_14270,N_11667);
or U17541 (N_17541,N_13962,N_11412);
and U17542 (N_17542,N_11673,N_10532);
and U17543 (N_17543,N_13695,N_10368);
nor U17544 (N_17544,N_14101,N_14325);
xor U17545 (N_17545,N_14212,N_10019);
nand U17546 (N_17546,N_10698,N_10234);
nand U17547 (N_17547,N_13936,N_12239);
nor U17548 (N_17548,N_11937,N_11644);
nor U17549 (N_17549,N_13535,N_12056);
and U17550 (N_17550,N_14835,N_14623);
nand U17551 (N_17551,N_10220,N_11244);
nor U17552 (N_17552,N_12779,N_10142);
or U17553 (N_17553,N_14397,N_12190);
or U17554 (N_17554,N_12143,N_11497);
nand U17555 (N_17555,N_10619,N_14861);
nand U17556 (N_17556,N_11799,N_11580);
nand U17557 (N_17557,N_13454,N_11465);
or U17558 (N_17558,N_14892,N_14403);
nor U17559 (N_17559,N_13445,N_10607);
nor U17560 (N_17560,N_13281,N_10188);
nand U17561 (N_17561,N_11425,N_13991);
or U17562 (N_17562,N_10508,N_14514);
nand U17563 (N_17563,N_13964,N_10264);
nor U17564 (N_17564,N_10215,N_10553);
nor U17565 (N_17565,N_12431,N_12711);
nor U17566 (N_17566,N_14848,N_11828);
or U17567 (N_17567,N_12560,N_14555);
and U17568 (N_17568,N_12392,N_11289);
nor U17569 (N_17569,N_11984,N_13944);
nand U17570 (N_17570,N_10425,N_14382);
nor U17571 (N_17571,N_10634,N_11559);
and U17572 (N_17572,N_11874,N_12089);
nand U17573 (N_17573,N_10249,N_13539);
nor U17574 (N_17574,N_11015,N_10914);
nor U17575 (N_17575,N_13524,N_12455);
and U17576 (N_17576,N_11018,N_13154);
or U17577 (N_17577,N_11012,N_12387);
or U17578 (N_17578,N_14797,N_13075);
and U17579 (N_17579,N_14225,N_12721);
or U17580 (N_17580,N_10643,N_10404);
and U17581 (N_17581,N_14834,N_11241);
nor U17582 (N_17582,N_14831,N_14646);
and U17583 (N_17583,N_14192,N_13251);
nor U17584 (N_17584,N_12232,N_14739);
nor U17585 (N_17585,N_10171,N_14532);
nand U17586 (N_17586,N_10092,N_11369);
nand U17587 (N_17587,N_12570,N_12429);
nand U17588 (N_17588,N_12356,N_12220);
nor U17589 (N_17589,N_10443,N_10042);
nand U17590 (N_17590,N_13821,N_13122);
or U17591 (N_17591,N_14625,N_13073);
nor U17592 (N_17592,N_14698,N_10965);
nor U17593 (N_17593,N_13471,N_13368);
or U17594 (N_17594,N_14093,N_12601);
and U17595 (N_17595,N_10870,N_12120);
xor U17596 (N_17596,N_10687,N_12535);
and U17597 (N_17597,N_14865,N_12977);
or U17598 (N_17598,N_11152,N_14865);
xnor U17599 (N_17599,N_10701,N_10114);
and U17600 (N_17600,N_12365,N_11480);
nor U17601 (N_17601,N_12200,N_11262);
nor U17602 (N_17602,N_12363,N_11202);
and U17603 (N_17603,N_10029,N_11491);
nor U17604 (N_17604,N_13093,N_14128);
and U17605 (N_17605,N_11005,N_10762);
nor U17606 (N_17606,N_10331,N_14872);
nand U17607 (N_17607,N_10573,N_10977);
and U17608 (N_17608,N_11557,N_11278);
or U17609 (N_17609,N_12600,N_11344);
nand U17610 (N_17610,N_12797,N_10554);
nand U17611 (N_17611,N_12031,N_13676);
xor U17612 (N_17612,N_14263,N_10469);
xnor U17613 (N_17613,N_12630,N_13594);
nand U17614 (N_17614,N_13775,N_14506);
nand U17615 (N_17615,N_14036,N_14051);
nand U17616 (N_17616,N_10172,N_13883);
or U17617 (N_17617,N_13571,N_11951);
or U17618 (N_17618,N_14061,N_10854);
or U17619 (N_17619,N_13215,N_12508);
xor U17620 (N_17620,N_13266,N_13647);
and U17621 (N_17621,N_11990,N_14565);
nand U17622 (N_17622,N_10224,N_12375);
and U17623 (N_17623,N_14416,N_13474);
nor U17624 (N_17624,N_13085,N_13477);
nand U17625 (N_17625,N_13214,N_12774);
xor U17626 (N_17626,N_13614,N_10142);
nor U17627 (N_17627,N_12826,N_12891);
or U17628 (N_17628,N_14046,N_14094);
nand U17629 (N_17629,N_13096,N_10628);
or U17630 (N_17630,N_11761,N_13005);
and U17631 (N_17631,N_10720,N_10713);
and U17632 (N_17632,N_12726,N_12467);
nor U17633 (N_17633,N_10411,N_12182);
nand U17634 (N_17634,N_11779,N_13224);
or U17635 (N_17635,N_11599,N_12771);
and U17636 (N_17636,N_12138,N_12418);
nand U17637 (N_17637,N_14042,N_10070);
nand U17638 (N_17638,N_14349,N_13163);
nor U17639 (N_17639,N_12384,N_10676);
and U17640 (N_17640,N_10183,N_11297);
and U17641 (N_17641,N_12945,N_11148);
and U17642 (N_17642,N_13994,N_11169);
and U17643 (N_17643,N_12440,N_11024);
and U17644 (N_17644,N_11672,N_11755);
or U17645 (N_17645,N_11768,N_12169);
and U17646 (N_17646,N_11738,N_11407);
nand U17647 (N_17647,N_10510,N_10844);
nor U17648 (N_17648,N_12252,N_11847);
or U17649 (N_17649,N_13688,N_14270);
or U17650 (N_17650,N_11680,N_12529);
nor U17651 (N_17651,N_10941,N_12762);
or U17652 (N_17652,N_11047,N_13205);
or U17653 (N_17653,N_12780,N_10556);
and U17654 (N_17654,N_14139,N_12008);
or U17655 (N_17655,N_14660,N_11817);
nand U17656 (N_17656,N_14763,N_14411);
nand U17657 (N_17657,N_10215,N_14845);
and U17658 (N_17658,N_11980,N_11924);
or U17659 (N_17659,N_14548,N_13496);
nand U17660 (N_17660,N_10268,N_11928);
xnor U17661 (N_17661,N_13823,N_12397);
and U17662 (N_17662,N_13298,N_12515);
or U17663 (N_17663,N_10304,N_11829);
or U17664 (N_17664,N_14728,N_12935);
nand U17665 (N_17665,N_14303,N_12169);
nor U17666 (N_17666,N_13398,N_10328);
and U17667 (N_17667,N_10278,N_12522);
and U17668 (N_17668,N_13564,N_11849);
xor U17669 (N_17669,N_13493,N_12528);
nor U17670 (N_17670,N_12616,N_12942);
nand U17671 (N_17671,N_10704,N_13764);
nand U17672 (N_17672,N_14823,N_10668);
nor U17673 (N_17673,N_13116,N_11725);
or U17674 (N_17674,N_10249,N_14473);
or U17675 (N_17675,N_10073,N_10110);
or U17676 (N_17676,N_10895,N_14076);
and U17677 (N_17677,N_14158,N_10103);
nor U17678 (N_17678,N_14975,N_12102);
nor U17679 (N_17679,N_11653,N_14446);
nor U17680 (N_17680,N_10884,N_10461);
nor U17681 (N_17681,N_11880,N_12823);
and U17682 (N_17682,N_10238,N_12636);
xnor U17683 (N_17683,N_12733,N_10028);
or U17684 (N_17684,N_14859,N_14755);
or U17685 (N_17685,N_10503,N_13349);
nand U17686 (N_17686,N_14006,N_14305);
xnor U17687 (N_17687,N_12234,N_12283);
and U17688 (N_17688,N_14483,N_14816);
or U17689 (N_17689,N_11234,N_14333);
xor U17690 (N_17690,N_12473,N_12584);
or U17691 (N_17691,N_11851,N_14153);
nand U17692 (N_17692,N_12169,N_10511);
or U17693 (N_17693,N_12407,N_14178);
nand U17694 (N_17694,N_10958,N_11315);
and U17695 (N_17695,N_12751,N_12798);
xor U17696 (N_17696,N_11121,N_10327);
nor U17697 (N_17697,N_12239,N_12350);
and U17698 (N_17698,N_14113,N_12612);
and U17699 (N_17699,N_14405,N_12875);
nand U17700 (N_17700,N_11026,N_12149);
nor U17701 (N_17701,N_11312,N_12054);
or U17702 (N_17702,N_14730,N_11028);
nand U17703 (N_17703,N_14437,N_11884);
and U17704 (N_17704,N_13773,N_12045);
nor U17705 (N_17705,N_13559,N_13852);
and U17706 (N_17706,N_14059,N_14825);
xor U17707 (N_17707,N_12339,N_11952);
nand U17708 (N_17708,N_13372,N_11469);
nor U17709 (N_17709,N_13222,N_12170);
or U17710 (N_17710,N_11789,N_12924);
and U17711 (N_17711,N_11731,N_10072);
or U17712 (N_17712,N_10184,N_13743);
nor U17713 (N_17713,N_13498,N_11315);
and U17714 (N_17714,N_14367,N_11576);
xnor U17715 (N_17715,N_10735,N_10396);
nor U17716 (N_17716,N_14598,N_10541);
nor U17717 (N_17717,N_10823,N_13895);
and U17718 (N_17718,N_12403,N_13556);
nand U17719 (N_17719,N_14509,N_13427);
or U17720 (N_17720,N_11889,N_11237);
nor U17721 (N_17721,N_11630,N_10079);
or U17722 (N_17722,N_13592,N_14363);
xor U17723 (N_17723,N_10867,N_12411);
or U17724 (N_17724,N_10025,N_11445);
or U17725 (N_17725,N_12570,N_12694);
nand U17726 (N_17726,N_14287,N_10026);
nor U17727 (N_17727,N_14306,N_11208);
and U17728 (N_17728,N_13810,N_12617);
nand U17729 (N_17729,N_11783,N_10027);
and U17730 (N_17730,N_10290,N_10613);
and U17731 (N_17731,N_14712,N_10269);
xor U17732 (N_17732,N_10748,N_10274);
nor U17733 (N_17733,N_11496,N_13484);
and U17734 (N_17734,N_12122,N_13121);
and U17735 (N_17735,N_13568,N_12239);
nand U17736 (N_17736,N_13918,N_10323);
nor U17737 (N_17737,N_10144,N_14232);
or U17738 (N_17738,N_12879,N_13256);
nor U17739 (N_17739,N_10797,N_12012);
nand U17740 (N_17740,N_13566,N_11003);
or U17741 (N_17741,N_11214,N_11100);
nand U17742 (N_17742,N_13063,N_14631);
or U17743 (N_17743,N_13862,N_13175);
or U17744 (N_17744,N_11479,N_14959);
or U17745 (N_17745,N_13804,N_13353);
xnor U17746 (N_17746,N_10635,N_12766);
and U17747 (N_17747,N_11685,N_14372);
or U17748 (N_17748,N_12160,N_13984);
nand U17749 (N_17749,N_11992,N_12206);
nand U17750 (N_17750,N_10147,N_14053);
or U17751 (N_17751,N_10880,N_13436);
or U17752 (N_17752,N_10742,N_10005);
xnor U17753 (N_17753,N_14588,N_14591);
or U17754 (N_17754,N_10215,N_12556);
nor U17755 (N_17755,N_11547,N_11644);
nand U17756 (N_17756,N_10900,N_13392);
nand U17757 (N_17757,N_11752,N_13268);
and U17758 (N_17758,N_13265,N_14064);
xor U17759 (N_17759,N_11873,N_14559);
nand U17760 (N_17760,N_11312,N_13686);
and U17761 (N_17761,N_13513,N_14434);
nand U17762 (N_17762,N_12289,N_11901);
nor U17763 (N_17763,N_13318,N_10775);
nand U17764 (N_17764,N_12053,N_14467);
nor U17765 (N_17765,N_10399,N_13170);
nor U17766 (N_17766,N_11371,N_10581);
and U17767 (N_17767,N_13103,N_13761);
xor U17768 (N_17768,N_14284,N_12682);
nand U17769 (N_17769,N_13282,N_13354);
or U17770 (N_17770,N_13028,N_11624);
and U17771 (N_17771,N_10125,N_10803);
xor U17772 (N_17772,N_13696,N_10340);
nand U17773 (N_17773,N_14566,N_10044);
xnor U17774 (N_17774,N_10097,N_12674);
nand U17775 (N_17775,N_11291,N_11116);
nor U17776 (N_17776,N_14805,N_13363);
and U17777 (N_17777,N_10867,N_10653);
xnor U17778 (N_17778,N_13470,N_11422);
and U17779 (N_17779,N_11924,N_13751);
nand U17780 (N_17780,N_13156,N_13559);
nand U17781 (N_17781,N_11606,N_13549);
or U17782 (N_17782,N_13334,N_13870);
or U17783 (N_17783,N_11705,N_14295);
nor U17784 (N_17784,N_10351,N_12870);
nand U17785 (N_17785,N_13078,N_12470);
and U17786 (N_17786,N_11099,N_13736);
and U17787 (N_17787,N_11182,N_11741);
nand U17788 (N_17788,N_10204,N_11600);
nand U17789 (N_17789,N_14654,N_11065);
nand U17790 (N_17790,N_10182,N_13984);
nor U17791 (N_17791,N_10895,N_12726);
and U17792 (N_17792,N_14590,N_13065);
nand U17793 (N_17793,N_11422,N_13607);
or U17794 (N_17794,N_12379,N_12369);
and U17795 (N_17795,N_13180,N_14718);
nand U17796 (N_17796,N_11534,N_14171);
xor U17797 (N_17797,N_11384,N_12598);
and U17798 (N_17798,N_13755,N_10333);
nor U17799 (N_17799,N_13251,N_10407);
xnor U17800 (N_17800,N_13660,N_13707);
nand U17801 (N_17801,N_12493,N_12034);
and U17802 (N_17802,N_11720,N_12030);
nor U17803 (N_17803,N_11563,N_11858);
or U17804 (N_17804,N_12102,N_14276);
nand U17805 (N_17805,N_10436,N_13076);
and U17806 (N_17806,N_10823,N_10852);
nand U17807 (N_17807,N_12138,N_14955);
and U17808 (N_17808,N_13137,N_14886);
or U17809 (N_17809,N_11559,N_13517);
nand U17810 (N_17810,N_14276,N_11167);
nand U17811 (N_17811,N_12110,N_14305);
and U17812 (N_17812,N_12045,N_12098);
xor U17813 (N_17813,N_13261,N_12149);
nand U17814 (N_17814,N_11957,N_13214);
nor U17815 (N_17815,N_14574,N_11903);
nand U17816 (N_17816,N_12843,N_12357);
nand U17817 (N_17817,N_14105,N_14230);
and U17818 (N_17818,N_11875,N_14413);
nor U17819 (N_17819,N_12156,N_10475);
nor U17820 (N_17820,N_14130,N_12069);
xnor U17821 (N_17821,N_13017,N_13132);
or U17822 (N_17822,N_13991,N_11042);
or U17823 (N_17823,N_11925,N_14562);
nor U17824 (N_17824,N_11101,N_12966);
and U17825 (N_17825,N_12933,N_10343);
and U17826 (N_17826,N_11662,N_11979);
or U17827 (N_17827,N_11783,N_10296);
nor U17828 (N_17828,N_12630,N_13316);
and U17829 (N_17829,N_11523,N_13834);
or U17830 (N_17830,N_12577,N_12277);
nor U17831 (N_17831,N_11616,N_13465);
nor U17832 (N_17832,N_12665,N_13813);
and U17833 (N_17833,N_13810,N_14305);
and U17834 (N_17834,N_14586,N_12517);
nor U17835 (N_17835,N_10971,N_14465);
nor U17836 (N_17836,N_11731,N_11061);
xor U17837 (N_17837,N_13266,N_13195);
and U17838 (N_17838,N_12024,N_14678);
and U17839 (N_17839,N_11272,N_10728);
or U17840 (N_17840,N_11433,N_12847);
or U17841 (N_17841,N_14009,N_13007);
or U17842 (N_17842,N_12795,N_13057);
nand U17843 (N_17843,N_12499,N_13766);
nor U17844 (N_17844,N_13217,N_10418);
nand U17845 (N_17845,N_10347,N_12760);
nand U17846 (N_17846,N_11737,N_11086);
and U17847 (N_17847,N_11136,N_14781);
nand U17848 (N_17848,N_14968,N_14099);
or U17849 (N_17849,N_13095,N_10602);
xor U17850 (N_17850,N_10706,N_14989);
nor U17851 (N_17851,N_13072,N_12833);
nand U17852 (N_17852,N_10374,N_13608);
xnor U17853 (N_17853,N_14726,N_13916);
and U17854 (N_17854,N_14442,N_14764);
nor U17855 (N_17855,N_11900,N_14501);
or U17856 (N_17856,N_10621,N_13382);
nand U17857 (N_17857,N_11135,N_11278);
and U17858 (N_17858,N_12702,N_10851);
or U17859 (N_17859,N_13253,N_14828);
nor U17860 (N_17860,N_12666,N_12264);
nor U17861 (N_17861,N_10497,N_12068);
nand U17862 (N_17862,N_11727,N_10362);
nand U17863 (N_17863,N_11108,N_13806);
and U17864 (N_17864,N_10739,N_12917);
or U17865 (N_17865,N_11056,N_10852);
and U17866 (N_17866,N_12950,N_13380);
nand U17867 (N_17867,N_12282,N_10893);
or U17868 (N_17868,N_12566,N_11417);
and U17869 (N_17869,N_11894,N_13934);
nor U17870 (N_17870,N_11027,N_14282);
nand U17871 (N_17871,N_13805,N_14533);
and U17872 (N_17872,N_10997,N_13289);
nor U17873 (N_17873,N_14101,N_14133);
or U17874 (N_17874,N_14204,N_11904);
nand U17875 (N_17875,N_11496,N_10385);
and U17876 (N_17876,N_13301,N_13855);
or U17877 (N_17877,N_13945,N_10913);
nand U17878 (N_17878,N_12639,N_14742);
nand U17879 (N_17879,N_10127,N_11983);
nand U17880 (N_17880,N_10145,N_10633);
xnor U17881 (N_17881,N_13043,N_12239);
and U17882 (N_17882,N_11846,N_11789);
and U17883 (N_17883,N_10402,N_11133);
nor U17884 (N_17884,N_14457,N_13506);
nand U17885 (N_17885,N_10463,N_11502);
or U17886 (N_17886,N_11600,N_11701);
or U17887 (N_17887,N_13886,N_12313);
xnor U17888 (N_17888,N_10327,N_13530);
nor U17889 (N_17889,N_13004,N_13399);
nand U17890 (N_17890,N_13346,N_12645);
nand U17891 (N_17891,N_10237,N_13532);
nand U17892 (N_17892,N_13609,N_10087);
nor U17893 (N_17893,N_12284,N_10843);
and U17894 (N_17894,N_13991,N_11246);
nor U17895 (N_17895,N_13982,N_14045);
or U17896 (N_17896,N_11394,N_12086);
nor U17897 (N_17897,N_10036,N_12842);
nor U17898 (N_17898,N_10012,N_10829);
or U17899 (N_17899,N_12312,N_14139);
nor U17900 (N_17900,N_14066,N_10600);
and U17901 (N_17901,N_12826,N_14522);
nor U17902 (N_17902,N_13687,N_14009);
nand U17903 (N_17903,N_11200,N_14277);
nand U17904 (N_17904,N_12785,N_12121);
nor U17905 (N_17905,N_12116,N_12349);
or U17906 (N_17906,N_11650,N_13534);
nand U17907 (N_17907,N_12461,N_11762);
nand U17908 (N_17908,N_14799,N_13615);
or U17909 (N_17909,N_12364,N_12236);
or U17910 (N_17910,N_13289,N_10978);
or U17911 (N_17911,N_14304,N_13173);
nor U17912 (N_17912,N_14239,N_12927);
nand U17913 (N_17913,N_14515,N_10609);
or U17914 (N_17914,N_11184,N_14000);
nor U17915 (N_17915,N_11538,N_10992);
and U17916 (N_17916,N_13259,N_14491);
and U17917 (N_17917,N_14244,N_10516);
nand U17918 (N_17918,N_14925,N_10397);
xnor U17919 (N_17919,N_12638,N_14891);
nor U17920 (N_17920,N_11382,N_11100);
nor U17921 (N_17921,N_10052,N_13091);
nor U17922 (N_17922,N_12339,N_14969);
nor U17923 (N_17923,N_10848,N_10156);
and U17924 (N_17924,N_12643,N_11611);
or U17925 (N_17925,N_12473,N_13356);
nand U17926 (N_17926,N_13438,N_14253);
and U17927 (N_17927,N_11567,N_10283);
or U17928 (N_17928,N_13848,N_14047);
and U17929 (N_17929,N_11104,N_14099);
or U17930 (N_17930,N_10723,N_12963);
nand U17931 (N_17931,N_13951,N_14252);
and U17932 (N_17932,N_12880,N_10816);
or U17933 (N_17933,N_14203,N_12388);
nand U17934 (N_17934,N_11012,N_11014);
nand U17935 (N_17935,N_12592,N_14964);
and U17936 (N_17936,N_11131,N_10117);
nor U17937 (N_17937,N_10122,N_10298);
nor U17938 (N_17938,N_10758,N_11519);
nor U17939 (N_17939,N_10062,N_11495);
nand U17940 (N_17940,N_14446,N_13358);
xor U17941 (N_17941,N_11030,N_10337);
and U17942 (N_17942,N_12334,N_12676);
or U17943 (N_17943,N_10042,N_12152);
nor U17944 (N_17944,N_13387,N_11037);
and U17945 (N_17945,N_10816,N_12306);
or U17946 (N_17946,N_14592,N_12442);
xnor U17947 (N_17947,N_12082,N_11084);
nor U17948 (N_17948,N_14657,N_12127);
and U17949 (N_17949,N_10403,N_10814);
nor U17950 (N_17950,N_10408,N_14686);
nor U17951 (N_17951,N_10288,N_13137);
and U17952 (N_17952,N_10906,N_14668);
or U17953 (N_17953,N_14404,N_12922);
or U17954 (N_17954,N_14229,N_12512);
and U17955 (N_17955,N_12585,N_10012);
nand U17956 (N_17956,N_12763,N_11807);
nor U17957 (N_17957,N_14485,N_14165);
or U17958 (N_17958,N_12243,N_14147);
xnor U17959 (N_17959,N_12503,N_14742);
and U17960 (N_17960,N_11670,N_12907);
or U17961 (N_17961,N_10996,N_10178);
or U17962 (N_17962,N_12099,N_13415);
or U17963 (N_17963,N_11703,N_11451);
or U17964 (N_17964,N_13675,N_11101);
and U17965 (N_17965,N_10116,N_13820);
and U17966 (N_17966,N_10266,N_10609);
and U17967 (N_17967,N_14233,N_14783);
or U17968 (N_17968,N_14220,N_11835);
xor U17969 (N_17969,N_12651,N_10129);
or U17970 (N_17970,N_12053,N_10867);
and U17971 (N_17971,N_10013,N_11198);
nand U17972 (N_17972,N_12269,N_12586);
nor U17973 (N_17973,N_12695,N_11494);
or U17974 (N_17974,N_13205,N_12271);
and U17975 (N_17975,N_11590,N_11555);
nor U17976 (N_17976,N_14469,N_12519);
and U17977 (N_17977,N_13483,N_12240);
nor U17978 (N_17978,N_11767,N_10107);
xor U17979 (N_17979,N_10215,N_12406);
xnor U17980 (N_17980,N_12940,N_13829);
xor U17981 (N_17981,N_13015,N_12544);
xnor U17982 (N_17982,N_13317,N_10908);
xor U17983 (N_17983,N_14476,N_10864);
nand U17984 (N_17984,N_14773,N_14365);
xnor U17985 (N_17985,N_14311,N_10216);
nand U17986 (N_17986,N_10717,N_12598);
nand U17987 (N_17987,N_14595,N_13317);
xor U17988 (N_17988,N_13379,N_14416);
nor U17989 (N_17989,N_10941,N_10588);
xnor U17990 (N_17990,N_12577,N_14646);
nand U17991 (N_17991,N_13307,N_14517);
or U17992 (N_17992,N_14618,N_12828);
or U17993 (N_17993,N_13622,N_12502);
or U17994 (N_17994,N_13333,N_10340);
xor U17995 (N_17995,N_14848,N_11263);
nor U17996 (N_17996,N_11968,N_11678);
nor U17997 (N_17997,N_10740,N_13031);
and U17998 (N_17998,N_11660,N_11798);
nor U17999 (N_17999,N_11008,N_13035);
or U18000 (N_18000,N_14383,N_10269);
and U18001 (N_18001,N_13047,N_13783);
nand U18002 (N_18002,N_14541,N_13541);
or U18003 (N_18003,N_14945,N_13381);
nor U18004 (N_18004,N_12742,N_13761);
nand U18005 (N_18005,N_14897,N_11393);
or U18006 (N_18006,N_10330,N_12636);
and U18007 (N_18007,N_12342,N_11081);
xnor U18008 (N_18008,N_14201,N_11782);
nor U18009 (N_18009,N_13056,N_14753);
and U18010 (N_18010,N_10146,N_11539);
and U18011 (N_18011,N_10446,N_10385);
xnor U18012 (N_18012,N_12206,N_13942);
nor U18013 (N_18013,N_12829,N_11381);
and U18014 (N_18014,N_13362,N_12931);
nor U18015 (N_18015,N_12729,N_10442);
nor U18016 (N_18016,N_12320,N_12457);
nor U18017 (N_18017,N_13952,N_14851);
nor U18018 (N_18018,N_14413,N_10849);
nand U18019 (N_18019,N_12731,N_13810);
nor U18020 (N_18020,N_11045,N_11059);
and U18021 (N_18021,N_14246,N_12510);
nand U18022 (N_18022,N_11408,N_10791);
xnor U18023 (N_18023,N_13289,N_13421);
nand U18024 (N_18024,N_12145,N_12390);
or U18025 (N_18025,N_13149,N_10613);
and U18026 (N_18026,N_14941,N_12222);
and U18027 (N_18027,N_13991,N_12579);
or U18028 (N_18028,N_10487,N_11578);
nor U18029 (N_18029,N_10105,N_11755);
or U18030 (N_18030,N_14395,N_11989);
and U18031 (N_18031,N_13667,N_10805);
nor U18032 (N_18032,N_12726,N_13783);
or U18033 (N_18033,N_11645,N_14726);
or U18034 (N_18034,N_12233,N_11951);
nand U18035 (N_18035,N_14204,N_11583);
xor U18036 (N_18036,N_13886,N_14498);
and U18037 (N_18037,N_12056,N_10418);
nor U18038 (N_18038,N_11041,N_12897);
nand U18039 (N_18039,N_11438,N_14566);
nand U18040 (N_18040,N_14323,N_11804);
xnor U18041 (N_18041,N_11775,N_12699);
nand U18042 (N_18042,N_10125,N_14300);
nand U18043 (N_18043,N_14323,N_12137);
and U18044 (N_18044,N_12613,N_10158);
or U18045 (N_18045,N_13327,N_14893);
or U18046 (N_18046,N_12023,N_11081);
nand U18047 (N_18047,N_11949,N_13468);
or U18048 (N_18048,N_12199,N_14258);
and U18049 (N_18049,N_12036,N_12039);
or U18050 (N_18050,N_11628,N_10975);
nand U18051 (N_18051,N_11180,N_11269);
or U18052 (N_18052,N_14406,N_13946);
or U18053 (N_18053,N_10150,N_12909);
nor U18054 (N_18054,N_14421,N_10737);
or U18055 (N_18055,N_13973,N_13044);
or U18056 (N_18056,N_13501,N_14747);
nand U18057 (N_18057,N_14410,N_11041);
nand U18058 (N_18058,N_11457,N_12218);
nor U18059 (N_18059,N_13358,N_12868);
nor U18060 (N_18060,N_11951,N_13185);
or U18061 (N_18061,N_14424,N_10690);
and U18062 (N_18062,N_11759,N_14066);
nand U18063 (N_18063,N_10158,N_11571);
nand U18064 (N_18064,N_14495,N_12208);
nand U18065 (N_18065,N_13735,N_10357);
and U18066 (N_18066,N_10655,N_13111);
or U18067 (N_18067,N_13478,N_10756);
nor U18068 (N_18068,N_10125,N_14904);
and U18069 (N_18069,N_13686,N_13659);
nand U18070 (N_18070,N_10136,N_12789);
or U18071 (N_18071,N_11562,N_10329);
nand U18072 (N_18072,N_13293,N_12604);
nor U18073 (N_18073,N_11498,N_10219);
nand U18074 (N_18074,N_13724,N_10765);
nand U18075 (N_18075,N_12062,N_14881);
nand U18076 (N_18076,N_13656,N_13795);
nor U18077 (N_18077,N_10168,N_14418);
and U18078 (N_18078,N_11571,N_10423);
nor U18079 (N_18079,N_12624,N_13430);
and U18080 (N_18080,N_10624,N_14441);
and U18081 (N_18081,N_12112,N_13817);
xnor U18082 (N_18082,N_14069,N_11103);
xor U18083 (N_18083,N_14536,N_12021);
and U18084 (N_18084,N_13531,N_13346);
and U18085 (N_18085,N_10936,N_10490);
and U18086 (N_18086,N_14595,N_10284);
or U18087 (N_18087,N_12910,N_14173);
nand U18088 (N_18088,N_12076,N_12956);
nor U18089 (N_18089,N_11023,N_10837);
and U18090 (N_18090,N_10255,N_13916);
nor U18091 (N_18091,N_12576,N_13433);
nand U18092 (N_18092,N_12309,N_14196);
nor U18093 (N_18093,N_13627,N_13043);
xor U18094 (N_18094,N_13198,N_10729);
or U18095 (N_18095,N_10925,N_13759);
and U18096 (N_18096,N_13652,N_12920);
or U18097 (N_18097,N_11230,N_11706);
nor U18098 (N_18098,N_14362,N_12060);
and U18099 (N_18099,N_13404,N_12021);
and U18100 (N_18100,N_14591,N_12507);
nand U18101 (N_18101,N_12796,N_11345);
nor U18102 (N_18102,N_10416,N_10222);
nand U18103 (N_18103,N_14729,N_14325);
and U18104 (N_18104,N_11232,N_10581);
nand U18105 (N_18105,N_10158,N_13894);
nor U18106 (N_18106,N_10124,N_11032);
nand U18107 (N_18107,N_13887,N_14118);
nor U18108 (N_18108,N_12232,N_14341);
nand U18109 (N_18109,N_11342,N_10737);
nor U18110 (N_18110,N_13738,N_12885);
nor U18111 (N_18111,N_12134,N_13374);
nand U18112 (N_18112,N_12023,N_11181);
or U18113 (N_18113,N_12961,N_13930);
nand U18114 (N_18114,N_11013,N_10457);
and U18115 (N_18115,N_14353,N_13528);
and U18116 (N_18116,N_14376,N_12730);
nor U18117 (N_18117,N_14857,N_13602);
nand U18118 (N_18118,N_10295,N_11515);
nand U18119 (N_18119,N_12897,N_10351);
nor U18120 (N_18120,N_11301,N_12061);
nor U18121 (N_18121,N_11981,N_10235);
nor U18122 (N_18122,N_14678,N_12630);
or U18123 (N_18123,N_10911,N_10319);
or U18124 (N_18124,N_11595,N_14819);
nand U18125 (N_18125,N_14029,N_13561);
or U18126 (N_18126,N_13940,N_10928);
and U18127 (N_18127,N_12022,N_12751);
nor U18128 (N_18128,N_14207,N_10398);
and U18129 (N_18129,N_13110,N_12297);
and U18130 (N_18130,N_11596,N_13087);
or U18131 (N_18131,N_13524,N_12950);
nand U18132 (N_18132,N_11978,N_13439);
and U18133 (N_18133,N_11890,N_13359);
nand U18134 (N_18134,N_12659,N_14304);
and U18135 (N_18135,N_13899,N_10707);
nand U18136 (N_18136,N_13806,N_10548);
and U18137 (N_18137,N_12577,N_14581);
nor U18138 (N_18138,N_10906,N_13918);
or U18139 (N_18139,N_14799,N_10637);
and U18140 (N_18140,N_11405,N_10268);
or U18141 (N_18141,N_12542,N_11919);
nor U18142 (N_18142,N_11824,N_14986);
and U18143 (N_18143,N_12390,N_11999);
nand U18144 (N_18144,N_12011,N_13043);
xor U18145 (N_18145,N_10670,N_14293);
and U18146 (N_18146,N_13816,N_13206);
xor U18147 (N_18147,N_13299,N_13993);
nor U18148 (N_18148,N_11906,N_13654);
and U18149 (N_18149,N_13772,N_13613);
or U18150 (N_18150,N_11182,N_11085);
nand U18151 (N_18151,N_12218,N_14072);
or U18152 (N_18152,N_12478,N_11562);
or U18153 (N_18153,N_10742,N_11798);
or U18154 (N_18154,N_11891,N_12579);
nor U18155 (N_18155,N_12532,N_11532);
nor U18156 (N_18156,N_10021,N_13815);
or U18157 (N_18157,N_10500,N_10468);
or U18158 (N_18158,N_11437,N_11530);
or U18159 (N_18159,N_13265,N_10570);
or U18160 (N_18160,N_10142,N_13069);
nand U18161 (N_18161,N_14391,N_11414);
xnor U18162 (N_18162,N_14748,N_14254);
and U18163 (N_18163,N_11308,N_13520);
nor U18164 (N_18164,N_13745,N_14198);
nand U18165 (N_18165,N_11944,N_11755);
nand U18166 (N_18166,N_14697,N_14322);
and U18167 (N_18167,N_14925,N_14538);
or U18168 (N_18168,N_10894,N_10365);
nor U18169 (N_18169,N_12233,N_10610);
nor U18170 (N_18170,N_11864,N_12520);
nand U18171 (N_18171,N_13723,N_11467);
and U18172 (N_18172,N_10273,N_11644);
nor U18173 (N_18173,N_12297,N_14634);
xor U18174 (N_18174,N_14425,N_13328);
nand U18175 (N_18175,N_11239,N_14512);
and U18176 (N_18176,N_12836,N_11188);
nor U18177 (N_18177,N_11685,N_12455);
or U18178 (N_18178,N_11361,N_12522);
or U18179 (N_18179,N_10301,N_12411);
or U18180 (N_18180,N_10505,N_12487);
or U18181 (N_18181,N_12734,N_14418);
nor U18182 (N_18182,N_13547,N_13632);
or U18183 (N_18183,N_12222,N_10722);
or U18184 (N_18184,N_14270,N_12019);
nor U18185 (N_18185,N_12471,N_10596);
nand U18186 (N_18186,N_12468,N_12019);
and U18187 (N_18187,N_13993,N_12851);
nor U18188 (N_18188,N_13345,N_13812);
nand U18189 (N_18189,N_12045,N_13852);
nand U18190 (N_18190,N_11226,N_12691);
nor U18191 (N_18191,N_14938,N_14176);
nand U18192 (N_18192,N_10000,N_10514);
or U18193 (N_18193,N_14094,N_12153);
nand U18194 (N_18194,N_12134,N_13272);
or U18195 (N_18195,N_10501,N_14232);
nand U18196 (N_18196,N_11993,N_14200);
or U18197 (N_18197,N_13648,N_13278);
nor U18198 (N_18198,N_11477,N_13175);
and U18199 (N_18199,N_10360,N_12750);
or U18200 (N_18200,N_14589,N_12392);
and U18201 (N_18201,N_10621,N_13679);
or U18202 (N_18202,N_14679,N_10491);
nand U18203 (N_18203,N_13263,N_10369);
and U18204 (N_18204,N_11333,N_11124);
nand U18205 (N_18205,N_11681,N_11456);
or U18206 (N_18206,N_14420,N_13841);
and U18207 (N_18207,N_11800,N_11472);
nand U18208 (N_18208,N_14934,N_13190);
nand U18209 (N_18209,N_10309,N_14864);
or U18210 (N_18210,N_12617,N_12161);
nand U18211 (N_18211,N_13480,N_13598);
xor U18212 (N_18212,N_10454,N_11809);
or U18213 (N_18213,N_11900,N_12793);
nand U18214 (N_18214,N_11562,N_13292);
nor U18215 (N_18215,N_13108,N_12997);
nand U18216 (N_18216,N_12070,N_10108);
and U18217 (N_18217,N_11846,N_11443);
nand U18218 (N_18218,N_10799,N_10188);
xor U18219 (N_18219,N_13101,N_10349);
or U18220 (N_18220,N_14350,N_10188);
xnor U18221 (N_18221,N_10628,N_12555);
nor U18222 (N_18222,N_10400,N_13323);
xor U18223 (N_18223,N_11984,N_10098);
nand U18224 (N_18224,N_13522,N_13795);
nand U18225 (N_18225,N_10257,N_12136);
xor U18226 (N_18226,N_10582,N_12809);
or U18227 (N_18227,N_10345,N_10334);
and U18228 (N_18228,N_12511,N_12123);
nand U18229 (N_18229,N_13983,N_10245);
and U18230 (N_18230,N_12760,N_12484);
nand U18231 (N_18231,N_11533,N_12157);
nor U18232 (N_18232,N_12527,N_10544);
and U18233 (N_18233,N_11012,N_14878);
nor U18234 (N_18234,N_14900,N_14312);
or U18235 (N_18235,N_14020,N_14805);
nor U18236 (N_18236,N_14704,N_14118);
xor U18237 (N_18237,N_10945,N_12434);
nor U18238 (N_18238,N_14824,N_12386);
nor U18239 (N_18239,N_12531,N_14094);
nand U18240 (N_18240,N_13134,N_10339);
nand U18241 (N_18241,N_11387,N_11717);
nor U18242 (N_18242,N_11040,N_12880);
nor U18243 (N_18243,N_12207,N_14142);
xnor U18244 (N_18244,N_14838,N_12085);
and U18245 (N_18245,N_10179,N_13589);
xnor U18246 (N_18246,N_14079,N_12974);
or U18247 (N_18247,N_12120,N_13313);
and U18248 (N_18248,N_11663,N_13349);
nor U18249 (N_18249,N_10072,N_11291);
and U18250 (N_18250,N_14861,N_10769);
or U18251 (N_18251,N_14425,N_14075);
xnor U18252 (N_18252,N_10807,N_12082);
or U18253 (N_18253,N_14480,N_13994);
or U18254 (N_18254,N_12270,N_14577);
or U18255 (N_18255,N_12354,N_12563);
nand U18256 (N_18256,N_14693,N_13509);
and U18257 (N_18257,N_11542,N_11311);
nand U18258 (N_18258,N_10601,N_14598);
or U18259 (N_18259,N_12344,N_12138);
and U18260 (N_18260,N_14503,N_11519);
nor U18261 (N_18261,N_11701,N_14818);
nor U18262 (N_18262,N_13035,N_10335);
or U18263 (N_18263,N_10256,N_11009);
and U18264 (N_18264,N_11124,N_12688);
nand U18265 (N_18265,N_13932,N_14058);
nand U18266 (N_18266,N_14183,N_13627);
and U18267 (N_18267,N_14429,N_10177);
nand U18268 (N_18268,N_14631,N_10271);
and U18269 (N_18269,N_12800,N_14484);
nand U18270 (N_18270,N_14162,N_13675);
nand U18271 (N_18271,N_10463,N_10006);
nand U18272 (N_18272,N_11188,N_14519);
and U18273 (N_18273,N_12481,N_10073);
nor U18274 (N_18274,N_10077,N_11473);
or U18275 (N_18275,N_12619,N_13574);
nor U18276 (N_18276,N_11951,N_14116);
or U18277 (N_18277,N_11423,N_11276);
nor U18278 (N_18278,N_10512,N_14488);
xor U18279 (N_18279,N_11070,N_14171);
and U18280 (N_18280,N_12693,N_14336);
or U18281 (N_18281,N_13404,N_12489);
or U18282 (N_18282,N_14322,N_13912);
nor U18283 (N_18283,N_13593,N_12144);
nor U18284 (N_18284,N_10052,N_13280);
and U18285 (N_18285,N_14355,N_14726);
nand U18286 (N_18286,N_11279,N_10703);
xor U18287 (N_18287,N_10778,N_13830);
nand U18288 (N_18288,N_13973,N_13318);
xnor U18289 (N_18289,N_11787,N_12227);
nand U18290 (N_18290,N_11454,N_11559);
nand U18291 (N_18291,N_14418,N_13305);
nor U18292 (N_18292,N_10536,N_12077);
and U18293 (N_18293,N_12126,N_11077);
nand U18294 (N_18294,N_13238,N_10647);
xor U18295 (N_18295,N_12946,N_14349);
and U18296 (N_18296,N_14896,N_12152);
xor U18297 (N_18297,N_13197,N_10073);
nor U18298 (N_18298,N_13121,N_10270);
nor U18299 (N_18299,N_11318,N_10428);
nor U18300 (N_18300,N_14897,N_12003);
and U18301 (N_18301,N_10672,N_12958);
and U18302 (N_18302,N_11388,N_13638);
nor U18303 (N_18303,N_13229,N_11510);
or U18304 (N_18304,N_13281,N_11228);
or U18305 (N_18305,N_14508,N_11153);
nand U18306 (N_18306,N_12627,N_14295);
and U18307 (N_18307,N_12366,N_10873);
xnor U18308 (N_18308,N_10254,N_11193);
and U18309 (N_18309,N_13988,N_10675);
and U18310 (N_18310,N_12769,N_10622);
nor U18311 (N_18311,N_10751,N_10509);
nor U18312 (N_18312,N_14142,N_11077);
or U18313 (N_18313,N_12118,N_12679);
nand U18314 (N_18314,N_11324,N_14165);
and U18315 (N_18315,N_14855,N_10076);
and U18316 (N_18316,N_11965,N_12603);
nand U18317 (N_18317,N_13791,N_12706);
or U18318 (N_18318,N_14559,N_13826);
nor U18319 (N_18319,N_12044,N_14968);
xnor U18320 (N_18320,N_12916,N_10817);
or U18321 (N_18321,N_12633,N_11235);
or U18322 (N_18322,N_13461,N_13348);
nand U18323 (N_18323,N_10700,N_10440);
xnor U18324 (N_18324,N_12530,N_10900);
and U18325 (N_18325,N_11595,N_12498);
and U18326 (N_18326,N_13393,N_10450);
nand U18327 (N_18327,N_14181,N_12398);
or U18328 (N_18328,N_13273,N_10968);
nor U18329 (N_18329,N_11111,N_14554);
or U18330 (N_18330,N_10138,N_14282);
nand U18331 (N_18331,N_11082,N_11214);
or U18332 (N_18332,N_11377,N_11317);
nand U18333 (N_18333,N_13993,N_14959);
or U18334 (N_18334,N_13988,N_13554);
nand U18335 (N_18335,N_14424,N_10352);
nor U18336 (N_18336,N_13292,N_13346);
nand U18337 (N_18337,N_10118,N_13122);
nor U18338 (N_18338,N_13934,N_13207);
nor U18339 (N_18339,N_12163,N_10015);
xnor U18340 (N_18340,N_14529,N_14945);
and U18341 (N_18341,N_14690,N_10664);
or U18342 (N_18342,N_10014,N_12626);
or U18343 (N_18343,N_11984,N_11019);
and U18344 (N_18344,N_12517,N_10012);
or U18345 (N_18345,N_13483,N_13886);
xnor U18346 (N_18346,N_14871,N_11679);
nand U18347 (N_18347,N_11894,N_14693);
xnor U18348 (N_18348,N_11702,N_11131);
and U18349 (N_18349,N_10456,N_11487);
and U18350 (N_18350,N_12620,N_11087);
or U18351 (N_18351,N_12583,N_12271);
nor U18352 (N_18352,N_13211,N_11354);
xor U18353 (N_18353,N_14311,N_11118);
nand U18354 (N_18354,N_13515,N_11808);
nor U18355 (N_18355,N_10695,N_12823);
nor U18356 (N_18356,N_12699,N_12164);
nand U18357 (N_18357,N_12143,N_14820);
or U18358 (N_18358,N_12962,N_14014);
xor U18359 (N_18359,N_10096,N_10988);
nand U18360 (N_18360,N_13911,N_14325);
or U18361 (N_18361,N_14271,N_10636);
nor U18362 (N_18362,N_10927,N_11062);
nand U18363 (N_18363,N_13705,N_14817);
xnor U18364 (N_18364,N_11336,N_13807);
xnor U18365 (N_18365,N_14382,N_11207);
and U18366 (N_18366,N_11359,N_12709);
or U18367 (N_18367,N_12363,N_14461);
nand U18368 (N_18368,N_10411,N_11759);
or U18369 (N_18369,N_12422,N_11390);
nand U18370 (N_18370,N_11953,N_13394);
nand U18371 (N_18371,N_14588,N_12150);
xnor U18372 (N_18372,N_14556,N_11520);
nand U18373 (N_18373,N_13005,N_10721);
and U18374 (N_18374,N_10876,N_11551);
nor U18375 (N_18375,N_11870,N_12340);
and U18376 (N_18376,N_14426,N_10163);
nor U18377 (N_18377,N_12731,N_10162);
nor U18378 (N_18378,N_12528,N_10124);
nor U18379 (N_18379,N_14127,N_10450);
nor U18380 (N_18380,N_12993,N_14045);
nand U18381 (N_18381,N_11693,N_12693);
nand U18382 (N_18382,N_11688,N_14114);
xor U18383 (N_18383,N_13215,N_14651);
nand U18384 (N_18384,N_11103,N_12114);
nor U18385 (N_18385,N_13094,N_12810);
nand U18386 (N_18386,N_12412,N_14049);
nor U18387 (N_18387,N_12521,N_12995);
and U18388 (N_18388,N_12517,N_13065);
or U18389 (N_18389,N_13472,N_10994);
or U18390 (N_18390,N_11348,N_10775);
and U18391 (N_18391,N_11949,N_11048);
nand U18392 (N_18392,N_12000,N_13247);
nor U18393 (N_18393,N_10601,N_13658);
and U18394 (N_18394,N_10952,N_14395);
nand U18395 (N_18395,N_10648,N_10719);
and U18396 (N_18396,N_10815,N_13826);
and U18397 (N_18397,N_14641,N_12793);
nand U18398 (N_18398,N_14544,N_10224);
nor U18399 (N_18399,N_13897,N_13221);
and U18400 (N_18400,N_11828,N_11498);
nor U18401 (N_18401,N_13763,N_12155);
nand U18402 (N_18402,N_14255,N_13386);
or U18403 (N_18403,N_11069,N_11950);
nand U18404 (N_18404,N_12869,N_14097);
nor U18405 (N_18405,N_13593,N_14360);
nor U18406 (N_18406,N_13758,N_11521);
or U18407 (N_18407,N_13729,N_14876);
or U18408 (N_18408,N_13998,N_14488);
nand U18409 (N_18409,N_14037,N_12794);
nand U18410 (N_18410,N_10009,N_10611);
and U18411 (N_18411,N_11509,N_11160);
nor U18412 (N_18412,N_13043,N_13567);
nand U18413 (N_18413,N_13792,N_11400);
nand U18414 (N_18414,N_12895,N_12819);
and U18415 (N_18415,N_11199,N_14471);
nand U18416 (N_18416,N_11569,N_11861);
xnor U18417 (N_18417,N_10093,N_12028);
nand U18418 (N_18418,N_11823,N_12934);
and U18419 (N_18419,N_11894,N_11462);
or U18420 (N_18420,N_10745,N_13933);
nand U18421 (N_18421,N_12829,N_13186);
nor U18422 (N_18422,N_10456,N_11802);
nor U18423 (N_18423,N_12094,N_11779);
nand U18424 (N_18424,N_10689,N_13808);
nor U18425 (N_18425,N_11493,N_11491);
and U18426 (N_18426,N_13903,N_13643);
xnor U18427 (N_18427,N_14281,N_10601);
nor U18428 (N_18428,N_11507,N_10702);
nand U18429 (N_18429,N_14240,N_12640);
or U18430 (N_18430,N_13950,N_10528);
and U18431 (N_18431,N_10960,N_14317);
nor U18432 (N_18432,N_10593,N_11555);
xnor U18433 (N_18433,N_12043,N_13020);
or U18434 (N_18434,N_12900,N_14896);
nor U18435 (N_18435,N_12633,N_12351);
or U18436 (N_18436,N_10966,N_12260);
xor U18437 (N_18437,N_10512,N_14861);
and U18438 (N_18438,N_11354,N_10228);
xor U18439 (N_18439,N_10881,N_10291);
xnor U18440 (N_18440,N_12534,N_10855);
and U18441 (N_18441,N_13298,N_10741);
nor U18442 (N_18442,N_11911,N_12022);
nor U18443 (N_18443,N_12837,N_12532);
nand U18444 (N_18444,N_13604,N_13104);
and U18445 (N_18445,N_11076,N_12480);
nor U18446 (N_18446,N_10001,N_11286);
nand U18447 (N_18447,N_12784,N_11716);
xnor U18448 (N_18448,N_14561,N_13607);
and U18449 (N_18449,N_13976,N_13570);
nor U18450 (N_18450,N_12184,N_14013);
and U18451 (N_18451,N_13517,N_14018);
or U18452 (N_18452,N_14553,N_13394);
and U18453 (N_18453,N_10092,N_12123);
and U18454 (N_18454,N_11049,N_11490);
nor U18455 (N_18455,N_12032,N_13744);
nor U18456 (N_18456,N_14676,N_11699);
nand U18457 (N_18457,N_11577,N_13124);
nand U18458 (N_18458,N_12236,N_11542);
or U18459 (N_18459,N_11758,N_12454);
nand U18460 (N_18460,N_11326,N_13726);
nor U18461 (N_18461,N_11345,N_12299);
nand U18462 (N_18462,N_14867,N_11909);
xnor U18463 (N_18463,N_10673,N_10511);
or U18464 (N_18464,N_13833,N_11278);
xor U18465 (N_18465,N_14911,N_11263);
nand U18466 (N_18466,N_12746,N_14301);
and U18467 (N_18467,N_14585,N_11990);
and U18468 (N_18468,N_10430,N_13449);
nand U18469 (N_18469,N_12256,N_10526);
and U18470 (N_18470,N_12335,N_14498);
or U18471 (N_18471,N_10422,N_13285);
nand U18472 (N_18472,N_14811,N_11105);
or U18473 (N_18473,N_10121,N_10186);
and U18474 (N_18474,N_12950,N_10456);
nor U18475 (N_18475,N_14598,N_14382);
and U18476 (N_18476,N_13295,N_10090);
or U18477 (N_18477,N_11062,N_13136);
nor U18478 (N_18478,N_13768,N_10397);
and U18479 (N_18479,N_13240,N_12165);
nand U18480 (N_18480,N_13639,N_14451);
nor U18481 (N_18481,N_10659,N_11036);
or U18482 (N_18482,N_11137,N_13462);
or U18483 (N_18483,N_14924,N_12528);
and U18484 (N_18484,N_11121,N_11581);
nor U18485 (N_18485,N_14129,N_13242);
nand U18486 (N_18486,N_10077,N_14038);
or U18487 (N_18487,N_11041,N_14467);
nor U18488 (N_18488,N_14175,N_12826);
or U18489 (N_18489,N_12523,N_10994);
xnor U18490 (N_18490,N_11366,N_13336);
and U18491 (N_18491,N_14263,N_10543);
nand U18492 (N_18492,N_11941,N_12401);
or U18493 (N_18493,N_14791,N_10824);
xnor U18494 (N_18494,N_10858,N_10996);
nor U18495 (N_18495,N_12945,N_12701);
and U18496 (N_18496,N_13628,N_11943);
or U18497 (N_18497,N_10274,N_12324);
nor U18498 (N_18498,N_11338,N_12883);
nor U18499 (N_18499,N_14437,N_11400);
or U18500 (N_18500,N_13572,N_12741);
and U18501 (N_18501,N_13779,N_14971);
or U18502 (N_18502,N_11473,N_14102);
and U18503 (N_18503,N_13208,N_11013);
xor U18504 (N_18504,N_13231,N_13238);
or U18505 (N_18505,N_13687,N_14001);
nor U18506 (N_18506,N_12897,N_12060);
nand U18507 (N_18507,N_11593,N_10308);
nand U18508 (N_18508,N_10711,N_12546);
xnor U18509 (N_18509,N_10266,N_14806);
or U18510 (N_18510,N_13194,N_10582);
and U18511 (N_18511,N_13403,N_10692);
and U18512 (N_18512,N_12204,N_11832);
nand U18513 (N_18513,N_10500,N_14436);
and U18514 (N_18514,N_12133,N_12725);
or U18515 (N_18515,N_11281,N_11145);
or U18516 (N_18516,N_13841,N_14064);
xor U18517 (N_18517,N_12055,N_12335);
nand U18518 (N_18518,N_11692,N_13170);
nor U18519 (N_18519,N_12944,N_13941);
and U18520 (N_18520,N_10160,N_12098);
nor U18521 (N_18521,N_12219,N_14032);
and U18522 (N_18522,N_11062,N_14388);
nor U18523 (N_18523,N_14932,N_13662);
nand U18524 (N_18524,N_12556,N_10184);
nand U18525 (N_18525,N_12149,N_13479);
or U18526 (N_18526,N_11327,N_13314);
nand U18527 (N_18527,N_11436,N_11565);
nor U18528 (N_18528,N_11324,N_12518);
nor U18529 (N_18529,N_12244,N_10757);
or U18530 (N_18530,N_12778,N_13309);
and U18531 (N_18531,N_10419,N_11750);
nor U18532 (N_18532,N_13473,N_14579);
nand U18533 (N_18533,N_10857,N_12582);
nor U18534 (N_18534,N_12837,N_14780);
and U18535 (N_18535,N_13870,N_11286);
nor U18536 (N_18536,N_14474,N_11422);
or U18537 (N_18537,N_13261,N_14079);
xnor U18538 (N_18538,N_12638,N_11658);
nand U18539 (N_18539,N_11498,N_10993);
nor U18540 (N_18540,N_11036,N_13380);
or U18541 (N_18541,N_10843,N_10985);
nand U18542 (N_18542,N_10218,N_12119);
nor U18543 (N_18543,N_11682,N_14480);
nand U18544 (N_18544,N_12042,N_10904);
and U18545 (N_18545,N_13326,N_12040);
xor U18546 (N_18546,N_10514,N_11656);
and U18547 (N_18547,N_14710,N_12262);
nand U18548 (N_18548,N_10900,N_13978);
and U18549 (N_18549,N_14099,N_13458);
and U18550 (N_18550,N_11840,N_11496);
or U18551 (N_18551,N_10266,N_12746);
and U18552 (N_18552,N_14680,N_10920);
nor U18553 (N_18553,N_10014,N_13759);
nand U18554 (N_18554,N_12203,N_11654);
or U18555 (N_18555,N_14007,N_13610);
xor U18556 (N_18556,N_14496,N_12662);
nand U18557 (N_18557,N_12255,N_12062);
nand U18558 (N_18558,N_11982,N_11302);
xor U18559 (N_18559,N_13543,N_10362);
and U18560 (N_18560,N_12963,N_12413);
nand U18561 (N_18561,N_12372,N_12716);
and U18562 (N_18562,N_12991,N_12885);
or U18563 (N_18563,N_13443,N_13081);
or U18564 (N_18564,N_13315,N_14008);
nand U18565 (N_18565,N_12087,N_14245);
nor U18566 (N_18566,N_12794,N_11547);
or U18567 (N_18567,N_10570,N_13988);
nor U18568 (N_18568,N_12552,N_10276);
nor U18569 (N_18569,N_11793,N_11116);
nand U18570 (N_18570,N_10575,N_11543);
and U18571 (N_18571,N_11886,N_10775);
nand U18572 (N_18572,N_11467,N_10798);
nand U18573 (N_18573,N_14751,N_13959);
nor U18574 (N_18574,N_13323,N_12787);
or U18575 (N_18575,N_14276,N_11581);
and U18576 (N_18576,N_11663,N_10843);
and U18577 (N_18577,N_13018,N_11290);
and U18578 (N_18578,N_11813,N_11261);
and U18579 (N_18579,N_11398,N_10127);
or U18580 (N_18580,N_11653,N_12618);
nand U18581 (N_18581,N_12263,N_12966);
nand U18582 (N_18582,N_12911,N_13954);
nand U18583 (N_18583,N_11592,N_10207);
xor U18584 (N_18584,N_10344,N_11203);
and U18585 (N_18585,N_11689,N_13615);
nor U18586 (N_18586,N_11936,N_13024);
or U18587 (N_18587,N_14356,N_14091);
and U18588 (N_18588,N_10398,N_13663);
xnor U18589 (N_18589,N_14875,N_12551);
nand U18590 (N_18590,N_11902,N_12400);
and U18591 (N_18591,N_10700,N_12349);
nor U18592 (N_18592,N_12478,N_11369);
and U18593 (N_18593,N_14363,N_14715);
and U18594 (N_18594,N_14204,N_12216);
nor U18595 (N_18595,N_11967,N_11993);
nand U18596 (N_18596,N_11722,N_13091);
and U18597 (N_18597,N_11668,N_11242);
nand U18598 (N_18598,N_13695,N_13474);
nand U18599 (N_18599,N_14262,N_10462);
or U18600 (N_18600,N_12180,N_10959);
nand U18601 (N_18601,N_10376,N_14485);
xor U18602 (N_18602,N_11861,N_14261);
or U18603 (N_18603,N_13127,N_14418);
xor U18604 (N_18604,N_11955,N_12197);
and U18605 (N_18605,N_10325,N_10092);
and U18606 (N_18606,N_12171,N_12560);
nor U18607 (N_18607,N_11817,N_11031);
or U18608 (N_18608,N_14942,N_14477);
nor U18609 (N_18609,N_10172,N_13876);
xnor U18610 (N_18610,N_14918,N_11666);
nor U18611 (N_18611,N_12044,N_11896);
nand U18612 (N_18612,N_13957,N_12179);
nand U18613 (N_18613,N_14950,N_14406);
nand U18614 (N_18614,N_14132,N_10784);
nor U18615 (N_18615,N_10532,N_10067);
or U18616 (N_18616,N_14282,N_14506);
or U18617 (N_18617,N_12475,N_10637);
nor U18618 (N_18618,N_14672,N_13779);
or U18619 (N_18619,N_10746,N_12041);
and U18620 (N_18620,N_14141,N_10620);
or U18621 (N_18621,N_12135,N_11540);
xor U18622 (N_18622,N_14338,N_12528);
and U18623 (N_18623,N_14149,N_10568);
nand U18624 (N_18624,N_11580,N_14648);
nor U18625 (N_18625,N_12214,N_11582);
or U18626 (N_18626,N_11728,N_13414);
and U18627 (N_18627,N_14999,N_12044);
nand U18628 (N_18628,N_13914,N_11694);
or U18629 (N_18629,N_10593,N_14326);
nand U18630 (N_18630,N_14339,N_10594);
xnor U18631 (N_18631,N_12801,N_10440);
nand U18632 (N_18632,N_10624,N_14652);
and U18633 (N_18633,N_11925,N_14290);
and U18634 (N_18634,N_14012,N_12043);
nand U18635 (N_18635,N_13172,N_10005);
xnor U18636 (N_18636,N_13998,N_12953);
and U18637 (N_18637,N_13338,N_12064);
or U18638 (N_18638,N_13334,N_12422);
xor U18639 (N_18639,N_14258,N_11874);
xor U18640 (N_18640,N_14728,N_11997);
and U18641 (N_18641,N_14651,N_13167);
or U18642 (N_18642,N_12902,N_10188);
and U18643 (N_18643,N_14949,N_13026);
and U18644 (N_18644,N_12795,N_13885);
nand U18645 (N_18645,N_10623,N_14333);
and U18646 (N_18646,N_10683,N_11596);
nor U18647 (N_18647,N_13204,N_14195);
nor U18648 (N_18648,N_14351,N_11004);
nor U18649 (N_18649,N_10011,N_13154);
and U18650 (N_18650,N_13081,N_13591);
nor U18651 (N_18651,N_13807,N_10544);
nand U18652 (N_18652,N_13694,N_11363);
nor U18653 (N_18653,N_14994,N_14973);
and U18654 (N_18654,N_14145,N_10603);
and U18655 (N_18655,N_13466,N_11922);
and U18656 (N_18656,N_12860,N_10350);
nor U18657 (N_18657,N_14126,N_11699);
or U18658 (N_18658,N_14364,N_14394);
or U18659 (N_18659,N_12344,N_12254);
nand U18660 (N_18660,N_11694,N_14392);
nor U18661 (N_18661,N_12661,N_14020);
and U18662 (N_18662,N_13110,N_11892);
nand U18663 (N_18663,N_11940,N_14161);
and U18664 (N_18664,N_11905,N_12717);
or U18665 (N_18665,N_14372,N_11273);
nor U18666 (N_18666,N_12481,N_12367);
nor U18667 (N_18667,N_14406,N_14706);
xnor U18668 (N_18668,N_11324,N_13774);
or U18669 (N_18669,N_13800,N_11801);
nor U18670 (N_18670,N_14935,N_12914);
or U18671 (N_18671,N_14686,N_14512);
or U18672 (N_18672,N_13351,N_13942);
nor U18673 (N_18673,N_11425,N_12131);
or U18674 (N_18674,N_14503,N_10658);
and U18675 (N_18675,N_14905,N_14848);
or U18676 (N_18676,N_11271,N_14543);
or U18677 (N_18677,N_14737,N_13608);
or U18678 (N_18678,N_10250,N_11184);
and U18679 (N_18679,N_14703,N_12024);
nand U18680 (N_18680,N_14421,N_12114);
or U18681 (N_18681,N_14957,N_10791);
nor U18682 (N_18682,N_13755,N_14823);
and U18683 (N_18683,N_11545,N_12919);
nand U18684 (N_18684,N_12611,N_12063);
and U18685 (N_18685,N_12797,N_12267);
nor U18686 (N_18686,N_14094,N_10749);
or U18687 (N_18687,N_11925,N_11515);
or U18688 (N_18688,N_11323,N_13631);
or U18689 (N_18689,N_14866,N_14377);
or U18690 (N_18690,N_13601,N_13881);
nand U18691 (N_18691,N_12187,N_14684);
nor U18692 (N_18692,N_12998,N_14757);
nor U18693 (N_18693,N_10502,N_11084);
or U18694 (N_18694,N_11066,N_14410);
nand U18695 (N_18695,N_10407,N_14031);
and U18696 (N_18696,N_11076,N_13562);
nand U18697 (N_18697,N_14654,N_11021);
nor U18698 (N_18698,N_12137,N_12874);
and U18699 (N_18699,N_10428,N_13343);
and U18700 (N_18700,N_14873,N_14488);
nand U18701 (N_18701,N_12762,N_10703);
or U18702 (N_18702,N_13977,N_11651);
and U18703 (N_18703,N_11402,N_10828);
nor U18704 (N_18704,N_12433,N_12374);
or U18705 (N_18705,N_12026,N_12136);
and U18706 (N_18706,N_10350,N_11970);
or U18707 (N_18707,N_10244,N_13389);
nand U18708 (N_18708,N_10175,N_10694);
nand U18709 (N_18709,N_14412,N_14037);
or U18710 (N_18710,N_14871,N_12083);
nand U18711 (N_18711,N_13964,N_10948);
xnor U18712 (N_18712,N_11181,N_11572);
xnor U18713 (N_18713,N_13853,N_11705);
and U18714 (N_18714,N_13601,N_10603);
or U18715 (N_18715,N_10195,N_11522);
nand U18716 (N_18716,N_14106,N_13083);
nand U18717 (N_18717,N_14481,N_11851);
and U18718 (N_18718,N_12792,N_10225);
or U18719 (N_18719,N_13085,N_13394);
xnor U18720 (N_18720,N_13927,N_10776);
nand U18721 (N_18721,N_14626,N_12737);
and U18722 (N_18722,N_12758,N_14440);
xnor U18723 (N_18723,N_14330,N_14008);
nand U18724 (N_18724,N_13966,N_11039);
or U18725 (N_18725,N_11315,N_10262);
nor U18726 (N_18726,N_13135,N_12940);
or U18727 (N_18727,N_11668,N_12674);
or U18728 (N_18728,N_10102,N_12616);
and U18729 (N_18729,N_10253,N_11652);
nand U18730 (N_18730,N_14026,N_11930);
nor U18731 (N_18731,N_13493,N_10641);
or U18732 (N_18732,N_10466,N_10352);
nor U18733 (N_18733,N_12298,N_11670);
nand U18734 (N_18734,N_13144,N_10476);
and U18735 (N_18735,N_13545,N_10353);
and U18736 (N_18736,N_11414,N_14602);
or U18737 (N_18737,N_14745,N_11139);
nand U18738 (N_18738,N_13197,N_13315);
xnor U18739 (N_18739,N_12409,N_14690);
nand U18740 (N_18740,N_11253,N_12448);
xor U18741 (N_18741,N_12313,N_14672);
and U18742 (N_18742,N_14847,N_13887);
or U18743 (N_18743,N_11998,N_13527);
nor U18744 (N_18744,N_10313,N_13148);
nand U18745 (N_18745,N_11621,N_10638);
nor U18746 (N_18746,N_13147,N_13111);
nand U18747 (N_18747,N_14419,N_13056);
nor U18748 (N_18748,N_13378,N_13983);
xor U18749 (N_18749,N_14221,N_10290);
and U18750 (N_18750,N_14454,N_12159);
or U18751 (N_18751,N_10310,N_14606);
nor U18752 (N_18752,N_14574,N_11815);
or U18753 (N_18753,N_13418,N_11414);
or U18754 (N_18754,N_10341,N_10254);
nor U18755 (N_18755,N_14203,N_13307);
nor U18756 (N_18756,N_13422,N_13238);
nand U18757 (N_18757,N_12966,N_10058);
or U18758 (N_18758,N_12107,N_12386);
nor U18759 (N_18759,N_14212,N_11570);
or U18760 (N_18760,N_12880,N_14624);
nor U18761 (N_18761,N_14719,N_11888);
or U18762 (N_18762,N_12086,N_10139);
nand U18763 (N_18763,N_10525,N_12224);
or U18764 (N_18764,N_13190,N_11515);
and U18765 (N_18765,N_14689,N_11069);
nor U18766 (N_18766,N_13246,N_10842);
nand U18767 (N_18767,N_10157,N_14944);
xnor U18768 (N_18768,N_10058,N_10064);
nand U18769 (N_18769,N_14456,N_11730);
nor U18770 (N_18770,N_13544,N_14366);
nor U18771 (N_18771,N_13549,N_10852);
and U18772 (N_18772,N_13507,N_11753);
nor U18773 (N_18773,N_10705,N_13010);
and U18774 (N_18774,N_10121,N_10659);
nand U18775 (N_18775,N_14618,N_10726);
and U18776 (N_18776,N_10376,N_11864);
nor U18777 (N_18777,N_14489,N_13833);
nand U18778 (N_18778,N_13198,N_10755);
or U18779 (N_18779,N_13071,N_14322);
nor U18780 (N_18780,N_10274,N_12813);
nor U18781 (N_18781,N_10028,N_14757);
and U18782 (N_18782,N_12093,N_10055);
or U18783 (N_18783,N_12113,N_14521);
or U18784 (N_18784,N_14693,N_10375);
nor U18785 (N_18785,N_14318,N_14786);
nor U18786 (N_18786,N_11507,N_10777);
or U18787 (N_18787,N_13679,N_10870);
and U18788 (N_18788,N_11497,N_12487);
nand U18789 (N_18789,N_12062,N_12478);
xor U18790 (N_18790,N_11907,N_11216);
nand U18791 (N_18791,N_14530,N_14012);
nor U18792 (N_18792,N_12027,N_14213);
nand U18793 (N_18793,N_11965,N_10016);
nor U18794 (N_18794,N_12053,N_11681);
and U18795 (N_18795,N_14656,N_12875);
nor U18796 (N_18796,N_11974,N_14800);
and U18797 (N_18797,N_12024,N_11905);
and U18798 (N_18798,N_12185,N_12816);
and U18799 (N_18799,N_11321,N_10533);
nor U18800 (N_18800,N_13845,N_12730);
nand U18801 (N_18801,N_12715,N_12767);
xor U18802 (N_18802,N_13733,N_10261);
nand U18803 (N_18803,N_11943,N_13270);
or U18804 (N_18804,N_14262,N_11917);
or U18805 (N_18805,N_10923,N_14240);
or U18806 (N_18806,N_12556,N_10315);
nor U18807 (N_18807,N_11644,N_10912);
or U18808 (N_18808,N_10714,N_12059);
nand U18809 (N_18809,N_11114,N_12977);
and U18810 (N_18810,N_11498,N_13498);
or U18811 (N_18811,N_10535,N_10368);
and U18812 (N_18812,N_13732,N_12456);
and U18813 (N_18813,N_10825,N_10567);
nand U18814 (N_18814,N_11023,N_11130);
xnor U18815 (N_18815,N_14636,N_13152);
or U18816 (N_18816,N_14688,N_12862);
or U18817 (N_18817,N_12869,N_14950);
nand U18818 (N_18818,N_12379,N_13037);
nand U18819 (N_18819,N_10152,N_14696);
nand U18820 (N_18820,N_10029,N_14900);
nor U18821 (N_18821,N_10177,N_13701);
nand U18822 (N_18822,N_12667,N_10840);
or U18823 (N_18823,N_13059,N_12956);
nand U18824 (N_18824,N_14391,N_13496);
or U18825 (N_18825,N_13224,N_13059);
nor U18826 (N_18826,N_13395,N_12054);
or U18827 (N_18827,N_14121,N_13233);
or U18828 (N_18828,N_10502,N_12794);
or U18829 (N_18829,N_10091,N_12433);
xnor U18830 (N_18830,N_10852,N_13113);
nor U18831 (N_18831,N_12924,N_11410);
nand U18832 (N_18832,N_13171,N_11628);
xor U18833 (N_18833,N_11242,N_13916);
xor U18834 (N_18834,N_12511,N_12835);
nand U18835 (N_18835,N_11939,N_10672);
and U18836 (N_18836,N_11103,N_10808);
and U18837 (N_18837,N_11865,N_13049);
nand U18838 (N_18838,N_10367,N_14459);
nor U18839 (N_18839,N_12079,N_10127);
nand U18840 (N_18840,N_11406,N_11176);
and U18841 (N_18841,N_14968,N_14122);
and U18842 (N_18842,N_14774,N_12009);
nor U18843 (N_18843,N_10557,N_10120);
nand U18844 (N_18844,N_12254,N_12695);
nand U18845 (N_18845,N_12010,N_12443);
and U18846 (N_18846,N_13582,N_12554);
and U18847 (N_18847,N_14305,N_10855);
xnor U18848 (N_18848,N_10641,N_14878);
and U18849 (N_18849,N_12390,N_10997);
xor U18850 (N_18850,N_10699,N_11041);
nor U18851 (N_18851,N_14882,N_14080);
or U18852 (N_18852,N_10900,N_10212);
nand U18853 (N_18853,N_11838,N_11653);
and U18854 (N_18854,N_13062,N_13970);
xnor U18855 (N_18855,N_12169,N_13755);
or U18856 (N_18856,N_14893,N_13691);
nor U18857 (N_18857,N_13480,N_11343);
nor U18858 (N_18858,N_12830,N_14784);
and U18859 (N_18859,N_11676,N_11467);
or U18860 (N_18860,N_11094,N_11212);
xor U18861 (N_18861,N_13583,N_14955);
nand U18862 (N_18862,N_12207,N_14516);
nand U18863 (N_18863,N_13115,N_13908);
or U18864 (N_18864,N_14926,N_10976);
nand U18865 (N_18865,N_11453,N_10891);
nand U18866 (N_18866,N_12350,N_13663);
nor U18867 (N_18867,N_13475,N_14075);
nor U18868 (N_18868,N_11534,N_11282);
nor U18869 (N_18869,N_10181,N_11735);
nor U18870 (N_18870,N_13028,N_12010);
xnor U18871 (N_18871,N_10349,N_10316);
and U18872 (N_18872,N_11158,N_11730);
nor U18873 (N_18873,N_12394,N_12089);
nor U18874 (N_18874,N_13691,N_14405);
or U18875 (N_18875,N_10322,N_13461);
xnor U18876 (N_18876,N_12119,N_13956);
nand U18877 (N_18877,N_12654,N_12365);
nor U18878 (N_18878,N_11727,N_12688);
or U18879 (N_18879,N_12472,N_11947);
and U18880 (N_18880,N_10515,N_14841);
and U18881 (N_18881,N_14647,N_11868);
nor U18882 (N_18882,N_10994,N_13958);
or U18883 (N_18883,N_10193,N_11718);
and U18884 (N_18884,N_12843,N_13229);
nor U18885 (N_18885,N_10116,N_14959);
nor U18886 (N_18886,N_11713,N_11523);
and U18887 (N_18887,N_14362,N_13254);
nor U18888 (N_18888,N_12371,N_10224);
nor U18889 (N_18889,N_10141,N_14044);
or U18890 (N_18890,N_12675,N_13177);
or U18891 (N_18891,N_13765,N_14731);
xor U18892 (N_18892,N_14550,N_12260);
nor U18893 (N_18893,N_12655,N_14036);
nand U18894 (N_18894,N_14097,N_13502);
and U18895 (N_18895,N_14578,N_10084);
or U18896 (N_18896,N_14731,N_10575);
or U18897 (N_18897,N_14707,N_12415);
nor U18898 (N_18898,N_10825,N_14515);
and U18899 (N_18899,N_10145,N_12403);
or U18900 (N_18900,N_10027,N_12992);
or U18901 (N_18901,N_14650,N_12685);
or U18902 (N_18902,N_14171,N_11305);
nand U18903 (N_18903,N_11060,N_10448);
nor U18904 (N_18904,N_11739,N_12996);
or U18905 (N_18905,N_12595,N_12984);
and U18906 (N_18906,N_13254,N_10610);
and U18907 (N_18907,N_11878,N_12534);
nor U18908 (N_18908,N_10990,N_13740);
xnor U18909 (N_18909,N_14630,N_13005);
nor U18910 (N_18910,N_11969,N_12122);
nand U18911 (N_18911,N_10107,N_10301);
nor U18912 (N_18912,N_14214,N_11882);
nand U18913 (N_18913,N_14461,N_12329);
nor U18914 (N_18914,N_11630,N_10396);
nor U18915 (N_18915,N_12885,N_12660);
nor U18916 (N_18916,N_12458,N_14151);
nor U18917 (N_18917,N_11582,N_12966);
or U18918 (N_18918,N_10290,N_11811);
or U18919 (N_18919,N_12279,N_11812);
and U18920 (N_18920,N_12578,N_12564);
nor U18921 (N_18921,N_11872,N_11907);
nor U18922 (N_18922,N_14160,N_10259);
or U18923 (N_18923,N_11992,N_13877);
nor U18924 (N_18924,N_12094,N_11311);
xor U18925 (N_18925,N_14821,N_11585);
nor U18926 (N_18926,N_12575,N_14664);
nor U18927 (N_18927,N_14058,N_12704);
nand U18928 (N_18928,N_12787,N_10940);
and U18929 (N_18929,N_14005,N_13011);
or U18930 (N_18930,N_11823,N_13252);
xor U18931 (N_18931,N_14149,N_13651);
nand U18932 (N_18932,N_11760,N_14592);
nor U18933 (N_18933,N_11516,N_12372);
or U18934 (N_18934,N_13913,N_12327);
xor U18935 (N_18935,N_12886,N_14902);
nor U18936 (N_18936,N_10049,N_11998);
nand U18937 (N_18937,N_13897,N_10662);
or U18938 (N_18938,N_14053,N_13880);
nor U18939 (N_18939,N_13801,N_10335);
nor U18940 (N_18940,N_10461,N_14841);
nor U18941 (N_18941,N_14998,N_10205);
xor U18942 (N_18942,N_12539,N_14387);
and U18943 (N_18943,N_11617,N_14021);
nand U18944 (N_18944,N_12913,N_11348);
nand U18945 (N_18945,N_10347,N_12212);
nand U18946 (N_18946,N_12236,N_12562);
and U18947 (N_18947,N_10589,N_12430);
or U18948 (N_18948,N_10936,N_10820);
nand U18949 (N_18949,N_13295,N_10342);
nor U18950 (N_18950,N_12985,N_13561);
or U18951 (N_18951,N_12086,N_11551);
and U18952 (N_18952,N_12679,N_12860);
or U18953 (N_18953,N_11615,N_11900);
or U18954 (N_18954,N_12859,N_14428);
and U18955 (N_18955,N_14219,N_14845);
xnor U18956 (N_18956,N_10184,N_11057);
nor U18957 (N_18957,N_14832,N_10760);
nand U18958 (N_18958,N_11457,N_12814);
or U18959 (N_18959,N_11793,N_14409);
nand U18960 (N_18960,N_14816,N_11568);
or U18961 (N_18961,N_11133,N_11703);
nand U18962 (N_18962,N_10139,N_11059);
and U18963 (N_18963,N_13508,N_14357);
or U18964 (N_18964,N_12250,N_13360);
xnor U18965 (N_18965,N_12323,N_12449);
nor U18966 (N_18966,N_13344,N_14455);
and U18967 (N_18967,N_13167,N_14231);
or U18968 (N_18968,N_14685,N_14319);
nand U18969 (N_18969,N_13727,N_10901);
nand U18970 (N_18970,N_14604,N_10891);
nand U18971 (N_18971,N_12220,N_13858);
or U18972 (N_18972,N_13005,N_13197);
nor U18973 (N_18973,N_10150,N_14553);
nor U18974 (N_18974,N_13965,N_14724);
nand U18975 (N_18975,N_14327,N_13123);
nand U18976 (N_18976,N_12897,N_13772);
nor U18977 (N_18977,N_11575,N_14670);
or U18978 (N_18978,N_14845,N_12066);
nor U18979 (N_18979,N_13777,N_14746);
nand U18980 (N_18980,N_12340,N_11096);
and U18981 (N_18981,N_12770,N_11097);
or U18982 (N_18982,N_11057,N_11294);
nor U18983 (N_18983,N_13141,N_11766);
and U18984 (N_18984,N_10887,N_10337);
or U18985 (N_18985,N_11720,N_13628);
xor U18986 (N_18986,N_13016,N_10453);
or U18987 (N_18987,N_12345,N_10457);
nand U18988 (N_18988,N_10868,N_10431);
nand U18989 (N_18989,N_11872,N_11838);
xor U18990 (N_18990,N_12904,N_13931);
nor U18991 (N_18991,N_12285,N_12178);
nor U18992 (N_18992,N_13925,N_13415);
or U18993 (N_18993,N_10917,N_11625);
nor U18994 (N_18994,N_14055,N_13913);
or U18995 (N_18995,N_14444,N_14969);
nor U18996 (N_18996,N_10814,N_12774);
nor U18997 (N_18997,N_11147,N_10726);
or U18998 (N_18998,N_12867,N_13924);
nand U18999 (N_18999,N_13307,N_13372);
nor U19000 (N_19000,N_14984,N_13370);
or U19001 (N_19001,N_14908,N_14657);
nor U19002 (N_19002,N_12863,N_13501);
and U19003 (N_19003,N_13025,N_14593);
and U19004 (N_19004,N_10691,N_12825);
and U19005 (N_19005,N_12723,N_14108);
nor U19006 (N_19006,N_14099,N_14026);
nor U19007 (N_19007,N_12095,N_10954);
and U19008 (N_19008,N_10713,N_11434);
xnor U19009 (N_19009,N_10226,N_10966);
or U19010 (N_19010,N_12239,N_11914);
xor U19011 (N_19011,N_13172,N_10700);
xor U19012 (N_19012,N_13466,N_10737);
nand U19013 (N_19013,N_14468,N_11945);
nor U19014 (N_19014,N_12918,N_14160);
or U19015 (N_19015,N_12189,N_10910);
and U19016 (N_19016,N_14552,N_13573);
xor U19017 (N_19017,N_12137,N_14297);
and U19018 (N_19018,N_14632,N_13201);
nor U19019 (N_19019,N_14662,N_10316);
nor U19020 (N_19020,N_11008,N_12553);
nor U19021 (N_19021,N_11045,N_13310);
and U19022 (N_19022,N_13641,N_12820);
nor U19023 (N_19023,N_10641,N_12157);
nand U19024 (N_19024,N_13482,N_14940);
or U19025 (N_19025,N_14999,N_11967);
or U19026 (N_19026,N_13784,N_14443);
and U19027 (N_19027,N_14059,N_12526);
xor U19028 (N_19028,N_10711,N_10540);
nand U19029 (N_19029,N_13828,N_11385);
nand U19030 (N_19030,N_14789,N_11165);
nand U19031 (N_19031,N_12680,N_13403);
and U19032 (N_19032,N_11578,N_14254);
nor U19033 (N_19033,N_10944,N_14799);
and U19034 (N_19034,N_14460,N_10767);
and U19035 (N_19035,N_13526,N_14814);
nor U19036 (N_19036,N_13749,N_14244);
and U19037 (N_19037,N_10952,N_11081);
nand U19038 (N_19038,N_11518,N_13822);
or U19039 (N_19039,N_11446,N_11803);
nor U19040 (N_19040,N_13306,N_14376);
or U19041 (N_19041,N_14155,N_14495);
or U19042 (N_19042,N_13929,N_13942);
and U19043 (N_19043,N_14110,N_11842);
and U19044 (N_19044,N_13118,N_11023);
xor U19045 (N_19045,N_10861,N_13941);
nor U19046 (N_19046,N_12722,N_14990);
or U19047 (N_19047,N_10551,N_10695);
nand U19048 (N_19048,N_11576,N_12313);
or U19049 (N_19049,N_12701,N_10481);
xor U19050 (N_19050,N_11634,N_10938);
or U19051 (N_19051,N_11934,N_10960);
or U19052 (N_19052,N_10925,N_10240);
or U19053 (N_19053,N_14420,N_10643);
and U19054 (N_19054,N_10563,N_12883);
nor U19055 (N_19055,N_14565,N_12124);
and U19056 (N_19056,N_11674,N_11224);
nand U19057 (N_19057,N_13799,N_13795);
and U19058 (N_19058,N_13622,N_13115);
and U19059 (N_19059,N_12059,N_11331);
nor U19060 (N_19060,N_10880,N_10813);
xnor U19061 (N_19061,N_12117,N_13820);
and U19062 (N_19062,N_12027,N_13879);
and U19063 (N_19063,N_10767,N_12965);
nand U19064 (N_19064,N_13965,N_10042);
nor U19065 (N_19065,N_10048,N_13787);
nand U19066 (N_19066,N_12652,N_12228);
nand U19067 (N_19067,N_12815,N_12664);
or U19068 (N_19068,N_11897,N_12385);
or U19069 (N_19069,N_13381,N_11453);
nand U19070 (N_19070,N_11341,N_12253);
nand U19071 (N_19071,N_10065,N_11468);
nor U19072 (N_19072,N_14318,N_13485);
nand U19073 (N_19073,N_13568,N_13220);
nand U19074 (N_19074,N_13957,N_14558);
nand U19075 (N_19075,N_12332,N_13965);
and U19076 (N_19076,N_10353,N_10290);
and U19077 (N_19077,N_13355,N_12964);
and U19078 (N_19078,N_12070,N_10460);
or U19079 (N_19079,N_12838,N_11930);
nor U19080 (N_19080,N_14230,N_14034);
and U19081 (N_19081,N_14393,N_13469);
nand U19082 (N_19082,N_11421,N_14366);
nand U19083 (N_19083,N_14064,N_11109);
and U19084 (N_19084,N_10719,N_10420);
nor U19085 (N_19085,N_14201,N_13274);
nor U19086 (N_19086,N_11032,N_13370);
nand U19087 (N_19087,N_14054,N_11973);
or U19088 (N_19088,N_10863,N_12417);
nor U19089 (N_19089,N_12198,N_10144);
nor U19090 (N_19090,N_13251,N_12380);
or U19091 (N_19091,N_10678,N_12123);
nand U19092 (N_19092,N_12018,N_14606);
nand U19093 (N_19093,N_13155,N_10539);
or U19094 (N_19094,N_13854,N_12955);
nor U19095 (N_19095,N_11381,N_10815);
or U19096 (N_19096,N_12472,N_13524);
nor U19097 (N_19097,N_14739,N_11154);
xnor U19098 (N_19098,N_11065,N_12764);
and U19099 (N_19099,N_12632,N_13150);
or U19100 (N_19100,N_12401,N_14100);
or U19101 (N_19101,N_13760,N_10405);
or U19102 (N_19102,N_11774,N_10128);
nand U19103 (N_19103,N_13614,N_14768);
xor U19104 (N_19104,N_11899,N_13241);
and U19105 (N_19105,N_12800,N_11906);
or U19106 (N_19106,N_13662,N_14411);
nor U19107 (N_19107,N_13485,N_10883);
or U19108 (N_19108,N_10143,N_13111);
nand U19109 (N_19109,N_10714,N_12185);
or U19110 (N_19110,N_12769,N_11500);
or U19111 (N_19111,N_11411,N_10577);
or U19112 (N_19112,N_10029,N_11975);
and U19113 (N_19113,N_10338,N_10973);
nor U19114 (N_19114,N_10325,N_10988);
nand U19115 (N_19115,N_12178,N_13179);
nand U19116 (N_19116,N_13716,N_11922);
nor U19117 (N_19117,N_12536,N_12484);
nand U19118 (N_19118,N_10927,N_14572);
or U19119 (N_19119,N_11188,N_12855);
nor U19120 (N_19120,N_13484,N_10910);
or U19121 (N_19121,N_12551,N_11423);
and U19122 (N_19122,N_11199,N_13612);
nor U19123 (N_19123,N_14056,N_12629);
or U19124 (N_19124,N_11511,N_10353);
nand U19125 (N_19125,N_13466,N_12263);
xnor U19126 (N_19126,N_13783,N_12235);
nand U19127 (N_19127,N_10474,N_10412);
nor U19128 (N_19128,N_14136,N_14437);
nor U19129 (N_19129,N_13745,N_11492);
nor U19130 (N_19130,N_12023,N_13321);
and U19131 (N_19131,N_11585,N_11193);
nor U19132 (N_19132,N_10581,N_13676);
and U19133 (N_19133,N_11892,N_10380);
and U19134 (N_19134,N_13509,N_12556);
nor U19135 (N_19135,N_10967,N_14827);
or U19136 (N_19136,N_12732,N_12430);
nor U19137 (N_19137,N_14994,N_10803);
nand U19138 (N_19138,N_13363,N_13843);
nand U19139 (N_19139,N_10396,N_13895);
or U19140 (N_19140,N_13710,N_10765);
nor U19141 (N_19141,N_11306,N_10838);
and U19142 (N_19142,N_12850,N_10509);
xor U19143 (N_19143,N_12297,N_14924);
xnor U19144 (N_19144,N_10442,N_12742);
nor U19145 (N_19145,N_13960,N_11801);
or U19146 (N_19146,N_11367,N_13300);
and U19147 (N_19147,N_12869,N_13144);
and U19148 (N_19148,N_10205,N_12241);
xor U19149 (N_19149,N_12788,N_12990);
nand U19150 (N_19150,N_12119,N_12180);
or U19151 (N_19151,N_14224,N_12440);
and U19152 (N_19152,N_12316,N_13508);
and U19153 (N_19153,N_11419,N_10137);
and U19154 (N_19154,N_11188,N_11877);
or U19155 (N_19155,N_10769,N_13266);
nor U19156 (N_19156,N_10928,N_14187);
nand U19157 (N_19157,N_14327,N_12001);
and U19158 (N_19158,N_10149,N_11670);
and U19159 (N_19159,N_14296,N_10391);
or U19160 (N_19160,N_13491,N_11101);
nand U19161 (N_19161,N_13453,N_11072);
nand U19162 (N_19162,N_11938,N_10901);
and U19163 (N_19163,N_13151,N_12053);
and U19164 (N_19164,N_14243,N_13090);
nor U19165 (N_19165,N_10183,N_14995);
nor U19166 (N_19166,N_14251,N_14862);
and U19167 (N_19167,N_14228,N_14641);
and U19168 (N_19168,N_14218,N_11034);
nor U19169 (N_19169,N_11328,N_13277);
and U19170 (N_19170,N_11513,N_11396);
xnor U19171 (N_19171,N_10060,N_11828);
nand U19172 (N_19172,N_14052,N_10501);
and U19173 (N_19173,N_11176,N_14324);
nand U19174 (N_19174,N_13189,N_12279);
nand U19175 (N_19175,N_10346,N_11298);
nor U19176 (N_19176,N_10237,N_13753);
nor U19177 (N_19177,N_14586,N_14436);
nor U19178 (N_19178,N_11355,N_13487);
xnor U19179 (N_19179,N_10610,N_11349);
or U19180 (N_19180,N_14775,N_10497);
or U19181 (N_19181,N_13260,N_14419);
nand U19182 (N_19182,N_11752,N_14749);
nor U19183 (N_19183,N_14699,N_11858);
nand U19184 (N_19184,N_12455,N_10897);
nand U19185 (N_19185,N_11879,N_10299);
xor U19186 (N_19186,N_14862,N_14115);
and U19187 (N_19187,N_10973,N_12340);
nor U19188 (N_19188,N_13471,N_10910);
or U19189 (N_19189,N_12989,N_14233);
nand U19190 (N_19190,N_11166,N_13563);
nor U19191 (N_19191,N_10796,N_13598);
and U19192 (N_19192,N_11649,N_11267);
nor U19193 (N_19193,N_12323,N_12767);
nor U19194 (N_19194,N_14197,N_12727);
nand U19195 (N_19195,N_11887,N_10731);
nor U19196 (N_19196,N_14446,N_10265);
or U19197 (N_19197,N_12031,N_11111);
and U19198 (N_19198,N_14087,N_13214);
and U19199 (N_19199,N_14343,N_13781);
nor U19200 (N_19200,N_10008,N_13230);
nand U19201 (N_19201,N_14868,N_10050);
nand U19202 (N_19202,N_10958,N_12407);
nor U19203 (N_19203,N_14072,N_12913);
nor U19204 (N_19204,N_14770,N_14125);
or U19205 (N_19205,N_13434,N_14289);
nand U19206 (N_19206,N_11214,N_11793);
nand U19207 (N_19207,N_13855,N_11697);
nand U19208 (N_19208,N_12170,N_12607);
or U19209 (N_19209,N_12745,N_14915);
nand U19210 (N_19210,N_11594,N_11397);
and U19211 (N_19211,N_12800,N_10104);
nand U19212 (N_19212,N_10004,N_11969);
or U19213 (N_19213,N_14810,N_13205);
nand U19214 (N_19214,N_10302,N_14090);
xnor U19215 (N_19215,N_12080,N_14394);
nor U19216 (N_19216,N_14275,N_10797);
nor U19217 (N_19217,N_11890,N_10373);
nor U19218 (N_19218,N_11529,N_11650);
or U19219 (N_19219,N_10227,N_14793);
nor U19220 (N_19220,N_10544,N_13753);
nor U19221 (N_19221,N_11324,N_10421);
nor U19222 (N_19222,N_13568,N_14455);
nor U19223 (N_19223,N_12226,N_10468);
nand U19224 (N_19224,N_14883,N_14357);
or U19225 (N_19225,N_11718,N_13112);
and U19226 (N_19226,N_12472,N_11859);
nand U19227 (N_19227,N_14218,N_12810);
or U19228 (N_19228,N_11605,N_10889);
nand U19229 (N_19229,N_10934,N_11376);
and U19230 (N_19230,N_14942,N_10203);
and U19231 (N_19231,N_14998,N_14207);
xnor U19232 (N_19232,N_14267,N_10285);
and U19233 (N_19233,N_11539,N_11810);
and U19234 (N_19234,N_11309,N_13877);
and U19235 (N_19235,N_12652,N_13658);
nor U19236 (N_19236,N_14626,N_10723);
and U19237 (N_19237,N_11002,N_14345);
nor U19238 (N_19238,N_14385,N_11023);
or U19239 (N_19239,N_13877,N_10402);
or U19240 (N_19240,N_12067,N_10094);
or U19241 (N_19241,N_11243,N_12234);
nand U19242 (N_19242,N_13630,N_13940);
nor U19243 (N_19243,N_12957,N_14457);
nor U19244 (N_19244,N_11739,N_11227);
nor U19245 (N_19245,N_12092,N_10351);
xor U19246 (N_19246,N_13773,N_14190);
or U19247 (N_19247,N_14042,N_12758);
and U19248 (N_19248,N_12171,N_14773);
xor U19249 (N_19249,N_14333,N_12802);
or U19250 (N_19250,N_13995,N_12086);
nand U19251 (N_19251,N_14573,N_14078);
xor U19252 (N_19252,N_12776,N_10986);
nor U19253 (N_19253,N_14037,N_14035);
or U19254 (N_19254,N_10781,N_10229);
and U19255 (N_19255,N_12219,N_10347);
or U19256 (N_19256,N_14266,N_13585);
or U19257 (N_19257,N_10328,N_10615);
or U19258 (N_19258,N_14656,N_12577);
nor U19259 (N_19259,N_12219,N_11651);
nand U19260 (N_19260,N_14256,N_13781);
xor U19261 (N_19261,N_14340,N_13071);
nor U19262 (N_19262,N_13955,N_12695);
nand U19263 (N_19263,N_10989,N_14673);
nor U19264 (N_19264,N_11211,N_14376);
or U19265 (N_19265,N_13568,N_10091);
nor U19266 (N_19266,N_13789,N_11299);
nor U19267 (N_19267,N_10111,N_12871);
nor U19268 (N_19268,N_12070,N_13059);
or U19269 (N_19269,N_11561,N_12738);
or U19270 (N_19270,N_13287,N_11003);
and U19271 (N_19271,N_12535,N_10729);
and U19272 (N_19272,N_14040,N_10102);
and U19273 (N_19273,N_13005,N_11741);
and U19274 (N_19274,N_13612,N_11686);
or U19275 (N_19275,N_11268,N_13451);
or U19276 (N_19276,N_11769,N_12035);
nand U19277 (N_19277,N_14390,N_10543);
nor U19278 (N_19278,N_10501,N_13656);
xnor U19279 (N_19279,N_12628,N_12929);
nor U19280 (N_19280,N_13307,N_13460);
xnor U19281 (N_19281,N_11237,N_14107);
and U19282 (N_19282,N_11253,N_10040);
nor U19283 (N_19283,N_12451,N_14791);
and U19284 (N_19284,N_14875,N_14531);
nand U19285 (N_19285,N_14390,N_13932);
xnor U19286 (N_19286,N_14657,N_12280);
nor U19287 (N_19287,N_11243,N_11864);
or U19288 (N_19288,N_14250,N_13919);
nor U19289 (N_19289,N_11597,N_14938);
and U19290 (N_19290,N_13157,N_13438);
and U19291 (N_19291,N_12814,N_11868);
and U19292 (N_19292,N_11722,N_12846);
nand U19293 (N_19293,N_11692,N_12978);
nor U19294 (N_19294,N_12664,N_13991);
xnor U19295 (N_19295,N_13891,N_12779);
or U19296 (N_19296,N_10691,N_10072);
nand U19297 (N_19297,N_12947,N_10538);
nor U19298 (N_19298,N_10093,N_13990);
nor U19299 (N_19299,N_14254,N_11007);
nand U19300 (N_19300,N_10200,N_14028);
nor U19301 (N_19301,N_13199,N_10279);
nand U19302 (N_19302,N_11028,N_11405);
and U19303 (N_19303,N_10888,N_11532);
xor U19304 (N_19304,N_13549,N_12197);
nor U19305 (N_19305,N_13973,N_13416);
or U19306 (N_19306,N_10725,N_11282);
nand U19307 (N_19307,N_13499,N_13011);
and U19308 (N_19308,N_13266,N_10944);
or U19309 (N_19309,N_10279,N_10686);
and U19310 (N_19310,N_14999,N_11481);
nand U19311 (N_19311,N_12327,N_13635);
nor U19312 (N_19312,N_11771,N_13745);
nor U19313 (N_19313,N_12413,N_13536);
nand U19314 (N_19314,N_14503,N_12456);
xor U19315 (N_19315,N_11245,N_13286);
and U19316 (N_19316,N_11841,N_13282);
or U19317 (N_19317,N_11292,N_13502);
or U19318 (N_19318,N_14479,N_11462);
nand U19319 (N_19319,N_13828,N_13612);
nand U19320 (N_19320,N_10974,N_11813);
and U19321 (N_19321,N_10189,N_13429);
or U19322 (N_19322,N_13461,N_12109);
nor U19323 (N_19323,N_13258,N_12513);
or U19324 (N_19324,N_14400,N_14452);
nand U19325 (N_19325,N_12423,N_13194);
or U19326 (N_19326,N_13126,N_14734);
nor U19327 (N_19327,N_12076,N_11677);
and U19328 (N_19328,N_10002,N_11467);
or U19329 (N_19329,N_10063,N_12103);
nor U19330 (N_19330,N_10089,N_12875);
or U19331 (N_19331,N_10500,N_14354);
nor U19332 (N_19332,N_11485,N_13892);
or U19333 (N_19333,N_12717,N_10389);
nor U19334 (N_19334,N_14338,N_11581);
and U19335 (N_19335,N_14376,N_11912);
xor U19336 (N_19336,N_12566,N_10172);
xnor U19337 (N_19337,N_11978,N_10680);
nor U19338 (N_19338,N_13701,N_12729);
nor U19339 (N_19339,N_11995,N_12887);
nor U19340 (N_19340,N_10008,N_14469);
or U19341 (N_19341,N_10583,N_11375);
nand U19342 (N_19342,N_13707,N_13023);
xor U19343 (N_19343,N_11854,N_14528);
or U19344 (N_19344,N_13176,N_13093);
nand U19345 (N_19345,N_12667,N_14991);
nand U19346 (N_19346,N_13706,N_10380);
nor U19347 (N_19347,N_12321,N_14145);
nor U19348 (N_19348,N_13218,N_13418);
xnor U19349 (N_19349,N_11802,N_10367);
nand U19350 (N_19350,N_10148,N_12633);
nand U19351 (N_19351,N_14998,N_13507);
and U19352 (N_19352,N_13689,N_11651);
nand U19353 (N_19353,N_10420,N_14770);
or U19354 (N_19354,N_11870,N_11635);
or U19355 (N_19355,N_13786,N_10165);
and U19356 (N_19356,N_12574,N_10715);
and U19357 (N_19357,N_12555,N_10643);
and U19358 (N_19358,N_14718,N_13236);
nand U19359 (N_19359,N_13213,N_14234);
and U19360 (N_19360,N_14792,N_14506);
and U19361 (N_19361,N_11532,N_14693);
nor U19362 (N_19362,N_14260,N_11943);
and U19363 (N_19363,N_10984,N_14542);
nand U19364 (N_19364,N_12706,N_13316);
nand U19365 (N_19365,N_12100,N_12511);
nand U19366 (N_19366,N_10112,N_11286);
or U19367 (N_19367,N_11293,N_14189);
or U19368 (N_19368,N_11516,N_10222);
nand U19369 (N_19369,N_10689,N_11051);
nand U19370 (N_19370,N_14502,N_10240);
and U19371 (N_19371,N_11408,N_13570);
or U19372 (N_19372,N_14350,N_12777);
or U19373 (N_19373,N_10161,N_12950);
and U19374 (N_19374,N_14843,N_11731);
and U19375 (N_19375,N_13238,N_12021);
and U19376 (N_19376,N_13624,N_11025);
and U19377 (N_19377,N_11259,N_13035);
xor U19378 (N_19378,N_10235,N_10310);
or U19379 (N_19379,N_14325,N_14487);
nand U19380 (N_19380,N_14722,N_14338);
or U19381 (N_19381,N_14662,N_12776);
or U19382 (N_19382,N_10802,N_13613);
nor U19383 (N_19383,N_10921,N_14096);
xnor U19384 (N_19384,N_14438,N_14784);
nor U19385 (N_19385,N_12084,N_11151);
or U19386 (N_19386,N_14702,N_12631);
nor U19387 (N_19387,N_14738,N_10824);
and U19388 (N_19388,N_11826,N_13163);
or U19389 (N_19389,N_12066,N_14876);
or U19390 (N_19390,N_12821,N_14376);
and U19391 (N_19391,N_14879,N_10629);
and U19392 (N_19392,N_10558,N_10580);
and U19393 (N_19393,N_10230,N_13458);
and U19394 (N_19394,N_13564,N_14962);
and U19395 (N_19395,N_10392,N_12276);
nand U19396 (N_19396,N_10126,N_14719);
nor U19397 (N_19397,N_14209,N_11524);
nand U19398 (N_19398,N_13640,N_10704);
or U19399 (N_19399,N_12880,N_10021);
xnor U19400 (N_19400,N_14670,N_14680);
nand U19401 (N_19401,N_13637,N_11951);
and U19402 (N_19402,N_12273,N_13386);
nand U19403 (N_19403,N_14585,N_12681);
and U19404 (N_19404,N_14355,N_11750);
or U19405 (N_19405,N_13785,N_13190);
and U19406 (N_19406,N_10492,N_14281);
nor U19407 (N_19407,N_11800,N_14671);
nand U19408 (N_19408,N_14382,N_10128);
xnor U19409 (N_19409,N_11043,N_11673);
nand U19410 (N_19410,N_14636,N_11374);
and U19411 (N_19411,N_12457,N_13383);
and U19412 (N_19412,N_10490,N_12447);
nand U19413 (N_19413,N_11572,N_12051);
or U19414 (N_19414,N_11177,N_13048);
nand U19415 (N_19415,N_11963,N_10008);
and U19416 (N_19416,N_11932,N_11269);
nor U19417 (N_19417,N_13362,N_12706);
nand U19418 (N_19418,N_14823,N_10635);
xor U19419 (N_19419,N_12380,N_11692);
and U19420 (N_19420,N_13666,N_13369);
nor U19421 (N_19421,N_13102,N_12495);
or U19422 (N_19422,N_13049,N_13203);
or U19423 (N_19423,N_12426,N_13681);
and U19424 (N_19424,N_13722,N_11739);
and U19425 (N_19425,N_12676,N_12933);
nor U19426 (N_19426,N_14254,N_11803);
or U19427 (N_19427,N_10628,N_13896);
nand U19428 (N_19428,N_11605,N_10182);
and U19429 (N_19429,N_13132,N_12912);
and U19430 (N_19430,N_10051,N_12226);
nor U19431 (N_19431,N_12052,N_12234);
nand U19432 (N_19432,N_11486,N_10455);
nor U19433 (N_19433,N_13360,N_11319);
xor U19434 (N_19434,N_14906,N_12567);
nand U19435 (N_19435,N_14686,N_14493);
nor U19436 (N_19436,N_10273,N_13517);
xnor U19437 (N_19437,N_10262,N_12118);
nor U19438 (N_19438,N_11116,N_14562);
and U19439 (N_19439,N_14777,N_14259);
nor U19440 (N_19440,N_10619,N_12136);
nor U19441 (N_19441,N_10048,N_10382);
nor U19442 (N_19442,N_11632,N_10181);
xnor U19443 (N_19443,N_12581,N_10280);
and U19444 (N_19444,N_11168,N_12671);
or U19445 (N_19445,N_11220,N_10858);
and U19446 (N_19446,N_10110,N_11348);
xnor U19447 (N_19447,N_11001,N_14399);
xnor U19448 (N_19448,N_12122,N_13815);
and U19449 (N_19449,N_12629,N_10974);
and U19450 (N_19450,N_11600,N_12440);
nor U19451 (N_19451,N_13528,N_11006);
or U19452 (N_19452,N_13940,N_13261);
nor U19453 (N_19453,N_11915,N_13963);
xnor U19454 (N_19454,N_11967,N_14077);
nand U19455 (N_19455,N_11444,N_12214);
and U19456 (N_19456,N_14097,N_10854);
and U19457 (N_19457,N_13961,N_11245);
and U19458 (N_19458,N_10696,N_14794);
nor U19459 (N_19459,N_14352,N_12148);
nor U19460 (N_19460,N_12058,N_11719);
nand U19461 (N_19461,N_12207,N_12506);
xor U19462 (N_19462,N_10474,N_11988);
nand U19463 (N_19463,N_10075,N_11240);
nor U19464 (N_19464,N_14956,N_12273);
xor U19465 (N_19465,N_10016,N_11710);
xor U19466 (N_19466,N_13215,N_14334);
xor U19467 (N_19467,N_13288,N_11456);
nor U19468 (N_19468,N_13367,N_12556);
and U19469 (N_19469,N_11423,N_14831);
nor U19470 (N_19470,N_13757,N_10187);
nand U19471 (N_19471,N_12591,N_12061);
nand U19472 (N_19472,N_10585,N_10267);
and U19473 (N_19473,N_11650,N_13631);
xor U19474 (N_19474,N_13206,N_11736);
nor U19475 (N_19475,N_13844,N_12510);
or U19476 (N_19476,N_11251,N_12792);
nand U19477 (N_19477,N_13278,N_14715);
nand U19478 (N_19478,N_10154,N_10781);
or U19479 (N_19479,N_14800,N_12203);
nor U19480 (N_19480,N_13033,N_11202);
nor U19481 (N_19481,N_13091,N_10184);
and U19482 (N_19482,N_13626,N_14764);
xnor U19483 (N_19483,N_14510,N_11767);
and U19484 (N_19484,N_10728,N_10915);
nand U19485 (N_19485,N_12968,N_13762);
and U19486 (N_19486,N_10662,N_11223);
nor U19487 (N_19487,N_12471,N_12610);
or U19488 (N_19488,N_11120,N_10322);
nand U19489 (N_19489,N_10404,N_10842);
nor U19490 (N_19490,N_11605,N_10946);
nor U19491 (N_19491,N_11683,N_10453);
and U19492 (N_19492,N_12578,N_10306);
nand U19493 (N_19493,N_10971,N_14036);
or U19494 (N_19494,N_13488,N_14409);
or U19495 (N_19495,N_10140,N_10176);
nor U19496 (N_19496,N_10391,N_12392);
nand U19497 (N_19497,N_10672,N_11391);
nand U19498 (N_19498,N_10666,N_11414);
nor U19499 (N_19499,N_12721,N_10409);
and U19500 (N_19500,N_13341,N_14063);
and U19501 (N_19501,N_10765,N_14247);
xnor U19502 (N_19502,N_11256,N_12612);
or U19503 (N_19503,N_12902,N_10148);
or U19504 (N_19504,N_11116,N_10765);
nor U19505 (N_19505,N_11941,N_12970);
nand U19506 (N_19506,N_11000,N_12565);
nand U19507 (N_19507,N_11374,N_12110);
and U19508 (N_19508,N_10797,N_10075);
and U19509 (N_19509,N_14463,N_10059);
or U19510 (N_19510,N_13004,N_11383);
nand U19511 (N_19511,N_10906,N_11547);
nor U19512 (N_19512,N_14321,N_13627);
nor U19513 (N_19513,N_13522,N_14798);
and U19514 (N_19514,N_14270,N_14937);
nand U19515 (N_19515,N_11659,N_12448);
nor U19516 (N_19516,N_13435,N_14768);
or U19517 (N_19517,N_14771,N_14351);
nor U19518 (N_19518,N_12569,N_11811);
or U19519 (N_19519,N_12458,N_14789);
xor U19520 (N_19520,N_14311,N_14101);
nor U19521 (N_19521,N_14838,N_11006);
xnor U19522 (N_19522,N_14386,N_14556);
nor U19523 (N_19523,N_14918,N_13050);
or U19524 (N_19524,N_14470,N_12372);
or U19525 (N_19525,N_10465,N_12890);
nor U19526 (N_19526,N_11325,N_13229);
nand U19527 (N_19527,N_11812,N_13576);
nor U19528 (N_19528,N_14804,N_11764);
and U19529 (N_19529,N_11738,N_10256);
or U19530 (N_19530,N_12471,N_10087);
and U19531 (N_19531,N_10042,N_13183);
or U19532 (N_19532,N_14763,N_13822);
nor U19533 (N_19533,N_14514,N_11523);
nand U19534 (N_19534,N_11509,N_14751);
and U19535 (N_19535,N_11488,N_12625);
nand U19536 (N_19536,N_13720,N_11517);
or U19537 (N_19537,N_14502,N_13363);
and U19538 (N_19538,N_11024,N_12871);
nand U19539 (N_19539,N_14085,N_14887);
or U19540 (N_19540,N_12411,N_13689);
nand U19541 (N_19541,N_10222,N_11664);
and U19542 (N_19542,N_11550,N_14402);
nand U19543 (N_19543,N_14752,N_10638);
nor U19544 (N_19544,N_14653,N_13026);
nand U19545 (N_19545,N_11399,N_13860);
nand U19546 (N_19546,N_13162,N_10132);
nor U19547 (N_19547,N_13220,N_10833);
nand U19548 (N_19548,N_14874,N_11879);
xnor U19549 (N_19549,N_10277,N_13688);
nand U19550 (N_19550,N_14565,N_11664);
xor U19551 (N_19551,N_13665,N_13144);
and U19552 (N_19552,N_10371,N_12266);
or U19553 (N_19553,N_14776,N_12797);
nand U19554 (N_19554,N_11720,N_12542);
nand U19555 (N_19555,N_14418,N_12430);
nand U19556 (N_19556,N_11981,N_11081);
and U19557 (N_19557,N_11529,N_11757);
nor U19558 (N_19558,N_11918,N_14421);
nor U19559 (N_19559,N_10804,N_13487);
or U19560 (N_19560,N_11248,N_10400);
nand U19561 (N_19561,N_14423,N_11648);
or U19562 (N_19562,N_13234,N_11995);
or U19563 (N_19563,N_11860,N_12245);
nand U19564 (N_19564,N_10340,N_11846);
nand U19565 (N_19565,N_12443,N_14501);
or U19566 (N_19566,N_11618,N_11814);
nand U19567 (N_19567,N_10184,N_14742);
xor U19568 (N_19568,N_14820,N_13093);
or U19569 (N_19569,N_12418,N_12671);
or U19570 (N_19570,N_11613,N_14894);
xor U19571 (N_19571,N_13652,N_11102);
and U19572 (N_19572,N_11703,N_11481);
and U19573 (N_19573,N_14789,N_13565);
nand U19574 (N_19574,N_10078,N_13193);
and U19575 (N_19575,N_12509,N_11449);
or U19576 (N_19576,N_13081,N_14175);
nor U19577 (N_19577,N_13856,N_13943);
xnor U19578 (N_19578,N_13430,N_12866);
nand U19579 (N_19579,N_13490,N_12986);
nand U19580 (N_19580,N_14400,N_12942);
or U19581 (N_19581,N_10303,N_12590);
or U19582 (N_19582,N_14430,N_13093);
nand U19583 (N_19583,N_10993,N_14302);
nor U19584 (N_19584,N_14287,N_10638);
and U19585 (N_19585,N_12264,N_13800);
nand U19586 (N_19586,N_14725,N_11196);
xnor U19587 (N_19587,N_14228,N_10331);
nor U19588 (N_19588,N_13442,N_13144);
and U19589 (N_19589,N_13902,N_12694);
or U19590 (N_19590,N_13555,N_11028);
xor U19591 (N_19591,N_10943,N_13340);
nand U19592 (N_19592,N_10191,N_11727);
nor U19593 (N_19593,N_12201,N_14018);
or U19594 (N_19594,N_14438,N_13920);
nand U19595 (N_19595,N_13662,N_12234);
or U19596 (N_19596,N_10269,N_10053);
nand U19597 (N_19597,N_11564,N_14653);
or U19598 (N_19598,N_10310,N_12326);
nand U19599 (N_19599,N_12729,N_10252);
and U19600 (N_19600,N_14797,N_13757);
nor U19601 (N_19601,N_12336,N_12050);
nand U19602 (N_19602,N_10164,N_14728);
xnor U19603 (N_19603,N_14868,N_11506);
nor U19604 (N_19604,N_11513,N_14314);
and U19605 (N_19605,N_10399,N_11287);
and U19606 (N_19606,N_14494,N_13287);
and U19607 (N_19607,N_14121,N_10392);
nor U19608 (N_19608,N_14704,N_13159);
or U19609 (N_19609,N_10493,N_14173);
nand U19610 (N_19610,N_11828,N_10102);
xor U19611 (N_19611,N_12506,N_11520);
xnor U19612 (N_19612,N_13790,N_12645);
or U19613 (N_19613,N_13047,N_13558);
nor U19614 (N_19614,N_11108,N_11731);
and U19615 (N_19615,N_13335,N_14579);
xnor U19616 (N_19616,N_13386,N_11838);
and U19617 (N_19617,N_10175,N_12045);
and U19618 (N_19618,N_12689,N_11484);
nor U19619 (N_19619,N_13905,N_13096);
or U19620 (N_19620,N_10927,N_10283);
nand U19621 (N_19621,N_11464,N_10468);
nor U19622 (N_19622,N_13976,N_13167);
nor U19623 (N_19623,N_14910,N_11367);
and U19624 (N_19624,N_11078,N_14732);
nand U19625 (N_19625,N_13248,N_13851);
and U19626 (N_19626,N_13931,N_14501);
nor U19627 (N_19627,N_13779,N_13784);
nor U19628 (N_19628,N_14038,N_10927);
and U19629 (N_19629,N_11488,N_10491);
or U19630 (N_19630,N_14762,N_14056);
nor U19631 (N_19631,N_11804,N_11231);
nand U19632 (N_19632,N_12760,N_11302);
xor U19633 (N_19633,N_13666,N_10935);
nand U19634 (N_19634,N_11015,N_11643);
nor U19635 (N_19635,N_11191,N_12212);
or U19636 (N_19636,N_14852,N_14653);
and U19637 (N_19637,N_10997,N_13005);
nor U19638 (N_19638,N_11346,N_10344);
nand U19639 (N_19639,N_13554,N_12506);
or U19640 (N_19640,N_10630,N_11014);
nor U19641 (N_19641,N_13459,N_11029);
and U19642 (N_19642,N_14603,N_14441);
xor U19643 (N_19643,N_12068,N_13367);
and U19644 (N_19644,N_14057,N_12517);
or U19645 (N_19645,N_13720,N_13822);
and U19646 (N_19646,N_13162,N_13715);
and U19647 (N_19647,N_13362,N_10934);
nor U19648 (N_19648,N_12044,N_10313);
or U19649 (N_19649,N_14385,N_11739);
xor U19650 (N_19650,N_10434,N_14414);
nor U19651 (N_19651,N_14378,N_11764);
xor U19652 (N_19652,N_13883,N_10323);
and U19653 (N_19653,N_14770,N_12381);
or U19654 (N_19654,N_12165,N_12416);
nor U19655 (N_19655,N_12077,N_10427);
or U19656 (N_19656,N_11022,N_11883);
and U19657 (N_19657,N_11085,N_14806);
or U19658 (N_19658,N_14321,N_12909);
nand U19659 (N_19659,N_11175,N_12623);
or U19660 (N_19660,N_10071,N_12205);
nor U19661 (N_19661,N_12036,N_13951);
xnor U19662 (N_19662,N_11770,N_11569);
or U19663 (N_19663,N_10548,N_11771);
nor U19664 (N_19664,N_12497,N_10779);
nor U19665 (N_19665,N_13075,N_10454);
or U19666 (N_19666,N_12925,N_12157);
nor U19667 (N_19667,N_10849,N_12096);
or U19668 (N_19668,N_14873,N_13026);
nand U19669 (N_19669,N_11506,N_12918);
xnor U19670 (N_19670,N_10887,N_10614);
nor U19671 (N_19671,N_13456,N_11991);
and U19672 (N_19672,N_12376,N_12014);
xnor U19673 (N_19673,N_11770,N_10845);
nand U19674 (N_19674,N_12485,N_14452);
nor U19675 (N_19675,N_11051,N_14808);
xor U19676 (N_19676,N_11794,N_11271);
nand U19677 (N_19677,N_13298,N_10604);
xnor U19678 (N_19678,N_14595,N_14914);
nor U19679 (N_19679,N_12626,N_10816);
nor U19680 (N_19680,N_14552,N_10903);
and U19681 (N_19681,N_13451,N_10391);
nand U19682 (N_19682,N_11107,N_11953);
or U19683 (N_19683,N_14863,N_13980);
and U19684 (N_19684,N_10859,N_13752);
and U19685 (N_19685,N_12261,N_13060);
and U19686 (N_19686,N_14396,N_11570);
nor U19687 (N_19687,N_13188,N_10560);
nand U19688 (N_19688,N_13508,N_12665);
or U19689 (N_19689,N_10954,N_12139);
or U19690 (N_19690,N_12478,N_12397);
nand U19691 (N_19691,N_10611,N_13551);
nand U19692 (N_19692,N_11107,N_13191);
and U19693 (N_19693,N_11992,N_14735);
xor U19694 (N_19694,N_12396,N_12802);
nor U19695 (N_19695,N_13130,N_11352);
and U19696 (N_19696,N_12145,N_10606);
and U19697 (N_19697,N_11150,N_14571);
and U19698 (N_19698,N_11919,N_12701);
or U19699 (N_19699,N_12853,N_13054);
nor U19700 (N_19700,N_13110,N_13801);
or U19701 (N_19701,N_11427,N_10783);
nand U19702 (N_19702,N_14429,N_10961);
and U19703 (N_19703,N_13508,N_11941);
nand U19704 (N_19704,N_13078,N_11177);
nor U19705 (N_19705,N_12017,N_13461);
and U19706 (N_19706,N_10721,N_12892);
or U19707 (N_19707,N_10999,N_13651);
or U19708 (N_19708,N_14872,N_10600);
nor U19709 (N_19709,N_10902,N_11970);
nor U19710 (N_19710,N_11856,N_11738);
or U19711 (N_19711,N_10966,N_11171);
and U19712 (N_19712,N_14288,N_14308);
nor U19713 (N_19713,N_13066,N_12951);
xnor U19714 (N_19714,N_11321,N_14859);
nor U19715 (N_19715,N_11643,N_12425);
and U19716 (N_19716,N_14727,N_10618);
or U19717 (N_19717,N_11031,N_14474);
nor U19718 (N_19718,N_10110,N_14717);
nand U19719 (N_19719,N_12637,N_10504);
xnor U19720 (N_19720,N_11130,N_11241);
or U19721 (N_19721,N_14531,N_12019);
nor U19722 (N_19722,N_10409,N_12503);
or U19723 (N_19723,N_12592,N_13360);
xnor U19724 (N_19724,N_13412,N_10454);
nor U19725 (N_19725,N_13447,N_12713);
nand U19726 (N_19726,N_11930,N_10708);
xnor U19727 (N_19727,N_10608,N_12840);
or U19728 (N_19728,N_12552,N_11801);
nor U19729 (N_19729,N_10229,N_13576);
nor U19730 (N_19730,N_12556,N_11175);
nand U19731 (N_19731,N_12969,N_11524);
nor U19732 (N_19732,N_14488,N_11884);
nand U19733 (N_19733,N_11961,N_12444);
or U19734 (N_19734,N_10255,N_13858);
nand U19735 (N_19735,N_12051,N_13023);
nand U19736 (N_19736,N_13602,N_10484);
and U19737 (N_19737,N_10914,N_14394);
or U19738 (N_19738,N_10728,N_10952);
xor U19739 (N_19739,N_11162,N_12087);
nor U19740 (N_19740,N_14818,N_11454);
or U19741 (N_19741,N_12352,N_14804);
nor U19742 (N_19742,N_14804,N_14580);
nand U19743 (N_19743,N_11503,N_10396);
nor U19744 (N_19744,N_12800,N_14664);
and U19745 (N_19745,N_11817,N_11018);
or U19746 (N_19746,N_12465,N_11046);
xor U19747 (N_19747,N_12287,N_14843);
and U19748 (N_19748,N_11710,N_11608);
xor U19749 (N_19749,N_10744,N_10707);
or U19750 (N_19750,N_14641,N_12634);
nand U19751 (N_19751,N_13070,N_14431);
or U19752 (N_19752,N_14043,N_14759);
nor U19753 (N_19753,N_12585,N_10137);
nand U19754 (N_19754,N_14142,N_11344);
and U19755 (N_19755,N_12601,N_10028);
and U19756 (N_19756,N_14390,N_13110);
nand U19757 (N_19757,N_12922,N_11586);
and U19758 (N_19758,N_13961,N_14094);
nor U19759 (N_19759,N_10832,N_13432);
or U19760 (N_19760,N_12290,N_14177);
nand U19761 (N_19761,N_14737,N_12946);
nor U19762 (N_19762,N_12364,N_11763);
nor U19763 (N_19763,N_12750,N_14601);
xnor U19764 (N_19764,N_11930,N_14659);
and U19765 (N_19765,N_11274,N_11665);
nand U19766 (N_19766,N_12328,N_14758);
nor U19767 (N_19767,N_14493,N_13363);
or U19768 (N_19768,N_12292,N_10594);
xnor U19769 (N_19769,N_14510,N_12940);
xor U19770 (N_19770,N_13933,N_13426);
nor U19771 (N_19771,N_14300,N_10195);
nor U19772 (N_19772,N_10910,N_14579);
or U19773 (N_19773,N_14401,N_12700);
xor U19774 (N_19774,N_13067,N_11341);
nand U19775 (N_19775,N_13871,N_12844);
nand U19776 (N_19776,N_11682,N_10224);
and U19777 (N_19777,N_12897,N_13566);
and U19778 (N_19778,N_12485,N_12282);
and U19779 (N_19779,N_11175,N_12483);
nor U19780 (N_19780,N_13791,N_11663);
xnor U19781 (N_19781,N_10709,N_11527);
nand U19782 (N_19782,N_13006,N_10193);
nor U19783 (N_19783,N_12545,N_13427);
nand U19784 (N_19784,N_12962,N_11169);
nor U19785 (N_19785,N_12209,N_10956);
and U19786 (N_19786,N_12375,N_13362);
or U19787 (N_19787,N_14903,N_13442);
or U19788 (N_19788,N_11715,N_10890);
nand U19789 (N_19789,N_14636,N_10854);
or U19790 (N_19790,N_10494,N_10749);
xor U19791 (N_19791,N_10295,N_10232);
nor U19792 (N_19792,N_10469,N_14582);
and U19793 (N_19793,N_10527,N_14130);
nor U19794 (N_19794,N_11959,N_12288);
xor U19795 (N_19795,N_13998,N_14498);
xnor U19796 (N_19796,N_10869,N_14078);
or U19797 (N_19797,N_10677,N_14801);
xnor U19798 (N_19798,N_14494,N_14251);
nand U19799 (N_19799,N_10536,N_14946);
nand U19800 (N_19800,N_10023,N_10155);
nor U19801 (N_19801,N_14115,N_11029);
xnor U19802 (N_19802,N_10960,N_13184);
nand U19803 (N_19803,N_14245,N_13997);
or U19804 (N_19804,N_10897,N_11412);
nor U19805 (N_19805,N_14185,N_10254);
nand U19806 (N_19806,N_14389,N_12020);
or U19807 (N_19807,N_11860,N_10914);
or U19808 (N_19808,N_10678,N_10109);
nor U19809 (N_19809,N_10989,N_12846);
nor U19810 (N_19810,N_12829,N_12650);
and U19811 (N_19811,N_10441,N_11991);
nor U19812 (N_19812,N_12073,N_14724);
or U19813 (N_19813,N_11192,N_12089);
and U19814 (N_19814,N_12854,N_10965);
and U19815 (N_19815,N_10429,N_10123);
or U19816 (N_19816,N_11473,N_12575);
nor U19817 (N_19817,N_11328,N_11074);
nor U19818 (N_19818,N_10053,N_11478);
or U19819 (N_19819,N_10635,N_13051);
or U19820 (N_19820,N_14479,N_13476);
xnor U19821 (N_19821,N_10411,N_10562);
nor U19822 (N_19822,N_12522,N_13630);
and U19823 (N_19823,N_10671,N_14944);
or U19824 (N_19824,N_11148,N_13950);
nor U19825 (N_19825,N_12922,N_11347);
or U19826 (N_19826,N_10518,N_11436);
nand U19827 (N_19827,N_14775,N_14277);
or U19828 (N_19828,N_14933,N_10156);
and U19829 (N_19829,N_11158,N_13417);
xor U19830 (N_19830,N_11349,N_13434);
nor U19831 (N_19831,N_11750,N_10948);
nor U19832 (N_19832,N_13690,N_10466);
nand U19833 (N_19833,N_10744,N_14161);
and U19834 (N_19834,N_13497,N_14964);
and U19835 (N_19835,N_13152,N_13954);
and U19836 (N_19836,N_11609,N_14132);
and U19837 (N_19837,N_11872,N_10528);
xnor U19838 (N_19838,N_10725,N_14492);
nor U19839 (N_19839,N_10610,N_14732);
nor U19840 (N_19840,N_12891,N_13889);
or U19841 (N_19841,N_13684,N_12002);
or U19842 (N_19842,N_11173,N_11118);
nor U19843 (N_19843,N_13921,N_12233);
nand U19844 (N_19844,N_13126,N_11975);
or U19845 (N_19845,N_10812,N_14168);
nand U19846 (N_19846,N_12559,N_11480);
or U19847 (N_19847,N_10048,N_13175);
and U19848 (N_19848,N_13290,N_14438);
nand U19849 (N_19849,N_11885,N_13074);
or U19850 (N_19850,N_13372,N_10611);
nor U19851 (N_19851,N_11260,N_14912);
or U19852 (N_19852,N_12375,N_11362);
and U19853 (N_19853,N_11165,N_11927);
nor U19854 (N_19854,N_11086,N_14068);
nand U19855 (N_19855,N_10963,N_14008);
and U19856 (N_19856,N_13118,N_13350);
xnor U19857 (N_19857,N_14518,N_11422);
nor U19858 (N_19858,N_10349,N_13387);
or U19859 (N_19859,N_12920,N_12241);
and U19860 (N_19860,N_12468,N_12375);
nand U19861 (N_19861,N_13145,N_14349);
nor U19862 (N_19862,N_12063,N_11875);
nand U19863 (N_19863,N_11899,N_14995);
nand U19864 (N_19864,N_13199,N_14170);
xor U19865 (N_19865,N_13199,N_12087);
nor U19866 (N_19866,N_10357,N_12483);
or U19867 (N_19867,N_14110,N_14672);
nor U19868 (N_19868,N_14533,N_14816);
and U19869 (N_19869,N_11705,N_14833);
nand U19870 (N_19870,N_14973,N_10328);
nor U19871 (N_19871,N_10859,N_11678);
nand U19872 (N_19872,N_13237,N_11390);
nor U19873 (N_19873,N_12279,N_11797);
nor U19874 (N_19874,N_12052,N_14174);
nor U19875 (N_19875,N_11247,N_11086);
nand U19876 (N_19876,N_13029,N_14174);
and U19877 (N_19877,N_13874,N_12567);
nand U19878 (N_19878,N_10600,N_11183);
nor U19879 (N_19879,N_14307,N_13092);
nand U19880 (N_19880,N_14385,N_12096);
or U19881 (N_19881,N_14109,N_13594);
or U19882 (N_19882,N_14802,N_10437);
and U19883 (N_19883,N_13261,N_14297);
or U19884 (N_19884,N_11883,N_12875);
nand U19885 (N_19885,N_11590,N_12419);
nor U19886 (N_19886,N_13699,N_11461);
or U19887 (N_19887,N_11162,N_13133);
xnor U19888 (N_19888,N_10306,N_14403);
and U19889 (N_19889,N_12219,N_11162);
nor U19890 (N_19890,N_14775,N_10829);
or U19891 (N_19891,N_13743,N_12325);
and U19892 (N_19892,N_12404,N_12254);
nand U19893 (N_19893,N_14838,N_13534);
nand U19894 (N_19894,N_14934,N_10790);
nand U19895 (N_19895,N_13636,N_12617);
nor U19896 (N_19896,N_11882,N_14407);
nand U19897 (N_19897,N_11605,N_11984);
nand U19898 (N_19898,N_12729,N_13850);
or U19899 (N_19899,N_12289,N_13029);
and U19900 (N_19900,N_13063,N_10370);
and U19901 (N_19901,N_13428,N_10929);
and U19902 (N_19902,N_11674,N_12561);
or U19903 (N_19903,N_11608,N_10752);
or U19904 (N_19904,N_13368,N_12241);
nor U19905 (N_19905,N_12376,N_11130);
nand U19906 (N_19906,N_14368,N_14796);
and U19907 (N_19907,N_13570,N_13013);
xnor U19908 (N_19908,N_12847,N_13171);
nand U19909 (N_19909,N_12571,N_13924);
xnor U19910 (N_19910,N_12229,N_13221);
nand U19911 (N_19911,N_11865,N_12062);
or U19912 (N_19912,N_10542,N_12823);
or U19913 (N_19913,N_10169,N_10886);
and U19914 (N_19914,N_12387,N_11229);
or U19915 (N_19915,N_14181,N_10584);
and U19916 (N_19916,N_10676,N_14699);
or U19917 (N_19917,N_10911,N_13614);
nand U19918 (N_19918,N_10141,N_10678);
or U19919 (N_19919,N_12107,N_14357);
nor U19920 (N_19920,N_14405,N_14856);
or U19921 (N_19921,N_11161,N_12328);
nor U19922 (N_19922,N_12321,N_13307);
xnor U19923 (N_19923,N_13682,N_10495);
and U19924 (N_19924,N_14218,N_12581);
or U19925 (N_19925,N_11050,N_14537);
nor U19926 (N_19926,N_14153,N_10378);
nor U19927 (N_19927,N_10014,N_10887);
or U19928 (N_19928,N_12730,N_14332);
or U19929 (N_19929,N_14224,N_13693);
nand U19930 (N_19930,N_14969,N_12325);
or U19931 (N_19931,N_12767,N_12859);
nor U19932 (N_19932,N_14950,N_14739);
nand U19933 (N_19933,N_13363,N_12402);
and U19934 (N_19934,N_11129,N_14236);
nand U19935 (N_19935,N_14527,N_13411);
or U19936 (N_19936,N_14973,N_11731);
and U19937 (N_19937,N_12319,N_10316);
xnor U19938 (N_19938,N_12873,N_12088);
or U19939 (N_19939,N_11657,N_11066);
and U19940 (N_19940,N_11835,N_13722);
and U19941 (N_19941,N_12993,N_11701);
nor U19942 (N_19942,N_10847,N_10235);
or U19943 (N_19943,N_14711,N_12361);
nor U19944 (N_19944,N_12411,N_14725);
nand U19945 (N_19945,N_11470,N_13325);
or U19946 (N_19946,N_12664,N_14286);
and U19947 (N_19947,N_14596,N_12093);
and U19948 (N_19948,N_11996,N_10360);
nor U19949 (N_19949,N_12471,N_12350);
and U19950 (N_19950,N_10840,N_10825);
nor U19951 (N_19951,N_11079,N_10715);
xnor U19952 (N_19952,N_11652,N_10344);
nor U19953 (N_19953,N_12019,N_12383);
nand U19954 (N_19954,N_12984,N_12239);
nand U19955 (N_19955,N_14918,N_14955);
nor U19956 (N_19956,N_12519,N_12552);
nor U19957 (N_19957,N_14832,N_12125);
or U19958 (N_19958,N_14096,N_11256);
or U19959 (N_19959,N_12839,N_12391);
or U19960 (N_19960,N_11695,N_12913);
nand U19961 (N_19961,N_10781,N_14930);
nand U19962 (N_19962,N_10542,N_11622);
and U19963 (N_19963,N_12392,N_11219);
or U19964 (N_19964,N_13086,N_10013);
xnor U19965 (N_19965,N_13338,N_14870);
nand U19966 (N_19966,N_14626,N_14199);
or U19967 (N_19967,N_10496,N_14419);
or U19968 (N_19968,N_11141,N_13801);
nor U19969 (N_19969,N_12543,N_11271);
nor U19970 (N_19970,N_11255,N_12009);
nand U19971 (N_19971,N_12949,N_10812);
nand U19972 (N_19972,N_11083,N_13394);
nand U19973 (N_19973,N_11672,N_11148);
or U19974 (N_19974,N_14904,N_13884);
nor U19975 (N_19975,N_14557,N_14896);
and U19976 (N_19976,N_11719,N_10122);
and U19977 (N_19977,N_11346,N_12690);
or U19978 (N_19978,N_14120,N_13173);
nand U19979 (N_19979,N_10334,N_12264);
nor U19980 (N_19980,N_11128,N_12289);
nand U19981 (N_19981,N_12748,N_11833);
and U19982 (N_19982,N_12663,N_10553);
or U19983 (N_19983,N_11336,N_14753);
nor U19984 (N_19984,N_11279,N_14313);
and U19985 (N_19985,N_10723,N_10365);
nor U19986 (N_19986,N_10367,N_14327);
or U19987 (N_19987,N_14082,N_11146);
and U19988 (N_19988,N_10816,N_10436);
and U19989 (N_19989,N_14382,N_12984);
xor U19990 (N_19990,N_10718,N_13163);
nor U19991 (N_19991,N_14497,N_13025);
or U19992 (N_19992,N_12340,N_11052);
and U19993 (N_19993,N_14649,N_10124);
nand U19994 (N_19994,N_13207,N_14183);
xor U19995 (N_19995,N_12011,N_13530);
nor U19996 (N_19996,N_12978,N_14395);
nand U19997 (N_19997,N_14530,N_13466);
and U19998 (N_19998,N_11251,N_13301);
nand U19999 (N_19999,N_10808,N_14402);
nand U20000 (N_20000,N_17213,N_16005);
and U20001 (N_20001,N_17734,N_16776);
nor U20002 (N_20002,N_18736,N_18142);
nor U20003 (N_20003,N_19616,N_16113);
or U20004 (N_20004,N_18241,N_19599);
nor U20005 (N_20005,N_19308,N_15477);
nand U20006 (N_20006,N_18308,N_18845);
or U20007 (N_20007,N_16421,N_17441);
nor U20008 (N_20008,N_17295,N_17283);
nor U20009 (N_20009,N_19327,N_18115);
nor U20010 (N_20010,N_19958,N_19809);
or U20011 (N_20011,N_15028,N_19148);
nor U20012 (N_20012,N_17942,N_18776);
nand U20013 (N_20013,N_16168,N_15607);
or U20014 (N_20014,N_18791,N_19498);
or U20015 (N_20015,N_15990,N_16226);
and U20016 (N_20016,N_17586,N_16112);
nor U20017 (N_20017,N_18177,N_18723);
and U20018 (N_20018,N_15219,N_19807);
nand U20019 (N_20019,N_15122,N_15094);
or U20020 (N_20020,N_15237,N_16433);
nand U20021 (N_20021,N_18541,N_17845);
or U20022 (N_20022,N_16396,N_15698);
nor U20023 (N_20023,N_19310,N_19132);
nand U20024 (N_20024,N_19014,N_16809);
or U20025 (N_20025,N_15846,N_18163);
nor U20026 (N_20026,N_15820,N_17137);
or U20027 (N_20027,N_15913,N_18173);
nor U20028 (N_20028,N_18051,N_19411);
xnor U20029 (N_20029,N_19403,N_16467);
nor U20030 (N_20030,N_18273,N_19072);
or U20031 (N_20031,N_15352,N_15433);
nand U20032 (N_20032,N_18571,N_17450);
or U20033 (N_20033,N_15946,N_16419);
nand U20034 (N_20034,N_15241,N_15210);
nor U20035 (N_20035,N_16294,N_15183);
nor U20036 (N_20036,N_19993,N_19284);
and U20037 (N_20037,N_19622,N_19100);
or U20038 (N_20038,N_18014,N_18963);
or U20039 (N_20039,N_19042,N_18487);
nor U20040 (N_20040,N_19026,N_18888);
xnor U20041 (N_20041,N_17689,N_16652);
or U20042 (N_20042,N_15144,N_18456);
and U20043 (N_20043,N_15888,N_18225);
or U20044 (N_20044,N_15484,N_16766);
nor U20045 (N_20045,N_19409,N_16637);
and U20046 (N_20046,N_15822,N_16519);
or U20047 (N_20047,N_16430,N_17403);
and U20048 (N_20048,N_17716,N_16574);
and U20049 (N_20049,N_15106,N_15960);
nand U20050 (N_20050,N_17397,N_17454);
and U20051 (N_20051,N_18559,N_18580);
nor U20052 (N_20052,N_17219,N_16784);
xnor U20053 (N_20053,N_17470,N_19111);
and U20054 (N_20054,N_16447,N_19768);
and U20055 (N_20055,N_18777,N_15032);
and U20056 (N_20056,N_17132,N_16144);
nand U20057 (N_20057,N_18378,N_17872);
or U20058 (N_20058,N_15489,N_19707);
nand U20059 (N_20059,N_15542,N_15162);
nand U20060 (N_20060,N_19461,N_19377);
nand U20061 (N_20061,N_18140,N_16432);
xor U20062 (N_20062,N_19523,N_15998);
and U20063 (N_20063,N_15713,N_18203);
nor U20064 (N_20064,N_17810,N_18459);
nand U20065 (N_20065,N_17077,N_15936);
and U20066 (N_20066,N_17147,N_15430);
or U20067 (N_20067,N_16231,N_18762);
nor U20068 (N_20068,N_16987,N_16427);
or U20069 (N_20069,N_18884,N_16928);
nand U20070 (N_20070,N_19397,N_19511);
or U20071 (N_20071,N_19580,N_16371);
nand U20072 (N_20072,N_15573,N_16364);
nor U20073 (N_20073,N_17442,N_16462);
or U20074 (N_20074,N_18620,N_18090);
or U20075 (N_20075,N_18385,N_18625);
or U20076 (N_20076,N_16331,N_19080);
nand U20077 (N_20077,N_17495,N_15073);
and U20078 (N_20078,N_19277,N_16358);
and U20079 (N_20079,N_19812,N_16434);
or U20080 (N_20080,N_15864,N_18712);
nor U20081 (N_20081,N_15858,N_19683);
nor U20082 (N_20082,N_18549,N_15746);
or U20083 (N_20083,N_19486,N_18169);
or U20084 (N_20084,N_17852,N_16448);
nor U20085 (N_20085,N_19475,N_18186);
and U20086 (N_20086,N_16191,N_16520);
and U20087 (N_20087,N_19384,N_18619);
nor U20088 (N_20088,N_15506,N_16444);
or U20089 (N_20089,N_16835,N_16667);
nor U20090 (N_20090,N_19542,N_19820);
or U20091 (N_20091,N_19399,N_19151);
xnor U20092 (N_20092,N_16913,N_15728);
nor U20093 (N_20093,N_15581,N_18413);
nor U20094 (N_20094,N_17879,N_19764);
or U20095 (N_20095,N_16681,N_16295);
nand U20096 (N_20096,N_17404,N_16536);
or U20097 (N_20097,N_15070,N_16685);
or U20098 (N_20098,N_18015,N_17655);
nor U20099 (N_20099,N_17264,N_16644);
or U20100 (N_20100,N_18281,N_17656);
nand U20101 (N_20101,N_15344,N_16618);
xnor U20102 (N_20102,N_18248,N_17573);
or U20103 (N_20103,N_19472,N_17739);
or U20104 (N_20104,N_18836,N_15103);
nand U20105 (N_20105,N_18893,N_18997);
nor U20106 (N_20106,N_19601,N_15969);
and U20107 (N_20107,N_17416,N_18697);
and U20108 (N_20108,N_18563,N_17850);
nand U20109 (N_20109,N_19126,N_15751);
nand U20110 (N_20110,N_16587,N_16834);
nor U20111 (N_20111,N_17233,N_18815);
or U20112 (N_20112,N_15035,N_15838);
nor U20113 (N_20113,N_19389,N_19861);
or U20114 (N_20114,N_17374,N_15526);
and U20115 (N_20115,N_19602,N_18551);
or U20116 (N_20116,N_15499,N_15608);
nand U20117 (N_20117,N_15671,N_17224);
or U20118 (N_20118,N_15686,N_15901);
nor U20119 (N_20119,N_17317,N_16489);
nand U20120 (N_20120,N_19655,N_15656);
nor U20121 (N_20121,N_16490,N_18605);
nand U20122 (N_20122,N_17535,N_17747);
nor U20123 (N_20123,N_18566,N_17697);
xor U20124 (N_20124,N_17835,N_17856);
nor U20125 (N_20125,N_15923,N_15668);
or U20126 (N_20126,N_19125,N_16951);
or U20127 (N_20127,N_17510,N_16334);
xnor U20128 (N_20128,N_19445,N_16690);
or U20129 (N_20129,N_18767,N_18759);
nand U20130 (N_20130,N_17136,N_18309);
nand U20131 (N_20131,N_17630,N_17103);
and U20132 (N_20132,N_15365,N_16515);
nor U20133 (N_20133,N_15918,N_18164);
nor U20134 (N_20134,N_16104,N_18363);
and U20135 (N_20135,N_16407,N_16084);
or U20136 (N_20136,N_16125,N_19033);
nand U20137 (N_20137,N_19496,N_19468);
or U20138 (N_20138,N_16418,N_17309);
xor U20139 (N_20139,N_19907,N_17173);
or U20140 (N_20140,N_17844,N_18264);
nand U20141 (N_20141,N_18584,N_17038);
xor U20142 (N_20142,N_17434,N_15112);
xnor U20143 (N_20143,N_17139,N_18381);
nor U20144 (N_20144,N_16038,N_17190);
nor U20145 (N_20145,N_18489,N_17811);
xor U20146 (N_20146,N_15143,N_16260);
nand U20147 (N_20147,N_19973,N_19423);
or U20148 (N_20148,N_15777,N_18864);
nand U20149 (N_20149,N_16968,N_17994);
and U20150 (N_20150,N_16789,N_18665);
or U20151 (N_20151,N_17800,N_16127);
xor U20152 (N_20152,N_19329,N_15222);
or U20153 (N_20153,N_15745,N_17271);
and U20154 (N_20154,N_18301,N_17832);
nand U20155 (N_20155,N_19871,N_17609);
and U20156 (N_20156,N_18906,N_17105);
or U20157 (N_20157,N_17154,N_18262);
or U20158 (N_20158,N_16889,N_19331);
nand U20159 (N_20159,N_19375,N_18590);
or U20160 (N_20160,N_16454,N_19909);
nand U20161 (N_20161,N_16623,N_15235);
xnor U20162 (N_20162,N_19571,N_18195);
or U20163 (N_20163,N_18856,N_18054);
or U20164 (N_20164,N_17830,N_15218);
or U20165 (N_20165,N_18480,N_16428);
and U20166 (N_20166,N_19699,N_17569);
or U20167 (N_20167,N_17731,N_17242);
and U20168 (N_20168,N_17097,N_15984);
xor U20169 (N_20169,N_18517,N_15709);
nor U20170 (N_20170,N_16000,N_18843);
nand U20171 (N_20171,N_17461,N_17071);
nor U20172 (N_20172,N_17414,N_18303);
nand U20173 (N_20173,N_17003,N_15059);
nor U20174 (N_20174,N_19674,N_16582);
and U20175 (N_20175,N_15599,N_16881);
nor U20176 (N_20176,N_19902,N_18438);
or U20177 (N_20177,N_19653,N_16675);
or U20178 (N_20178,N_18630,N_15973);
or U20179 (N_20179,N_18387,N_19893);
or U20180 (N_20180,N_18131,N_16500);
nor U20181 (N_20181,N_15253,N_18391);
and U20182 (N_20182,N_15403,N_19933);
or U20183 (N_20183,N_19345,N_18276);
nand U20184 (N_20184,N_16254,N_17983);
xnor U20185 (N_20185,N_15940,N_19049);
nand U20186 (N_20186,N_18465,N_17817);
nor U20187 (N_20187,N_19235,N_17289);
or U20188 (N_20188,N_17333,N_16716);
nand U20189 (N_20189,N_15481,N_16458);
or U20190 (N_20190,N_18933,N_15322);
or U20191 (N_20191,N_16341,N_19165);
nand U20192 (N_20192,N_16643,N_19927);
and U20193 (N_20193,N_19695,N_19474);
or U20194 (N_20194,N_18356,N_17316);
and U20195 (N_20195,N_15287,N_16629);
nor U20196 (N_20196,N_16793,N_15125);
or U20197 (N_20197,N_15985,N_17758);
nand U20198 (N_20198,N_15232,N_16631);
nor U20199 (N_20199,N_18778,N_19478);
nand U20200 (N_20200,N_17669,N_17618);
xor U20201 (N_20201,N_17371,N_19766);
xnor U20202 (N_20202,N_19649,N_15999);
nor U20203 (N_20203,N_17914,N_16807);
or U20204 (N_20204,N_17590,N_15958);
nand U20205 (N_20205,N_17700,N_17883);
or U20206 (N_20206,N_19879,N_16514);
nand U20207 (N_20207,N_15342,N_15531);
nand U20208 (N_20208,N_15332,N_16128);
nor U20209 (N_20209,N_18831,N_15251);
or U20210 (N_20210,N_17318,N_15646);
nand U20211 (N_20211,N_16921,N_16734);
or U20212 (N_20212,N_19150,N_15680);
nor U20213 (N_20213,N_16501,N_15217);
and U20214 (N_20214,N_16981,N_19174);
nor U20215 (N_20215,N_17762,N_19913);
and U20216 (N_20216,N_19306,N_19037);
nor U20217 (N_20217,N_18467,N_17073);
nor U20218 (N_20218,N_17534,N_18020);
or U20219 (N_20219,N_18372,N_19328);
nand U20220 (N_20220,N_17964,N_19212);
or U20221 (N_20221,N_18261,N_19206);
nor U20222 (N_20222,N_18609,N_15691);
and U20223 (N_20223,N_19758,N_15610);
nand U20224 (N_20224,N_18875,N_15196);
nand U20225 (N_20225,N_17620,N_16692);
xor U20226 (N_20226,N_16126,N_16468);
nand U20227 (N_20227,N_19581,N_15429);
nand U20228 (N_20228,N_19057,N_19684);
nor U20229 (N_20229,N_18801,N_19842);
nor U20230 (N_20230,N_15245,N_15133);
nor U20231 (N_20231,N_18962,N_19263);
and U20232 (N_20232,N_17598,N_16062);
and U20233 (N_20233,N_17662,N_18497);
nand U20234 (N_20234,N_15571,N_16588);
or U20235 (N_20235,N_16886,N_18122);
or U20236 (N_20236,N_18932,N_17639);
and U20237 (N_20237,N_17388,N_18221);
and U20238 (N_20238,N_19662,N_17692);
xor U20239 (N_20239,N_19422,N_15426);
or U20240 (N_20240,N_18439,N_18038);
and U20241 (N_20241,N_17338,N_15009);
nand U20242 (N_20242,N_15464,N_16121);
xnor U20243 (N_20243,N_18857,N_16831);
xnor U20244 (N_20244,N_18855,N_18751);
nand U20245 (N_20245,N_15362,N_15509);
nand U20246 (N_20246,N_17702,N_18735);
or U20247 (N_20247,N_15712,N_18573);
and U20248 (N_20248,N_16336,N_19552);
nor U20249 (N_20249,N_17542,N_17650);
or U20250 (N_20250,N_17440,N_15215);
and U20251 (N_20251,N_18799,N_18501);
or U20252 (N_20252,N_16597,N_17214);
or U20253 (N_20253,N_15965,N_15694);
or U20254 (N_20254,N_18114,N_15749);
nor U20255 (N_20255,N_17140,N_18642);
nor U20256 (N_20256,N_16930,N_18041);
or U20257 (N_20257,N_15517,N_17538);
nor U20258 (N_20258,N_17917,N_18513);
nor U20259 (N_20259,N_19260,N_19210);
or U20260 (N_20260,N_17562,N_18505);
xor U20261 (N_20261,N_15737,N_17217);
nor U20262 (N_20262,N_16204,N_19387);
and U20263 (N_20263,N_17250,N_16552);
xnor U20264 (N_20264,N_15340,N_18327);
nor U20265 (N_20265,N_15769,N_16924);
nand U20266 (N_20266,N_17096,N_15663);
nand U20267 (N_20267,N_18398,N_17059);
nand U20268 (N_20268,N_18389,N_19005);
or U20269 (N_20269,N_19234,N_16978);
xnor U20270 (N_20270,N_15812,N_18362);
and U20271 (N_20271,N_19518,N_15229);
nor U20272 (N_20272,N_16292,N_19921);
and U20273 (N_20273,N_19429,N_15205);
nor U20274 (N_20274,N_19124,N_19681);
and U20275 (N_20275,N_16081,N_16954);
or U20276 (N_20276,N_16869,N_15598);
or U20277 (N_20277,N_15716,N_15213);
or U20278 (N_20278,N_18427,N_15800);
nor U20279 (N_20279,N_18616,N_15279);
nand U20280 (N_20280,N_18833,N_19245);
and U20281 (N_20281,N_16449,N_16155);
nand U20282 (N_20282,N_18253,N_17381);
xnor U20283 (N_20283,N_17089,N_16170);
or U20284 (N_20284,N_16586,N_16946);
xnor U20285 (N_20285,N_19962,N_19451);
and U20286 (N_20286,N_18190,N_19757);
or U20287 (N_20287,N_18556,N_15091);
nand U20288 (N_20288,N_17952,N_18271);
and U20289 (N_20289,N_19198,N_16083);
and U20290 (N_20290,N_16787,N_17505);
and U20291 (N_20291,N_18025,N_18560);
nor U20292 (N_20292,N_19597,N_15117);
nor U20293 (N_20293,N_17439,N_18539);
nor U20294 (N_20294,N_16518,N_19368);
and U20295 (N_20295,N_19173,N_18034);
xnor U20296 (N_20296,N_16939,N_18508);
and U20297 (N_20297,N_16306,N_18636);
and U20298 (N_20298,N_17298,N_17910);
and U20299 (N_20299,N_18550,N_19313);
xnor U20300 (N_20300,N_15078,N_16145);
nand U20301 (N_20301,N_19023,N_18087);
nand U20302 (N_20302,N_17429,N_18670);
nand U20303 (N_20303,N_19142,N_15977);
nand U20304 (N_20304,N_15718,N_16989);
nor U20305 (N_20305,N_16542,N_17592);
nor U20306 (N_20306,N_15095,N_15634);
nor U20307 (N_20307,N_15051,N_18939);
nand U20308 (N_20308,N_16510,N_15371);
or U20309 (N_20309,N_16122,N_19894);
and U20310 (N_20310,N_16699,N_18604);
nand U20311 (N_20311,N_18078,N_18468);
or U20312 (N_20312,N_18184,N_17045);
and U20313 (N_20313,N_16953,N_15620);
nand U20314 (N_20314,N_17902,N_15413);
or U20315 (N_20315,N_18204,N_18816);
and U20316 (N_20316,N_15184,N_15267);
and U20317 (N_20317,N_17972,N_16680);
or U20318 (N_20318,N_19860,N_17085);
or U20319 (N_20319,N_18607,N_19841);
nand U20320 (N_20320,N_17988,N_17194);
or U20321 (N_20321,N_16480,N_18804);
nand U20322 (N_20322,N_16821,N_15508);
nand U20323 (N_20323,N_18249,N_19529);
nor U20324 (N_20324,N_17130,N_15919);
nand U20325 (N_20325,N_17539,N_18355);
or U20326 (N_20326,N_17030,N_18237);
nor U20327 (N_20327,N_16992,N_17548);
and U20328 (N_20328,N_17612,N_18202);
nor U20329 (N_20329,N_16002,N_19742);
xor U20330 (N_20330,N_18229,N_15804);
nor U20331 (N_20331,N_18490,N_16949);
or U20332 (N_20332,N_19577,N_19904);
nand U20333 (N_20333,N_18943,N_18012);
nand U20334 (N_20334,N_17499,N_17978);
xnor U20335 (N_20335,N_17049,N_18082);
and U20336 (N_20336,N_16740,N_16641);
nand U20337 (N_20337,N_16197,N_18023);
nor U20338 (N_20338,N_17961,N_18265);
and U20339 (N_20339,N_15724,N_17325);
nand U20340 (N_20340,N_16134,N_17960);
or U20341 (N_20341,N_15040,N_17293);
nor U20342 (N_20342,N_15087,N_19781);
nor U20343 (N_20343,N_19554,N_19952);
or U20344 (N_20344,N_18294,N_18737);
and U20345 (N_20345,N_17476,N_19876);
and U20346 (N_20346,N_16980,N_18645);
and U20347 (N_20347,N_17890,N_15714);
nor U20348 (N_20348,N_16838,N_17710);
nand U20349 (N_20349,N_16232,N_16902);
xor U20350 (N_20350,N_15981,N_15136);
nor U20351 (N_20351,N_16705,N_16620);
and U20352 (N_20352,N_18311,N_17659);
xnor U20353 (N_20353,N_15052,N_15900);
and U20354 (N_20354,N_19532,N_18971);
xor U20355 (N_20355,N_18935,N_15808);
xnor U20356 (N_20356,N_19066,N_19382);
nor U20357 (N_20357,N_16103,N_18522);
or U20358 (N_20358,N_15453,N_16593);
nand U20359 (N_20359,N_15832,N_18315);
nor U20360 (N_20360,N_18805,N_17649);
and U20361 (N_20361,N_19538,N_15639);
xor U20362 (N_20362,N_19827,N_17080);
nand U20363 (N_20363,N_16193,N_18069);
xnor U20364 (N_20364,N_18111,N_17272);
and U20365 (N_20365,N_18384,N_15869);
or U20366 (N_20366,N_16321,N_17243);
or U20367 (N_20367,N_17435,N_17153);
and U20368 (N_20368,N_19324,N_19319);
xnor U20369 (N_20369,N_19546,N_18827);
nor U20370 (N_20370,N_16004,N_15932);
and U20371 (N_20371,N_17377,N_16516);
nor U20372 (N_20372,N_16325,N_15329);
nor U20373 (N_20373,N_17195,N_18710);
xnor U20374 (N_20374,N_17491,N_18651);
nor U20375 (N_20375,N_16309,N_16074);
or U20376 (N_20376,N_17232,N_17922);
nand U20377 (N_20377,N_15565,N_17492);
xnor U20378 (N_20378,N_15039,N_18344);
or U20379 (N_20379,N_15549,N_19143);
and U20380 (N_20380,N_17421,N_15283);
and U20381 (N_20381,N_19975,N_15443);
and U20382 (N_20382,N_15313,N_19394);
xnor U20383 (N_20383,N_15814,N_16267);
or U20384 (N_20384,N_16075,N_17806);
or U20385 (N_20385,N_16739,N_17965);
or U20386 (N_20386,N_16072,N_17009);
xor U20387 (N_20387,N_17544,N_16799);
nand U20388 (N_20388,N_16967,N_19706);
nor U20389 (N_20389,N_19633,N_17028);
and U20390 (N_20390,N_17768,N_19205);
xor U20391 (N_20391,N_16572,N_18416);
and U20392 (N_20392,N_17724,N_19054);
and U20393 (N_20393,N_19579,N_18085);
nor U20394 (N_20394,N_17876,N_19339);
xor U20395 (N_20395,N_15273,N_16042);
or U20396 (N_20396,N_18916,N_18088);
nor U20397 (N_20397,N_18904,N_19756);
nand U20398 (N_20398,N_16357,N_15991);
and U20399 (N_20399,N_19925,N_15816);
nor U20400 (N_20400,N_19795,N_19463);
xor U20401 (N_20401,N_19365,N_19901);
xor U20402 (N_20402,N_18162,N_17407);
nor U20403 (N_20403,N_15450,N_17340);
nor U20404 (N_20404,N_19223,N_19330);
or U20405 (N_20405,N_15881,N_18537);
and U20406 (N_20406,N_19318,N_15894);
nand U20407 (N_20407,N_19859,N_19116);
or U20408 (N_20408,N_15446,N_17726);
nand U20409 (N_20409,N_17935,N_15361);
and U20410 (N_20410,N_15711,N_16061);
xor U20411 (N_20411,N_16288,N_16340);
nand U20412 (N_20412,N_16366,N_16940);
or U20413 (N_20413,N_18320,N_15791);
nand U20414 (N_20414,N_15621,N_19469);
nand U20415 (N_20415,N_19122,N_18570);
nor U20416 (N_20416,N_19942,N_18101);
and U20417 (N_20417,N_16848,N_19018);
nor U20418 (N_20418,N_19686,N_19986);
nand U20419 (N_20419,N_15090,N_19340);
nor U20420 (N_20420,N_19715,N_17344);
nand U20421 (N_20421,N_15569,N_16669);
nand U20422 (N_20422,N_17522,N_18353);
or U20423 (N_20423,N_19976,N_17594);
and U20424 (N_20424,N_15725,N_15892);
and U20425 (N_20425,N_15418,N_17993);
nand U20426 (N_20426,N_16596,N_16132);
nand U20427 (N_20427,N_18157,N_19484);
nor U20428 (N_20428,N_19821,N_19385);
nor U20429 (N_20429,N_19296,N_19584);
or U20430 (N_20430,N_15314,N_15707);
nor U20431 (N_20431,N_18175,N_16355);
or U20432 (N_20432,N_16655,N_15425);
and U20433 (N_20433,N_19839,N_16849);
xnor U20434 (N_20434,N_16211,N_15911);
and U20435 (N_20435,N_15293,N_19883);
nor U20436 (N_20436,N_15319,N_19572);
and U20437 (N_20437,N_18821,N_19374);
xor U20438 (N_20438,N_17300,N_18510);
nand U20439 (N_20439,N_15783,N_17711);
and U20440 (N_20440,N_19240,N_19863);
xnor U20441 (N_20441,N_17629,N_17842);
nor U20442 (N_20442,N_19275,N_19170);
or U20443 (N_20443,N_15114,N_18673);
nand U20444 (N_20444,N_15355,N_15645);
or U20445 (N_20445,N_16877,N_17012);
and U20446 (N_20446,N_18181,N_16818);
nor U20447 (N_20447,N_17525,N_17412);
xnor U20448 (N_20448,N_18639,N_15030);
nand U20449 (N_20449,N_18742,N_18252);
and U20450 (N_20450,N_18881,N_16408);
or U20451 (N_20451,N_16365,N_18703);
xnor U20452 (N_20452,N_15614,N_17392);
or U20453 (N_20453,N_18552,N_18614);
and U20454 (N_20454,N_19970,N_17670);
and U20455 (N_20455,N_19494,N_19104);
and U20456 (N_20456,N_18364,N_16386);
nor U20457 (N_20457,N_17991,N_18950);
and U20458 (N_20458,N_17694,N_19858);
and U20459 (N_20459,N_17064,N_19343);
and U20460 (N_20460,N_16811,N_19835);
xor U20461 (N_20461,N_18083,N_16673);
nand U20462 (N_20462,N_17368,N_19844);
or U20463 (N_20463,N_16639,N_19785);
nor U20464 (N_20464,N_15334,N_17123);
or U20465 (N_20465,N_17036,N_16162);
nor U20466 (N_20466,N_16617,N_16099);
nor U20467 (N_20467,N_17828,N_18366);
and U20468 (N_20468,N_17688,N_17164);
and U20469 (N_20469,N_18495,N_19522);
nand U20470 (N_20470,N_18464,N_16806);
xnor U20471 (N_20471,N_19888,N_16636);
nand U20472 (N_20472,N_19979,N_16106);
or U20473 (N_20473,N_16626,N_17120);
nand U20474 (N_20474,N_18841,N_19354);
nor U20475 (N_20475,N_16361,N_16014);
nor U20476 (N_20476,N_18008,N_17487);
nand U20477 (N_20477,N_16320,N_17322);
and U20478 (N_20478,N_18727,N_18530);
or U20479 (N_20479,N_16151,N_16303);
and U20480 (N_20480,N_18418,N_19433);
nand U20481 (N_20481,N_15843,N_19735);
or U20482 (N_20482,N_16863,N_18473);
or U20483 (N_20483,N_17905,N_19629);
or U20484 (N_20484,N_18455,N_16771);
or U20485 (N_20485,N_17751,N_17866);
nor U20486 (N_20486,N_18268,N_16815);
and U20487 (N_20487,N_16329,N_15448);
and U20488 (N_20488,N_16948,N_16892);
or U20489 (N_20489,N_15185,N_18089);
nor U20490 (N_20490,N_19246,N_18733);
nor U20491 (N_20491,N_16095,N_17924);
nor U20492 (N_20492,N_19039,N_18696);
and U20493 (N_20493,N_17446,N_16794);
nand U20494 (N_20494,N_15294,N_18167);
nand U20495 (N_20495,N_15891,N_17827);
nand U20496 (N_20496,N_19175,N_19344);
and U20497 (N_20497,N_17170,N_17033);
and U20498 (N_20498,N_18282,N_16308);
or U20499 (N_20499,N_19407,N_15240);
and U20500 (N_20500,N_18618,N_15105);
nand U20501 (N_20501,N_15770,N_17860);
nor U20502 (N_20502,N_15616,N_16141);
nor U20503 (N_20503,N_18374,N_16715);
or U20504 (N_20504,N_16965,N_16659);
or U20505 (N_20505,N_18137,N_16737);
xnor U20506 (N_20506,N_18341,N_17748);
and U20507 (N_20507,N_15049,N_18622);
nor U20508 (N_20508,N_18141,N_19797);
nand U20509 (N_20509,N_18870,N_15742);
nand U20510 (N_20510,N_18220,N_18756);
nand U20511 (N_20511,N_17472,N_16547);
xnor U20512 (N_20512,N_16833,N_17900);
nor U20513 (N_20513,N_15633,N_18685);
nand U20514 (N_20514,N_17501,N_18745);
and U20515 (N_20515,N_16654,N_18135);
or U20516 (N_20516,N_19378,N_19218);
nand U20517 (N_20517,N_18879,N_18409);
and U20518 (N_20518,N_16146,N_19227);
nand U20519 (N_20519,N_17305,N_16727);
nor U20520 (N_20520,N_15071,N_19563);
and U20521 (N_20521,N_19652,N_15422);
or U20522 (N_20522,N_17920,N_17216);
nor U20523 (N_20523,N_16240,N_15139);
or U20524 (N_20524,N_19444,N_15497);
nand U20525 (N_20525,N_19673,N_16741);
and U20526 (N_20526,N_19698,N_19931);
nor U20527 (N_20527,N_19065,N_18930);
nor U20528 (N_20528,N_18747,N_17849);
nor U20529 (N_20529,N_16098,N_18538);
xor U20530 (N_20530,N_16710,N_18424);
or U20531 (N_20531,N_19219,N_18451);
xor U20532 (N_20532,N_16595,N_19261);
xnor U20533 (N_20533,N_19818,N_17261);
nand U20534 (N_20534,N_19038,N_17366);
and U20535 (N_20535,N_15138,N_15873);
xnor U20536 (N_20536,N_15700,N_15098);
nor U20537 (N_20537,N_15524,N_15527);
or U20538 (N_20538,N_16161,N_17857);
nand U20539 (N_20539,N_19015,N_15930);
xnor U20540 (N_20540,N_19743,N_15895);
and U20541 (N_20541,N_17193,N_15016);
nor U20542 (N_20542,N_17483,N_19914);
or U20543 (N_20543,N_19421,N_17926);
nor U20544 (N_20544,N_17353,N_18231);
and U20545 (N_20545,N_16114,N_18178);
nand U20546 (N_20546,N_16638,N_18708);
nor U20547 (N_20547,N_18989,N_17347);
nor U20548 (N_20548,N_17868,N_15710);
and U20549 (N_20549,N_18867,N_19789);
nor U20550 (N_20550,N_17373,N_18773);
nor U20551 (N_20551,N_19201,N_15779);
or U20552 (N_20552,N_19321,N_17750);
or U20553 (N_20553,N_16250,N_16688);
or U20554 (N_20554,N_15950,N_15395);
xor U20555 (N_20555,N_15866,N_19916);
nor U20556 (N_20556,N_18102,N_17053);
nor U20557 (N_20557,N_16909,N_18212);
or U20558 (N_20558,N_15175,N_17658);
or U20559 (N_20559,N_17613,N_18478);
nor U20560 (N_20560,N_15957,N_17011);
or U20561 (N_20561,N_17545,N_15494);
nor U20562 (N_20562,N_16938,N_15297);
nand U20563 (N_20563,N_18994,N_18748);
nor U20564 (N_20564,N_17854,N_17129);
or U20565 (N_20565,N_15478,N_18689);
and U20566 (N_20566,N_17676,N_18535);
nand U20567 (N_20567,N_18000,N_18275);
and U20568 (N_20568,N_15910,N_15993);
nor U20569 (N_20569,N_19960,N_19846);
nor U20570 (N_20570,N_17415,N_17449);
or U20571 (N_20571,N_16663,N_16389);
nand U20572 (N_20572,N_15720,N_16936);
or U20573 (N_20573,N_19658,N_15255);
nor U20574 (N_20574,N_16060,N_19544);
or U20575 (N_20575,N_19297,N_16017);
nor U20576 (N_20576,N_16952,N_16410);
or U20577 (N_20577,N_16786,N_16651);
or U20578 (N_20578,N_15417,N_17098);
nand U20579 (N_20579,N_15131,N_16435);
and U20580 (N_20580,N_16749,N_17266);
nand U20581 (N_20581,N_17026,N_19322);
or U20582 (N_20582,N_18100,N_16369);
xnor U20583 (N_20583,N_18844,N_15301);
nand U20584 (N_20584,N_17804,N_15545);
and U20585 (N_20585,N_18976,N_18717);
and U20586 (N_20586,N_17732,N_19843);
nand U20587 (N_20587,N_15225,N_17228);
xnor U20588 (N_20588,N_18575,N_15584);
and U20589 (N_20589,N_19947,N_19643);
nand U20590 (N_20590,N_19404,N_15522);
or U20591 (N_20591,N_17941,N_18842);
and U20592 (N_20592,N_16290,N_19667);
and U20593 (N_20593,N_16350,N_19158);
and U20594 (N_20594,N_19528,N_19691);
nor U20595 (N_20595,N_18431,N_16660);
or U20596 (N_20596,N_16962,N_19615);
nor U20597 (N_20597,N_19505,N_15916);
nand U20598 (N_20598,N_17183,N_18149);
nand U20599 (N_20599,N_17599,N_16744);
nand U20600 (N_20600,N_19560,N_16843);
nand U20601 (N_20601,N_19853,N_17908);
xnor U20602 (N_20602,N_18880,N_17721);
or U20603 (N_20603,N_16379,N_15802);
or U20604 (N_20604,N_16565,N_15756);
nand U20605 (N_20605,N_17126,N_16411);
and U20606 (N_20606,N_17042,N_18232);
and U20607 (N_20607,N_19156,N_16495);
nor U20608 (N_20608,N_15915,N_16496);
and U20609 (N_20609,N_18059,N_15321);
and U20610 (N_20610,N_16852,N_18030);
and U20611 (N_20611,N_15795,N_16278);
nand U20612 (N_20612,N_15104,N_15258);
xnor U20613 (N_20613,N_16874,N_17722);
nor U20614 (N_20614,N_18985,N_15757);
and U20615 (N_20615,N_18172,N_19262);
nand U20616 (N_20616,N_16266,N_18240);
or U20617 (N_20617,N_19228,N_18274);
nor U20618 (N_20618,N_19183,N_18222);
nor U20619 (N_20619,N_17803,N_19770);
and U20620 (N_20620,N_17568,N_18348);
nor U20621 (N_20621,N_19059,N_18958);
or U20622 (N_20622,N_19369,N_18610);
nand U20623 (N_20623,N_18124,N_16384);
nor U20624 (N_20624,N_18491,N_15992);
or U20625 (N_20625,N_18840,N_18547);
and U20626 (N_20626,N_15559,N_15111);
nand U20627 (N_20627,N_18433,N_17646);
nand U20628 (N_20628,N_15424,N_18227);
and U20629 (N_20629,N_15941,N_18048);
or U20630 (N_20630,N_15060,N_15763);
or U20631 (N_20631,N_19281,N_15951);
and U20632 (N_20632,N_15582,N_15023);
nand U20633 (N_20633,N_16845,N_17529);
xnor U20634 (N_20634,N_15818,N_16717);
nand U20635 (N_20635,N_17115,N_17241);
xnor U20636 (N_20636,N_19694,N_18898);
or U20637 (N_20637,N_16762,N_17135);
nor U20638 (N_20638,N_18545,N_15160);
and U20639 (N_20639,N_17307,N_16376);
nor U20640 (N_20640,N_16917,N_16612);
nand U20641 (N_20641,N_18084,N_15796);
and U20642 (N_20642,N_18046,N_17387);
nand U20643 (N_20643,N_17199,N_16120);
nor U20644 (N_20644,N_19603,N_17088);
and U20645 (N_20645,N_17391,N_17060);
nand U20646 (N_20646,N_15819,N_17358);
or U20647 (N_20647,N_17644,N_17553);
nor U20648 (N_20648,N_16054,N_15462);
or U20649 (N_20649,N_15652,N_17356);
or U20650 (N_20650,N_15989,N_19314);
nor U20651 (N_20651,N_18127,N_17282);
nand U20652 (N_20652,N_19427,N_18257);
nand U20653 (N_20653,N_19929,N_17884);
or U20654 (N_20654,N_17311,N_18587);
and U20655 (N_20655,N_17660,N_15211);
nand U20656 (N_20656,N_15170,N_19270);
nor U20657 (N_20657,N_19500,N_16093);
nor U20658 (N_20658,N_15702,N_18367);
and U20659 (N_20659,N_19459,N_16769);
or U20660 (N_20660,N_19437,N_19750);
or U20661 (N_20661,N_18925,N_16910);
or U20662 (N_20662,N_17046,N_16022);
nand U20663 (N_20663,N_17578,N_16380);
or U20664 (N_20664,N_17477,N_16820);
and U20665 (N_20665,N_19166,N_17774);
nand U20666 (N_20666,N_15788,N_17359);
nor U20667 (N_20667,N_19031,N_18405);
and U20668 (N_20668,N_17114,N_19220);
nand U20669 (N_20669,N_16102,N_17863);
nand U20670 (N_20670,N_15420,N_19922);
or U20671 (N_20671,N_18500,N_19082);
or U20672 (N_20672,N_16459,N_18644);
or U20673 (N_20673,N_18965,N_18216);
and U20674 (N_20674,N_15552,N_19114);
nand U20675 (N_20675,N_18116,N_15659);
or U20676 (N_20676,N_18612,N_15739);
and U20677 (N_20677,N_17118,N_16632);
or U20678 (N_20678,N_15212,N_15188);
or U20679 (N_20679,N_18613,N_16363);
nand U20680 (N_20680,N_18536,N_19790);
nor U20681 (N_20681,N_16304,N_19386);
nor U20682 (N_20682,N_18097,N_19096);
and U20683 (N_20683,N_17222,N_16453);
or U20684 (N_20684,N_19977,N_17962);
nand U20685 (N_20685,N_16019,N_15860);
or U20686 (N_20686,N_17229,N_18369);
or U20687 (N_20687,N_19293,N_16840);
xnor U20688 (N_20688,N_19596,N_17781);
or U20689 (N_20689,N_19355,N_15441);
and U20690 (N_20690,N_16998,N_15026);
or U20691 (N_20691,N_16855,N_17719);
nand U20692 (N_20692,N_15664,N_18346);
or U20693 (N_20693,N_17675,N_18694);
nand U20694 (N_20694,N_16607,N_17186);
nor U20695 (N_20695,N_17201,N_17648);
and U20696 (N_20696,N_15475,N_17430);
nand U20697 (N_20697,N_17141,N_19833);
nor U20698 (N_20698,N_17526,N_19147);
or U20699 (N_20699,N_18546,N_17755);
and U20700 (N_20700,N_18959,N_19779);
or U20701 (N_20701,N_15252,N_18992);
nand U20702 (N_20702,N_19963,N_17677);
xnor U20703 (N_20703,N_16990,N_16941);
and U20704 (N_20704,N_16217,N_17257);
or U20705 (N_20705,N_16964,N_16763);
nand U20706 (N_20706,N_15747,N_16167);
nor U20707 (N_20707,N_19696,N_19971);
xnor U20708 (N_20708,N_16533,N_15172);
nand U20709 (N_20709,N_19793,N_19168);
xnor U20710 (N_20710,N_15893,N_19055);
or U20711 (N_20711,N_19915,N_19252);
or U20712 (N_20712,N_17203,N_18053);
nor U20713 (N_20713,N_15473,N_18627);
or U20714 (N_20714,N_19892,N_15166);
or U20715 (N_20715,N_18244,N_19852);
xor U20716 (N_20716,N_19388,N_19177);
or U20717 (N_20717,N_15370,N_17280);
nor U20718 (N_20718,N_18668,N_19672);
nor U20719 (N_20719,N_18287,N_18170);
and U20720 (N_20720,N_16722,N_15740);
nand U20721 (N_20721,N_19559,N_17083);
and U20722 (N_20722,N_19027,N_16282);
or U20723 (N_20723,N_18897,N_19086);
or U20724 (N_20724,N_18862,N_19619);
nor U20725 (N_20725,N_19021,N_18589);
xnor U20726 (N_20726,N_17310,N_16234);
nand U20727 (N_20727,N_19533,N_15591);
and U20728 (N_20728,N_16856,N_19108);
or U20729 (N_20729,N_19515,N_15851);
nor U20730 (N_20730,N_19535,N_15084);
nand U20731 (N_20731,N_17192,N_19441);
nor U20732 (N_20732,N_18663,N_15945);
or U20733 (N_20733,N_19588,N_19642);
and U20734 (N_20734,N_15061,N_17063);
xor U20735 (N_20735,N_15474,N_19719);
nand U20736 (N_20736,N_15471,N_16731);
nor U20737 (N_20737,N_18741,N_19231);
and U20738 (N_20738,N_19146,N_16100);
nor U20739 (N_20739,N_18404,N_18878);
or U20740 (N_20740,N_17110,N_17248);
or U20741 (N_20741,N_15730,N_19624);
nand U20742 (N_20742,N_15833,N_18542);
nand U20743 (N_20743,N_15515,N_17382);
and U20744 (N_20744,N_18337,N_18136);
and U20745 (N_20745,N_16695,N_16559);
nor U20746 (N_20746,N_15320,N_18153);
nor U20747 (N_20747,N_18482,N_16569);
or U20748 (N_20748,N_19832,N_19551);
nand U20749 (N_20749,N_19102,N_15300);
and U20750 (N_20750,N_18915,N_19413);
and U20751 (N_20751,N_15525,N_17509);
or U20752 (N_20752,N_18514,N_17438);
nor U20753 (N_20753,N_15924,N_18106);
xnor U20754 (N_20754,N_17321,N_15528);
nor U20755 (N_20755,N_15341,N_15952);
nand U20756 (N_20756,N_19834,N_18013);
nor U20757 (N_20757,N_15003,N_18182);
nor U20758 (N_20758,N_16920,N_16816);
or U20759 (N_20759,N_18984,N_18349);
or U20760 (N_20760,N_18076,N_15632);
nor U20761 (N_20761,N_18251,N_15387);
nor U20762 (N_20762,N_18719,N_16362);
and U20763 (N_20763,N_19507,N_15379);
and U20764 (N_20764,N_17107,N_15336);
nor U20765 (N_20765,N_17235,N_19714);
or U20766 (N_20766,N_15556,N_16873);
or U20767 (N_20767,N_18796,N_15823);
or U20768 (N_20768,N_16788,N_17682);
or U20769 (N_20769,N_16756,N_18938);
nor U20770 (N_20770,N_17666,N_17519);
and U20771 (N_20771,N_17532,N_17463);
xnor U20772 (N_20772,N_17423,N_18811);
or U20773 (N_20773,N_16166,N_18569);
nand U20774 (N_20774,N_19928,N_17466);
or U20775 (N_20775,N_19885,N_15223);
nand U20776 (N_20776,N_17119,N_19995);
nand U20777 (N_20777,N_19782,N_16298);
or U20778 (N_20778,N_15576,N_16342);
nor U20779 (N_20779,N_19783,N_19088);
or U20780 (N_20780,N_15703,N_17744);
and U20781 (N_20781,N_19969,N_17899);
and U20782 (N_20782,N_18147,N_18223);
or U20783 (N_20783,N_17494,N_17869);
xnor U20784 (N_20784,N_18611,N_15244);
and U20785 (N_20785,N_16056,N_18057);
nand U20786 (N_20786,N_18434,N_19145);
nor U20787 (N_20787,N_19824,N_19557);
or U20788 (N_20788,N_19945,N_17693);
or U20789 (N_20789,N_17798,N_18518);
nor U20790 (N_20790,N_17819,N_18246);
nand U20791 (N_20791,N_18488,N_18907);
nand U20792 (N_20792,N_17484,N_15067);
or U20793 (N_20793,N_16602,N_16461);
nor U20794 (N_20794,N_18718,N_16517);
xnor U20795 (N_20795,N_19091,N_19051);
nand U20796 (N_20796,N_19233,N_19336);
and U20797 (N_20797,N_18621,N_19836);
and U20798 (N_20798,N_19483,N_19008);
or U20799 (N_20799,N_15767,N_17196);
nand U20800 (N_20800,N_18877,N_16752);
and U20801 (N_20801,N_17826,N_16018);
nand U20802 (N_20802,N_16284,N_17843);
nor U20803 (N_20803,N_15179,N_16301);
nand U20804 (N_20804,N_17507,N_15961);
nor U20805 (N_20805,N_16525,N_15909);
xor U20806 (N_20806,N_18033,N_19810);
xor U20807 (N_20807,N_19711,N_15053);
or U20808 (N_20808,N_17871,N_19489);
nor U20809 (N_20809,N_17684,N_17764);
nand U20810 (N_20810,N_19869,N_19391);
or U20811 (N_20811,N_16929,N_19604);
nor U20812 (N_20812,N_17823,N_19121);
nor U20813 (N_20813,N_17162,N_15844);
or U20814 (N_20814,N_19521,N_18144);
or U20815 (N_20815,N_18335,N_19360);
or U20816 (N_20816,N_15886,N_15914);
xnor U20817 (N_20817,N_18098,N_15583);
or U20818 (N_20818,N_15109,N_16390);
nor U20819 (N_20819,N_15415,N_18637);
xnor U20820 (N_20820,N_19716,N_16943);
xor U20821 (N_20821,N_16801,N_17680);
and U20822 (N_20822,N_15292,N_19119);
or U20823 (N_20823,N_17198,N_19083);
and U20824 (N_20824,N_15360,N_17623);
xnor U20825 (N_20825,N_15020,N_16318);
or U20826 (N_20826,N_18280,N_16589);
and U20827 (N_20827,N_17163,N_17607);
nand U20828 (N_20828,N_17807,N_19592);
or U20829 (N_20829,N_16630,N_18432);
nor U20830 (N_20830,N_19325,N_19357);
nor U20831 (N_20831,N_16378,N_18908);
nor U20832 (N_20832,N_15752,N_16222);
or U20833 (N_20833,N_15529,N_19561);
or U20834 (N_20834,N_17017,N_16252);
or U20835 (N_20835,N_17919,N_18370);
xnor U20836 (N_20836,N_15452,N_17839);
nand U20837 (N_20837,N_18396,N_16438);
and U20838 (N_20838,N_16925,N_15953);
and U20839 (N_20839,N_16876,N_16150);
and U20840 (N_20840,N_16333,N_15626);
xnor U20841 (N_20841,N_19341,N_15538);
xnor U20842 (N_20842,N_19333,N_19501);
nor U20843 (N_20843,N_16247,N_17363);
and U20844 (N_20844,N_16927,N_16828);
nand U20845 (N_20845,N_19193,N_15177);
nor U20846 (N_20846,N_18931,N_17636);
or U20847 (N_20847,N_18047,N_18080);
nand U20848 (N_20848,N_18753,N_19406);
or U20849 (N_20849,N_18732,N_15887);
or U20850 (N_20850,N_16347,N_17537);
and U20851 (N_20851,N_17308,N_17427);
nand U20852 (N_20852,N_16860,N_17306);
xnor U20853 (N_20853,N_17950,N_15590);
or U20854 (N_20854,N_15760,N_19607);
nand U20855 (N_20855,N_15054,N_15612);
and U20856 (N_20856,N_17372,N_17558);
nor U20857 (N_20857,N_16322,N_16571);
xor U20858 (N_20858,N_18940,N_18698);
xnor U20859 (N_20859,N_19047,N_19796);
nand U20860 (N_20860,N_15325,N_19733);
and U20861 (N_20861,N_16416,N_16944);
nand U20862 (N_20862,N_19752,N_19727);
nand U20863 (N_20863,N_15762,N_19583);
and U20864 (N_20864,N_18123,N_18218);
nor U20865 (N_20865,N_18603,N_17836);
and U20866 (N_20866,N_17290,N_15784);
nand U20867 (N_20867,N_17025,N_19738);
and U20868 (N_20868,N_16482,N_17174);
or U20869 (N_20869,N_19420,N_17622);
nor U20870 (N_20870,N_16212,N_16257);
or U20871 (N_20871,N_17002,N_18330);
nor U20872 (N_20872,N_17018,N_16352);
nand U20873 (N_20873,N_17733,N_18507);
or U20874 (N_20874,N_19548,N_18107);
nand U20875 (N_20875,N_15705,N_16697);
and U20876 (N_20876,N_17474,N_18926);
nor U20877 (N_20877,N_18449,N_18238);
nor U20878 (N_20878,N_19002,N_19910);
or U20879 (N_20879,N_17390,N_19787);
nand U20880 (N_20880,N_16445,N_17380);
nor U20881 (N_20881,N_19530,N_18110);
or U20882 (N_20882,N_19747,N_17995);
nor U20883 (N_20883,N_18035,N_18437);
nor U20884 (N_20884,N_18674,N_15047);
nor U20885 (N_20885,N_19857,N_17600);
and U20886 (N_20886,N_18492,N_18450);
nor U20887 (N_20887,N_18474,N_19393);
or U20888 (N_20888,N_19801,N_16774);
nor U20889 (N_20889,N_16725,N_18873);
and U20890 (N_20890,N_15119,N_19103);
nor U20891 (N_20891,N_17150,N_17615);
nand U20892 (N_20892,N_18561,N_19753);
nand U20893 (N_20893,N_15988,N_17954);
nand U20894 (N_20894,N_17263,N_15057);
nand U20895 (N_20895,N_17247,N_19516);
or U20896 (N_20896,N_16479,N_15034);
nor U20897 (N_20897,N_16906,N_17789);
nand U20898 (N_20898,N_18011,N_15872);
and U20899 (N_20899,N_15147,N_19991);
nand U20900 (N_20900,N_17771,N_15758);
or U20901 (N_20901,N_19432,N_18004);
or U20902 (N_20902,N_18528,N_16550);
or U20903 (N_20903,N_15794,N_15507);
nand U20904 (N_20904,N_15384,N_15701);
or U20905 (N_20905,N_17848,N_19813);
or U20906 (N_20906,N_16698,N_17498);
and U20907 (N_20907,N_17113,N_19084);
nand U20908 (N_20908,N_19666,N_15848);
and U20909 (N_20909,N_16314,N_19582);
and U20910 (N_20910,N_17645,N_15638);
xor U20911 (N_20911,N_19115,N_19455);
and U20912 (N_20912,N_15773,N_18105);
nor U20913 (N_20913,N_16983,N_18475);
or U20914 (N_20914,N_15163,N_19965);
and U20915 (N_20915,N_18829,N_17379);
or U20916 (N_20916,N_19802,N_16394);
nand U20917 (N_20917,N_17155,N_17533);
nor U20918 (N_20918,N_15906,N_15019);
and U20919 (N_20919,N_16723,N_16899);
and U20920 (N_20920,N_15504,N_17287);
or U20921 (N_20921,N_15406,N_16275);
and U20922 (N_20922,N_19182,N_15363);
or U20923 (N_20923,N_16176,N_15976);
and U20924 (N_20924,N_19274,N_17133);
or U20925 (N_20925,N_15001,N_15513);
nor U20926 (N_20926,N_19867,N_16265);
and U20927 (N_20927,N_17706,N_15080);
or U20928 (N_20928,N_15262,N_17445);
or U20929 (N_20929,N_17350,N_17209);
nand U20930 (N_20930,N_15904,N_19636);
and U20931 (N_20931,N_15727,N_18990);
nor U20932 (N_20932,N_16116,N_17979);
nand U20933 (N_20933,N_18006,N_15956);
or U20934 (N_20934,N_19216,N_17685);
and U20935 (N_20935,N_16105,N_17020);
or U20936 (N_20936,N_19668,N_19074);
and U20937 (N_20937,N_19414,N_18236);
or U20938 (N_20938,N_18032,N_16557);
nand U20939 (N_20939,N_16558,N_18338);
xor U20940 (N_20940,N_19076,N_16033);
nor U20941 (N_20941,N_16898,N_19936);
nor U20942 (N_20942,N_17517,N_16315);
or U20943 (N_20943,N_17904,N_16812);
nand U20944 (N_20944,N_18623,N_16139);
and U20945 (N_20945,N_15890,N_19739);
nor U20946 (N_20946,N_15676,N_19614);
xor U20947 (N_20947,N_18224,N_15574);
nor U20948 (N_20948,N_16891,N_15877);
or U20949 (N_20949,N_15378,N_17144);
nand U20950 (N_20950,N_18417,N_18125);
and U20951 (N_20951,N_17749,N_18155);
and U20952 (N_20952,N_15345,N_18039);
or U20953 (N_20953,N_19309,N_16931);
nor U20954 (N_20954,N_18928,N_19870);
nor U20955 (N_20955,N_19020,N_19638);
and U20956 (N_20956,N_16351,N_16273);
xnor U20957 (N_20957,N_16836,N_18574);
or U20958 (N_20958,N_17547,N_19266);
nand U20959 (N_20959,N_15679,N_19645);
or U20960 (N_20960,N_18399,N_19203);
and U20961 (N_20961,N_15089,N_19428);
and U20962 (N_20962,N_19265,N_19988);
or U20963 (N_20963,N_17055,N_16109);
nand U20964 (N_20964,N_17717,N_17086);
nor U20965 (N_20965,N_16847,N_19191);
and U20966 (N_20966,N_17953,N_16932);
nand U20967 (N_20967,N_15380,N_16779);
and U20968 (N_20968,N_17502,N_16661);
nor U20969 (N_20969,N_19644,N_19512);
and U20970 (N_20970,N_18104,N_15837);
xor U20971 (N_20971,N_15330,N_18838);
or U20972 (N_20972,N_15640,N_18109);
nand U20973 (N_20973,N_15726,N_18401);
or U20974 (N_20974,N_19258,N_18531);
or U20975 (N_20975,N_16417,N_17015);
and U20976 (N_20976,N_17455,N_15787);
and U20977 (N_20977,N_19688,N_15642);
nand U20978 (N_20978,N_16184,N_17791);
nor U20979 (N_20979,N_15250,N_17571);
nand U20980 (N_20980,N_17227,N_17109);
nand U20981 (N_20981,N_19278,N_18072);
nor U20982 (N_20982,N_17332,N_18192);
nor U20983 (N_20983,N_16460,N_15978);
nor U20984 (N_20984,N_16272,N_18918);
nand U20985 (N_20985,N_18070,N_18998);
nor U20986 (N_20986,N_19079,N_17408);
nor U20987 (N_20987,N_18839,N_17478);
and U20988 (N_20988,N_18126,N_16058);
and U20989 (N_20989,N_18094,N_16576);
nor U20990 (N_20990,N_18213,N_18453);
nand U20991 (N_20991,N_19291,N_16509);
xnor U20992 (N_20992,N_19610,N_19651);
nand U20993 (N_20993,N_17334,N_15600);
and U20994 (N_20994,N_19961,N_17078);
nor U20995 (N_20995,N_18407,N_15208);
nand U20996 (N_20996,N_17299,N_16409);
xnor U20997 (N_20997,N_15282,N_18640);
or U20998 (N_20998,N_16110,N_17788);
and U20999 (N_20999,N_18657,N_17275);
or U21000 (N_21000,N_17777,N_16908);
xor U21001 (N_21001,N_17236,N_18134);
nor U21002 (N_21002,N_18477,N_19197);
xnor U21003 (N_21003,N_16452,N_16914);
nor U21004 (N_21004,N_18436,N_19851);
nor U21005 (N_21005,N_16012,N_16823);
nand U21006 (N_21006,N_15434,N_17584);
nor U21007 (N_21007,N_15922,N_18284);
or U21008 (N_21008,N_19734,N_16404);
nand U21009 (N_21009,N_17337,N_18496);
xor U21010 (N_21010,N_18360,N_19396);
nor U21011 (N_21011,N_15404,N_18676);
xnor U21012 (N_21012,N_15847,N_18686);
and U21013 (N_21013,N_16893,N_17376);
nand U21014 (N_21014,N_19157,N_19509);
nand U21015 (N_21015,N_15242,N_19458);
nand U21016 (N_21016,N_18677,N_17128);
nor U21017 (N_21017,N_19286,N_15683);
nor U21018 (N_21018,N_18909,N_15220);
nand U21019 (N_21019,N_16382,N_19457);
nor U21020 (N_21020,N_17124,N_18351);
or U21021 (N_21021,N_18891,N_17554);
xor U21022 (N_21022,N_16498,N_19028);
or U21023 (N_21023,N_18649,N_18197);
or U21024 (N_21024,N_19912,N_18752);
or U21025 (N_21025,N_18065,N_18375);
xor U21026 (N_21026,N_19830,N_19221);
or U21027 (N_21027,N_19417,N_18412);
or U21028 (N_21028,N_17016,N_16634);
nand U21029 (N_21029,N_18691,N_15627);
xor U21030 (N_21030,N_15980,N_15810);
nand U21031 (N_21031,N_15031,N_19823);
and U21032 (N_21032,N_16159,N_16960);
nand U21033 (N_21033,N_15127,N_18152);
nand U21034 (N_21034,N_15004,N_18631);
or U21035 (N_21035,N_17776,N_18558);
nor U21036 (N_21036,N_18313,N_19438);
nand U21037 (N_21037,N_19301,N_17364);
nand U21038 (N_21038,N_16702,N_18300);
nor U21039 (N_21039,N_19510,N_19748);
nand U21040 (N_21040,N_15027,N_15882);
and U21041 (N_21041,N_18168,N_18198);
and U21042 (N_21042,N_16189,N_18007);
and U21043 (N_21043,N_15488,N_18562);
and U21044 (N_21044,N_19209,N_19905);
and U21045 (N_21045,N_17223,N_17031);
nand U21046 (N_21046,N_17265,N_19964);
or U21047 (N_21047,N_15409,N_18470);
nor U21048 (N_21048,N_19460,N_16628);
or U21049 (N_21049,N_15811,N_17980);
nand U21050 (N_21050,N_16147,N_16826);
and U21051 (N_21051,N_18869,N_17652);
nand U21052 (N_21052,N_19138,N_17389);
nor U21053 (N_21053,N_16894,N_19828);
xor U21054 (N_21054,N_18794,N_16079);
nor U21055 (N_21055,N_19401,N_19575);
nand U21056 (N_21056,N_16915,N_18675);
and U21057 (N_21057,N_18941,N_15265);
nand U21058 (N_21058,N_16359,N_16556);
or U21059 (N_21059,N_17577,N_15311);
nand U21060 (N_21060,N_16757,N_17587);
and U21061 (N_21061,N_17262,N_18982);
nor U21062 (N_21062,N_17221,N_19524);
nor U21063 (N_21063,N_19920,N_19664);
nor U21064 (N_21064,N_15729,N_18325);
nor U21065 (N_21065,N_16721,N_16160);
xnor U21066 (N_21066,N_17365,N_18828);
nor U21067 (N_21067,N_19013,N_18081);
nand U21068 (N_21068,N_15492,N_19957);
and U21069 (N_21069,N_18555,N_18702);
or U21070 (N_21070,N_17936,N_15772);
and U21071 (N_21071,N_15979,N_15625);
or U21072 (N_21072,N_19771,N_17990);
nor U21073 (N_21073,N_16531,N_15118);
xor U21074 (N_21074,N_17593,N_17249);
or U21075 (N_21075,N_16817,N_15721);
nor U21076 (N_21076,N_16575,N_17759);
and U21077 (N_21077,N_16696,N_15826);
nand U21078 (N_21078,N_15038,N_16653);
nor U21079 (N_21079,N_19363,N_16259);
and U21080 (N_21080,N_16157,N_19732);
and U21081 (N_21081,N_15629,N_18286);
nor U21082 (N_21082,N_17549,N_17171);
and U21083 (N_21083,N_15029,N_17651);
and U21084 (N_21084,N_17870,N_16068);
or U21085 (N_21085,N_15206,N_18797);
nand U21086 (N_21086,N_19776,N_18781);
xnor U21087 (N_21087,N_19878,N_18593);
xor U21088 (N_21088,N_19620,N_18858);
and U21089 (N_21089,N_17268,N_16761);
or U21090 (N_21090,N_17515,N_15855);
xor U21091 (N_21091,N_15908,N_16003);
xor U21092 (N_21092,N_19184,N_19440);
or U21093 (N_21093,N_17740,N_17795);
and U21094 (N_21094,N_19160,N_19134);
nor U21095 (N_21095,N_16001,N_15115);
and U21096 (N_21096,N_18812,N_18886);
xor U21097 (N_21097,N_15377,N_16406);
or U21098 (N_21098,N_19751,N_17375);
nand U21099 (N_21099,N_17766,N_18503);
nand U21100 (N_21100,N_15102,N_17514);
xor U21101 (N_21101,N_15134,N_15761);
xor U21102 (N_21102,N_19849,N_15005);
nor U21103 (N_21103,N_15077,N_17930);
nor U21104 (N_21104,N_17001,N_19012);
and U21105 (N_21105,N_17840,N_16999);
nor U21106 (N_21106,N_15630,N_18598);
nor U21107 (N_21107,N_16323,N_19332);
or U21108 (N_21108,N_16173,N_15312);
and U21109 (N_21109,N_17127,N_15968);
and U21110 (N_21110,N_18334,N_19069);
nand U21111 (N_21111,N_19009,N_16142);
nor U21112 (N_21112,N_17887,N_16511);
and U21113 (N_21113,N_15926,N_19954);
or U21114 (N_21114,N_16844,N_15385);
or U21115 (N_21115,N_18800,N_16241);
nand U21116 (N_21116,N_17000,N_15343);
nand U21117 (N_21117,N_17745,N_18103);
and U21118 (N_21118,N_15708,N_19093);
nor U21119 (N_21119,N_19682,N_15544);
and U21120 (N_21120,N_19352,N_16491);
nor U21121 (N_21121,N_18761,N_17273);
nor U21122 (N_21122,N_15151,N_16878);
or U21123 (N_21123,N_17730,N_18077);
nor U21124 (N_21124,N_17746,N_18058);
nand U21125 (N_21125,N_15955,N_18108);
or U21126 (N_21126,N_15315,N_18543);
nand U21127 (N_21127,N_16055,N_18586);
and U21128 (N_21128,N_16137,N_18986);
and U21129 (N_21129,N_18730,N_19946);
and U21130 (N_21130,N_17206,N_15641);
nor U21131 (N_21131,N_17022,N_15182);
or U21132 (N_21132,N_17465,N_17058);
nand U21133 (N_21133,N_15809,N_16783);
nor U21134 (N_21134,N_16872,N_18329);
or U21135 (N_21135,N_18428,N_19848);
nand U21136 (N_21136,N_17032,N_18318);
nor U21137 (N_21137,N_17775,N_18302);
nand U21138 (N_21138,N_17270,N_16772);
nor U21139 (N_21139,N_18945,N_16566);
xor U21140 (N_21140,N_16825,N_19939);
nor U21141 (N_21141,N_19190,N_19346);
nand U21142 (N_21142,N_19959,N_15140);
or U21143 (N_21143,N_18707,N_19367);
or U21144 (N_21144,N_15521,N_17985);
nor U21145 (N_21145,N_15199,N_18972);
nor U21146 (N_21146,N_18577,N_15817);
nand U21147 (N_21147,N_17348,N_18435);
nor U21148 (N_21148,N_16375,N_16158);
and U21149 (N_21149,N_15781,N_17184);
nor U21150 (N_21150,N_18452,N_16471);
or U21151 (N_21151,N_18117,N_15239);
and U21152 (N_21152,N_19452,N_18226);
nand U21153 (N_21153,N_19854,N_19447);
xnor U21154 (N_21154,N_17360,N_15339);
and U21155 (N_21155,N_18245,N_19746);
and U21156 (N_21156,N_16345,N_19724);
and U21157 (N_21157,N_16537,N_17285);
or U21158 (N_21158,N_17467,N_15017);
and U21159 (N_21159,N_16420,N_17893);
and U21160 (N_21160,N_18290,N_15660);
or U21161 (N_21161,N_15852,N_15706);
nor U21162 (N_21162,N_19364,N_15228);
nor U21163 (N_21163,N_16689,N_15192);
nor U21164 (N_21164,N_17099,N_18960);
and U21165 (N_21165,N_15839,N_16625);
nand U21166 (N_21166,N_15290,N_17004);
nor U21167 (N_21167,N_17027,N_17881);
xnor U21168 (N_21168,N_18952,N_18889);
nand U21169 (N_21169,N_19608,N_15657);
and U21170 (N_21170,N_17605,N_19948);
nor U21171 (N_21171,N_17760,N_19425);
nor U21172 (N_21172,N_15503,N_17065);
xor U21173 (N_21173,N_17829,N_18692);
nor U21174 (N_21174,N_17328,N_17786);
nand U21175 (N_21175,N_15502,N_19159);
xnor U21176 (N_21176,N_19017,N_17614);
or U21177 (N_21177,N_15076,N_17253);
and U21178 (N_21178,N_17932,N_19896);
nand U21179 (N_21179,N_15635,N_15690);
nor U21180 (N_21180,N_18896,N_16650);
nand U21181 (N_21181,N_18016,N_19351);
nor U21182 (N_21182,N_19568,N_15750);
nor U21183 (N_21183,N_15514,N_15438);
xor U21184 (N_21184,N_16604,N_16238);
or U21185 (N_21185,N_15423,N_17220);
nand U21186 (N_21186,N_15797,N_19117);
or U21187 (N_21187,N_17813,N_15130);
nor U21188 (N_21188,N_15209,N_15295);
xor U21189 (N_21189,N_18242,N_15256);
or U21190 (N_21190,N_19195,N_15025);
nor U21191 (N_21191,N_17054,N_19934);
nor U21192 (N_21192,N_18347,N_17276);
xnor U21193 (N_21193,N_17812,N_18721);
or U21194 (N_21194,N_17921,N_17191);
xnor U21195 (N_21195,N_17531,N_17143);
and U21196 (N_21196,N_17148,N_19983);
nand U21197 (N_21197,N_15666,N_17330);
and U21198 (N_21198,N_19630,N_17320);
or U21199 (N_21199,N_15567,N_19930);
and U21200 (N_21200,N_19850,N_19481);
or U21201 (N_21201,N_15398,N_15878);
xor U21202 (N_21202,N_17940,N_16554);
nor U21203 (N_21203,N_19032,N_19323);
nor U21204 (N_21204,N_19760,N_17891);
nor U21205 (N_21205,N_19884,N_19874);
nor U21206 (N_21206,N_17024,N_15096);
xnor U21207 (N_21207,N_16436,N_15064);
and U21208 (N_21208,N_19941,N_16682);
and U21209 (N_21209,N_15435,N_16082);
or U21210 (N_21210,N_15948,N_18043);
nor U21211 (N_21211,N_19482,N_17122);
nand U21212 (N_21212,N_18092,N_18188);
and U21213 (N_21213,N_15929,N_17051);
nor U21214 (N_21214,N_17948,N_16814);
xnor U21215 (N_21215,N_19144,N_17989);
or U21216 (N_21216,N_15259,N_18579);
or U21217 (N_21217,N_17934,N_19179);
nand U21218 (N_21218,N_16051,N_17197);
nor U21219 (N_21219,N_19294,N_16684);
nor U21220 (N_21220,N_18298,N_16486);
nor U21221 (N_21221,N_15142,N_19094);
nor U21222 (N_21222,N_15364,N_17277);
or U21223 (N_21223,N_15386,N_16397);
and U21224 (N_21224,N_15414,N_19431);
and U21225 (N_21225,N_15296,N_19935);
or U21226 (N_21226,N_18380,N_18835);
nor U21227 (N_21227,N_15214,N_15248);
and U21228 (N_21228,N_17780,N_15692);
and U21229 (N_21229,N_16441,N_16819);
or U21230 (N_21230,N_18750,N_17231);
nor U21231 (N_21231,N_18557,N_16841);
and U21232 (N_21232,N_18112,N_18554);
or U21233 (N_21233,N_17244,N_19989);
and U21234 (N_21234,N_16305,N_18128);
nor U21235 (N_21235,N_16958,N_19418);
and U21236 (N_21236,N_15622,N_18903);
xnor U21237 (N_21237,N_18787,N_17410);
and U21238 (N_21238,N_16181,N_19761);
nand U21239 (N_21239,N_18895,N_18017);
nor U21240 (N_21240,N_17482,N_18254);
or U21241 (N_21241,N_16671,N_16154);
nor U21242 (N_21242,N_19736,N_19334);
and U21243 (N_21243,N_16707,N_16319);
xor U21244 (N_21244,N_16023,N_16403);
or U21245 (N_21245,N_16264,N_19349);
or U21246 (N_21246,N_16080,N_16041);
nor U21247 (N_21247,N_15681,N_17653);
nor U21248 (N_21248,N_16568,N_17696);
xnor U21249 (N_21249,N_19439,N_16668);
nor U21250 (N_21250,N_15128,N_17411);
and U21251 (N_21251,N_18948,N_18628);
and U21252 (N_21252,N_15665,N_18209);
nand U21253 (N_21253,N_18585,N_16709);
nand U21254 (N_21254,N_17061,N_16670);
nor U21255 (N_21255,N_16773,N_18096);
or U21256 (N_21256,N_15307,N_15670);
and U21257 (N_21257,N_16832,N_15421);
or U21258 (N_21258,N_16244,N_15236);
or U21259 (N_21259,N_18892,N_19704);
or U21260 (N_21260,N_16530,N_18420);
and U21261 (N_21261,N_17496,N_19811);
nand U21262 (N_21262,N_19670,N_16674);
xnor U21263 (N_21263,N_19024,N_18183);
or U21264 (N_21264,N_16635,N_18523);
or U21265 (N_21265,N_17251,N_18429);
nand U21266 (N_21266,N_18230,N_17035);
nand U21267 (N_21267,N_16683,N_16299);
nor U21268 (N_21268,N_16047,N_17457);
xor U21269 (N_21269,N_16463,N_17274);
xnor U21270 (N_21270,N_19257,N_18392);
nand U21271 (N_21271,N_15619,N_18872);
and U21272 (N_21272,N_15113,N_17034);
nand U21273 (N_21273,N_19186,N_17068);
xor U21274 (N_21274,N_18208,N_16747);
xor U21275 (N_21275,N_15390,N_18296);
or U21276 (N_21276,N_17176,N_16578);
nand U21277 (N_21277,N_17142,N_15124);
or U21278 (N_21278,N_15126,N_17149);
or U21279 (N_21279,N_15854,N_15835);
and U21280 (N_21280,N_16854,N_15516);
or U21281 (N_21281,N_18243,N_16726);
and U21282 (N_21282,N_19075,N_19099);
nand U21283 (N_21283,N_19831,N_18646);
nor U21284 (N_21284,N_18852,N_17638);
nand U21285 (N_21285,N_15902,N_17947);
or U21286 (N_21286,N_18684,N_18026);
or U21287 (N_21287,N_15428,N_15548);
or U21288 (N_21288,N_19061,N_15485);
nor U21289 (N_21289,N_17601,N_15350);
or U21290 (N_21290,N_18705,N_16178);
and U21291 (N_21291,N_15533,N_18462);
and U21292 (N_21292,N_18947,N_17524);
and U21293 (N_21293,N_18044,N_16645);
or U21294 (N_21294,N_19490,N_19701);
nor U21295 (N_21295,N_19657,N_17864);
nor U21296 (N_21296,N_16163,N_18292);
or U21297 (N_21297,N_15519,N_15606);
nor U21298 (N_21298,N_16859,N_15191);
nand U21299 (N_21299,N_15785,N_17489);
xor U21300 (N_21300,N_17383,N_16337);
nor U21301 (N_21301,N_17386,N_15308);
and U21302 (N_21302,N_15674,N_19098);
nand U21303 (N_21303,N_16994,N_17820);
nand U21304 (N_21304,N_18634,N_17970);
nor U21305 (N_21305,N_16136,N_16367);
and U21306 (N_21306,N_16401,N_15367);
or U21307 (N_21307,N_18373,N_19029);
nor U21308 (N_21308,N_16724,N_19889);
nor U21309 (N_21309,N_17117,N_17708);
or U21310 (N_21310,N_15338,N_16897);
and U21311 (N_21311,N_19137,N_16268);
nor U21312 (N_21312,N_19372,N_18754);
xor U21313 (N_21313,N_16092,N_15407);
and U21314 (N_21314,N_18359,N_19078);
or U21315 (N_21315,N_16025,N_16977);
nand U21316 (N_21316,N_19659,N_16090);
nand U21317 (N_21317,N_17158,N_17686);
or U21318 (N_21318,N_17862,N_18578);
nand U21319 (N_21319,N_16248,N_17160);
and U21320 (N_21320,N_19966,N_18062);
nor U21321 (N_21321,N_17048,N_17784);
or U21322 (N_21322,N_16870,N_18967);
nand U21323 (N_21323,N_18394,N_19675);
nand U21324 (N_21324,N_19605,N_15825);
and U21325 (N_21325,N_15351,N_17345);
or U21326 (N_21326,N_16719,N_16228);
and U21327 (N_21327,N_17763,N_18476);
nand U21328 (N_21328,N_16429,N_16224);
xor U21329 (N_21329,N_15337,N_15586);
nor U21330 (N_21330,N_18615,N_15200);
nor U21331 (N_21331,N_17976,N_17631);
xnor U21332 (N_21332,N_15505,N_16901);
and U21333 (N_21333,N_15967,N_18156);
xnor U21334 (N_21334,N_19141,N_19728);
and U21335 (N_21335,N_17673,N_18576);
nand U21336 (N_21336,N_19503,N_19129);
or U21337 (N_21337,N_19940,N_18421);
nand U21338 (N_21338,N_17738,N_19689);
nand U21339 (N_21339,N_16888,N_17818);
and U21340 (N_21340,N_16974,N_19229);
nand U21341 (N_21341,N_18914,N_16640);
nand U21342 (N_21342,N_19984,N_18299);
and U21343 (N_21343,N_18321,N_18883);
nor U21344 (N_21344,N_19506,N_19722);
and U21345 (N_21345,N_18148,N_18323);
or U21346 (N_21346,N_15883,N_19890);
and U21347 (N_21347,N_17010,N_17327);
or U21348 (N_21348,N_17713,N_16175);
xor U21349 (N_21349,N_17851,N_15782);
and U21350 (N_21350,N_17256,N_18233);
nand U21351 (N_21351,N_16414,N_17395);
or U21352 (N_21352,N_15856,N_16398);
nand U21353 (N_21353,N_18666,N_19467);
or U21354 (N_21354,N_15304,N_18158);
or U21355 (N_21355,N_17667,N_18516);
and U21356 (N_21356,N_16765,N_17837);
and U21357 (N_21357,N_19188,N_16775);
nor U21358 (N_21358,N_19517,N_16328);
nor U21359 (N_21359,N_18368,N_17082);
nor U21360 (N_21360,N_16579,N_18052);
or U21361 (N_21361,N_17394,N_18365);
nand U21362 (N_21362,N_19817,N_15801);
nor U21363 (N_21363,N_16904,N_19395);
nor U21364 (N_21364,N_17714,N_15821);
and U21365 (N_21365,N_15348,N_16470);
nor U21366 (N_21366,N_15198,N_15359);
and U21367 (N_21367,N_16280,N_19640);
xnor U21368 (N_21368,N_16312,N_16475);
nand U21369 (N_21369,N_17037,N_19737);
xnor U21370 (N_21370,N_19585,N_17873);
and U21371 (N_21371,N_15879,N_16646);
and U21372 (N_21372,N_18390,N_16527);
and U21373 (N_21373,N_18269,N_16555);
nand U21374 (N_21374,N_16180,N_19647);
xor U21375 (N_21375,N_15934,N_16522);
nand U21376 (N_21376,N_16214,N_19273);
or U21377 (N_21377,N_15862,N_15636);
and U21378 (N_21378,N_18448,N_15555);
xnor U21379 (N_21379,N_15353,N_16223);
and U21380 (N_21380,N_15316,N_18956);
nand U21381 (N_21381,N_16236,N_15460);
and U21382 (N_21382,N_16297,N_16896);
xnor U21383 (N_21383,N_19492,N_16594);
and U21384 (N_21384,N_16455,N_18746);
or U21385 (N_21385,N_19232,N_18808);
nor U21386 (N_21386,N_18743,N_19700);
nor U21387 (N_21387,N_17095,N_17969);
and U21388 (N_21388,N_15454,N_16986);
or U21389 (N_21389,N_19825,N_18028);
and U21390 (N_21390,N_16203,N_18352);
nor U21391 (N_21391,N_17292,N_18779);
nor U21392 (N_21392,N_17480,N_15093);
nand U21393 (N_21393,N_16402,N_19215);
xnor U21394 (N_21394,N_17657,N_17814);
and U21395 (N_21395,N_18825,N_19128);
or U21396 (N_21396,N_19628,N_16286);
and U21397 (N_21397,N_15532,N_19718);
nand U21398 (N_21398,N_15966,N_17469);
nand U21399 (N_21399,N_18285,N_16529);
or U21400 (N_21400,N_17084,N_18185);
or U21401 (N_21401,N_15546,N_19493);
or U21402 (N_21402,N_18446,N_15274);
nor U21403 (N_21403,N_19895,N_15044);
nor U21404 (N_21404,N_15150,N_15108);
or U21405 (N_21405,N_18923,N_18768);
nand U21406 (N_21406,N_17595,N_16391);
nand U21407 (N_21407,N_17628,N_19804);
and U21408 (N_21408,N_16862,N_17237);
or U21409 (N_21409,N_16400,N_18951);
and U21410 (N_21410,N_18763,N_16465);
nand U21411 (N_21411,N_19968,N_17075);
and U21412 (N_21412,N_19053,N_15075);
and U21413 (N_21413,N_18724,N_19660);
nor U21414 (N_21414,N_19338,N_17992);
or U21415 (N_21415,N_15927,N_15479);
and U21416 (N_21416,N_17557,N_15637);
nor U21417 (N_21417,N_15309,N_19149);
and U21418 (N_21418,N_17453,N_15303);
nor U21419 (N_21419,N_15234,N_15579);
nand U21420 (N_21420,N_18073,N_19019);
or U21421 (N_21421,N_19370,N_18151);
nor U21422 (N_21422,N_19003,N_18912);
nor U21423 (N_21423,N_15775,N_15792);
nor U21424 (N_21424,N_15828,N_19663);
and U21425 (N_21425,N_18206,N_16156);
and U21426 (N_21426,N_15347,N_19777);
nand U21427 (N_21427,N_15480,N_18672);
nand U21428 (N_21428,N_17559,N_16466);
nor U21429 (N_21429,N_19626,N_19497);
or U21430 (N_21430,N_17100,N_16067);
xnor U21431 (N_21431,N_18425,N_19044);
xnor U21432 (N_21432,N_18771,N_19767);
or U21433 (N_21433,N_16481,N_19665);
and U21434 (N_21434,N_17323,N_19241);
or U21435 (N_21435,N_18063,N_18772);
and U21436 (N_21436,N_17591,N_16887);
xor U21437 (N_21437,N_15667,N_19176);
nor U21438 (N_21438,N_17349,N_18690);
and U21439 (N_21439,N_18461,N_18306);
nand U21440 (N_21440,N_16528,N_17070);
and U21441 (N_21441,N_19276,N_18291);
and U21442 (N_21442,N_16494,N_15050);
nor U21443 (N_21443,N_16945,N_16094);
or U21444 (N_21444,N_17975,N_15699);
or U21445 (N_21445,N_18260,N_15540);
or U21446 (N_21446,N_18256,N_19011);
and U21447 (N_21447,N_18180,N_16287);
xor U21448 (N_21448,N_18317,N_17909);
xnor U21449 (N_21449,N_16169,N_19573);
or U21450 (N_21450,N_18890,N_18874);
or U21451 (N_21451,N_15302,N_15550);
and U21452 (N_21452,N_15539,N_16353);
xor U21453 (N_21453,N_16885,N_15107);
and U21454 (N_21454,N_16890,N_16686);
and U21455 (N_21455,N_19161,N_18460);
and U21456 (N_21456,N_19316,N_18749);
nand U21457 (N_21457,N_15291,N_15618);
nor U21458 (N_21458,N_17178,N_16768);
nand U21459 (N_21459,N_18328,N_17425);
nor U21460 (N_21460,N_16219,N_19107);
and U21461 (N_21461,N_17169,N_15734);
or U21462 (N_21462,N_16313,N_18074);
or U21463 (N_21463,N_18682,N_16346);
and U21464 (N_21464,N_17413,N_16622);
and U21465 (N_21465,N_15158,N_16615);
and U21466 (N_21466,N_18293,N_19712);
or U21467 (N_21467,N_15437,N_17718);
or U21468 (N_21468,N_16642,N_18996);
nor U21469 (N_21469,N_18853,N_17451);
nand U21470 (N_21470,N_16138,N_19272);
nor U21471 (N_21471,N_16437,N_15845);
or U21472 (N_21472,N_17029,N_16601);
or U21473 (N_21473,N_18656,N_18139);
nor U21474 (N_21474,N_16487,N_15677);
nand U21475 (N_21475,N_18822,N_16097);
and U21476 (N_21476,N_15286,N_15554);
xnor U21477 (N_21477,N_17362,N_19488);
nor U21478 (N_21478,N_16508,N_18731);
and U21479 (N_21479,N_16678,N_19268);
nor U21480 (N_21480,N_16485,N_16119);
nor U21481 (N_21481,N_19167,N_17286);
nor U21482 (N_21482,N_15644,N_18515);
or U21483 (N_21483,N_16413,N_16714);
nand U21484 (N_21484,N_17896,N_16549);
nor U21485 (N_21485,N_16919,N_17741);
or U21486 (N_21486,N_19392,N_19886);
or U21487 (N_21487,N_15416,N_15857);
and U21488 (N_21488,N_15410,N_18395);
or U21489 (N_21489,N_16326,N_15202);
nor U21490 (N_21490,N_18977,N_17112);
and U21491 (N_21491,N_18738,N_17200);
and U21492 (N_21492,N_18339,N_19264);
nor U21493 (N_21493,N_18342,N_18525);
or U21494 (N_21494,N_16750,N_16171);
nand U21495 (N_21495,N_17937,N_18481);
and U21496 (N_21496,N_19547,N_18207);
or U21497 (N_21497,N_18809,N_16348);
or U21498 (N_21498,N_16846,N_19586);
xor U21499 (N_21499,N_17269,N_17471);
nand U21500 (N_21500,N_18472,N_19000);
nand U21501 (N_21501,N_18770,N_16966);
xnor U21502 (N_21502,N_19908,N_19990);
xor U21503 (N_21503,N_15898,N_16803);
nand U21504 (N_21504,N_17695,N_17865);
nor U21505 (N_21505,N_17479,N_17901);
xor U21506 (N_21506,N_19199,N_15512);
nand U21507 (N_21507,N_18174,N_15765);
and U21508 (N_21508,N_18093,N_18121);
nor U21509 (N_21509,N_18200,N_17773);
and U21510 (N_21510,N_15717,N_18031);
nand U21511 (N_21511,N_16089,N_17588);
and U21512 (N_21512,N_17013,N_19606);
nand U21513 (N_21513,N_18146,N_16335);
nor U21514 (N_21514,N_16457,N_18790);
nand U21515 (N_21515,N_15662,N_19539);
and U21516 (N_21516,N_19006,N_18711);
or U21517 (N_21517,N_15373,N_19997);
or U21518 (N_21518,N_19462,N_19499);
xnor U21519 (N_21519,N_17398,N_19725);
nand U21520 (N_21520,N_17131,N_18988);
or U21521 (N_21521,N_18632,N_17966);
or U21522 (N_21522,N_17335,N_19676);
or U21523 (N_21523,N_17824,N_16349);
nor U21524 (N_21524,N_19609,N_19085);
and U21525 (N_21525,N_16202,N_16269);
nor U21526 (N_21526,N_18086,N_17815);
and U21527 (N_21527,N_18196,N_17409);
nand U21528 (N_21528,N_18410,N_17874);
and U21529 (N_21529,N_19840,N_18040);
xnor U21530 (N_21530,N_18980,N_19172);
and U21531 (N_21531,N_19052,N_15088);
or U21532 (N_21532,N_19127,N_15518);
or U21533 (N_21533,N_16274,N_18648);
or U21534 (N_21534,N_18594,N_15022);
nor U21535 (N_21535,N_18154,N_15830);
or U21536 (N_21536,N_15431,N_16996);
or U21537 (N_21537,N_19202,N_16703);
or U21538 (N_21538,N_19550,N_15201);
xor U21539 (N_21539,N_19112,N_16392);
nand U21540 (N_21540,N_15655,N_16923);
nor U21541 (N_21541,N_18295,N_19949);
nor U21542 (N_21542,N_15097,N_19611);
and U21543 (N_21543,N_16532,N_16580);
or U21544 (N_21544,N_15405,N_19133);
nor U21545 (N_21545,N_16755,N_15964);
or U21546 (N_21546,N_18524,N_17861);
and U21547 (N_21547,N_19282,N_17853);
nor U21548 (N_21548,N_15577,N_16469);
or U21549 (N_21549,N_15834,N_19687);
nor U21550 (N_21550,N_18826,N_17284);
nor U21551 (N_21551,N_16796,N_16207);
and U21552 (N_21552,N_15468,N_19769);
xnor U21553 (N_21553,N_15928,N_19089);
or U21554 (N_21554,N_15931,N_19326);
and U21555 (N_21555,N_16011,N_19242);
nor U21556 (N_21556,N_15776,N_16971);
and U21557 (N_21557,N_15278,N_16013);
nor U21558 (N_21558,N_16237,N_19200);
nor U21559 (N_21559,N_19720,N_16882);
nand U21560 (N_21560,N_17050,N_15153);
nor U21561 (N_21561,N_16069,N_19537);
nand U21562 (N_21562,N_16188,N_16956);
and U21563 (N_21563,N_19288,N_19967);
and U21564 (N_21564,N_15079,N_16656);
and U21565 (N_21565,N_19254,N_17215);
or U21566 (N_21566,N_19446,N_15141);
nor U21567 (N_21567,N_19480,N_18010);
xor U21568 (N_21568,N_15588,N_17987);
and U21569 (N_21569,N_17172,N_17617);
or U21570 (N_21570,N_18150,N_17166);
nor U21571 (N_21571,N_17808,N_18803);
nand U21572 (N_21572,N_17146,N_17226);
and U21573 (N_21573,N_16770,N_15173);
and U21574 (N_21574,N_15596,N_17833);
or U21575 (N_21575,N_17346,N_16997);
or U21576 (N_21576,N_16233,N_15010);
and U21577 (N_21577,N_19068,N_18430);
and U21578 (N_21578,N_17417,N_17632);
nor U21579 (N_21579,N_15917,N_16186);
and U21580 (N_21580,N_19123,N_15482);
nor U21581 (N_21581,N_16474,N_19410);
or U21582 (N_21582,N_18919,N_17999);
and U21583 (N_21583,N_15447,N_18215);
nor U21584 (N_21584,N_15689,N_19152);
xor U21585 (N_21585,N_16664,N_15658);
nor U21586 (N_21586,N_18987,N_17816);
or U21587 (N_21587,N_15326,N_15442);
xnor U21588 (N_21588,N_19565,N_17342);
nand U21589 (N_21589,N_17260,N_16385);
nor U21590 (N_21590,N_17460,N_18699);
and U21591 (N_21591,N_16198,N_17894);
xor U21592 (N_21592,N_15786,N_19070);
or U21593 (N_21593,N_19987,N_16657);
xor U21594 (N_21594,N_15015,N_18851);
nor U21595 (N_21595,N_19903,N_17252);
and U21596 (N_21596,N_15449,N_17396);
nand U21597 (N_21597,N_17069,N_16736);
nor U21598 (N_21598,N_17765,N_19466);
nand U21599 (N_21599,N_19943,N_15624);
nor U21600 (N_21600,N_16526,N_17493);
nor U21601 (N_21601,N_19454,N_16864);
nand U21602 (N_21602,N_19717,N_15402);
nor U21603 (N_21603,N_19255,N_19317);
nor U21604 (N_21604,N_17564,N_15161);
and U21605 (N_21605,N_16289,N_17125);
or U21606 (N_21606,N_16111,N_19230);
and U21607 (N_21607,N_17431,N_16543);
or U21608 (N_21608,N_16911,N_16694);
nand U21609 (N_21609,N_17949,N_16036);
or U21610 (N_21610,N_17116,N_19416);
nand U21611 (N_21611,N_16492,N_17361);
or U21612 (N_21612,N_19999,N_17938);
nand U21613 (N_21613,N_18567,N_15458);
xor U21614 (N_21614,N_18386,N_19612);
xnor U21615 (N_21615,N_17072,N_16344);
nand U21616 (N_21616,N_17674,N_18045);
and U21617 (N_21617,N_15651,N_16279);
and U21618 (N_21618,N_15137,N_16616);
nand U21619 (N_21619,N_18924,N_18848);
or U21620 (N_21620,N_19259,N_16343);
nor U21621 (N_21621,N_17021,N_16781);
or U21622 (N_21622,N_16708,N_17202);
xnor U21623 (N_21623,N_15233,N_18376);
and U21624 (N_21624,N_18247,N_15033);
nor U21625 (N_21625,N_18806,N_18075);
and U21626 (N_21626,N_16015,N_16679);
xnor U21627 (N_21627,N_19856,N_18601);
or U21628 (N_21628,N_18937,N_19648);
or U21629 (N_21629,N_16609,N_17508);
nor U21630 (N_21630,N_18744,N_15880);
nand U21631 (N_21631,N_18027,N_16598);
nand U21632 (N_21632,N_19081,N_16270);
and U21633 (N_21633,N_16423,N_18526);
and U21634 (N_21634,N_16044,N_18345);
or U21635 (N_21635,N_15180,N_17296);
and U21636 (N_21636,N_18442,N_15695);
or U21637 (N_21637,N_18540,N_19541);
nand U21638 (N_21638,N_15875,N_15937);
nor U21639 (N_21639,N_15327,N_16795);
nor U21640 (N_21640,N_16071,N_19595);
or U21641 (N_21641,N_15176,N_19348);
nor U21642 (N_21642,N_19347,N_16477);
nand U21643 (N_21643,N_16961,N_17401);
and U21644 (N_21644,N_17875,N_18957);
nor U21645 (N_21645,N_16276,N_15263);
nand U21646 (N_21646,N_18340,N_19110);
nor U21647 (N_21647,N_17906,N_18974);
and U21648 (N_21648,N_17023,N_19872);
xnor U21649 (N_21649,N_16210,N_16871);
or U21650 (N_21650,N_17767,N_16194);
and U21651 (N_21651,N_16785,N_16753);
nand U21652 (N_21652,N_16253,N_19745);
xnor U21653 (N_21653,N_16021,N_17014);
nand U21654 (N_21654,N_15006,N_19730);
and U21655 (N_21655,N_16192,N_19136);
xor U21656 (N_21656,N_16614,N_17145);
nor U21657 (N_21657,N_15687,N_17291);
nor U21658 (N_21658,N_19315,N_15557);
nand U21659 (N_21659,N_15346,N_16088);
nor U21660 (N_21660,N_15601,N_19477);
or U21661 (N_21661,N_19381,N_19692);
or U21662 (N_21662,N_15203,N_16245);
and U21663 (N_21663,N_18316,N_17886);
and U21664 (N_21664,N_18458,N_17589);
or U21665 (N_21665,N_18929,N_18060);
or U21666 (N_21666,N_15085,N_17288);
or U21667 (N_21667,N_16857,N_15643);
nand U21668 (N_21668,N_16412,N_17663);
xnor U21669 (N_21669,N_17475,N_16200);
or U21670 (N_21670,N_17604,N_17723);
nor U21671 (N_21671,N_19713,N_18485);
and U21672 (N_21672,N_16149,N_16101);
nor U21673 (N_21673,N_17369,N_18278);
nand U21674 (N_21674,N_15167,N_15008);
xor U21675 (N_21675,N_15081,N_18239);
or U21676 (N_21676,N_17452,N_15281);
or U21677 (N_21677,N_18018,N_15943);
nand U21678 (N_21678,N_16368,N_17681);
nand U21679 (N_21679,N_18406,N_17419);
nand U21680 (N_21680,N_15836,N_15439);
nor U21681 (N_21681,N_16164,N_17052);
and U21682 (N_21682,N_17462,N_16091);
nor U21683 (N_21683,N_17556,N_18792);
xnor U21684 (N_21684,N_19016,N_19868);
and U21685 (N_21685,N_16330,N_15799);
nor U21686 (N_21686,N_18789,N_18263);
xnor U21687 (N_21687,N_15174,N_19792);
nor U21688 (N_21688,N_16605,N_18819);
and U21689 (N_21689,N_17877,N_17778);
nand U21690 (N_21690,N_19690,N_17281);
nor U21691 (N_21691,N_19071,N_19847);
and U21692 (N_21692,N_17769,N_17074);
or U21693 (N_21693,N_19627,N_18361);
or U21694 (N_21694,N_18596,N_15063);
nor U21695 (N_21695,N_19805,N_16443);
nor U21696 (N_21696,N_15135,N_19569);
nor U21697 (N_21697,N_15275,N_18498);
and U21698 (N_21698,N_19164,N_15261);
xnor U21699 (N_21699,N_19169,N_17516);
and U21700 (N_21700,N_19171,N_16540);
xnor U21701 (N_21701,N_16926,N_16415);
xnor U21702 (N_21702,N_15216,N_16563);
or U21703 (N_21703,N_17911,N_16377);
or U21704 (N_21704,N_15563,N_15066);
or U21705 (N_21705,N_15007,N_17378);
xnor U21706 (N_21706,N_15046,N_17834);
nor U21707 (N_21707,N_17664,N_19073);
nand U21708 (N_21708,N_15257,N_15903);
and U21709 (N_21709,N_16087,N_15204);
nor U21710 (N_21710,N_16190,N_17736);
nand U21711 (N_21711,N_18466,N_18597);
nand U21712 (N_21712,N_15493,N_18704);
and U21713 (N_21713,N_15272,N_19784);
or U21714 (N_21714,N_18860,N_19267);
and U21715 (N_21715,N_17090,N_16007);
xor U21716 (N_21716,N_17402,N_19519);
xor U21717 (N_21717,N_17151,N_16973);
nand U21718 (N_21718,N_19680,N_15815);
nor U21719 (N_21719,N_17643,N_19415);
and U21720 (N_21720,N_17712,N_18336);
nand U21721 (N_21721,N_17897,N_18445);
and U21722 (N_21722,N_18865,N_15723);
and U21723 (N_21723,N_19120,N_16979);
or U21724 (N_21724,N_18653,N_19845);
nand U21725 (N_21725,N_15149,N_15271);
or U21726 (N_21726,N_15754,N_18993);
nand U21727 (N_21727,N_18629,N_17671);
nand U21728 (N_21728,N_15486,N_16942);
and U21729 (N_21729,N_18199,N_16199);
xnor U21730 (N_21730,N_19556,N_15498);
xnor U21731 (N_21731,N_19800,N_17157);
or U21732 (N_21732,N_16837,N_15260);
nand U21733 (N_21733,N_17703,N_19010);
nand U21734 (N_21734,N_15043,N_16024);
and U21735 (N_21735,N_17570,N_17621);
or U21736 (N_21736,N_16053,N_17351);
nor U21737 (N_21737,N_19778,N_17944);
or U21738 (N_21738,N_19956,N_17794);
nor U21739 (N_21739,N_16743,N_17279);
or U21740 (N_21740,N_18818,N_16118);
or U21741 (N_21741,N_18942,N_15842);
nor U21742 (N_21742,N_16255,N_19917);
nand U21743 (N_21743,N_17560,N_15072);
nand U21744 (N_21744,N_15456,N_18807);
or U21745 (N_21745,N_15186,N_15536);
nand U21746 (N_21746,N_16179,N_18118);
nand U21747 (N_21747,N_17567,N_19829);
nor U21748 (N_21748,N_18661,N_19578);
or U21749 (N_21749,N_18354,N_16866);
nand U21750 (N_21750,N_19786,N_17189);
or U21751 (N_21751,N_16300,N_17303);
and U21752 (N_21752,N_15171,N_18310);
or U21753 (N_21753,N_19932,N_18332);
nor U21754 (N_21754,N_18534,N_16063);
nor U21755 (N_21755,N_15083,N_19034);
or U21756 (N_21756,N_16043,N_19822);
and U21757 (N_21757,N_16153,N_18055);
and U21758 (N_21758,N_16778,N_15850);
and U21759 (N_21759,N_19998,N_18953);
nor U21760 (N_21760,N_16086,N_15693);
nor U21761 (N_21761,N_16677,N_17929);
or U21762 (N_21762,N_18305,N_19424);
and U21763 (N_21763,N_17138,N_18171);
nor U21764 (N_21764,N_19816,N_17757);
nor U21765 (N_21765,N_16215,N_17331);
nand U21766 (N_21766,N_19163,N_15036);
and U21767 (N_21767,N_15092,N_18382);
and U21768 (N_21768,N_17576,N_16798);
and U21769 (N_21769,N_19982,N_16124);
and U21770 (N_21770,N_19058,N_16957);
nor U21771 (N_21771,N_18267,N_18471);
xnor U21772 (N_21772,N_17743,N_15154);
nand U21773 (N_21773,N_19808,N_18863);
and U21774 (N_21774,N_18635,N_17297);
xnor U21775 (N_21775,N_16209,N_17406);
nand U21776 (N_21776,N_16476,N_16425);
nand U21777 (N_21777,N_18383,N_16545);
nor U21778 (N_21778,N_18687,N_16548);
and U21779 (N_21779,N_19359,N_19269);
nor U21780 (N_21780,N_15397,N_19862);
or U21781 (N_21781,N_17506,N_15831);
nand U21782 (N_21782,N_15678,N_16172);
nor U21783 (N_21783,N_19755,N_17005);
or U21784 (N_21784,N_16246,N_18258);
nand U21785 (N_21785,N_18143,N_19866);
or U21786 (N_21786,N_16767,N_15181);
and U21787 (N_21787,N_19287,N_18120);
and U21788 (N_21788,N_16608,N_16249);
and U21789 (N_21789,N_17846,N_17859);
nand U21790 (N_21790,N_17437,N_19749);
xnor U21791 (N_21791,N_16032,N_19589);
and U21792 (N_21792,N_19036,N_18899);
nor U21793 (N_21793,N_18037,N_17998);
and U21794 (N_21794,N_15333,N_15382);
nor U21795 (N_21795,N_19570,N_15647);
nand U21796 (N_21796,N_17384,N_15921);
and U21797 (N_21797,N_17878,N_15623);
and U21798 (N_21798,N_16195,N_16672);
nor U21799 (N_21799,N_19380,N_19911);
nor U21800 (N_21800,N_18991,N_15318);
nor U21801 (N_21801,N_19060,N_18995);
and U21802 (N_21802,N_15759,N_16478);
and U21803 (N_21803,N_15920,N_17121);
or U21804 (N_21804,N_15564,N_15768);
nor U21805 (N_21805,N_16281,N_16728);
nor U21806 (N_21806,N_19118,N_17040);
xor U21807 (N_21807,N_17581,N_16220);
nand U21808 (N_21808,N_15491,N_19919);
or U21809 (N_21809,N_18966,N_19419);
and U21810 (N_21810,N_18211,N_17665);
or U21811 (N_21811,N_19476,N_17057);
nor U21812 (N_21812,N_19587,N_17521);
nand U21813 (N_21813,N_16627,N_19705);
and U21814 (N_21814,N_18343,N_19087);
nor U21815 (N_21815,N_19217,N_19178);
and U21816 (N_21816,N_15249,N_15396);
xor U21817 (N_21817,N_19621,N_15451);
or U21818 (N_21818,N_15935,N_18720);
nor U21819 (N_21819,N_16317,N_17473);
nor U21820 (N_21820,N_15164,N_16905);
nand U21821 (N_21821,N_16581,N_18064);
nor U21822 (N_21822,N_18887,N_16129);
nor U21823 (N_21823,N_18795,N_19985);
xnor U21824 (N_21824,N_15594,N_15391);
and U21825 (N_21825,N_18572,N_19754);
nand U21826 (N_21826,N_16583,N_16165);
and U21827 (N_21827,N_17903,N_15306);
and U21828 (N_21828,N_16225,N_17304);
and U21829 (N_21829,N_15807,N_17915);
nor U21830 (N_21830,N_17585,N_18219);
nand U21831 (N_21831,N_19305,N_18161);
nand U21832 (N_21832,N_17925,N_18493);
nand U21833 (N_21833,N_18734,N_15732);
or U21834 (N_21834,N_15520,N_18617);
xnor U21835 (N_21835,N_16205,N_15243);
nand U21836 (N_21836,N_18726,N_16738);
nand U21837 (N_21837,N_16360,N_15938);
and U21838 (N_21838,N_17957,N_19600);
or U21839 (N_21839,N_18944,N_17211);
nand U21840 (N_21840,N_18954,N_19045);
and U21841 (N_21841,N_17278,N_15227);
xnor U21842 (N_21842,N_19307,N_18920);
nand U21843 (N_21843,N_15595,N_17087);
and U21844 (N_21844,N_15899,N_18414);
nor U21845 (N_21845,N_15056,N_17982);
or U21846 (N_21846,N_15609,N_19697);
xnor U21847 (N_21847,N_16442,N_17019);
and U21848 (N_21848,N_19153,N_19448);
nand U21849 (N_21849,N_19775,N_17805);
nor U21850 (N_21850,N_16701,N_19944);
or U21851 (N_21851,N_16174,N_17094);
nand U21852 (N_21852,N_17606,N_17458);
or U21853 (N_21853,N_15511,N_19237);
nand U21854 (N_21854,N_15476,N_17168);
nand U21855 (N_21855,N_19534,N_17512);
or U21856 (N_21856,N_17481,N_15912);
or U21857 (N_21857,N_18066,N_18970);
nand U21858 (N_21858,N_16049,N_17892);
nor U21859 (N_21859,N_15997,N_17727);
or U21860 (N_21860,N_16751,N_15445);
nor U21861 (N_21861,N_17313,N_19479);
and U21862 (N_21862,N_18548,N_18760);
or U21863 (N_21863,N_17927,N_19598);
or U21864 (N_21864,N_19358,N_19899);
nand U21865 (N_21865,N_16229,N_18647);
xnor U21866 (N_21866,N_15349,N_18331);
and U21867 (N_21867,N_18403,N_19525);
nand U21868 (N_21868,N_17540,N_16034);
nand U21869 (N_21869,N_18210,N_17039);
and U21870 (N_21870,N_17802,N_17367);
nand U21871 (N_21871,N_17500,N_19631);
nand U21872 (N_21872,N_15467,N_19453);
nor U21873 (N_21873,N_19189,N_16665);
and U21874 (N_21874,N_19487,N_15603);
nor U21875 (N_21875,N_15276,N_16206);
or U21876 (N_21876,N_17687,N_16883);
nor U21877 (N_21877,N_16143,N_18900);
nand U21878 (N_21878,N_16115,N_19043);
xor U21879 (N_21879,N_15148,N_16792);
nor U21880 (N_21880,N_18824,N_15247);
or U21881 (N_21881,N_16560,N_16373);
nor U21882 (N_21882,N_16020,N_19207);
or U21883 (N_21883,N_19625,N_15002);
or U21884 (N_21884,N_16073,N_15042);
and U21885 (N_21885,N_17787,N_15024);
nor U21886 (N_21886,N_19618,N_17047);
and U21887 (N_21887,N_17218,N_15356);
nor U21888 (N_21888,N_17602,N_16296);
and U21889 (N_21889,N_17647,N_19562);
and U21890 (N_21890,N_19256,N_16332);
xor U21891 (N_21891,N_17161,N_15585);
or U21892 (N_21892,N_17225,N_19837);
nor U21893 (N_21893,N_18846,N_17797);
and U21894 (N_21894,N_17527,N_15357);
or U21895 (N_21895,N_19135,N_16456);
nor U21896 (N_21896,N_16285,N_15764);
and U21897 (N_21897,N_17563,N_18894);
nand U21898 (N_21898,N_17619,N_19390);
and U21899 (N_21899,N_16483,N_17770);
and U21900 (N_21900,N_15501,N_17385);
and U21901 (N_21901,N_16523,N_18441);
or U21902 (N_21902,N_15572,N_19526);
nor U21903 (N_21903,N_18934,N_17977);
nand U21904 (N_21904,N_17541,N_18713);
nor U21905 (N_21905,N_15535,N_18350);
nor U21906 (N_21906,N_19311,N_17081);
or U21907 (N_21907,N_16619,N_15530);
xnor U21908 (N_21908,N_15459,N_16907);
and U21909 (N_21909,N_18832,N_18288);
nand U21910 (N_21910,N_17691,N_15738);
and U21911 (N_21911,N_16472,N_18729);
nor U21912 (N_21912,N_16006,N_18255);
xnor U21913 (N_21913,N_15959,N_17255);
or U21914 (N_21914,N_18067,N_15537);
xor U21915 (N_21915,N_18664,N_17551);
and U21916 (N_21916,N_18913,N_18658);
nor U21917 (N_21917,N_15305,N_18850);
nand U21918 (N_21918,N_19677,N_17885);
nor U21919 (N_21919,N_16451,N_19740);
xor U21920 (N_21920,N_16963,N_19196);
nor U21921 (N_21921,N_16208,N_19791);
and U21922 (N_21922,N_15383,N_18486);
nor U21923 (N_21923,N_16027,N_18679);
nand U21924 (N_21924,N_17958,N_19996);
and U21925 (N_21925,N_18160,N_17867);
and U21926 (N_21926,N_16648,N_19877);
and U21927 (N_21927,N_18502,N_19744);
nand U21928 (N_21928,N_19077,N_16008);
or U21929 (N_21929,N_17523,N_17610);
and U21930 (N_21930,N_16040,N_17729);
or U21931 (N_21931,N_15146,N_15650);
xor U21932 (N_21932,N_19379,N_18600);
and U21933 (N_21933,N_18716,N_16567);
or U21934 (N_21934,N_16995,N_15562);
and U21935 (N_21935,N_19900,N_16693);
and U21936 (N_21936,N_17761,N_15741);
and U21937 (N_21937,N_19025,N_15673);
or U21938 (N_21938,N_18042,N_15905);
xor U21939 (N_21939,N_15975,N_18758);
or U21940 (N_21940,N_18638,N_19514);
or U21941 (N_21941,N_15840,N_15487);
or U21942 (N_21942,N_16035,N_16839);
xor U21943 (N_21943,N_16316,N_18652);
nand U21944 (N_21944,N_18608,N_17608);
and U21945 (N_21945,N_18521,N_16512);
nand U21946 (N_21946,N_19450,N_19236);
nand U21947 (N_21947,N_19095,N_15983);
and U21948 (N_21948,N_19464,N_16307);
or U21949 (N_21949,N_16030,N_15058);
nor U21950 (N_21950,N_17207,N_18194);
nor U21951 (N_21951,N_16577,N_17705);
nor U21952 (N_21952,N_15685,N_19485);
xnor U21953 (N_21953,N_17422,N_16706);
nand U21954 (N_21954,N_17067,N_19926);
or U21955 (N_21955,N_19661,N_16538);
or U21956 (N_21956,N_17267,N_15152);
and U21957 (N_21957,N_16662,N_16800);
nand U21958 (N_21958,N_18975,N_19918);
nand U21959 (N_21959,N_18483,N_17424);
xnor U21960 (N_21960,N_19335,N_16243);
xor U21961 (N_21961,N_15195,N_16291);
xnor U21962 (N_21962,N_18005,N_17513);
xor U21963 (N_21963,N_16603,N_15558);
nand U21964 (N_21964,N_18145,N_15189);
or U21965 (N_21965,N_18949,N_18823);
nor U21966 (N_21966,N_15466,N_15432);
xnor U21967 (N_21967,N_16108,N_19040);
or U21968 (N_21968,N_15285,N_16399);
nand U21969 (N_21969,N_18009,N_15495);
and U21970 (N_21970,N_16327,N_19244);
nand U21971 (N_21971,N_16850,N_18595);
or U21972 (N_21972,N_17008,N_15197);
and U21973 (N_21973,N_17945,N_15697);
xor U21974 (N_21974,N_16970,N_16405);
or U21975 (N_21975,N_17447,N_18314);
nor U21976 (N_21976,N_17102,N_18786);
nor U21977 (N_21977,N_19891,N_19140);
nor U21978 (N_21978,N_18936,N_15715);
nor U21979 (N_21979,N_15284,N_16950);
nor U21980 (N_21980,N_17782,N_17302);
nand U21981 (N_21981,N_18667,N_16691);
or U21982 (N_21982,N_19204,N_18484);
nand U21983 (N_21983,N_16666,N_19067);
and U21984 (N_21984,N_16780,N_18765);
nand U21985 (N_21985,N_18527,N_19950);
or U21986 (N_21986,N_19855,N_19430);
or U21987 (N_21987,N_18469,N_18633);
and U21988 (N_21988,N_15238,N_18377);
or U21989 (N_21989,N_19937,N_16687);
or U21990 (N_21990,N_19154,N_15323);
nor U21991 (N_21991,N_17704,N_16076);
nand U21992 (N_21992,N_19101,N_15372);
xor U21993 (N_21993,N_17104,N_15266);
and U21994 (N_21994,N_18371,N_18868);
or U21995 (N_21995,N_17165,N_19353);
nand U21996 (N_21996,N_19710,N_15012);
and U21997 (N_21997,N_16064,N_16096);
nand U21998 (N_21998,N_17792,N_17239);
or U21999 (N_21999,N_19050,N_16791);
and U22000 (N_22000,N_17418,N_19304);
xnor U22001 (N_22001,N_15748,N_18444);
nand U22002 (N_22002,N_19035,N_15254);
nor U22003 (N_22003,N_16544,N_19536);
and U22004 (N_22004,N_15939,N_19564);
nor U22005 (N_22005,N_16808,N_16045);
and U22006 (N_22006,N_19632,N_15827);
and U22007 (N_22007,N_17329,N_19302);
nor U22008 (N_22008,N_16324,N_18659);
xnor U22009 (N_22009,N_16227,N_15230);
or U22010 (N_22010,N_17822,N_15605);
nor U22011 (N_22011,N_15696,N_15793);
nand U22012 (N_22012,N_15193,N_16046);
xor U22013 (N_22013,N_19865,N_19798);
and U22014 (N_22014,N_16777,N_18999);
nand U22015 (N_22015,N_17555,N_16133);
nand U22016 (N_22016,N_19224,N_16185);
and U22017 (N_22017,N_19289,N_19567);
or U22018 (N_22018,N_15613,N_16895);
xnor U22019 (N_22019,N_17159,N_17986);
and U22020 (N_22020,N_15074,N_18946);
or U22021 (N_22021,N_19549,N_16658);
nand U22022 (N_22022,N_19283,N_16959);
nor U22023 (N_22023,N_17943,N_16077);
nand U22024 (N_22024,N_16969,N_19763);
nand U22025 (N_22025,N_15684,N_18289);
and U22026 (N_22026,N_16450,N_15246);
nor U22027 (N_22027,N_18755,N_18095);
xnor U22028 (N_22028,N_18165,N_15602);
nor U22029 (N_22029,N_19361,N_18715);
xor U22030 (N_22030,N_16123,N_18968);
or U22031 (N_22031,N_15500,N_15299);
and U22032 (N_22032,N_18660,N_17880);
nand U22033 (N_22033,N_15560,N_15226);
nor U22034 (N_22034,N_15735,N_18671);
nand U22035 (N_22035,N_16446,N_15461);
or U22036 (N_22036,N_17187,N_18911);
or U22037 (N_22037,N_15744,N_18830);
xor U22038 (N_22038,N_17672,N_18049);
nor U22039 (N_22039,N_19048,N_15849);
or U22040 (N_22040,N_15392,N_15317);
nor U22041 (N_22041,N_15269,N_18591);
nand U22042 (N_22042,N_17951,N_15970);
nor U22043 (N_22043,N_19194,N_17062);
xnor U22044 (N_22044,N_18783,N_15805);
xnor U22045 (N_22045,N_17530,N_17679);
nor U22046 (N_22046,N_19001,N_19097);
nor U22047 (N_22047,N_15870,N_18866);
nand U22048 (N_22048,N_16140,N_15368);
and U22049 (N_22049,N_15798,N_16251);
and U22050 (N_22050,N_18266,N_15288);
or U22051 (N_22051,N_19162,N_17626);
xor U22052 (N_22052,N_15048,N_16016);
nand U22053 (N_22053,N_18725,N_18506);
or U22054 (N_22054,N_17889,N_15190);
and U22055 (N_22055,N_17661,N_17783);
nor U22056 (N_22056,N_15829,N_15593);
nand U22057 (N_22057,N_18722,N_17821);
nor U22058 (N_22058,N_18250,N_19139);
nand U22059 (N_22059,N_18166,N_17111);
nor U22060 (N_22060,N_16748,N_15389);
nand U22061 (N_22061,N_19299,N_19972);
or U22062 (N_22062,N_17546,N_18228);
nand U22063 (N_22063,N_15399,N_16239);
nor U22064 (N_22064,N_19594,N_18688);
nand U22065 (N_22065,N_16048,N_19250);
nand U22066 (N_22066,N_19063,N_16387);
or U22067 (N_22067,N_18624,N_17056);
nand U22068 (N_22068,N_15868,N_17167);
xor U22069 (N_22069,N_18071,N_15755);
and U22070 (N_22070,N_16760,N_18810);
or U22071 (N_22071,N_15121,N_18650);
nor U22072 (N_22072,N_17967,N_19729);
and U22073 (N_22073,N_18774,N_19974);
and U22074 (N_22074,N_17212,N_15731);
xnor U22075 (N_22075,N_19864,N_17503);
nand U22076 (N_22076,N_19155,N_19470);
or U22077 (N_22077,N_18457,N_16733);
xor U22078 (N_22078,N_15653,N_18179);
and U22079 (N_22079,N_19826,N_15675);
nor U22080 (N_22080,N_18511,N_15086);
nor U22081 (N_22081,N_19709,N_19881);
nor U22082 (N_22082,N_15328,N_17079);
nand U22083 (N_22083,N_17968,N_17939);
or U22084 (N_22084,N_19679,N_19398);
and U22085 (N_22085,N_16867,N_16858);
or U22086 (N_22086,N_16600,N_17043);
and U22087 (N_22087,N_16742,N_16984);
nand U22088 (N_22088,N_15874,N_19650);
nand U22089 (N_22089,N_19443,N_16066);
or U22090 (N_22090,N_17997,N_19880);
xnor U22091 (N_22091,N_15472,N_17838);
and U22092 (N_22092,N_16972,N_17642);
and U22093 (N_22093,N_17405,N_19819);
nand U22094 (N_22094,N_15611,N_19814);
nor U22095 (N_22095,N_16277,N_17259);
nor U22096 (N_22096,N_19875,N_19214);
or U22097 (N_22097,N_17044,N_16152);
or U22098 (N_22098,N_17701,N_17580);
nor U22099 (N_22099,N_15000,N_17698);
and U22100 (N_22100,N_18193,N_16218);
nand U22101 (N_22101,N_18509,N_17185);
or U22102 (N_22102,N_18973,N_16759);
and U22103 (N_22103,N_19105,N_15947);
nor U22104 (N_22104,N_16829,N_18969);
and U22105 (N_22105,N_19062,N_15419);
or U22106 (N_22106,N_18532,N_17486);
nor U22107 (N_22107,N_16842,N_15159);
or U22108 (N_22108,N_17301,N_16148);
and U22109 (N_22109,N_17735,N_17456);
and U22110 (N_22110,N_18921,N_15021);
nor U22111 (N_22111,N_16130,N_16440);
xor U22112 (N_22112,N_15933,N_15962);
xor U22113 (N_22113,N_18602,N_19243);
xnor U22114 (N_22114,N_18419,N_16827);
and U22115 (N_22115,N_15682,N_15523);
or U22116 (N_22116,N_19654,N_17582);
nand U22117 (N_22117,N_16395,N_19924);
or U22118 (N_22118,N_16196,N_17955);
xor U22119 (N_22119,N_15440,N_16187);
and U22120 (N_22120,N_15231,N_17238);
nor U22121 (N_22121,N_19371,N_16599);
nand U22122 (N_22122,N_17152,N_16649);
nand U22123 (N_22123,N_17205,N_18129);
nor U22124 (N_22124,N_19591,N_19773);
nor U22125 (N_22125,N_17715,N_15324);
or U22126 (N_22126,N_19703,N_18669);
and U22127 (N_22127,N_19980,N_15587);
nor U22128 (N_22128,N_15401,N_19794);
nor U22129 (N_22129,N_18519,N_17354);
nor U22130 (N_22130,N_19788,N_17341);
xnor U22131 (N_22131,N_16177,N_16261);
or U22132 (N_22132,N_17928,N_19456);
or U22133 (N_22133,N_17603,N_18782);
and U22134 (N_22134,N_15510,N_16822);
nand U22135 (N_22135,N_19806,N_19545);
nor U22136 (N_22136,N_16221,N_19376);
nor U22137 (N_22137,N_19495,N_18564);
and U22138 (N_22138,N_17841,N_18641);
nor U22139 (N_22139,N_19774,N_18654);
and U22140 (N_22140,N_18861,N_18769);
or U22141 (N_22141,N_18297,N_18019);
nor U22142 (N_22142,N_19004,N_16037);
xor U22143 (N_22143,N_19617,N_18393);
and U22144 (N_22144,N_18259,N_15055);
and U22145 (N_22145,N_15264,N_16052);
xor U22146 (N_22146,N_17959,N_19400);
and U22147 (N_22147,N_15277,N_15648);
nand U22148 (N_22148,N_17490,N_17754);
or U22149 (N_22149,N_19131,N_18788);
and U22150 (N_22150,N_17634,N_16935);
and U22151 (N_22151,N_19222,N_19741);
nor U22152 (N_22152,N_15194,N_17566);
or U22153 (N_22153,N_18905,N_18029);
or U22154 (N_22154,N_18379,N_17156);
or U22155 (N_22155,N_16271,N_15018);
nand U22156 (N_22156,N_17399,N_17041);
and U22157 (N_22157,N_16302,N_17633);
and U22158 (N_22158,N_17076,N_16573);
nor U22159 (N_22159,N_16730,N_19951);
or U22160 (N_22160,N_15280,N_17210);
nand U22161 (N_22161,N_19279,N_18454);
or U22162 (N_22162,N_16711,N_18217);
or U22163 (N_22163,N_17974,N_18626);
nor U22164 (N_22164,N_19897,N_15436);
and U22165 (N_22165,N_18544,N_17825);
or U22166 (N_22166,N_18785,N_17093);
or U22167 (N_22167,N_18728,N_17204);
nand U22168 (N_22168,N_15771,N_17683);
or U22169 (N_22169,N_15045,N_17912);
nand U22170 (N_22170,N_16372,N_17996);
and U22171 (N_22171,N_19113,N_16880);
and U22172 (N_22172,N_18581,N_17528);
nor U22173 (N_22173,N_16085,N_18319);
or U22174 (N_22174,N_18002,N_15974);
or U22175 (N_22175,N_17616,N_18176);
and U22176 (N_22176,N_18113,N_17918);
or U22177 (N_22177,N_18927,N_15982);
or U22178 (N_22178,N_19473,N_18739);
and U22179 (N_22179,N_18854,N_18447);
or U22180 (N_22180,N_18277,N_16505);
nand U22181 (N_22181,N_15889,N_16439);
or U22182 (N_22182,N_17831,N_19064);
and U22183 (N_22183,N_16797,N_18091);
or U22184 (N_22184,N_18333,N_15268);
and U22185 (N_22185,N_19726,N_18422);
nand U22186 (N_22186,N_16564,N_19041);
or U22187 (N_22187,N_19442,N_16824);
and U22188 (N_22188,N_19981,N_16507);
xnor U22189 (N_22189,N_18678,N_19312);
nor U22190 (N_22190,N_17579,N_19558);
nand U22191 (N_22191,N_16647,N_15444);
and U22192 (N_22192,N_15944,N_19342);
and U22193 (N_22193,N_15270,N_18655);
or U22194 (N_22194,N_15896,N_15298);
xor U22195 (N_22195,N_18910,N_17627);
nand U22196 (N_22196,N_18022,N_16258);
or U22197 (N_22197,N_19356,N_17181);
nor U22198 (N_22198,N_18205,N_19295);
nor U22199 (N_22199,N_15604,N_16534);
nand U22200 (N_22200,N_18961,N_18443);
nand U22201 (N_22201,N_16633,N_17796);
nor U22202 (N_22202,N_19527,N_16993);
or U22203 (N_22203,N_17637,N_18312);
or U22204 (N_22204,N_16553,N_15543);
or U22205 (N_22205,N_17597,N_15841);
xnor U22206 (N_22206,N_16937,N_18061);
and U22207 (N_22207,N_19030,N_16551);
and U22208 (N_22208,N_15455,N_17690);
or U22209 (N_22209,N_16370,N_19249);
or U22210 (N_22210,N_16293,N_17772);
nor U22211 (N_22211,N_16339,N_18326);
nor U22212 (N_22212,N_16611,N_15566);
and U22213 (N_22213,N_17518,N_16606);
nor U22214 (N_22214,N_18036,N_19383);
or U22215 (N_22215,N_15463,N_16713);
nor U22216 (N_22216,N_15884,N_16868);
nor U22217 (N_22217,N_19185,N_16354);
and U22218 (N_22218,N_16585,N_18001);
or U22219 (N_22219,N_19540,N_16916);
nor U22220 (N_22220,N_16879,N_19022);
nor U22221 (N_22221,N_18700,N_18701);
nand U22222 (N_22222,N_19685,N_16383);
or U22223 (N_22223,N_16853,N_18662);
or U22224 (N_22224,N_17888,N_15289);
nand U22225 (N_22225,N_16078,N_16503);
nor U22226 (N_22226,N_16497,N_15971);
or U22227 (N_22227,N_18820,N_19678);
or U22228 (N_22228,N_17426,N_15069);
and U22229 (N_22229,N_18695,N_16546);
nor U22230 (N_22230,N_15065,N_17234);
or U22231 (N_22231,N_15863,N_16592);
nor U22232 (N_22232,N_15013,N_19637);
nor U22233 (N_22233,N_19838,N_18214);
nand U22234 (N_22234,N_17520,N_15110);
and U22235 (N_22235,N_15457,N_15766);
or U22236 (N_22236,N_19978,N_15100);
or U22237 (N_22237,N_16735,N_16947);
and U22238 (N_22238,N_18201,N_17575);
nor U22239 (N_22239,N_17428,N_16933);
xor U22240 (N_22240,N_18922,N_15400);
nor U22241 (N_22241,N_18599,N_19574);
or U22242 (N_22242,N_15388,N_19772);
nand U22243 (N_22243,N_17511,N_15589);
and U22244 (N_22244,N_17433,N_16991);
nor U22245 (N_22245,N_17707,N_15132);
or U22246 (N_22246,N_16504,N_15631);
xor U22247 (N_22247,N_15972,N_15169);
nand U22248 (N_22248,N_19247,N_17258);
and U22249 (N_22249,N_18606,N_17779);
and U22250 (N_22250,N_17611,N_18408);
nand U22251 (N_22251,N_15722,N_17799);
and U22252 (N_22252,N_19531,N_19555);
or U22253 (N_22253,N_17907,N_15876);
nand U22254 (N_22254,N_16764,N_15561);
and U22255 (N_22255,N_16754,N_19211);
and U22256 (N_22256,N_16502,N_16065);
or U22257 (N_22257,N_18582,N_18680);
nor U22258 (N_22258,N_18130,N_16201);
and U22259 (N_22259,N_17793,N_16976);
nand U22260 (N_22260,N_16539,N_18068);
nand U22261 (N_22261,N_17913,N_15068);
nor U22262 (N_22262,N_17809,N_15987);
nand U22263 (N_22263,N_16070,N_17134);
or U22264 (N_22264,N_17066,N_17753);
or U22265 (N_22265,N_17188,N_18499);
and U22266 (N_22266,N_15789,N_19641);
nor U22267 (N_22267,N_15570,N_17725);
nand U22268 (N_22268,N_18981,N_16310);
nor U22269 (N_22269,N_18132,N_19906);
nor U22270 (N_22270,N_19187,N_17956);
nor U22271 (N_22271,N_16988,N_19669);
or U22272 (N_22272,N_16584,N_16613);
nand U22273 (N_22273,N_18187,N_16431);
or U22274 (N_22274,N_16484,N_19449);
xor U22275 (N_22275,N_16562,N_15719);
nand U22276 (N_22276,N_15101,N_18964);
or U22277 (N_22277,N_19248,N_18793);
or U22278 (N_22278,N_17468,N_18766);
or U22279 (N_22279,N_17464,N_15394);
and U22280 (N_22280,N_18917,N_19426);
nor U22281 (N_22281,N_16790,N_19402);
or U22282 (N_22282,N_17946,N_15813);
nor U22283 (N_22283,N_19239,N_19955);
or U22284 (N_22284,N_16031,N_19046);
and U22285 (N_22285,N_15496,N_15547);
or U22286 (N_22286,N_15778,N_17312);
or U22287 (N_22287,N_16338,N_15871);
and U22288 (N_22288,N_17339,N_16059);
nand U22289 (N_22289,N_17572,N_19435);
nand U22290 (N_22290,N_18885,N_18565);
and U22291 (N_22291,N_19225,N_18798);
or U22292 (N_22292,N_15470,N_17355);
nand U22293 (N_22293,N_17294,N_19887);
or U22294 (N_22294,N_15803,N_18955);
nor U22295 (N_22295,N_15986,N_16183);
and U22296 (N_22296,N_18784,N_15411);
and U22297 (N_22297,N_18978,N_19731);
and U22298 (N_22298,N_18757,N_15123);
nor U22299 (N_22299,N_19815,N_16356);
nor U22300 (N_22300,N_19671,N_16506);
or U22301 (N_22301,N_18415,N_16182);
or U22302 (N_22302,N_19765,N_18133);
nand U22303 (N_22303,N_16242,N_16621);
nor U22304 (N_22304,N_18400,N_19513);
xnor U22305 (N_22305,N_15736,N_15824);
or U22306 (N_22306,N_19320,N_19303);
xor U22307 (N_22307,N_18056,N_15469);
and U22308 (N_22308,N_16985,N_19271);
or U22309 (N_22309,N_15865,N_18189);
nor U22310 (N_22310,N_15963,N_17504);
or U22311 (N_22311,N_18358,N_17448);
nor U22312 (N_22312,N_16922,N_19300);
nor U22313 (N_22313,N_19799,N_17400);
or U22314 (N_22314,N_19226,N_15178);
or U22315 (N_22315,N_16975,N_15753);
or U22316 (N_22316,N_17641,N_16039);
and U22317 (N_22317,N_16524,N_17246);
nor U22318 (N_22318,N_18388,N_19693);
and U22319 (N_22319,N_19056,N_17785);
and U22320 (N_22320,N_17720,N_19090);
nor U22321 (N_22321,N_18304,N_17314);
nand U22322 (N_22322,N_17625,N_18520);
and U22323 (N_22323,N_19007,N_15187);
nand U22324 (N_22324,N_18693,N_17640);
nand U22325 (N_22325,N_15907,N_19465);
nand U22326 (N_22326,N_19590,N_15116);
nand U22327 (N_22327,N_18533,N_17971);
or U22328 (N_22328,N_17737,N_18003);
or U22329 (N_22329,N_18871,N_15672);
or U22330 (N_22330,N_16493,N_18504);
nor U22331 (N_22331,N_18119,N_15168);
or U22332 (N_22332,N_15661,N_19623);
nor U22333 (N_22333,N_16712,N_18024);
and U22334 (N_22334,N_15551,N_16884);
or U22335 (N_22335,N_18849,N_18882);
and U22336 (N_22336,N_15867,N_18235);
and U22337 (N_22337,N_16131,N_16746);
nor U22338 (N_22338,N_18764,N_17668);
or U22339 (N_22339,N_19520,N_16535);
or U22340 (N_22340,N_15578,N_19350);
or U22341 (N_22341,N_16028,N_18817);
nand U22342 (N_22342,N_15774,N_17357);
nor U22343 (N_22343,N_19280,N_19180);
and U22344 (N_22344,N_17336,N_17459);
nand U22345 (N_22345,N_17436,N_17497);
nor U22346 (N_22346,N_17550,N_15861);
nand U22347 (N_22347,N_16422,N_18272);
nand U22348 (N_22348,N_19092,N_19708);
nor U22349 (N_22349,N_17709,N_16624);
or U22350 (N_22350,N_15427,N_19298);
and U22351 (N_22351,N_15374,N_19408);
nand U22352 (N_22352,N_17443,N_15575);
nand U22353 (N_22353,N_17370,N_15335);
xor U22354 (N_22354,N_19656,N_17984);
and U22355 (N_22355,N_17855,N_16050);
and U22356 (N_22356,N_17752,N_17324);
or U22357 (N_22357,N_19923,N_18159);
and U22358 (N_22358,N_15885,N_16610);
and U22359 (N_22359,N_19251,N_15954);
xor U22360 (N_22360,N_18780,N_15897);
nor U22361 (N_22361,N_15568,N_15654);
or U22362 (N_22362,N_17728,N_15704);
xnor U22363 (N_22363,N_15925,N_15120);
and U22364 (N_22364,N_17007,N_18902);
and U22365 (N_22365,N_17343,N_15145);
xnor U22366 (N_22366,N_16473,N_15376);
nor U22367 (N_22367,N_16955,N_17678);
and U22368 (N_22368,N_17536,N_19366);
nand U22369 (N_22369,N_18512,N_19106);
or U22370 (N_22370,N_15733,N_15994);
nor U22371 (N_22371,N_16865,N_18324);
nor U22372 (N_22372,N_17091,N_16426);
nand U22373 (N_22373,N_16745,N_16720);
nor U22374 (N_22374,N_16903,N_16590);
or U22375 (N_22375,N_18847,N_15628);
and U22376 (N_22376,N_15949,N_17654);
nand U22377 (N_22377,N_15615,N_18279);
nor U22378 (N_22378,N_17790,N_19576);
and U22379 (N_22379,N_19898,N_19634);
nand U22380 (N_22380,N_19639,N_17180);
and U22381 (N_22381,N_18050,N_15553);
nand U22382 (N_22382,N_18463,N_16424);
and U22383 (N_22383,N_18423,N_16676);
or U22384 (N_22384,N_16782,N_18099);
nor U22385 (N_22385,N_17108,N_18813);
and U22386 (N_22386,N_18859,N_17175);
and U22387 (N_22387,N_17635,N_17933);
and U22388 (N_22388,N_15129,N_18079);
nor U22389 (N_22389,N_15853,N_18681);
or U22390 (N_22390,N_16283,N_16311);
nor U22391 (N_22391,N_19613,N_16499);
nor U22392 (N_22392,N_19436,N_16861);
xor U22393 (N_22393,N_17574,N_15806);
or U22394 (N_22394,N_15688,N_18479);
or U22395 (N_22395,N_16235,N_18709);
and U22396 (N_22396,N_17240,N_18357);
and U22397 (N_22397,N_19109,N_16830);
nor U22398 (N_22398,N_17858,N_16591);
nand U22399 (N_22399,N_17981,N_18876);
nand U22400 (N_22400,N_16216,N_19543);
or U22401 (N_22401,N_17543,N_17565);
xor U22402 (N_22402,N_16804,N_15310);
nor U22403 (N_22403,N_16057,N_15996);
nand U22404 (N_22404,N_16393,N_17801);
nor U22405 (N_22405,N_15412,N_15369);
and U22406 (N_22406,N_15224,N_19593);
nand U22407 (N_22407,N_19759,N_15366);
or U22408 (N_22408,N_19702,N_16718);
or U22409 (N_22409,N_17756,N_16135);
nand U22410 (N_22410,N_19253,N_19412);
nor U22411 (N_22411,N_19337,N_17006);
nor U22412 (N_22412,N_16813,N_18592);
or U22413 (N_22413,N_19192,N_15221);
nand U22414 (N_22414,N_16570,N_15381);
or U22415 (N_22415,N_17847,N_15541);
nor U22416 (N_22416,N_15331,N_18901);
and U22417 (N_22417,N_16851,N_17092);
nand U22418 (N_22418,N_16758,N_18021);
nand U22419 (N_22419,N_16875,N_17106);
xnor U22420 (N_22420,N_18983,N_16810);
xor U22421 (N_22421,N_18494,N_18529);
or U22422 (N_22422,N_18837,N_15534);
nand U22423 (N_22423,N_16704,N_16488);
nand U22424 (N_22424,N_17208,N_17177);
nand U22425 (N_22425,N_16729,N_15859);
nand U22426 (N_22426,N_19362,N_15995);
and U22427 (N_22427,N_16464,N_17742);
nor U22428 (N_22428,N_17596,N_18775);
nand U22429 (N_22429,N_19646,N_16561);
nand U22430 (N_22430,N_15580,N_19992);
xnor U22431 (N_22431,N_16900,N_17420);
xnor U22432 (N_22432,N_17432,N_18440);
nor U22433 (N_22433,N_16388,N_16513);
or U22434 (N_22434,N_15669,N_17916);
nand U22435 (N_22435,N_16230,N_19130);
and U22436 (N_22436,N_16381,N_18740);
nand U22437 (N_22437,N_19208,N_17101);
nand U22438 (N_22438,N_15157,N_19373);
nand U22439 (N_22439,N_18979,N_17485);
and U22440 (N_22440,N_16918,N_19285);
nand U22441 (N_22441,N_19938,N_19873);
or U22442 (N_22442,N_19491,N_16805);
nor U22443 (N_22443,N_18802,N_15375);
or U22444 (N_22444,N_18568,N_17319);
or U22445 (N_22445,N_17393,N_15156);
nand U22446 (N_22446,N_16700,N_19803);
and U22447 (N_22447,N_18588,N_18191);
or U22448 (N_22448,N_15358,N_19994);
xnor U22449 (N_22449,N_16521,N_19502);
xnor U22450 (N_22450,N_15207,N_15155);
nor U22451 (N_22451,N_15037,N_15597);
nand U22452 (N_22452,N_16802,N_18426);
nand U22453 (N_22453,N_15942,N_17315);
and U22454 (N_22454,N_16541,N_15062);
xnor U22455 (N_22455,N_17488,N_19723);
or U22456 (N_22456,N_19780,N_16256);
or U22457 (N_22457,N_16029,N_16010);
or U22458 (N_22458,N_16213,N_17230);
nand U22459 (N_22459,N_18643,N_17326);
and U22460 (N_22460,N_16912,N_15490);
nand U22461 (N_22461,N_16934,N_19508);
nor U22462 (N_22462,N_15790,N_15617);
and U22463 (N_22463,N_19290,N_16263);
xor U22464 (N_22464,N_16117,N_17583);
and U22465 (N_22465,N_19635,N_19566);
or U22466 (N_22466,N_18234,N_15099);
nor U22467 (N_22467,N_16107,N_16982);
or U22468 (N_22468,N_18683,N_19292);
and U22469 (N_22469,N_19213,N_18553);
nand U22470 (N_22470,N_15483,N_18397);
or U22471 (N_22471,N_18714,N_19405);
nand U22472 (N_22472,N_15014,N_15780);
or U22473 (N_22473,N_17973,N_17182);
and U22474 (N_22474,N_15592,N_18583);
nor U22475 (N_22475,N_17561,N_17552);
nand U22476 (N_22476,N_18307,N_17245);
or U22477 (N_22477,N_19504,N_19471);
and U22478 (N_22478,N_18411,N_15743);
or U22479 (N_22479,N_17882,N_18814);
and U22480 (N_22480,N_18706,N_17923);
and U22481 (N_22481,N_15165,N_16374);
nor U22482 (N_22482,N_17179,N_16026);
or U22483 (N_22483,N_19553,N_19238);
xor U22484 (N_22484,N_18322,N_17898);
nor U22485 (N_22485,N_15041,N_18834);
or U22486 (N_22486,N_16009,N_19181);
nand U22487 (N_22487,N_15649,N_15354);
and U22488 (N_22488,N_17444,N_17895);
and U22489 (N_22489,N_19721,N_19882);
xnor U22490 (N_22490,N_17254,N_17624);
xnor U22491 (N_22491,N_16732,N_15082);
nand U22492 (N_22492,N_19953,N_17352);
nor U22493 (N_22493,N_17963,N_15011);
nor U22494 (N_22494,N_15393,N_15408);
or U22495 (N_22495,N_15465,N_17931);
or U22496 (N_22496,N_17699,N_18283);
xor U22497 (N_22497,N_18402,N_18270);
or U22498 (N_22498,N_16262,N_19762);
or U22499 (N_22499,N_18138,N_19434);
nand U22500 (N_22500,N_15463,N_17882);
and U22501 (N_22501,N_19017,N_16359);
or U22502 (N_22502,N_18603,N_15532);
nand U22503 (N_22503,N_18075,N_19885);
or U22504 (N_22504,N_16340,N_17208);
and U22505 (N_22505,N_18241,N_17810);
and U22506 (N_22506,N_18737,N_15289);
nand U22507 (N_22507,N_15365,N_16138);
nand U22508 (N_22508,N_15501,N_16157);
nand U22509 (N_22509,N_18721,N_18405);
and U22510 (N_22510,N_16739,N_19828);
xnor U22511 (N_22511,N_19052,N_17555);
or U22512 (N_22512,N_15933,N_19563);
and U22513 (N_22513,N_16440,N_18148);
nor U22514 (N_22514,N_15837,N_16053);
and U22515 (N_22515,N_17981,N_15287);
and U22516 (N_22516,N_15956,N_15656);
or U22517 (N_22517,N_18548,N_17457);
nand U22518 (N_22518,N_17063,N_15309);
or U22519 (N_22519,N_17901,N_19296);
nor U22520 (N_22520,N_15946,N_19579);
or U22521 (N_22521,N_18430,N_17918);
and U22522 (N_22522,N_15752,N_18064);
nand U22523 (N_22523,N_19877,N_16267);
or U22524 (N_22524,N_15993,N_19872);
nand U22525 (N_22525,N_18126,N_18411);
xnor U22526 (N_22526,N_18463,N_18753);
nor U22527 (N_22527,N_17048,N_17768);
nor U22528 (N_22528,N_19600,N_15383);
nand U22529 (N_22529,N_18513,N_16988);
nor U22530 (N_22530,N_18945,N_16751);
xnor U22531 (N_22531,N_17245,N_17598);
and U22532 (N_22532,N_16888,N_17375);
nand U22533 (N_22533,N_16229,N_16457);
nand U22534 (N_22534,N_19301,N_19465);
nand U22535 (N_22535,N_18052,N_16405);
xnor U22536 (N_22536,N_17161,N_15338);
nand U22537 (N_22537,N_15880,N_15700);
nor U22538 (N_22538,N_18728,N_16429);
or U22539 (N_22539,N_15136,N_17900);
nor U22540 (N_22540,N_17079,N_19669);
nor U22541 (N_22541,N_19397,N_17211);
and U22542 (N_22542,N_17619,N_18895);
and U22543 (N_22543,N_17119,N_17006);
or U22544 (N_22544,N_19520,N_18501);
and U22545 (N_22545,N_15104,N_16888);
or U22546 (N_22546,N_16608,N_17240);
nor U22547 (N_22547,N_16301,N_18942);
and U22548 (N_22548,N_19709,N_15312);
and U22549 (N_22549,N_18067,N_17938);
nand U22550 (N_22550,N_15132,N_15861);
nor U22551 (N_22551,N_17763,N_19136);
nand U22552 (N_22552,N_15881,N_16538);
nor U22553 (N_22553,N_19976,N_15385);
and U22554 (N_22554,N_16005,N_19214);
or U22555 (N_22555,N_17088,N_18333);
or U22556 (N_22556,N_16337,N_15582);
or U22557 (N_22557,N_17720,N_16199);
nand U22558 (N_22558,N_19229,N_15868);
nor U22559 (N_22559,N_18589,N_15085);
or U22560 (N_22560,N_19323,N_18063);
nand U22561 (N_22561,N_18146,N_18345);
and U22562 (N_22562,N_19367,N_15637);
or U22563 (N_22563,N_15956,N_19954);
and U22564 (N_22564,N_16143,N_18495);
and U22565 (N_22565,N_15283,N_16645);
nand U22566 (N_22566,N_16114,N_18937);
nand U22567 (N_22567,N_18620,N_17392);
nand U22568 (N_22568,N_18662,N_15225);
nand U22569 (N_22569,N_18244,N_18005);
nor U22570 (N_22570,N_19949,N_17707);
nand U22571 (N_22571,N_17197,N_18247);
and U22572 (N_22572,N_19265,N_16252);
and U22573 (N_22573,N_19910,N_17336);
nor U22574 (N_22574,N_18230,N_19360);
and U22575 (N_22575,N_17042,N_19748);
and U22576 (N_22576,N_19176,N_15675);
nor U22577 (N_22577,N_19697,N_15804);
nor U22578 (N_22578,N_15397,N_16255);
nor U22579 (N_22579,N_19652,N_17459);
or U22580 (N_22580,N_16289,N_15880);
nand U22581 (N_22581,N_19108,N_16418);
nor U22582 (N_22582,N_15294,N_19238);
nor U22583 (N_22583,N_15112,N_15682);
or U22584 (N_22584,N_18137,N_17006);
nor U22585 (N_22585,N_19511,N_19092);
or U22586 (N_22586,N_15022,N_17975);
nor U22587 (N_22587,N_19956,N_16063);
nand U22588 (N_22588,N_17038,N_18446);
and U22589 (N_22589,N_16843,N_16575);
or U22590 (N_22590,N_16175,N_17481);
and U22591 (N_22591,N_19857,N_17958);
nand U22592 (N_22592,N_17179,N_15343);
or U22593 (N_22593,N_18633,N_16476);
nand U22594 (N_22594,N_19632,N_17114);
or U22595 (N_22595,N_16356,N_19599);
or U22596 (N_22596,N_19096,N_16614);
nand U22597 (N_22597,N_16842,N_15399);
xor U22598 (N_22598,N_16302,N_17539);
and U22599 (N_22599,N_15615,N_16970);
or U22600 (N_22600,N_15979,N_16383);
or U22601 (N_22601,N_19265,N_17921);
or U22602 (N_22602,N_15868,N_17032);
nand U22603 (N_22603,N_16492,N_17349);
nand U22604 (N_22604,N_15673,N_19363);
or U22605 (N_22605,N_16017,N_17493);
nor U22606 (N_22606,N_18124,N_17801);
or U22607 (N_22607,N_17306,N_18324);
or U22608 (N_22608,N_15493,N_19801);
xnor U22609 (N_22609,N_18097,N_15320);
and U22610 (N_22610,N_15266,N_18479);
nand U22611 (N_22611,N_16362,N_17381);
nand U22612 (N_22612,N_18468,N_18926);
xor U22613 (N_22613,N_19175,N_15589);
nor U22614 (N_22614,N_18010,N_16874);
or U22615 (N_22615,N_18853,N_19011);
and U22616 (N_22616,N_15001,N_16015);
nand U22617 (N_22617,N_19989,N_17701);
xor U22618 (N_22618,N_16885,N_18595);
nor U22619 (N_22619,N_16005,N_17724);
or U22620 (N_22620,N_19607,N_18768);
nor U22621 (N_22621,N_15069,N_16594);
nand U22622 (N_22622,N_16044,N_17523);
and U22623 (N_22623,N_17418,N_18650);
nand U22624 (N_22624,N_16680,N_19107);
nor U22625 (N_22625,N_16413,N_17568);
xnor U22626 (N_22626,N_15221,N_17475);
or U22627 (N_22627,N_15452,N_15973);
nand U22628 (N_22628,N_17368,N_18582);
or U22629 (N_22629,N_15290,N_18360);
xor U22630 (N_22630,N_18604,N_15756);
or U22631 (N_22631,N_19342,N_15618);
or U22632 (N_22632,N_18695,N_15795);
nor U22633 (N_22633,N_18689,N_19192);
and U22634 (N_22634,N_15358,N_18211);
xnor U22635 (N_22635,N_18442,N_18617);
nand U22636 (N_22636,N_17274,N_18426);
nand U22637 (N_22637,N_16200,N_18276);
nand U22638 (N_22638,N_17960,N_17586);
nor U22639 (N_22639,N_15991,N_18797);
or U22640 (N_22640,N_15250,N_19650);
nand U22641 (N_22641,N_16698,N_17163);
or U22642 (N_22642,N_17799,N_16076);
nor U22643 (N_22643,N_18133,N_19658);
xnor U22644 (N_22644,N_19446,N_17340);
nand U22645 (N_22645,N_15429,N_18983);
nand U22646 (N_22646,N_15121,N_18835);
nor U22647 (N_22647,N_18302,N_17000);
or U22648 (N_22648,N_16980,N_19154);
and U22649 (N_22649,N_15105,N_15315);
or U22650 (N_22650,N_16674,N_17779);
and U22651 (N_22651,N_15274,N_15522);
nand U22652 (N_22652,N_15368,N_17033);
or U22653 (N_22653,N_17643,N_18432);
and U22654 (N_22654,N_17442,N_18223);
xnor U22655 (N_22655,N_17230,N_16352);
and U22656 (N_22656,N_15011,N_17465);
and U22657 (N_22657,N_19283,N_16700);
and U22658 (N_22658,N_15642,N_16533);
xor U22659 (N_22659,N_19948,N_17819);
and U22660 (N_22660,N_16376,N_15156);
or U22661 (N_22661,N_19397,N_18084);
nor U22662 (N_22662,N_15760,N_15329);
nand U22663 (N_22663,N_18389,N_17969);
and U22664 (N_22664,N_15612,N_18651);
or U22665 (N_22665,N_16752,N_17459);
or U22666 (N_22666,N_17024,N_18107);
and U22667 (N_22667,N_16453,N_19419);
nor U22668 (N_22668,N_17278,N_17450);
or U22669 (N_22669,N_18417,N_18770);
nor U22670 (N_22670,N_18829,N_18871);
nor U22671 (N_22671,N_17120,N_19472);
or U22672 (N_22672,N_15127,N_16271);
and U22673 (N_22673,N_17068,N_18444);
or U22674 (N_22674,N_16371,N_15788);
nand U22675 (N_22675,N_19179,N_19983);
or U22676 (N_22676,N_18624,N_15889);
and U22677 (N_22677,N_19721,N_18136);
and U22678 (N_22678,N_16152,N_16338);
and U22679 (N_22679,N_18464,N_17702);
or U22680 (N_22680,N_17541,N_18423);
or U22681 (N_22681,N_16525,N_17742);
or U22682 (N_22682,N_19962,N_16604);
or U22683 (N_22683,N_18379,N_16760);
or U22684 (N_22684,N_15369,N_19427);
or U22685 (N_22685,N_16453,N_15277);
nand U22686 (N_22686,N_19939,N_19305);
nor U22687 (N_22687,N_17947,N_18655);
nand U22688 (N_22688,N_17161,N_19296);
and U22689 (N_22689,N_17660,N_19339);
and U22690 (N_22690,N_16577,N_15415);
or U22691 (N_22691,N_18321,N_19401);
nand U22692 (N_22692,N_16117,N_19147);
nand U22693 (N_22693,N_17992,N_16020);
or U22694 (N_22694,N_16156,N_19646);
nor U22695 (N_22695,N_17713,N_18888);
nor U22696 (N_22696,N_18393,N_18279);
and U22697 (N_22697,N_17552,N_15293);
nand U22698 (N_22698,N_16314,N_15930);
or U22699 (N_22699,N_15594,N_15330);
nand U22700 (N_22700,N_18063,N_17259);
nor U22701 (N_22701,N_19505,N_18227);
nand U22702 (N_22702,N_18002,N_18447);
or U22703 (N_22703,N_18789,N_16914);
or U22704 (N_22704,N_16923,N_16254);
and U22705 (N_22705,N_15925,N_17178);
nor U22706 (N_22706,N_15129,N_15309);
and U22707 (N_22707,N_17663,N_15193);
or U22708 (N_22708,N_16193,N_16087);
and U22709 (N_22709,N_16196,N_16034);
and U22710 (N_22710,N_15424,N_19825);
nand U22711 (N_22711,N_17279,N_19257);
and U22712 (N_22712,N_18227,N_16846);
nand U22713 (N_22713,N_19934,N_16503);
nand U22714 (N_22714,N_18286,N_15961);
nand U22715 (N_22715,N_16720,N_17814);
nand U22716 (N_22716,N_19250,N_15422);
nor U22717 (N_22717,N_18400,N_17762);
or U22718 (N_22718,N_17049,N_19934);
xnor U22719 (N_22719,N_17989,N_16905);
nand U22720 (N_22720,N_17634,N_19106);
nand U22721 (N_22721,N_16191,N_19391);
nor U22722 (N_22722,N_16714,N_15082);
nand U22723 (N_22723,N_17655,N_19523);
nand U22724 (N_22724,N_18963,N_15696);
nand U22725 (N_22725,N_17671,N_16681);
and U22726 (N_22726,N_16682,N_16661);
or U22727 (N_22727,N_15813,N_16795);
or U22728 (N_22728,N_19070,N_15467);
nor U22729 (N_22729,N_15038,N_18545);
and U22730 (N_22730,N_18885,N_17853);
nand U22731 (N_22731,N_16811,N_18861);
or U22732 (N_22732,N_15290,N_17957);
nor U22733 (N_22733,N_15299,N_16371);
and U22734 (N_22734,N_18714,N_17096);
and U22735 (N_22735,N_19727,N_18944);
or U22736 (N_22736,N_16310,N_15360);
and U22737 (N_22737,N_15960,N_16743);
and U22738 (N_22738,N_18185,N_18306);
or U22739 (N_22739,N_19945,N_15594);
and U22740 (N_22740,N_17626,N_15963);
nor U22741 (N_22741,N_16243,N_19079);
or U22742 (N_22742,N_19746,N_19280);
and U22743 (N_22743,N_15680,N_16100);
nor U22744 (N_22744,N_15497,N_15354);
and U22745 (N_22745,N_17221,N_16349);
and U22746 (N_22746,N_15653,N_18996);
and U22747 (N_22747,N_16520,N_16544);
nor U22748 (N_22748,N_15428,N_15813);
xor U22749 (N_22749,N_16083,N_19808);
and U22750 (N_22750,N_17714,N_17370);
xor U22751 (N_22751,N_15890,N_18672);
nand U22752 (N_22752,N_18424,N_17446);
nor U22753 (N_22753,N_15456,N_16536);
nor U22754 (N_22754,N_17310,N_19755);
nor U22755 (N_22755,N_16335,N_18437);
nand U22756 (N_22756,N_19042,N_17312);
and U22757 (N_22757,N_15445,N_17799);
or U22758 (N_22758,N_17207,N_16339);
nor U22759 (N_22759,N_15754,N_18489);
or U22760 (N_22760,N_16770,N_16225);
and U22761 (N_22761,N_17598,N_15887);
nand U22762 (N_22762,N_16405,N_18879);
and U22763 (N_22763,N_17072,N_19114);
nor U22764 (N_22764,N_18361,N_18244);
or U22765 (N_22765,N_19160,N_17493);
nor U22766 (N_22766,N_16965,N_16745);
and U22767 (N_22767,N_18582,N_15937);
nand U22768 (N_22768,N_15853,N_16424);
nor U22769 (N_22769,N_19553,N_18889);
and U22770 (N_22770,N_16773,N_17442);
and U22771 (N_22771,N_16512,N_19960);
xor U22772 (N_22772,N_16613,N_15867);
nor U22773 (N_22773,N_17697,N_17199);
and U22774 (N_22774,N_17536,N_16313);
or U22775 (N_22775,N_15495,N_17645);
nor U22776 (N_22776,N_15538,N_18646);
nor U22777 (N_22777,N_16748,N_18213);
and U22778 (N_22778,N_18769,N_19536);
xor U22779 (N_22779,N_16234,N_18805);
nor U22780 (N_22780,N_17120,N_19918);
xor U22781 (N_22781,N_15038,N_19521);
nor U22782 (N_22782,N_16320,N_17580);
or U22783 (N_22783,N_15180,N_18689);
and U22784 (N_22784,N_19380,N_16194);
and U22785 (N_22785,N_18314,N_15749);
nand U22786 (N_22786,N_17193,N_19927);
and U22787 (N_22787,N_17865,N_15055);
and U22788 (N_22788,N_18329,N_15939);
or U22789 (N_22789,N_19679,N_19741);
xnor U22790 (N_22790,N_15313,N_15037);
and U22791 (N_22791,N_18386,N_18013);
or U22792 (N_22792,N_19918,N_18892);
nor U22793 (N_22793,N_15663,N_15136);
and U22794 (N_22794,N_16046,N_19796);
nand U22795 (N_22795,N_18336,N_17309);
nor U22796 (N_22796,N_16310,N_15871);
nand U22797 (N_22797,N_17588,N_15128);
nand U22798 (N_22798,N_16631,N_18706);
nor U22799 (N_22799,N_18235,N_18108);
nand U22800 (N_22800,N_15240,N_19885);
or U22801 (N_22801,N_16348,N_18676);
xnor U22802 (N_22802,N_15560,N_17079);
or U22803 (N_22803,N_17740,N_16047);
and U22804 (N_22804,N_17001,N_18038);
or U22805 (N_22805,N_15711,N_17627);
nor U22806 (N_22806,N_15658,N_17741);
nand U22807 (N_22807,N_18148,N_18445);
nand U22808 (N_22808,N_18069,N_17370);
nor U22809 (N_22809,N_16548,N_18586);
nand U22810 (N_22810,N_17878,N_16206);
or U22811 (N_22811,N_16307,N_16997);
nor U22812 (N_22812,N_17490,N_17004);
nand U22813 (N_22813,N_19056,N_16097);
nor U22814 (N_22814,N_17650,N_16672);
nand U22815 (N_22815,N_16289,N_15505);
or U22816 (N_22816,N_19525,N_15974);
xnor U22817 (N_22817,N_19894,N_15915);
and U22818 (N_22818,N_17688,N_16161);
and U22819 (N_22819,N_15200,N_16303);
or U22820 (N_22820,N_17321,N_19004);
nand U22821 (N_22821,N_15708,N_17145);
or U22822 (N_22822,N_15641,N_16697);
and U22823 (N_22823,N_15503,N_19029);
or U22824 (N_22824,N_19269,N_19239);
and U22825 (N_22825,N_16137,N_16070);
nor U22826 (N_22826,N_16263,N_16276);
nor U22827 (N_22827,N_18507,N_17947);
nand U22828 (N_22828,N_17052,N_19925);
nor U22829 (N_22829,N_18295,N_18164);
and U22830 (N_22830,N_19289,N_17945);
nand U22831 (N_22831,N_19475,N_17001);
nor U22832 (N_22832,N_17761,N_17882);
nor U22833 (N_22833,N_17623,N_16386);
nor U22834 (N_22834,N_18752,N_16795);
nand U22835 (N_22835,N_19939,N_19634);
and U22836 (N_22836,N_18371,N_18266);
xnor U22837 (N_22837,N_16441,N_18495);
and U22838 (N_22838,N_17635,N_17822);
nor U22839 (N_22839,N_15809,N_15102);
xor U22840 (N_22840,N_16369,N_18112);
nand U22841 (N_22841,N_16137,N_15851);
or U22842 (N_22842,N_18284,N_15165);
nor U22843 (N_22843,N_17718,N_17643);
and U22844 (N_22844,N_16151,N_17790);
nand U22845 (N_22845,N_15392,N_15437);
or U22846 (N_22846,N_17031,N_19535);
nand U22847 (N_22847,N_15212,N_16778);
xor U22848 (N_22848,N_16181,N_17196);
xor U22849 (N_22849,N_17061,N_19690);
or U22850 (N_22850,N_19371,N_16113);
nor U22851 (N_22851,N_19497,N_16982);
and U22852 (N_22852,N_15568,N_18325);
and U22853 (N_22853,N_19384,N_16228);
and U22854 (N_22854,N_18266,N_17743);
nand U22855 (N_22855,N_15887,N_15271);
nor U22856 (N_22856,N_18380,N_17015);
or U22857 (N_22857,N_19779,N_16457);
nand U22858 (N_22858,N_18573,N_18937);
nand U22859 (N_22859,N_18829,N_19482);
nor U22860 (N_22860,N_19599,N_17517);
nand U22861 (N_22861,N_15802,N_18327);
and U22862 (N_22862,N_16936,N_19503);
nor U22863 (N_22863,N_16266,N_15636);
and U22864 (N_22864,N_17649,N_19195);
and U22865 (N_22865,N_18422,N_19763);
and U22866 (N_22866,N_16182,N_19503);
nand U22867 (N_22867,N_17221,N_16689);
or U22868 (N_22868,N_15639,N_17023);
or U22869 (N_22869,N_17149,N_16515);
and U22870 (N_22870,N_19321,N_17111);
nor U22871 (N_22871,N_19013,N_17052);
or U22872 (N_22872,N_15625,N_15610);
nor U22873 (N_22873,N_18270,N_17660);
and U22874 (N_22874,N_18179,N_19848);
and U22875 (N_22875,N_18667,N_15647);
nor U22876 (N_22876,N_17178,N_19173);
nand U22877 (N_22877,N_16851,N_18222);
and U22878 (N_22878,N_15395,N_17533);
nor U22879 (N_22879,N_15688,N_15034);
or U22880 (N_22880,N_17411,N_15091);
nand U22881 (N_22881,N_15816,N_17523);
nor U22882 (N_22882,N_15249,N_15302);
nor U22883 (N_22883,N_16313,N_19703);
nand U22884 (N_22884,N_15502,N_17944);
and U22885 (N_22885,N_16637,N_15978);
and U22886 (N_22886,N_16701,N_15373);
or U22887 (N_22887,N_15122,N_19007);
or U22888 (N_22888,N_17219,N_16773);
or U22889 (N_22889,N_18550,N_19211);
nand U22890 (N_22890,N_15713,N_19134);
or U22891 (N_22891,N_18933,N_18700);
or U22892 (N_22892,N_16355,N_15844);
or U22893 (N_22893,N_17294,N_18769);
and U22894 (N_22894,N_19768,N_15055);
or U22895 (N_22895,N_18439,N_19227);
and U22896 (N_22896,N_18917,N_16158);
nor U22897 (N_22897,N_18873,N_19225);
or U22898 (N_22898,N_16307,N_17358);
nor U22899 (N_22899,N_16710,N_17174);
and U22900 (N_22900,N_19906,N_19673);
nand U22901 (N_22901,N_16236,N_18356);
xor U22902 (N_22902,N_19194,N_17242);
nand U22903 (N_22903,N_18549,N_15810);
or U22904 (N_22904,N_17145,N_19670);
or U22905 (N_22905,N_16945,N_18556);
or U22906 (N_22906,N_15448,N_16243);
and U22907 (N_22907,N_19545,N_15755);
and U22908 (N_22908,N_19311,N_16874);
nor U22909 (N_22909,N_17509,N_17031);
nor U22910 (N_22910,N_18222,N_15743);
xnor U22911 (N_22911,N_15115,N_16042);
nand U22912 (N_22912,N_17719,N_19511);
nand U22913 (N_22913,N_17023,N_16535);
or U22914 (N_22914,N_18356,N_16742);
nand U22915 (N_22915,N_19939,N_16769);
or U22916 (N_22916,N_19054,N_17114);
and U22917 (N_22917,N_15052,N_18911);
xnor U22918 (N_22918,N_16280,N_17399);
nor U22919 (N_22919,N_19095,N_19785);
and U22920 (N_22920,N_16539,N_15036);
nor U22921 (N_22921,N_15533,N_19922);
xnor U22922 (N_22922,N_15678,N_18243);
and U22923 (N_22923,N_19114,N_18224);
xnor U22924 (N_22924,N_15185,N_18549);
nor U22925 (N_22925,N_17263,N_16276);
or U22926 (N_22926,N_19940,N_18552);
or U22927 (N_22927,N_19905,N_17785);
nand U22928 (N_22928,N_16662,N_18879);
nand U22929 (N_22929,N_16095,N_17634);
xor U22930 (N_22930,N_18056,N_18832);
or U22931 (N_22931,N_18049,N_15701);
xnor U22932 (N_22932,N_19869,N_19337);
or U22933 (N_22933,N_15743,N_16042);
or U22934 (N_22934,N_18203,N_17884);
nor U22935 (N_22935,N_17902,N_17868);
and U22936 (N_22936,N_17477,N_17872);
nand U22937 (N_22937,N_19119,N_18119);
or U22938 (N_22938,N_18894,N_17043);
and U22939 (N_22939,N_19615,N_15991);
nor U22940 (N_22940,N_16345,N_18553);
and U22941 (N_22941,N_19456,N_16037);
xor U22942 (N_22942,N_15822,N_19155);
or U22943 (N_22943,N_16207,N_18079);
nor U22944 (N_22944,N_15739,N_18699);
and U22945 (N_22945,N_17826,N_17029);
nor U22946 (N_22946,N_16165,N_17313);
nand U22947 (N_22947,N_19758,N_18493);
nand U22948 (N_22948,N_16587,N_17679);
nor U22949 (N_22949,N_17682,N_19512);
or U22950 (N_22950,N_19084,N_17420);
nand U22951 (N_22951,N_19263,N_15828);
and U22952 (N_22952,N_17609,N_16691);
or U22953 (N_22953,N_16221,N_15427);
or U22954 (N_22954,N_18059,N_19462);
or U22955 (N_22955,N_19854,N_16115);
or U22956 (N_22956,N_17932,N_17148);
or U22957 (N_22957,N_19130,N_18145);
nand U22958 (N_22958,N_16335,N_15398);
or U22959 (N_22959,N_16446,N_19834);
and U22960 (N_22960,N_19357,N_18054);
nor U22961 (N_22961,N_18093,N_15349);
nor U22962 (N_22962,N_16706,N_19614);
nand U22963 (N_22963,N_15632,N_16123);
nor U22964 (N_22964,N_17775,N_18480);
and U22965 (N_22965,N_16599,N_18490);
nand U22966 (N_22966,N_18414,N_17312);
nor U22967 (N_22967,N_16155,N_16120);
xor U22968 (N_22968,N_18365,N_19552);
nor U22969 (N_22969,N_16175,N_18374);
nor U22970 (N_22970,N_15939,N_18937);
nor U22971 (N_22971,N_16459,N_15488);
and U22972 (N_22972,N_17970,N_18770);
nand U22973 (N_22973,N_16975,N_15887);
nor U22974 (N_22974,N_19033,N_19306);
or U22975 (N_22975,N_15774,N_18184);
nand U22976 (N_22976,N_15816,N_17026);
and U22977 (N_22977,N_15682,N_16440);
or U22978 (N_22978,N_17478,N_16388);
nand U22979 (N_22979,N_19869,N_15315);
and U22980 (N_22980,N_16259,N_17580);
nor U22981 (N_22981,N_17967,N_16406);
nor U22982 (N_22982,N_17100,N_18130);
and U22983 (N_22983,N_18606,N_15958);
nor U22984 (N_22984,N_19957,N_19041);
xnor U22985 (N_22985,N_15744,N_15497);
or U22986 (N_22986,N_17648,N_16489);
xor U22987 (N_22987,N_19028,N_19605);
xnor U22988 (N_22988,N_19666,N_17520);
nand U22989 (N_22989,N_15879,N_17636);
nor U22990 (N_22990,N_16459,N_19573);
nor U22991 (N_22991,N_16390,N_16807);
or U22992 (N_22992,N_16998,N_19201);
and U22993 (N_22993,N_15965,N_16972);
nor U22994 (N_22994,N_17068,N_15424);
and U22995 (N_22995,N_19090,N_16388);
and U22996 (N_22996,N_19676,N_16831);
nand U22997 (N_22997,N_19265,N_19781);
and U22998 (N_22998,N_15462,N_19355);
nand U22999 (N_22999,N_15962,N_18385);
and U23000 (N_23000,N_18473,N_16146);
or U23001 (N_23001,N_16596,N_18091);
and U23002 (N_23002,N_16564,N_18623);
nor U23003 (N_23003,N_19791,N_19943);
nand U23004 (N_23004,N_16862,N_16982);
and U23005 (N_23005,N_15042,N_18503);
nand U23006 (N_23006,N_17080,N_15520);
nand U23007 (N_23007,N_17142,N_19794);
and U23008 (N_23008,N_15391,N_17941);
or U23009 (N_23009,N_19330,N_17453);
nor U23010 (N_23010,N_19577,N_15159);
nand U23011 (N_23011,N_16773,N_18832);
xor U23012 (N_23012,N_15931,N_18889);
nor U23013 (N_23013,N_15402,N_16253);
nand U23014 (N_23014,N_19458,N_19331);
nand U23015 (N_23015,N_17711,N_18416);
nand U23016 (N_23016,N_16972,N_19203);
or U23017 (N_23017,N_19069,N_15718);
or U23018 (N_23018,N_17692,N_16865);
or U23019 (N_23019,N_16383,N_15844);
xor U23020 (N_23020,N_19323,N_16448);
nor U23021 (N_23021,N_18838,N_16635);
or U23022 (N_23022,N_19493,N_16599);
and U23023 (N_23023,N_15468,N_18882);
or U23024 (N_23024,N_18498,N_17691);
and U23025 (N_23025,N_17852,N_15243);
nor U23026 (N_23026,N_16981,N_17083);
nor U23027 (N_23027,N_15169,N_18412);
nand U23028 (N_23028,N_19821,N_15563);
or U23029 (N_23029,N_19682,N_15581);
or U23030 (N_23030,N_17093,N_19362);
and U23031 (N_23031,N_16672,N_19871);
nor U23032 (N_23032,N_19779,N_15173);
nand U23033 (N_23033,N_17133,N_18400);
or U23034 (N_23034,N_15274,N_16159);
nand U23035 (N_23035,N_17658,N_19196);
or U23036 (N_23036,N_16485,N_19964);
nor U23037 (N_23037,N_17504,N_18822);
and U23038 (N_23038,N_15163,N_19461);
nor U23039 (N_23039,N_15908,N_15196);
and U23040 (N_23040,N_18673,N_17410);
xor U23041 (N_23041,N_19736,N_18180);
nand U23042 (N_23042,N_18674,N_19090);
or U23043 (N_23043,N_17595,N_17152);
nor U23044 (N_23044,N_15468,N_15545);
nand U23045 (N_23045,N_15571,N_16538);
or U23046 (N_23046,N_15002,N_17699);
nor U23047 (N_23047,N_15243,N_19563);
and U23048 (N_23048,N_16329,N_17852);
or U23049 (N_23049,N_15213,N_15838);
or U23050 (N_23050,N_18828,N_17674);
or U23051 (N_23051,N_16999,N_19020);
nor U23052 (N_23052,N_18290,N_18715);
and U23053 (N_23053,N_17701,N_18442);
nand U23054 (N_23054,N_18434,N_18412);
and U23055 (N_23055,N_15861,N_18710);
and U23056 (N_23056,N_19904,N_15935);
or U23057 (N_23057,N_17616,N_17217);
and U23058 (N_23058,N_16148,N_17776);
and U23059 (N_23059,N_17515,N_15361);
nor U23060 (N_23060,N_18658,N_17332);
xor U23061 (N_23061,N_16076,N_18639);
nand U23062 (N_23062,N_19334,N_16605);
and U23063 (N_23063,N_18556,N_17652);
nand U23064 (N_23064,N_15590,N_15240);
and U23065 (N_23065,N_16341,N_16801);
and U23066 (N_23066,N_19613,N_19846);
and U23067 (N_23067,N_19339,N_18015);
nor U23068 (N_23068,N_15697,N_17852);
or U23069 (N_23069,N_18290,N_15228);
nand U23070 (N_23070,N_19739,N_17987);
and U23071 (N_23071,N_17088,N_15732);
nand U23072 (N_23072,N_15748,N_19971);
nor U23073 (N_23073,N_17879,N_15287);
xnor U23074 (N_23074,N_16012,N_17261);
and U23075 (N_23075,N_19221,N_19298);
or U23076 (N_23076,N_16634,N_16471);
nor U23077 (N_23077,N_19802,N_16878);
or U23078 (N_23078,N_17804,N_16422);
nor U23079 (N_23079,N_18498,N_17996);
nor U23080 (N_23080,N_16874,N_18004);
nand U23081 (N_23081,N_19322,N_19224);
nor U23082 (N_23082,N_15465,N_18647);
or U23083 (N_23083,N_17024,N_15793);
nand U23084 (N_23084,N_19939,N_17077);
nand U23085 (N_23085,N_19620,N_16006);
nand U23086 (N_23086,N_18552,N_15037);
and U23087 (N_23087,N_18861,N_15676);
and U23088 (N_23088,N_16198,N_17859);
and U23089 (N_23089,N_16185,N_18162);
nand U23090 (N_23090,N_19005,N_17548);
nor U23091 (N_23091,N_17284,N_16540);
nor U23092 (N_23092,N_18040,N_18283);
and U23093 (N_23093,N_18286,N_19418);
or U23094 (N_23094,N_15341,N_17886);
nor U23095 (N_23095,N_16239,N_15272);
nand U23096 (N_23096,N_15775,N_18841);
nand U23097 (N_23097,N_16200,N_17526);
and U23098 (N_23098,N_19759,N_15419);
or U23099 (N_23099,N_19911,N_19808);
and U23100 (N_23100,N_16382,N_15630);
or U23101 (N_23101,N_15189,N_17631);
nor U23102 (N_23102,N_15578,N_18247);
or U23103 (N_23103,N_19621,N_15481);
nand U23104 (N_23104,N_15889,N_17362);
xnor U23105 (N_23105,N_18596,N_17570);
and U23106 (N_23106,N_19495,N_16086);
nor U23107 (N_23107,N_17215,N_15857);
or U23108 (N_23108,N_19797,N_18263);
and U23109 (N_23109,N_15493,N_15963);
and U23110 (N_23110,N_18431,N_15917);
and U23111 (N_23111,N_17558,N_16069);
nor U23112 (N_23112,N_18535,N_17403);
nor U23113 (N_23113,N_15963,N_19363);
and U23114 (N_23114,N_15634,N_16842);
xor U23115 (N_23115,N_16274,N_19773);
nand U23116 (N_23116,N_17080,N_17952);
nand U23117 (N_23117,N_16492,N_16071);
or U23118 (N_23118,N_17277,N_15912);
or U23119 (N_23119,N_15141,N_19304);
nor U23120 (N_23120,N_18009,N_19310);
nand U23121 (N_23121,N_17563,N_18625);
nand U23122 (N_23122,N_17202,N_17452);
nor U23123 (N_23123,N_17142,N_15335);
and U23124 (N_23124,N_16089,N_17984);
nand U23125 (N_23125,N_15144,N_18032);
nand U23126 (N_23126,N_15929,N_17656);
nor U23127 (N_23127,N_17736,N_18227);
nand U23128 (N_23128,N_16294,N_15913);
or U23129 (N_23129,N_17551,N_16113);
nand U23130 (N_23130,N_19869,N_17233);
or U23131 (N_23131,N_15766,N_17053);
or U23132 (N_23132,N_17293,N_17394);
or U23133 (N_23133,N_15405,N_18357);
xor U23134 (N_23134,N_15488,N_15357);
nand U23135 (N_23135,N_15569,N_16863);
xor U23136 (N_23136,N_17169,N_19521);
or U23137 (N_23137,N_17495,N_15919);
nand U23138 (N_23138,N_16751,N_18494);
nor U23139 (N_23139,N_15499,N_17045);
nand U23140 (N_23140,N_18949,N_16592);
and U23141 (N_23141,N_17203,N_15115);
and U23142 (N_23142,N_15124,N_18282);
nand U23143 (N_23143,N_15487,N_17467);
nor U23144 (N_23144,N_16602,N_16944);
nand U23145 (N_23145,N_15896,N_16883);
nand U23146 (N_23146,N_19387,N_16642);
and U23147 (N_23147,N_15628,N_19407);
or U23148 (N_23148,N_19686,N_16527);
or U23149 (N_23149,N_16793,N_18850);
xnor U23150 (N_23150,N_18603,N_17489);
or U23151 (N_23151,N_18281,N_18016);
nor U23152 (N_23152,N_19191,N_17812);
and U23153 (N_23153,N_19443,N_19801);
nand U23154 (N_23154,N_19914,N_17995);
xor U23155 (N_23155,N_17618,N_18254);
nor U23156 (N_23156,N_17561,N_19069);
or U23157 (N_23157,N_16319,N_16077);
nand U23158 (N_23158,N_17550,N_16098);
nor U23159 (N_23159,N_16049,N_16316);
nor U23160 (N_23160,N_16465,N_19246);
or U23161 (N_23161,N_19056,N_18591);
or U23162 (N_23162,N_15343,N_17802);
nand U23163 (N_23163,N_15519,N_16287);
nand U23164 (N_23164,N_19564,N_17223);
nor U23165 (N_23165,N_18468,N_17526);
or U23166 (N_23166,N_18339,N_18189);
nand U23167 (N_23167,N_19098,N_19678);
or U23168 (N_23168,N_16043,N_19663);
and U23169 (N_23169,N_15066,N_19195);
nand U23170 (N_23170,N_19497,N_17378);
nand U23171 (N_23171,N_17674,N_18097);
and U23172 (N_23172,N_17031,N_16960);
or U23173 (N_23173,N_19592,N_16363);
nand U23174 (N_23174,N_16506,N_18058);
nor U23175 (N_23175,N_17036,N_15727);
nor U23176 (N_23176,N_15869,N_19237);
nor U23177 (N_23177,N_15059,N_19236);
nand U23178 (N_23178,N_16490,N_19486);
or U23179 (N_23179,N_16931,N_19726);
nor U23180 (N_23180,N_18048,N_16660);
or U23181 (N_23181,N_19549,N_18158);
nor U23182 (N_23182,N_15799,N_19732);
and U23183 (N_23183,N_16845,N_18098);
nor U23184 (N_23184,N_17442,N_18405);
or U23185 (N_23185,N_18361,N_19519);
and U23186 (N_23186,N_19613,N_17900);
nor U23187 (N_23187,N_18232,N_15243);
xnor U23188 (N_23188,N_15779,N_18841);
nor U23189 (N_23189,N_16977,N_19249);
and U23190 (N_23190,N_15713,N_16107);
nand U23191 (N_23191,N_16453,N_16160);
nand U23192 (N_23192,N_19645,N_18481);
xnor U23193 (N_23193,N_16426,N_19947);
and U23194 (N_23194,N_15433,N_19818);
or U23195 (N_23195,N_17207,N_19890);
nor U23196 (N_23196,N_19814,N_17549);
and U23197 (N_23197,N_19940,N_18637);
or U23198 (N_23198,N_17549,N_16353);
and U23199 (N_23199,N_19936,N_19721);
or U23200 (N_23200,N_16604,N_17093);
nor U23201 (N_23201,N_18947,N_16981);
and U23202 (N_23202,N_15255,N_19122);
nand U23203 (N_23203,N_16457,N_19916);
and U23204 (N_23204,N_15517,N_17019);
nor U23205 (N_23205,N_17452,N_17797);
nand U23206 (N_23206,N_18990,N_17755);
nor U23207 (N_23207,N_19544,N_18956);
nor U23208 (N_23208,N_17906,N_16867);
or U23209 (N_23209,N_17627,N_15223);
nand U23210 (N_23210,N_19236,N_18408);
and U23211 (N_23211,N_19630,N_18473);
and U23212 (N_23212,N_15495,N_19334);
nor U23213 (N_23213,N_15419,N_15005);
nor U23214 (N_23214,N_16173,N_19133);
xnor U23215 (N_23215,N_15325,N_17015);
nor U23216 (N_23216,N_17053,N_19691);
nand U23217 (N_23217,N_19524,N_17807);
and U23218 (N_23218,N_18972,N_16316);
and U23219 (N_23219,N_18302,N_18883);
nor U23220 (N_23220,N_15628,N_15517);
nor U23221 (N_23221,N_16889,N_15763);
xnor U23222 (N_23222,N_16284,N_19716);
or U23223 (N_23223,N_16990,N_18605);
xor U23224 (N_23224,N_15138,N_17911);
nor U23225 (N_23225,N_15368,N_15721);
nand U23226 (N_23226,N_15826,N_16510);
nand U23227 (N_23227,N_17586,N_15883);
nand U23228 (N_23228,N_18591,N_19847);
and U23229 (N_23229,N_18279,N_18476);
or U23230 (N_23230,N_18802,N_19307);
nand U23231 (N_23231,N_16084,N_19159);
nor U23232 (N_23232,N_15137,N_19863);
nor U23233 (N_23233,N_16404,N_18893);
and U23234 (N_23234,N_15655,N_15693);
nand U23235 (N_23235,N_19949,N_16967);
nand U23236 (N_23236,N_16944,N_16836);
nand U23237 (N_23237,N_19661,N_19174);
nor U23238 (N_23238,N_17178,N_16903);
nor U23239 (N_23239,N_17411,N_16874);
or U23240 (N_23240,N_16700,N_15741);
and U23241 (N_23241,N_16378,N_18097);
or U23242 (N_23242,N_15827,N_15083);
nand U23243 (N_23243,N_15945,N_18195);
nor U23244 (N_23244,N_18290,N_17821);
nor U23245 (N_23245,N_17520,N_17266);
nor U23246 (N_23246,N_17118,N_16738);
nor U23247 (N_23247,N_18025,N_16723);
or U23248 (N_23248,N_16020,N_15091);
xor U23249 (N_23249,N_17863,N_16045);
or U23250 (N_23250,N_18266,N_15406);
or U23251 (N_23251,N_19363,N_16588);
xnor U23252 (N_23252,N_18792,N_17347);
nor U23253 (N_23253,N_18526,N_19871);
nand U23254 (N_23254,N_18005,N_15676);
xnor U23255 (N_23255,N_18612,N_19171);
or U23256 (N_23256,N_16518,N_16845);
or U23257 (N_23257,N_18200,N_15007);
and U23258 (N_23258,N_19792,N_19136);
nand U23259 (N_23259,N_17945,N_19294);
and U23260 (N_23260,N_19762,N_17071);
nand U23261 (N_23261,N_18564,N_17555);
nand U23262 (N_23262,N_18675,N_16556);
or U23263 (N_23263,N_15893,N_17807);
nand U23264 (N_23264,N_15611,N_17094);
or U23265 (N_23265,N_17915,N_15102);
nand U23266 (N_23266,N_19737,N_15204);
or U23267 (N_23267,N_18038,N_16475);
nand U23268 (N_23268,N_16598,N_16578);
and U23269 (N_23269,N_15228,N_16341);
and U23270 (N_23270,N_16808,N_15418);
nor U23271 (N_23271,N_18423,N_18081);
and U23272 (N_23272,N_18830,N_15611);
xnor U23273 (N_23273,N_19293,N_18182);
and U23274 (N_23274,N_15652,N_18736);
or U23275 (N_23275,N_18014,N_15432);
nor U23276 (N_23276,N_19515,N_17999);
or U23277 (N_23277,N_19685,N_16566);
nand U23278 (N_23278,N_19581,N_19392);
nor U23279 (N_23279,N_19065,N_16721);
nor U23280 (N_23280,N_18330,N_15063);
or U23281 (N_23281,N_15090,N_18804);
and U23282 (N_23282,N_19263,N_17731);
nor U23283 (N_23283,N_18433,N_15193);
nand U23284 (N_23284,N_18537,N_18019);
xnor U23285 (N_23285,N_16622,N_15566);
nor U23286 (N_23286,N_18037,N_18800);
nor U23287 (N_23287,N_17123,N_16589);
nor U23288 (N_23288,N_18546,N_15401);
or U23289 (N_23289,N_16148,N_18087);
or U23290 (N_23290,N_15209,N_16848);
xor U23291 (N_23291,N_19014,N_17590);
and U23292 (N_23292,N_19561,N_19451);
nor U23293 (N_23293,N_18748,N_17890);
or U23294 (N_23294,N_15857,N_15081);
or U23295 (N_23295,N_19934,N_19737);
or U23296 (N_23296,N_18551,N_18293);
nand U23297 (N_23297,N_18396,N_19444);
and U23298 (N_23298,N_18956,N_15728);
nor U23299 (N_23299,N_16662,N_16646);
nand U23300 (N_23300,N_17394,N_15066);
or U23301 (N_23301,N_15295,N_18061);
or U23302 (N_23302,N_17685,N_17030);
nor U23303 (N_23303,N_16677,N_19595);
nand U23304 (N_23304,N_19987,N_16018);
and U23305 (N_23305,N_15649,N_19233);
and U23306 (N_23306,N_19489,N_17419);
nand U23307 (N_23307,N_19778,N_16930);
nand U23308 (N_23308,N_19573,N_19962);
nand U23309 (N_23309,N_15678,N_19843);
nor U23310 (N_23310,N_18070,N_15298);
and U23311 (N_23311,N_16296,N_18859);
xnor U23312 (N_23312,N_19389,N_15125);
xor U23313 (N_23313,N_15552,N_17832);
or U23314 (N_23314,N_18820,N_17514);
and U23315 (N_23315,N_17416,N_17418);
nand U23316 (N_23316,N_17849,N_17845);
or U23317 (N_23317,N_17328,N_16145);
nor U23318 (N_23318,N_18338,N_16248);
nor U23319 (N_23319,N_15717,N_15694);
or U23320 (N_23320,N_16495,N_19721);
or U23321 (N_23321,N_16437,N_17581);
and U23322 (N_23322,N_15934,N_16469);
and U23323 (N_23323,N_19833,N_16931);
nor U23324 (N_23324,N_17993,N_15959);
and U23325 (N_23325,N_19762,N_17274);
nor U23326 (N_23326,N_16223,N_15041);
nand U23327 (N_23327,N_16612,N_19438);
and U23328 (N_23328,N_15205,N_16874);
nor U23329 (N_23329,N_17751,N_15097);
nor U23330 (N_23330,N_16712,N_19916);
xor U23331 (N_23331,N_19865,N_19454);
or U23332 (N_23332,N_19458,N_19378);
or U23333 (N_23333,N_18955,N_16243);
or U23334 (N_23334,N_16680,N_16054);
nand U23335 (N_23335,N_19649,N_19183);
nand U23336 (N_23336,N_17185,N_18339);
and U23337 (N_23337,N_18765,N_17485);
nor U23338 (N_23338,N_19462,N_17033);
and U23339 (N_23339,N_19950,N_16816);
or U23340 (N_23340,N_15709,N_16804);
or U23341 (N_23341,N_17730,N_17193);
and U23342 (N_23342,N_16653,N_16960);
or U23343 (N_23343,N_15972,N_17038);
nand U23344 (N_23344,N_15837,N_16148);
and U23345 (N_23345,N_16491,N_18179);
or U23346 (N_23346,N_17018,N_19962);
nand U23347 (N_23347,N_16216,N_16138);
and U23348 (N_23348,N_18089,N_15629);
and U23349 (N_23349,N_17150,N_17749);
nand U23350 (N_23350,N_19586,N_17891);
or U23351 (N_23351,N_18788,N_19475);
and U23352 (N_23352,N_15127,N_17788);
nor U23353 (N_23353,N_16288,N_17462);
nand U23354 (N_23354,N_19479,N_17146);
or U23355 (N_23355,N_18645,N_18664);
and U23356 (N_23356,N_16485,N_16570);
nor U23357 (N_23357,N_17614,N_19751);
nor U23358 (N_23358,N_15254,N_16351);
or U23359 (N_23359,N_17762,N_18829);
nand U23360 (N_23360,N_16957,N_16669);
and U23361 (N_23361,N_19302,N_17379);
xnor U23362 (N_23362,N_19813,N_16714);
and U23363 (N_23363,N_15262,N_17354);
nor U23364 (N_23364,N_16184,N_17250);
xor U23365 (N_23365,N_19194,N_16229);
and U23366 (N_23366,N_18739,N_18524);
and U23367 (N_23367,N_15878,N_15533);
nand U23368 (N_23368,N_15909,N_16508);
nor U23369 (N_23369,N_18279,N_17695);
and U23370 (N_23370,N_16351,N_16081);
nor U23371 (N_23371,N_15780,N_17647);
nor U23372 (N_23372,N_17286,N_15842);
or U23373 (N_23373,N_19986,N_18048);
and U23374 (N_23374,N_15781,N_19422);
nor U23375 (N_23375,N_16851,N_15668);
or U23376 (N_23376,N_17743,N_15481);
nor U23377 (N_23377,N_15224,N_15046);
nand U23378 (N_23378,N_19701,N_17806);
and U23379 (N_23379,N_16081,N_19763);
nor U23380 (N_23380,N_15032,N_17958);
xor U23381 (N_23381,N_18458,N_18560);
nor U23382 (N_23382,N_15736,N_18181);
xnor U23383 (N_23383,N_16682,N_15478);
nand U23384 (N_23384,N_19356,N_16179);
and U23385 (N_23385,N_18606,N_17603);
nand U23386 (N_23386,N_19492,N_16402);
nand U23387 (N_23387,N_15006,N_18664);
nor U23388 (N_23388,N_17894,N_17953);
nand U23389 (N_23389,N_19321,N_16710);
nand U23390 (N_23390,N_19419,N_15413);
nand U23391 (N_23391,N_17882,N_16166);
xnor U23392 (N_23392,N_16779,N_17234);
and U23393 (N_23393,N_15485,N_19902);
or U23394 (N_23394,N_15629,N_19464);
or U23395 (N_23395,N_19678,N_17280);
nand U23396 (N_23396,N_16108,N_18172);
and U23397 (N_23397,N_19889,N_17857);
nand U23398 (N_23398,N_15466,N_17093);
and U23399 (N_23399,N_17743,N_15333);
nand U23400 (N_23400,N_16736,N_17206);
nor U23401 (N_23401,N_16527,N_15407);
or U23402 (N_23402,N_15544,N_17040);
nand U23403 (N_23403,N_17625,N_16033);
nor U23404 (N_23404,N_19364,N_19874);
or U23405 (N_23405,N_19471,N_16472);
and U23406 (N_23406,N_16880,N_18317);
and U23407 (N_23407,N_15463,N_18405);
nor U23408 (N_23408,N_19189,N_18076);
nand U23409 (N_23409,N_19251,N_19176);
or U23410 (N_23410,N_19862,N_18102);
nor U23411 (N_23411,N_18093,N_18789);
nand U23412 (N_23412,N_15859,N_19831);
xor U23413 (N_23413,N_16406,N_18295);
nand U23414 (N_23414,N_19716,N_18529);
or U23415 (N_23415,N_16476,N_17327);
nor U23416 (N_23416,N_16898,N_19993);
or U23417 (N_23417,N_17934,N_18870);
xnor U23418 (N_23418,N_16126,N_17592);
nor U23419 (N_23419,N_18731,N_16102);
nand U23420 (N_23420,N_16127,N_18581);
and U23421 (N_23421,N_18460,N_18644);
and U23422 (N_23422,N_17550,N_19374);
nor U23423 (N_23423,N_18630,N_19801);
nor U23424 (N_23424,N_19630,N_19326);
nand U23425 (N_23425,N_15281,N_16297);
and U23426 (N_23426,N_18967,N_15290);
and U23427 (N_23427,N_18030,N_19438);
nor U23428 (N_23428,N_16489,N_19827);
nor U23429 (N_23429,N_19046,N_15484);
and U23430 (N_23430,N_16449,N_18408);
xnor U23431 (N_23431,N_16374,N_18838);
nand U23432 (N_23432,N_17521,N_15785);
xor U23433 (N_23433,N_16443,N_15939);
nand U23434 (N_23434,N_18058,N_15104);
nand U23435 (N_23435,N_17613,N_19522);
and U23436 (N_23436,N_16628,N_15581);
nor U23437 (N_23437,N_15158,N_15786);
xor U23438 (N_23438,N_17465,N_18752);
and U23439 (N_23439,N_19222,N_19764);
and U23440 (N_23440,N_17595,N_19418);
nor U23441 (N_23441,N_17309,N_18595);
nor U23442 (N_23442,N_19530,N_15037);
nor U23443 (N_23443,N_15438,N_15989);
and U23444 (N_23444,N_17424,N_19906);
nand U23445 (N_23445,N_19468,N_18029);
or U23446 (N_23446,N_17525,N_15121);
xnor U23447 (N_23447,N_19506,N_19555);
nand U23448 (N_23448,N_15552,N_19190);
nand U23449 (N_23449,N_17691,N_18546);
nor U23450 (N_23450,N_15832,N_16275);
nor U23451 (N_23451,N_19825,N_19925);
or U23452 (N_23452,N_19316,N_16037);
nor U23453 (N_23453,N_17373,N_15236);
or U23454 (N_23454,N_16346,N_18330);
xnor U23455 (N_23455,N_18047,N_16563);
nand U23456 (N_23456,N_18599,N_17867);
or U23457 (N_23457,N_15783,N_19618);
nor U23458 (N_23458,N_18387,N_18332);
xor U23459 (N_23459,N_16816,N_18460);
or U23460 (N_23460,N_19392,N_16917);
nand U23461 (N_23461,N_16416,N_17263);
nand U23462 (N_23462,N_16561,N_19391);
and U23463 (N_23463,N_19056,N_17269);
xnor U23464 (N_23464,N_15467,N_17467);
and U23465 (N_23465,N_15190,N_15970);
nand U23466 (N_23466,N_15084,N_18520);
and U23467 (N_23467,N_16962,N_16876);
or U23468 (N_23468,N_18022,N_16732);
nor U23469 (N_23469,N_18223,N_18447);
and U23470 (N_23470,N_19786,N_18891);
nor U23471 (N_23471,N_19133,N_15593);
nand U23472 (N_23472,N_19817,N_17498);
nor U23473 (N_23473,N_18856,N_15903);
xor U23474 (N_23474,N_18905,N_16128);
nand U23475 (N_23475,N_17086,N_15061);
or U23476 (N_23476,N_15569,N_17624);
or U23477 (N_23477,N_16675,N_15863);
nor U23478 (N_23478,N_18804,N_15345);
nor U23479 (N_23479,N_15775,N_18970);
nand U23480 (N_23480,N_16772,N_18191);
xnor U23481 (N_23481,N_17469,N_19751);
nor U23482 (N_23482,N_18384,N_18634);
xor U23483 (N_23483,N_16502,N_19508);
nand U23484 (N_23484,N_18329,N_17568);
nor U23485 (N_23485,N_18240,N_19793);
and U23486 (N_23486,N_15630,N_15769);
or U23487 (N_23487,N_15711,N_17010);
nor U23488 (N_23488,N_18523,N_15537);
and U23489 (N_23489,N_16910,N_16252);
nand U23490 (N_23490,N_15383,N_16308);
and U23491 (N_23491,N_18807,N_17969);
or U23492 (N_23492,N_15932,N_16961);
and U23493 (N_23493,N_15535,N_15663);
or U23494 (N_23494,N_15088,N_17358);
nand U23495 (N_23495,N_16612,N_15854);
nor U23496 (N_23496,N_17752,N_15841);
and U23497 (N_23497,N_15977,N_16544);
nand U23498 (N_23498,N_17745,N_16104);
nand U23499 (N_23499,N_15250,N_15369);
nor U23500 (N_23500,N_18172,N_17603);
and U23501 (N_23501,N_18329,N_18228);
or U23502 (N_23502,N_17947,N_17396);
nor U23503 (N_23503,N_18637,N_18726);
and U23504 (N_23504,N_16849,N_19226);
nand U23505 (N_23505,N_17471,N_19153);
or U23506 (N_23506,N_15247,N_19463);
and U23507 (N_23507,N_15962,N_18085);
or U23508 (N_23508,N_18996,N_17505);
and U23509 (N_23509,N_19401,N_19830);
nand U23510 (N_23510,N_19783,N_18824);
nor U23511 (N_23511,N_19868,N_17583);
nor U23512 (N_23512,N_19080,N_15180);
or U23513 (N_23513,N_15208,N_16834);
nor U23514 (N_23514,N_15795,N_15875);
xor U23515 (N_23515,N_18102,N_16964);
xnor U23516 (N_23516,N_16317,N_18508);
or U23517 (N_23517,N_18981,N_15716);
and U23518 (N_23518,N_18525,N_16355);
and U23519 (N_23519,N_15958,N_17944);
or U23520 (N_23520,N_17353,N_16876);
nor U23521 (N_23521,N_18147,N_19339);
xnor U23522 (N_23522,N_17705,N_17148);
and U23523 (N_23523,N_17729,N_15289);
xnor U23524 (N_23524,N_16013,N_16054);
or U23525 (N_23525,N_16983,N_15673);
xnor U23526 (N_23526,N_16483,N_16349);
and U23527 (N_23527,N_15084,N_17048);
nand U23528 (N_23528,N_15957,N_19250);
xor U23529 (N_23529,N_17970,N_15500);
and U23530 (N_23530,N_19323,N_19342);
and U23531 (N_23531,N_19107,N_17413);
nor U23532 (N_23532,N_16398,N_18221);
and U23533 (N_23533,N_17616,N_18620);
nor U23534 (N_23534,N_19147,N_18141);
or U23535 (N_23535,N_16795,N_16721);
and U23536 (N_23536,N_19686,N_15158);
xnor U23537 (N_23537,N_16341,N_15738);
nor U23538 (N_23538,N_15276,N_17196);
nand U23539 (N_23539,N_18846,N_17151);
and U23540 (N_23540,N_16680,N_19719);
xnor U23541 (N_23541,N_18047,N_16920);
nor U23542 (N_23542,N_19267,N_17096);
nor U23543 (N_23543,N_16642,N_15708);
and U23544 (N_23544,N_16488,N_16472);
nor U23545 (N_23545,N_16098,N_15778);
or U23546 (N_23546,N_16118,N_18023);
nor U23547 (N_23547,N_19958,N_18950);
nand U23548 (N_23548,N_18123,N_18138);
and U23549 (N_23549,N_18539,N_18723);
and U23550 (N_23550,N_17505,N_16090);
or U23551 (N_23551,N_18120,N_16377);
nor U23552 (N_23552,N_15000,N_17254);
xor U23553 (N_23553,N_19019,N_18301);
nor U23554 (N_23554,N_17484,N_15384);
or U23555 (N_23555,N_17850,N_18006);
or U23556 (N_23556,N_17309,N_15917);
nor U23557 (N_23557,N_17115,N_18974);
nor U23558 (N_23558,N_17229,N_18232);
nor U23559 (N_23559,N_15253,N_17270);
nand U23560 (N_23560,N_17871,N_15370);
or U23561 (N_23561,N_19817,N_18312);
nand U23562 (N_23562,N_16272,N_15022);
and U23563 (N_23563,N_18963,N_18730);
and U23564 (N_23564,N_16085,N_19727);
or U23565 (N_23565,N_17040,N_16023);
nor U23566 (N_23566,N_17317,N_16134);
nor U23567 (N_23567,N_17241,N_15206);
and U23568 (N_23568,N_15316,N_15744);
nand U23569 (N_23569,N_16180,N_19377);
nor U23570 (N_23570,N_18355,N_18323);
or U23571 (N_23571,N_15020,N_16408);
and U23572 (N_23572,N_18453,N_19245);
nor U23573 (N_23573,N_16343,N_17867);
nor U23574 (N_23574,N_15511,N_16040);
nor U23575 (N_23575,N_16612,N_17685);
or U23576 (N_23576,N_16239,N_17168);
or U23577 (N_23577,N_19962,N_15803);
nand U23578 (N_23578,N_19700,N_16988);
and U23579 (N_23579,N_18580,N_16676);
nand U23580 (N_23580,N_17826,N_19505);
nor U23581 (N_23581,N_15196,N_16458);
or U23582 (N_23582,N_16157,N_18153);
nand U23583 (N_23583,N_17446,N_16203);
nor U23584 (N_23584,N_19633,N_15437);
nand U23585 (N_23585,N_19688,N_19401);
nor U23586 (N_23586,N_16609,N_19249);
and U23587 (N_23587,N_15324,N_16788);
xor U23588 (N_23588,N_18042,N_15082);
or U23589 (N_23589,N_16614,N_15135);
or U23590 (N_23590,N_15772,N_17467);
nor U23591 (N_23591,N_15192,N_15426);
or U23592 (N_23592,N_17537,N_18281);
nand U23593 (N_23593,N_17717,N_17136);
nor U23594 (N_23594,N_19781,N_18355);
nor U23595 (N_23595,N_17379,N_19059);
nand U23596 (N_23596,N_17796,N_16452);
or U23597 (N_23597,N_17330,N_16554);
xnor U23598 (N_23598,N_19144,N_18873);
nand U23599 (N_23599,N_18669,N_17315);
nor U23600 (N_23600,N_15222,N_16029);
and U23601 (N_23601,N_17100,N_18789);
nand U23602 (N_23602,N_19682,N_18263);
nand U23603 (N_23603,N_16567,N_18635);
or U23604 (N_23604,N_17809,N_16276);
and U23605 (N_23605,N_15107,N_19396);
nand U23606 (N_23606,N_19512,N_19407);
nand U23607 (N_23607,N_19039,N_17512);
or U23608 (N_23608,N_18177,N_19086);
nor U23609 (N_23609,N_16192,N_19295);
xnor U23610 (N_23610,N_19578,N_17416);
nand U23611 (N_23611,N_17883,N_19847);
nand U23612 (N_23612,N_17964,N_17412);
nand U23613 (N_23613,N_17090,N_16658);
xor U23614 (N_23614,N_16335,N_15407);
and U23615 (N_23615,N_18118,N_15746);
nor U23616 (N_23616,N_16065,N_18620);
nor U23617 (N_23617,N_19455,N_19734);
nand U23618 (N_23618,N_19072,N_17510);
nand U23619 (N_23619,N_19057,N_15234);
nand U23620 (N_23620,N_16574,N_15498);
nand U23621 (N_23621,N_15471,N_17575);
nor U23622 (N_23622,N_18995,N_18905);
or U23623 (N_23623,N_17041,N_15264);
or U23624 (N_23624,N_19055,N_19370);
or U23625 (N_23625,N_15374,N_16471);
or U23626 (N_23626,N_17455,N_15516);
nand U23627 (N_23627,N_16723,N_15293);
nor U23628 (N_23628,N_19671,N_19641);
nand U23629 (N_23629,N_17650,N_18376);
or U23630 (N_23630,N_17682,N_17766);
and U23631 (N_23631,N_18554,N_16619);
nor U23632 (N_23632,N_17129,N_16938);
or U23633 (N_23633,N_15708,N_16400);
and U23634 (N_23634,N_16401,N_17075);
nor U23635 (N_23635,N_16596,N_19598);
or U23636 (N_23636,N_18187,N_18032);
and U23637 (N_23637,N_18020,N_19976);
or U23638 (N_23638,N_18129,N_16948);
or U23639 (N_23639,N_15325,N_16065);
nand U23640 (N_23640,N_16273,N_17656);
xor U23641 (N_23641,N_18269,N_15519);
nor U23642 (N_23642,N_18809,N_16056);
xor U23643 (N_23643,N_16123,N_15388);
or U23644 (N_23644,N_18844,N_16292);
or U23645 (N_23645,N_18205,N_19338);
nor U23646 (N_23646,N_16163,N_18100);
or U23647 (N_23647,N_19192,N_16575);
and U23648 (N_23648,N_17071,N_18283);
nor U23649 (N_23649,N_16789,N_16017);
nor U23650 (N_23650,N_16223,N_18069);
nand U23651 (N_23651,N_16876,N_16730);
and U23652 (N_23652,N_18795,N_15414);
or U23653 (N_23653,N_16800,N_18288);
nand U23654 (N_23654,N_18679,N_17867);
nor U23655 (N_23655,N_19690,N_15491);
or U23656 (N_23656,N_17104,N_19218);
and U23657 (N_23657,N_16618,N_16716);
nor U23658 (N_23658,N_15044,N_17872);
and U23659 (N_23659,N_17817,N_19838);
and U23660 (N_23660,N_16495,N_16094);
nor U23661 (N_23661,N_18844,N_17691);
nor U23662 (N_23662,N_17340,N_18333);
or U23663 (N_23663,N_16961,N_19284);
and U23664 (N_23664,N_15734,N_16233);
nand U23665 (N_23665,N_19617,N_19818);
nor U23666 (N_23666,N_16928,N_15517);
or U23667 (N_23667,N_17292,N_16688);
and U23668 (N_23668,N_18995,N_19691);
nand U23669 (N_23669,N_16736,N_15200);
xor U23670 (N_23670,N_18845,N_16133);
and U23671 (N_23671,N_18414,N_17041);
or U23672 (N_23672,N_18053,N_15168);
nor U23673 (N_23673,N_16735,N_16640);
xnor U23674 (N_23674,N_19221,N_16146);
nand U23675 (N_23675,N_18626,N_19456);
or U23676 (N_23676,N_17824,N_17221);
xor U23677 (N_23677,N_15536,N_16084);
nand U23678 (N_23678,N_15780,N_17572);
xnor U23679 (N_23679,N_16267,N_15109);
nor U23680 (N_23680,N_18777,N_19710);
nor U23681 (N_23681,N_16750,N_19551);
or U23682 (N_23682,N_15862,N_18853);
nand U23683 (N_23683,N_19748,N_17588);
or U23684 (N_23684,N_16122,N_18847);
nor U23685 (N_23685,N_18707,N_17049);
or U23686 (N_23686,N_18762,N_17581);
or U23687 (N_23687,N_15529,N_15914);
and U23688 (N_23688,N_17672,N_19027);
xor U23689 (N_23689,N_19384,N_17466);
nor U23690 (N_23690,N_18120,N_15845);
and U23691 (N_23691,N_16151,N_16764);
nand U23692 (N_23692,N_17926,N_16847);
or U23693 (N_23693,N_16296,N_16618);
and U23694 (N_23694,N_17441,N_19832);
nand U23695 (N_23695,N_19250,N_17766);
nor U23696 (N_23696,N_15349,N_15108);
or U23697 (N_23697,N_15227,N_19350);
nor U23698 (N_23698,N_15260,N_18356);
and U23699 (N_23699,N_18088,N_16058);
nand U23700 (N_23700,N_16373,N_15347);
xor U23701 (N_23701,N_15278,N_19003);
and U23702 (N_23702,N_17213,N_16110);
or U23703 (N_23703,N_17518,N_16459);
nor U23704 (N_23704,N_15023,N_19507);
and U23705 (N_23705,N_18759,N_16507);
or U23706 (N_23706,N_18347,N_17910);
and U23707 (N_23707,N_15926,N_15869);
nand U23708 (N_23708,N_17671,N_17159);
xnor U23709 (N_23709,N_16314,N_17837);
or U23710 (N_23710,N_19776,N_15073);
xor U23711 (N_23711,N_16328,N_17320);
nor U23712 (N_23712,N_15581,N_15062);
nor U23713 (N_23713,N_15670,N_15257);
nor U23714 (N_23714,N_15654,N_16606);
and U23715 (N_23715,N_18849,N_17232);
nand U23716 (N_23716,N_15061,N_16026);
nor U23717 (N_23717,N_16787,N_15159);
nand U23718 (N_23718,N_16025,N_16401);
xnor U23719 (N_23719,N_15921,N_18046);
or U23720 (N_23720,N_18757,N_16407);
or U23721 (N_23721,N_19549,N_15008);
nor U23722 (N_23722,N_17978,N_18005);
nor U23723 (N_23723,N_19626,N_15674);
and U23724 (N_23724,N_18333,N_15694);
nor U23725 (N_23725,N_19450,N_17577);
nand U23726 (N_23726,N_15521,N_15382);
nand U23727 (N_23727,N_16366,N_19441);
or U23728 (N_23728,N_15335,N_17461);
nand U23729 (N_23729,N_17478,N_15425);
nand U23730 (N_23730,N_19236,N_18717);
xor U23731 (N_23731,N_17800,N_16177);
nand U23732 (N_23732,N_16014,N_16624);
nand U23733 (N_23733,N_15771,N_15765);
nor U23734 (N_23734,N_18796,N_17047);
xor U23735 (N_23735,N_15440,N_19799);
nor U23736 (N_23736,N_19936,N_16233);
and U23737 (N_23737,N_17646,N_19782);
nor U23738 (N_23738,N_16872,N_15494);
and U23739 (N_23739,N_16187,N_19970);
and U23740 (N_23740,N_19029,N_19972);
and U23741 (N_23741,N_19996,N_18506);
xor U23742 (N_23742,N_18325,N_17590);
or U23743 (N_23743,N_17426,N_15565);
nor U23744 (N_23744,N_16319,N_15217);
nand U23745 (N_23745,N_15508,N_15985);
nor U23746 (N_23746,N_15741,N_18237);
nor U23747 (N_23747,N_15573,N_16073);
nand U23748 (N_23748,N_18952,N_18029);
and U23749 (N_23749,N_17083,N_18767);
and U23750 (N_23750,N_18023,N_16783);
nor U23751 (N_23751,N_19717,N_19981);
nor U23752 (N_23752,N_16661,N_15875);
nand U23753 (N_23753,N_16156,N_17053);
nor U23754 (N_23754,N_15998,N_16294);
and U23755 (N_23755,N_17805,N_16588);
or U23756 (N_23756,N_19138,N_18838);
or U23757 (N_23757,N_15602,N_17282);
nand U23758 (N_23758,N_18011,N_19279);
nor U23759 (N_23759,N_19424,N_19704);
nand U23760 (N_23760,N_18437,N_17515);
and U23761 (N_23761,N_15319,N_18802);
xnor U23762 (N_23762,N_16717,N_15680);
nand U23763 (N_23763,N_16086,N_18387);
xor U23764 (N_23764,N_15124,N_18724);
and U23765 (N_23765,N_18896,N_19430);
nand U23766 (N_23766,N_18758,N_17443);
or U23767 (N_23767,N_19194,N_17772);
nand U23768 (N_23768,N_19382,N_19221);
nor U23769 (N_23769,N_17945,N_19182);
nand U23770 (N_23770,N_18480,N_16833);
nor U23771 (N_23771,N_15428,N_18382);
or U23772 (N_23772,N_17297,N_19675);
nor U23773 (N_23773,N_18166,N_18765);
nor U23774 (N_23774,N_18215,N_16677);
or U23775 (N_23775,N_17645,N_16899);
nor U23776 (N_23776,N_17770,N_16580);
and U23777 (N_23777,N_16251,N_17159);
or U23778 (N_23778,N_16265,N_16180);
nor U23779 (N_23779,N_15696,N_17335);
and U23780 (N_23780,N_19212,N_15472);
xnor U23781 (N_23781,N_17864,N_15751);
nand U23782 (N_23782,N_16430,N_17398);
and U23783 (N_23783,N_19073,N_16347);
nand U23784 (N_23784,N_17724,N_17441);
and U23785 (N_23785,N_16626,N_15785);
xor U23786 (N_23786,N_15233,N_18888);
nand U23787 (N_23787,N_18464,N_18761);
or U23788 (N_23788,N_16307,N_15254);
and U23789 (N_23789,N_18178,N_17814);
or U23790 (N_23790,N_17819,N_15493);
and U23791 (N_23791,N_18787,N_15428);
nand U23792 (N_23792,N_19586,N_19142);
nor U23793 (N_23793,N_19264,N_19486);
nand U23794 (N_23794,N_18619,N_18045);
or U23795 (N_23795,N_19240,N_15475);
or U23796 (N_23796,N_19651,N_15540);
nor U23797 (N_23797,N_16103,N_17655);
and U23798 (N_23798,N_18491,N_16851);
and U23799 (N_23799,N_16720,N_15442);
nand U23800 (N_23800,N_16742,N_15710);
nand U23801 (N_23801,N_16952,N_18250);
and U23802 (N_23802,N_16338,N_17489);
and U23803 (N_23803,N_18026,N_15110);
nand U23804 (N_23804,N_18092,N_17646);
or U23805 (N_23805,N_18067,N_18769);
or U23806 (N_23806,N_16843,N_16747);
and U23807 (N_23807,N_15450,N_19976);
nand U23808 (N_23808,N_15752,N_16493);
and U23809 (N_23809,N_19998,N_19609);
nor U23810 (N_23810,N_16549,N_19201);
or U23811 (N_23811,N_15659,N_18618);
nand U23812 (N_23812,N_18635,N_18614);
xnor U23813 (N_23813,N_15424,N_17228);
nor U23814 (N_23814,N_19913,N_17191);
nand U23815 (N_23815,N_18289,N_16773);
nand U23816 (N_23816,N_18088,N_18902);
and U23817 (N_23817,N_19227,N_15835);
nor U23818 (N_23818,N_16893,N_15922);
or U23819 (N_23819,N_15249,N_16445);
and U23820 (N_23820,N_16372,N_18038);
xor U23821 (N_23821,N_16272,N_18249);
nor U23822 (N_23822,N_18477,N_16000);
and U23823 (N_23823,N_15528,N_18055);
or U23824 (N_23824,N_18606,N_15165);
and U23825 (N_23825,N_18828,N_17574);
nand U23826 (N_23826,N_15929,N_18781);
nor U23827 (N_23827,N_19696,N_18072);
and U23828 (N_23828,N_18480,N_19958);
and U23829 (N_23829,N_15767,N_19462);
and U23830 (N_23830,N_15438,N_19845);
or U23831 (N_23831,N_16564,N_19071);
nand U23832 (N_23832,N_17896,N_17393);
nand U23833 (N_23833,N_16203,N_18112);
and U23834 (N_23834,N_16780,N_18810);
xor U23835 (N_23835,N_16170,N_16627);
nand U23836 (N_23836,N_16812,N_19249);
nand U23837 (N_23837,N_16695,N_17781);
and U23838 (N_23838,N_18750,N_16657);
and U23839 (N_23839,N_17684,N_16536);
and U23840 (N_23840,N_19551,N_18624);
and U23841 (N_23841,N_19487,N_17950);
nand U23842 (N_23842,N_17314,N_16613);
nor U23843 (N_23843,N_15889,N_15680);
and U23844 (N_23844,N_15683,N_17223);
and U23845 (N_23845,N_15182,N_15613);
or U23846 (N_23846,N_16199,N_19386);
or U23847 (N_23847,N_16671,N_17989);
nand U23848 (N_23848,N_17507,N_19465);
nand U23849 (N_23849,N_15488,N_19459);
and U23850 (N_23850,N_18457,N_16005);
and U23851 (N_23851,N_19891,N_19627);
nand U23852 (N_23852,N_18143,N_15069);
nand U23853 (N_23853,N_17156,N_16361);
nor U23854 (N_23854,N_18266,N_17134);
nor U23855 (N_23855,N_17653,N_17957);
or U23856 (N_23856,N_16235,N_16550);
xnor U23857 (N_23857,N_15443,N_15956);
and U23858 (N_23858,N_18219,N_16263);
nor U23859 (N_23859,N_16799,N_19253);
nand U23860 (N_23860,N_18569,N_19095);
nand U23861 (N_23861,N_17815,N_17027);
or U23862 (N_23862,N_19976,N_19666);
and U23863 (N_23863,N_15053,N_19028);
or U23864 (N_23864,N_18388,N_18995);
and U23865 (N_23865,N_15895,N_15078);
nor U23866 (N_23866,N_18966,N_19476);
nor U23867 (N_23867,N_18818,N_17368);
or U23868 (N_23868,N_15238,N_19985);
nand U23869 (N_23869,N_15092,N_15174);
and U23870 (N_23870,N_15156,N_18533);
nand U23871 (N_23871,N_19387,N_17699);
and U23872 (N_23872,N_15565,N_16366);
and U23873 (N_23873,N_18958,N_18521);
nand U23874 (N_23874,N_17652,N_17921);
or U23875 (N_23875,N_17962,N_18476);
or U23876 (N_23876,N_15381,N_15321);
or U23877 (N_23877,N_19986,N_19728);
nor U23878 (N_23878,N_15173,N_19146);
nor U23879 (N_23879,N_15016,N_15937);
nor U23880 (N_23880,N_17204,N_18251);
xor U23881 (N_23881,N_17909,N_19472);
nor U23882 (N_23882,N_15105,N_19244);
and U23883 (N_23883,N_16304,N_18037);
nor U23884 (N_23884,N_18708,N_16771);
nor U23885 (N_23885,N_18141,N_15168);
or U23886 (N_23886,N_18419,N_18273);
nor U23887 (N_23887,N_19499,N_16485);
or U23888 (N_23888,N_18639,N_16764);
and U23889 (N_23889,N_17702,N_16839);
nand U23890 (N_23890,N_17211,N_19986);
nor U23891 (N_23891,N_16229,N_16045);
or U23892 (N_23892,N_17976,N_19734);
nor U23893 (N_23893,N_17631,N_19597);
or U23894 (N_23894,N_17242,N_17109);
nor U23895 (N_23895,N_15374,N_18272);
nand U23896 (N_23896,N_16649,N_19847);
or U23897 (N_23897,N_17682,N_15929);
nor U23898 (N_23898,N_18715,N_19919);
nor U23899 (N_23899,N_17370,N_16548);
or U23900 (N_23900,N_16286,N_19237);
or U23901 (N_23901,N_15016,N_19470);
nor U23902 (N_23902,N_18944,N_16769);
and U23903 (N_23903,N_18374,N_16470);
or U23904 (N_23904,N_16626,N_18685);
or U23905 (N_23905,N_19936,N_18896);
nor U23906 (N_23906,N_17557,N_18682);
or U23907 (N_23907,N_15215,N_19730);
nand U23908 (N_23908,N_16411,N_19856);
and U23909 (N_23909,N_18639,N_17595);
nor U23910 (N_23910,N_18047,N_16754);
nand U23911 (N_23911,N_15669,N_16347);
and U23912 (N_23912,N_17970,N_15876);
nor U23913 (N_23913,N_16636,N_17104);
nand U23914 (N_23914,N_15412,N_16716);
nor U23915 (N_23915,N_15922,N_18559);
nor U23916 (N_23916,N_18683,N_15658);
nor U23917 (N_23917,N_17662,N_18708);
xnor U23918 (N_23918,N_19076,N_18423);
or U23919 (N_23919,N_16004,N_17125);
and U23920 (N_23920,N_15267,N_15172);
xnor U23921 (N_23921,N_18962,N_19406);
or U23922 (N_23922,N_15852,N_18298);
or U23923 (N_23923,N_16797,N_17558);
nor U23924 (N_23924,N_18770,N_19340);
xnor U23925 (N_23925,N_19733,N_19670);
and U23926 (N_23926,N_17769,N_16539);
nor U23927 (N_23927,N_16799,N_19627);
and U23928 (N_23928,N_19618,N_18402);
or U23929 (N_23929,N_18634,N_19623);
and U23930 (N_23930,N_17065,N_19766);
nor U23931 (N_23931,N_15469,N_19326);
and U23932 (N_23932,N_16836,N_16732);
and U23933 (N_23933,N_16055,N_16601);
or U23934 (N_23934,N_19442,N_18919);
and U23935 (N_23935,N_19633,N_18431);
and U23936 (N_23936,N_19440,N_17832);
and U23937 (N_23937,N_17512,N_18021);
nand U23938 (N_23938,N_17317,N_15529);
xnor U23939 (N_23939,N_15995,N_17546);
and U23940 (N_23940,N_19974,N_16550);
nand U23941 (N_23941,N_18497,N_19530);
and U23942 (N_23942,N_19095,N_15911);
and U23943 (N_23943,N_19835,N_17910);
xor U23944 (N_23944,N_15598,N_19117);
or U23945 (N_23945,N_19196,N_16045);
or U23946 (N_23946,N_17841,N_18119);
or U23947 (N_23947,N_17498,N_17137);
or U23948 (N_23948,N_19611,N_18292);
or U23949 (N_23949,N_15808,N_16608);
nand U23950 (N_23950,N_16693,N_15331);
xor U23951 (N_23951,N_16976,N_16897);
nor U23952 (N_23952,N_18280,N_16475);
nor U23953 (N_23953,N_18825,N_19854);
and U23954 (N_23954,N_18434,N_17470);
or U23955 (N_23955,N_15412,N_17310);
and U23956 (N_23956,N_16008,N_17770);
and U23957 (N_23957,N_17191,N_17084);
and U23958 (N_23958,N_18785,N_15000);
nand U23959 (N_23959,N_17469,N_18829);
and U23960 (N_23960,N_17037,N_17778);
or U23961 (N_23961,N_17311,N_18780);
nor U23962 (N_23962,N_17287,N_18231);
or U23963 (N_23963,N_16218,N_19810);
and U23964 (N_23964,N_18096,N_16213);
or U23965 (N_23965,N_16287,N_16074);
nor U23966 (N_23966,N_17213,N_16047);
and U23967 (N_23967,N_17856,N_18397);
xor U23968 (N_23968,N_19410,N_16467);
nand U23969 (N_23969,N_17253,N_15484);
nand U23970 (N_23970,N_15456,N_15659);
nor U23971 (N_23971,N_17975,N_17941);
or U23972 (N_23972,N_18902,N_18950);
nand U23973 (N_23973,N_16576,N_19623);
or U23974 (N_23974,N_18622,N_18800);
xor U23975 (N_23975,N_15181,N_19428);
nand U23976 (N_23976,N_15747,N_15663);
nand U23977 (N_23977,N_16365,N_19122);
and U23978 (N_23978,N_17528,N_17258);
nand U23979 (N_23979,N_16331,N_15297);
or U23980 (N_23980,N_19401,N_18132);
nor U23981 (N_23981,N_18494,N_17048);
nor U23982 (N_23982,N_17318,N_18400);
or U23983 (N_23983,N_17551,N_15975);
or U23984 (N_23984,N_16212,N_16997);
nand U23985 (N_23985,N_17084,N_16867);
and U23986 (N_23986,N_18085,N_15797);
xor U23987 (N_23987,N_18672,N_15485);
nand U23988 (N_23988,N_19434,N_19063);
and U23989 (N_23989,N_16189,N_17623);
or U23990 (N_23990,N_18284,N_17885);
and U23991 (N_23991,N_15433,N_16293);
or U23992 (N_23992,N_18686,N_15870);
nand U23993 (N_23993,N_18585,N_17407);
and U23994 (N_23994,N_18861,N_18710);
or U23995 (N_23995,N_15818,N_18869);
or U23996 (N_23996,N_17059,N_17713);
or U23997 (N_23997,N_16065,N_17108);
xnor U23998 (N_23998,N_16883,N_16189);
nor U23999 (N_23999,N_15138,N_16122);
nand U24000 (N_24000,N_17285,N_18533);
or U24001 (N_24001,N_15592,N_19262);
nand U24002 (N_24002,N_17391,N_18089);
and U24003 (N_24003,N_15707,N_19339);
or U24004 (N_24004,N_18142,N_18333);
or U24005 (N_24005,N_17663,N_16392);
nor U24006 (N_24006,N_18197,N_17715);
nor U24007 (N_24007,N_15988,N_18799);
nand U24008 (N_24008,N_16644,N_16380);
nand U24009 (N_24009,N_17401,N_19355);
nand U24010 (N_24010,N_19768,N_15602);
nand U24011 (N_24011,N_19559,N_16343);
and U24012 (N_24012,N_19157,N_17254);
or U24013 (N_24013,N_19588,N_19584);
nand U24014 (N_24014,N_18195,N_16073);
or U24015 (N_24015,N_18065,N_15048);
nor U24016 (N_24016,N_15126,N_19971);
xor U24017 (N_24017,N_16133,N_19372);
nor U24018 (N_24018,N_18501,N_18645);
and U24019 (N_24019,N_16142,N_16188);
and U24020 (N_24020,N_18001,N_19840);
nand U24021 (N_24021,N_18506,N_19232);
or U24022 (N_24022,N_19813,N_18213);
nand U24023 (N_24023,N_19372,N_18958);
or U24024 (N_24024,N_19095,N_17742);
and U24025 (N_24025,N_16016,N_19585);
nand U24026 (N_24026,N_18237,N_18993);
nand U24027 (N_24027,N_16276,N_15154);
and U24028 (N_24028,N_19891,N_17426);
nor U24029 (N_24029,N_15977,N_16865);
nand U24030 (N_24030,N_18104,N_16097);
or U24031 (N_24031,N_15738,N_17335);
nor U24032 (N_24032,N_15930,N_16464);
nor U24033 (N_24033,N_15456,N_16852);
and U24034 (N_24034,N_17500,N_17408);
nor U24035 (N_24035,N_16087,N_18986);
or U24036 (N_24036,N_17998,N_16387);
and U24037 (N_24037,N_16621,N_19217);
and U24038 (N_24038,N_15003,N_17475);
nand U24039 (N_24039,N_16194,N_17336);
nand U24040 (N_24040,N_17690,N_16743);
nor U24041 (N_24041,N_17554,N_17416);
or U24042 (N_24042,N_17922,N_15027);
nor U24043 (N_24043,N_18426,N_17004);
or U24044 (N_24044,N_16577,N_17258);
and U24045 (N_24045,N_19109,N_15971);
or U24046 (N_24046,N_15454,N_15184);
and U24047 (N_24047,N_16681,N_17446);
and U24048 (N_24048,N_19405,N_15934);
and U24049 (N_24049,N_15565,N_17139);
nor U24050 (N_24050,N_19411,N_18563);
nand U24051 (N_24051,N_19088,N_16313);
nor U24052 (N_24052,N_16000,N_15199);
and U24053 (N_24053,N_18255,N_16007);
nor U24054 (N_24054,N_16910,N_19237);
nand U24055 (N_24055,N_16177,N_16054);
and U24056 (N_24056,N_19646,N_18131);
and U24057 (N_24057,N_16886,N_16680);
nor U24058 (N_24058,N_19786,N_18200);
xor U24059 (N_24059,N_17413,N_17430);
or U24060 (N_24060,N_18254,N_19104);
or U24061 (N_24061,N_18293,N_18454);
and U24062 (N_24062,N_19508,N_16115);
and U24063 (N_24063,N_15632,N_16099);
nand U24064 (N_24064,N_16988,N_15606);
nand U24065 (N_24065,N_15884,N_18376);
or U24066 (N_24066,N_18911,N_15035);
xnor U24067 (N_24067,N_19760,N_19456);
nor U24068 (N_24068,N_15562,N_18670);
and U24069 (N_24069,N_17637,N_15842);
or U24070 (N_24070,N_17646,N_19775);
nand U24071 (N_24071,N_19139,N_16670);
xnor U24072 (N_24072,N_15490,N_16516);
or U24073 (N_24073,N_16847,N_15309);
nor U24074 (N_24074,N_19202,N_18724);
or U24075 (N_24075,N_17282,N_17497);
nor U24076 (N_24076,N_18604,N_16763);
nor U24077 (N_24077,N_18352,N_15547);
and U24078 (N_24078,N_16876,N_16537);
nor U24079 (N_24079,N_17877,N_15384);
and U24080 (N_24080,N_19252,N_17139);
nor U24081 (N_24081,N_19333,N_18299);
and U24082 (N_24082,N_15145,N_17370);
and U24083 (N_24083,N_19753,N_18913);
nand U24084 (N_24084,N_16210,N_18952);
and U24085 (N_24085,N_16812,N_18033);
nand U24086 (N_24086,N_16717,N_17629);
nand U24087 (N_24087,N_17318,N_19097);
nand U24088 (N_24088,N_16083,N_15350);
or U24089 (N_24089,N_18186,N_18476);
nand U24090 (N_24090,N_19812,N_17550);
or U24091 (N_24091,N_19652,N_18668);
xor U24092 (N_24092,N_15092,N_17819);
and U24093 (N_24093,N_16804,N_19273);
nor U24094 (N_24094,N_19294,N_18582);
or U24095 (N_24095,N_18747,N_15600);
or U24096 (N_24096,N_16698,N_15199);
nand U24097 (N_24097,N_15898,N_15447);
nand U24098 (N_24098,N_16862,N_18594);
nor U24099 (N_24099,N_17773,N_18260);
and U24100 (N_24100,N_17238,N_18388);
nor U24101 (N_24101,N_19192,N_15989);
nand U24102 (N_24102,N_19225,N_15225);
nor U24103 (N_24103,N_16591,N_15875);
nand U24104 (N_24104,N_15429,N_19213);
xor U24105 (N_24105,N_16237,N_18989);
nand U24106 (N_24106,N_17919,N_19002);
and U24107 (N_24107,N_17691,N_19753);
nor U24108 (N_24108,N_15352,N_15967);
nor U24109 (N_24109,N_16996,N_18059);
and U24110 (N_24110,N_16059,N_17750);
nor U24111 (N_24111,N_15245,N_15642);
and U24112 (N_24112,N_19475,N_16517);
and U24113 (N_24113,N_18987,N_16208);
and U24114 (N_24114,N_17826,N_16660);
and U24115 (N_24115,N_15417,N_15455);
nand U24116 (N_24116,N_15765,N_16613);
and U24117 (N_24117,N_16589,N_19835);
nor U24118 (N_24118,N_15155,N_18117);
nor U24119 (N_24119,N_17151,N_19337);
and U24120 (N_24120,N_18609,N_19540);
nor U24121 (N_24121,N_16145,N_15131);
nor U24122 (N_24122,N_15447,N_18170);
or U24123 (N_24123,N_17099,N_19609);
and U24124 (N_24124,N_19147,N_16103);
and U24125 (N_24125,N_18583,N_19776);
and U24126 (N_24126,N_19333,N_16852);
and U24127 (N_24127,N_19008,N_15055);
xnor U24128 (N_24128,N_17358,N_15239);
xor U24129 (N_24129,N_19958,N_18927);
nand U24130 (N_24130,N_17541,N_18636);
nand U24131 (N_24131,N_17125,N_17479);
or U24132 (N_24132,N_19849,N_15964);
and U24133 (N_24133,N_17085,N_15365);
nor U24134 (N_24134,N_15165,N_16249);
nand U24135 (N_24135,N_18324,N_19304);
and U24136 (N_24136,N_19374,N_17952);
nor U24137 (N_24137,N_18730,N_19208);
nor U24138 (N_24138,N_18032,N_15176);
or U24139 (N_24139,N_16390,N_17350);
nand U24140 (N_24140,N_19691,N_17701);
or U24141 (N_24141,N_19363,N_15645);
nor U24142 (N_24142,N_16415,N_18867);
and U24143 (N_24143,N_16356,N_19401);
nor U24144 (N_24144,N_16713,N_16727);
nand U24145 (N_24145,N_17546,N_19140);
xor U24146 (N_24146,N_16570,N_16097);
xor U24147 (N_24147,N_18426,N_17446);
and U24148 (N_24148,N_17979,N_16485);
and U24149 (N_24149,N_15162,N_19414);
xor U24150 (N_24150,N_19720,N_16750);
and U24151 (N_24151,N_18555,N_19631);
nand U24152 (N_24152,N_15206,N_19669);
nand U24153 (N_24153,N_15623,N_17018);
nor U24154 (N_24154,N_19309,N_17864);
nor U24155 (N_24155,N_16858,N_19928);
or U24156 (N_24156,N_15874,N_19501);
nor U24157 (N_24157,N_15237,N_16853);
and U24158 (N_24158,N_17056,N_15219);
nand U24159 (N_24159,N_16059,N_17796);
nand U24160 (N_24160,N_16002,N_19536);
or U24161 (N_24161,N_17373,N_18286);
and U24162 (N_24162,N_18805,N_16322);
and U24163 (N_24163,N_17929,N_15271);
xor U24164 (N_24164,N_18158,N_19963);
nand U24165 (N_24165,N_15236,N_16005);
or U24166 (N_24166,N_16665,N_16922);
nand U24167 (N_24167,N_16075,N_15790);
and U24168 (N_24168,N_19156,N_17711);
nand U24169 (N_24169,N_19744,N_15403);
and U24170 (N_24170,N_15951,N_17843);
nor U24171 (N_24171,N_17468,N_15666);
nor U24172 (N_24172,N_16051,N_19791);
and U24173 (N_24173,N_19857,N_19416);
nor U24174 (N_24174,N_16435,N_16713);
and U24175 (N_24175,N_17939,N_18967);
or U24176 (N_24176,N_16430,N_18902);
xnor U24177 (N_24177,N_19231,N_19468);
nand U24178 (N_24178,N_16901,N_15927);
nand U24179 (N_24179,N_18242,N_19826);
nor U24180 (N_24180,N_19037,N_17110);
nor U24181 (N_24181,N_15056,N_16816);
and U24182 (N_24182,N_15740,N_16307);
or U24183 (N_24183,N_18557,N_18535);
xnor U24184 (N_24184,N_19756,N_16170);
nand U24185 (N_24185,N_17793,N_17114);
or U24186 (N_24186,N_15814,N_19059);
nand U24187 (N_24187,N_18537,N_17375);
or U24188 (N_24188,N_18769,N_18790);
and U24189 (N_24189,N_15048,N_18477);
nand U24190 (N_24190,N_19544,N_16470);
nand U24191 (N_24191,N_18642,N_17820);
or U24192 (N_24192,N_15496,N_19340);
or U24193 (N_24193,N_18941,N_17505);
nor U24194 (N_24194,N_15372,N_15865);
and U24195 (N_24195,N_18967,N_16725);
nor U24196 (N_24196,N_15873,N_15441);
nand U24197 (N_24197,N_18765,N_19294);
and U24198 (N_24198,N_16675,N_17989);
nand U24199 (N_24199,N_17268,N_15386);
xor U24200 (N_24200,N_16243,N_18970);
nand U24201 (N_24201,N_19489,N_18344);
nor U24202 (N_24202,N_19790,N_17408);
or U24203 (N_24203,N_18248,N_19925);
and U24204 (N_24204,N_17101,N_19422);
xor U24205 (N_24205,N_17304,N_16495);
nor U24206 (N_24206,N_16181,N_17124);
nand U24207 (N_24207,N_15528,N_18623);
nor U24208 (N_24208,N_15499,N_15683);
nand U24209 (N_24209,N_16062,N_18979);
nor U24210 (N_24210,N_17543,N_15983);
nand U24211 (N_24211,N_17583,N_15797);
nand U24212 (N_24212,N_15053,N_16214);
and U24213 (N_24213,N_16428,N_19822);
nor U24214 (N_24214,N_17352,N_15333);
xor U24215 (N_24215,N_16907,N_19822);
nor U24216 (N_24216,N_15986,N_19512);
and U24217 (N_24217,N_19840,N_16345);
or U24218 (N_24218,N_17794,N_18695);
and U24219 (N_24219,N_17485,N_15006);
or U24220 (N_24220,N_17770,N_17771);
and U24221 (N_24221,N_15338,N_18988);
xnor U24222 (N_24222,N_18491,N_15049);
nand U24223 (N_24223,N_16816,N_16099);
nor U24224 (N_24224,N_15620,N_15690);
nor U24225 (N_24225,N_18151,N_18518);
nand U24226 (N_24226,N_19257,N_16345);
or U24227 (N_24227,N_19447,N_17145);
xor U24228 (N_24228,N_17018,N_18843);
xor U24229 (N_24229,N_18364,N_19985);
or U24230 (N_24230,N_17905,N_19225);
xor U24231 (N_24231,N_15542,N_19578);
and U24232 (N_24232,N_18256,N_18490);
xor U24233 (N_24233,N_17166,N_15974);
nand U24234 (N_24234,N_15288,N_15784);
nand U24235 (N_24235,N_15684,N_16458);
and U24236 (N_24236,N_15786,N_16581);
nor U24237 (N_24237,N_18382,N_17490);
nor U24238 (N_24238,N_15355,N_18635);
nor U24239 (N_24239,N_15942,N_19295);
and U24240 (N_24240,N_16815,N_18106);
and U24241 (N_24241,N_17736,N_15533);
nor U24242 (N_24242,N_16759,N_17235);
and U24243 (N_24243,N_17651,N_17632);
nand U24244 (N_24244,N_17341,N_18649);
nand U24245 (N_24245,N_17341,N_19885);
nand U24246 (N_24246,N_19447,N_17864);
nor U24247 (N_24247,N_19690,N_18817);
xnor U24248 (N_24248,N_16081,N_18741);
nor U24249 (N_24249,N_16043,N_15310);
nor U24250 (N_24250,N_15475,N_15101);
xnor U24251 (N_24251,N_17185,N_15921);
nor U24252 (N_24252,N_19895,N_16983);
or U24253 (N_24253,N_18444,N_19511);
nand U24254 (N_24254,N_18427,N_17578);
nor U24255 (N_24255,N_18100,N_18257);
nand U24256 (N_24256,N_17465,N_17468);
and U24257 (N_24257,N_17515,N_19503);
and U24258 (N_24258,N_15902,N_16648);
or U24259 (N_24259,N_19217,N_15158);
or U24260 (N_24260,N_19065,N_18215);
nand U24261 (N_24261,N_17905,N_17046);
and U24262 (N_24262,N_16572,N_19922);
nor U24263 (N_24263,N_15768,N_19309);
nor U24264 (N_24264,N_16801,N_19244);
nand U24265 (N_24265,N_18100,N_15944);
nand U24266 (N_24266,N_17107,N_16280);
xor U24267 (N_24267,N_16655,N_15442);
nor U24268 (N_24268,N_16860,N_17782);
and U24269 (N_24269,N_19993,N_18062);
nor U24270 (N_24270,N_17028,N_15399);
or U24271 (N_24271,N_18042,N_19100);
xnor U24272 (N_24272,N_15771,N_16447);
nor U24273 (N_24273,N_19412,N_15590);
xnor U24274 (N_24274,N_16241,N_15490);
and U24275 (N_24275,N_18464,N_19125);
nor U24276 (N_24276,N_17893,N_17871);
nand U24277 (N_24277,N_15912,N_16008);
nor U24278 (N_24278,N_17693,N_18373);
nand U24279 (N_24279,N_18328,N_17305);
nor U24280 (N_24280,N_18333,N_19333);
nand U24281 (N_24281,N_18024,N_16619);
xnor U24282 (N_24282,N_18782,N_17882);
nor U24283 (N_24283,N_17896,N_19922);
xor U24284 (N_24284,N_17940,N_16352);
nor U24285 (N_24285,N_17034,N_19033);
or U24286 (N_24286,N_19268,N_18052);
and U24287 (N_24287,N_17762,N_15262);
and U24288 (N_24288,N_17703,N_16775);
or U24289 (N_24289,N_17921,N_15671);
or U24290 (N_24290,N_18872,N_16761);
and U24291 (N_24291,N_16375,N_15210);
nand U24292 (N_24292,N_19669,N_15786);
nor U24293 (N_24293,N_18080,N_18857);
xnor U24294 (N_24294,N_17973,N_17084);
xnor U24295 (N_24295,N_16234,N_19145);
and U24296 (N_24296,N_16887,N_16789);
xnor U24297 (N_24297,N_15015,N_18555);
nand U24298 (N_24298,N_15618,N_18053);
and U24299 (N_24299,N_15413,N_16001);
and U24300 (N_24300,N_15328,N_17692);
nor U24301 (N_24301,N_15325,N_18224);
or U24302 (N_24302,N_17490,N_18537);
nand U24303 (N_24303,N_16682,N_16786);
nor U24304 (N_24304,N_19497,N_16236);
xnor U24305 (N_24305,N_15629,N_19112);
nor U24306 (N_24306,N_16056,N_17524);
or U24307 (N_24307,N_19950,N_18602);
xnor U24308 (N_24308,N_15666,N_16796);
nand U24309 (N_24309,N_18558,N_17175);
nand U24310 (N_24310,N_19702,N_19805);
and U24311 (N_24311,N_18305,N_16002);
or U24312 (N_24312,N_15321,N_19153);
nor U24313 (N_24313,N_15063,N_17884);
nand U24314 (N_24314,N_15257,N_16984);
and U24315 (N_24315,N_19342,N_15603);
nand U24316 (N_24316,N_17842,N_19605);
and U24317 (N_24317,N_17493,N_15697);
or U24318 (N_24318,N_18477,N_18156);
xnor U24319 (N_24319,N_16389,N_17577);
and U24320 (N_24320,N_17023,N_18187);
nor U24321 (N_24321,N_15299,N_15627);
and U24322 (N_24322,N_16696,N_19245);
nand U24323 (N_24323,N_17234,N_19021);
nand U24324 (N_24324,N_19911,N_16465);
or U24325 (N_24325,N_19983,N_19209);
and U24326 (N_24326,N_17801,N_18958);
or U24327 (N_24327,N_15999,N_16222);
xnor U24328 (N_24328,N_18646,N_16610);
and U24329 (N_24329,N_15025,N_18758);
or U24330 (N_24330,N_19890,N_17972);
xnor U24331 (N_24331,N_15678,N_17920);
nor U24332 (N_24332,N_16019,N_15121);
and U24333 (N_24333,N_17143,N_19327);
xnor U24334 (N_24334,N_15110,N_15572);
or U24335 (N_24335,N_18429,N_18581);
nor U24336 (N_24336,N_18732,N_19037);
nand U24337 (N_24337,N_15565,N_19669);
nand U24338 (N_24338,N_15935,N_15933);
nand U24339 (N_24339,N_18060,N_17671);
and U24340 (N_24340,N_18336,N_16641);
nand U24341 (N_24341,N_16552,N_17486);
or U24342 (N_24342,N_16540,N_16132);
nor U24343 (N_24343,N_15494,N_17134);
nor U24344 (N_24344,N_18802,N_17449);
or U24345 (N_24345,N_15921,N_16229);
or U24346 (N_24346,N_15054,N_18715);
nor U24347 (N_24347,N_16483,N_18332);
or U24348 (N_24348,N_17879,N_19661);
nor U24349 (N_24349,N_15957,N_18136);
xnor U24350 (N_24350,N_17057,N_17552);
and U24351 (N_24351,N_16973,N_17843);
xor U24352 (N_24352,N_18060,N_18065);
xnor U24353 (N_24353,N_17383,N_15109);
nand U24354 (N_24354,N_17800,N_17597);
or U24355 (N_24355,N_16037,N_18874);
or U24356 (N_24356,N_17581,N_15510);
and U24357 (N_24357,N_18127,N_18355);
nand U24358 (N_24358,N_17485,N_15963);
nor U24359 (N_24359,N_15062,N_16947);
nor U24360 (N_24360,N_19530,N_16798);
nand U24361 (N_24361,N_19705,N_19646);
and U24362 (N_24362,N_17843,N_16006);
nand U24363 (N_24363,N_19765,N_15978);
nand U24364 (N_24364,N_19453,N_17432);
and U24365 (N_24365,N_16364,N_16348);
xnor U24366 (N_24366,N_18028,N_16370);
and U24367 (N_24367,N_17295,N_17608);
xor U24368 (N_24368,N_16673,N_17397);
xnor U24369 (N_24369,N_18547,N_15289);
and U24370 (N_24370,N_16098,N_16073);
xnor U24371 (N_24371,N_15262,N_17359);
and U24372 (N_24372,N_17064,N_17988);
nand U24373 (N_24373,N_16835,N_16954);
or U24374 (N_24374,N_18961,N_17655);
and U24375 (N_24375,N_18591,N_17553);
and U24376 (N_24376,N_18685,N_17977);
nand U24377 (N_24377,N_19444,N_18149);
nor U24378 (N_24378,N_17184,N_17628);
nor U24379 (N_24379,N_17898,N_19929);
or U24380 (N_24380,N_17908,N_16077);
and U24381 (N_24381,N_17797,N_15662);
nand U24382 (N_24382,N_19766,N_16240);
nor U24383 (N_24383,N_18197,N_16228);
and U24384 (N_24384,N_15319,N_18330);
xnor U24385 (N_24385,N_15570,N_16303);
nor U24386 (N_24386,N_16511,N_19848);
or U24387 (N_24387,N_16344,N_15648);
nor U24388 (N_24388,N_16936,N_18381);
nand U24389 (N_24389,N_18468,N_16949);
and U24390 (N_24390,N_18829,N_19734);
nor U24391 (N_24391,N_17329,N_17596);
and U24392 (N_24392,N_18367,N_18536);
and U24393 (N_24393,N_17495,N_18879);
nand U24394 (N_24394,N_18923,N_18352);
nor U24395 (N_24395,N_19550,N_19393);
or U24396 (N_24396,N_16009,N_19635);
or U24397 (N_24397,N_19752,N_19988);
nand U24398 (N_24398,N_16057,N_17834);
or U24399 (N_24399,N_15614,N_18954);
and U24400 (N_24400,N_16085,N_18081);
and U24401 (N_24401,N_16681,N_16636);
and U24402 (N_24402,N_15087,N_19541);
xor U24403 (N_24403,N_18167,N_16451);
and U24404 (N_24404,N_17538,N_16402);
or U24405 (N_24405,N_18292,N_15240);
and U24406 (N_24406,N_15872,N_15276);
nor U24407 (N_24407,N_16693,N_18131);
xnor U24408 (N_24408,N_16439,N_15023);
nor U24409 (N_24409,N_15414,N_19778);
or U24410 (N_24410,N_15377,N_19042);
nand U24411 (N_24411,N_18895,N_16104);
or U24412 (N_24412,N_18743,N_19271);
or U24413 (N_24413,N_15269,N_17372);
nand U24414 (N_24414,N_17658,N_19950);
nor U24415 (N_24415,N_15049,N_16157);
xnor U24416 (N_24416,N_17041,N_17620);
and U24417 (N_24417,N_17229,N_17660);
or U24418 (N_24418,N_19723,N_16979);
nand U24419 (N_24419,N_19771,N_16230);
nand U24420 (N_24420,N_17166,N_16020);
nand U24421 (N_24421,N_16965,N_18485);
or U24422 (N_24422,N_17282,N_19942);
nor U24423 (N_24423,N_17367,N_17725);
nor U24424 (N_24424,N_17797,N_17959);
nand U24425 (N_24425,N_15047,N_15453);
nand U24426 (N_24426,N_15822,N_17682);
nor U24427 (N_24427,N_15320,N_19148);
or U24428 (N_24428,N_15700,N_15295);
xnor U24429 (N_24429,N_18595,N_15982);
or U24430 (N_24430,N_18439,N_18313);
nand U24431 (N_24431,N_16750,N_16756);
nand U24432 (N_24432,N_16206,N_16979);
and U24433 (N_24433,N_19344,N_17968);
or U24434 (N_24434,N_18250,N_19827);
nor U24435 (N_24435,N_16463,N_15111);
nor U24436 (N_24436,N_15868,N_19745);
and U24437 (N_24437,N_16377,N_15381);
nor U24438 (N_24438,N_18081,N_18898);
nand U24439 (N_24439,N_15243,N_17613);
nor U24440 (N_24440,N_15852,N_18304);
nor U24441 (N_24441,N_19863,N_16055);
xnor U24442 (N_24442,N_15893,N_15166);
and U24443 (N_24443,N_16239,N_18957);
nand U24444 (N_24444,N_15013,N_18659);
xnor U24445 (N_24445,N_16399,N_16107);
nand U24446 (N_24446,N_19433,N_16469);
nand U24447 (N_24447,N_15351,N_18109);
nor U24448 (N_24448,N_16732,N_15598);
nand U24449 (N_24449,N_16668,N_15660);
or U24450 (N_24450,N_15885,N_15318);
xnor U24451 (N_24451,N_17669,N_19148);
nor U24452 (N_24452,N_18464,N_18095);
and U24453 (N_24453,N_15007,N_16044);
and U24454 (N_24454,N_17314,N_17910);
xor U24455 (N_24455,N_16834,N_16274);
xnor U24456 (N_24456,N_19961,N_16914);
nand U24457 (N_24457,N_18272,N_16173);
nand U24458 (N_24458,N_19632,N_17254);
nor U24459 (N_24459,N_15028,N_19192);
or U24460 (N_24460,N_15113,N_19891);
xor U24461 (N_24461,N_15098,N_15731);
or U24462 (N_24462,N_19997,N_18677);
nor U24463 (N_24463,N_18937,N_18867);
xnor U24464 (N_24464,N_16037,N_18070);
nand U24465 (N_24465,N_19608,N_18534);
and U24466 (N_24466,N_19825,N_16128);
or U24467 (N_24467,N_19687,N_18244);
and U24468 (N_24468,N_17525,N_19432);
nand U24469 (N_24469,N_16904,N_15355);
and U24470 (N_24470,N_19742,N_16142);
nor U24471 (N_24471,N_18396,N_18943);
xnor U24472 (N_24472,N_15963,N_17499);
xnor U24473 (N_24473,N_15726,N_16230);
nand U24474 (N_24474,N_17556,N_18237);
and U24475 (N_24475,N_18410,N_18641);
nand U24476 (N_24476,N_19558,N_15729);
nor U24477 (N_24477,N_15534,N_17019);
nand U24478 (N_24478,N_18650,N_17467);
nand U24479 (N_24479,N_18709,N_17092);
xor U24480 (N_24480,N_15597,N_15755);
nand U24481 (N_24481,N_16395,N_17903);
or U24482 (N_24482,N_17956,N_16464);
nand U24483 (N_24483,N_15512,N_19328);
nand U24484 (N_24484,N_17615,N_18408);
nand U24485 (N_24485,N_18870,N_19436);
xnor U24486 (N_24486,N_15173,N_18828);
xnor U24487 (N_24487,N_16608,N_17174);
nand U24488 (N_24488,N_19777,N_16774);
nand U24489 (N_24489,N_19313,N_16875);
xnor U24490 (N_24490,N_17769,N_17938);
or U24491 (N_24491,N_16075,N_19598);
and U24492 (N_24492,N_18309,N_16502);
nand U24493 (N_24493,N_19570,N_19239);
or U24494 (N_24494,N_18944,N_17145);
and U24495 (N_24495,N_19580,N_15743);
or U24496 (N_24496,N_17074,N_16911);
and U24497 (N_24497,N_15888,N_15280);
nor U24498 (N_24498,N_17303,N_18840);
nand U24499 (N_24499,N_15427,N_15763);
or U24500 (N_24500,N_15918,N_19769);
and U24501 (N_24501,N_19687,N_19599);
nand U24502 (N_24502,N_15009,N_16309);
nor U24503 (N_24503,N_16281,N_16006);
nand U24504 (N_24504,N_17275,N_15187);
and U24505 (N_24505,N_18115,N_19771);
nand U24506 (N_24506,N_18194,N_19561);
nand U24507 (N_24507,N_19977,N_19662);
nand U24508 (N_24508,N_16568,N_19475);
nand U24509 (N_24509,N_15121,N_17567);
nor U24510 (N_24510,N_19261,N_17144);
nor U24511 (N_24511,N_15450,N_15610);
nand U24512 (N_24512,N_16599,N_15794);
xor U24513 (N_24513,N_15041,N_18782);
nor U24514 (N_24514,N_17740,N_17563);
xnor U24515 (N_24515,N_17032,N_16422);
xor U24516 (N_24516,N_15866,N_16442);
nor U24517 (N_24517,N_18230,N_19713);
nor U24518 (N_24518,N_15361,N_17395);
nor U24519 (N_24519,N_17451,N_15884);
and U24520 (N_24520,N_17455,N_17802);
nand U24521 (N_24521,N_19227,N_17651);
and U24522 (N_24522,N_18279,N_17855);
nor U24523 (N_24523,N_15722,N_18369);
nor U24524 (N_24524,N_19905,N_18248);
and U24525 (N_24525,N_18321,N_19449);
nor U24526 (N_24526,N_18634,N_17949);
nor U24527 (N_24527,N_15685,N_18648);
and U24528 (N_24528,N_17946,N_16713);
nand U24529 (N_24529,N_19188,N_18807);
and U24530 (N_24530,N_17209,N_19193);
or U24531 (N_24531,N_16772,N_17233);
nand U24532 (N_24532,N_18566,N_18768);
xnor U24533 (N_24533,N_15710,N_17019);
and U24534 (N_24534,N_18149,N_17438);
or U24535 (N_24535,N_15110,N_16563);
or U24536 (N_24536,N_17359,N_19818);
and U24537 (N_24537,N_16006,N_15427);
nor U24538 (N_24538,N_16424,N_15389);
nor U24539 (N_24539,N_15154,N_18709);
nor U24540 (N_24540,N_16665,N_19956);
or U24541 (N_24541,N_15443,N_19590);
nor U24542 (N_24542,N_18459,N_16265);
and U24543 (N_24543,N_17151,N_17668);
or U24544 (N_24544,N_16619,N_19364);
or U24545 (N_24545,N_19741,N_18697);
and U24546 (N_24546,N_18264,N_16582);
nand U24547 (N_24547,N_16763,N_16776);
nor U24548 (N_24548,N_16359,N_19001);
and U24549 (N_24549,N_16212,N_17615);
and U24550 (N_24550,N_15947,N_17707);
or U24551 (N_24551,N_19630,N_15993);
and U24552 (N_24552,N_18852,N_19055);
or U24553 (N_24553,N_17924,N_19905);
and U24554 (N_24554,N_16762,N_18101);
nor U24555 (N_24555,N_15359,N_16492);
or U24556 (N_24556,N_19094,N_17166);
nor U24557 (N_24557,N_16090,N_17068);
nand U24558 (N_24558,N_19234,N_16605);
xor U24559 (N_24559,N_19245,N_16380);
nor U24560 (N_24560,N_18110,N_18487);
or U24561 (N_24561,N_15223,N_18644);
xnor U24562 (N_24562,N_16220,N_18214);
or U24563 (N_24563,N_16258,N_18925);
nor U24564 (N_24564,N_18685,N_17024);
and U24565 (N_24565,N_19340,N_18007);
and U24566 (N_24566,N_18307,N_19339);
and U24567 (N_24567,N_15158,N_19957);
nand U24568 (N_24568,N_17117,N_17590);
nand U24569 (N_24569,N_18293,N_16321);
and U24570 (N_24570,N_16749,N_18883);
nor U24571 (N_24571,N_15671,N_19547);
nand U24572 (N_24572,N_15601,N_18451);
and U24573 (N_24573,N_15274,N_15587);
xor U24574 (N_24574,N_19324,N_17286);
and U24575 (N_24575,N_15277,N_15566);
and U24576 (N_24576,N_15794,N_17898);
nor U24577 (N_24577,N_17868,N_18845);
or U24578 (N_24578,N_17382,N_18373);
and U24579 (N_24579,N_17036,N_16520);
or U24580 (N_24580,N_19280,N_19636);
nand U24581 (N_24581,N_19301,N_17764);
xnor U24582 (N_24582,N_18919,N_18671);
nor U24583 (N_24583,N_17000,N_19248);
nand U24584 (N_24584,N_15998,N_16592);
nor U24585 (N_24585,N_15756,N_19790);
or U24586 (N_24586,N_17952,N_15606);
xor U24587 (N_24587,N_18768,N_19635);
and U24588 (N_24588,N_19593,N_17634);
nand U24589 (N_24589,N_17395,N_15453);
or U24590 (N_24590,N_16962,N_15456);
nor U24591 (N_24591,N_16172,N_16963);
nor U24592 (N_24592,N_18976,N_17158);
xor U24593 (N_24593,N_17094,N_15936);
and U24594 (N_24594,N_19835,N_19370);
and U24595 (N_24595,N_15500,N_15339);
nand U24596 (N_24596,N_17252,N_17314);
or U24597 (N_24597,N_18560,N_16873);
and U24598 (N_24598,N_19811,N_16815);
and U24599 (N_24599,N_17355,N_17461);
and U24600 (N_24600,N_16874,N_16216);
and U24601 (N_24601,N_18608,N_17156);
and U24602 (N_24602,N_16299,N_16437);
and U24603 (N_24603,N_19006,N_18321);
xnor U24604 (N_24604,N_15283,N_19048);
nand U24605 (N_24605,N_16415,N_16241);
nor U24606 (N_24606,N_19675,N_16471);
nor U24607 (N_24607,N_16529,N_19499);
nand U24608 (N_24608,N_17647,N_19513);
and U24609 (N_24609,N_16310,N_16164);
nand U24610 (N_24610,N_18318,N_19970);
xnor U24611 (N_24611,N_18956,N_16571);
or U24612 (N_24612,N_19071,N_17933);
or U24613 (N_24613,N_15282,N_18796);
or U24614 (N_24614,N_16497,N_17430);
and U24615 (N_24615,N_19069,N_16752);
or U24616 (N_24616,N_19046,N_17440);
xnor U24617 (N_24617,N_18574,N_18733);
xnor U24618 (N_24618,N_18076,N_18863);
and U24619 (N_24619,N_18586,N_19959);
and U24620 (N_24620,N_17138,N_19341);
or U24621 (N_24621,N_18697,N_15774);
xor U24622 (N_24622,N_16595,N_19446);
nand U24623 (N_24623,N_17623,N_15723);
or U24624 (N_24624,N_19470,N_16384);
and U24625 (N_24625,N_19806,N_16810);
and U24626 (N_24626,N_17283,N_18116);
nor U24627 (N_24627,N_19935,N_16089);
xnor U24628 (N_24628,N_17715,N_19714);
nand U24629 (N_24629,N_17417,N_15515);
and U24630 (N_24630,N_18335,N_16030);
nor U24631 (N_24631,N_16754,N_18642);
or U24632 (N_24632,N_18530,N_15179);
and U24633 (N_24633,N_15069,N_19586);
nand U24634 (N_24634,N_19247,N_16713);
nand U24635 (N_24635,N_16830,N_19219);
and U24636 (N_24636,N_19085,N_16565);
nand U24637 (N_24637,N_19652,N_19058);
nand U24638 (N_24638,N_16034,N_17026);
and U24639 (N_24639,N_19487,N_18645);
or U24640 (N_24640,N_19730,N_18980);
or U24641 (N_24641,N_15310,N_19512);
nor U24642 (N_24642,N_17340,N_16100);
xor U24643 (N_24643,N_16376,N_19133);
or U24644 (N_24644,N_15225,N_17381);
or U24645 (N_24645,N_16683,N_18759);
nand U24646 (N_24646,N_17590,N_17973);
or U24647 (N_24647,N_18735,N_17222);
nor U24648 (N_24648,N_16524,N_16064);
or U24649 (N_24649,N_18167,N_15763);
xnor U24650 (N_24650,N_18420,N_19968);
xor U24651 (N_24651,N_18713,N_16932);
nand U24652 (N_24652,N_18239,N_16926);
nand U24653 (N_24653,N_17999,N_18715);
and U24654 (N_24654,N_18366,N_15424);
or U24655 (N_24655,N_18494,N_16112);
or U24656 (N_24656,N_18197,N_17844);
or U24657 (N_24657,N_17813,N_19645);
nand U24658 (N_24658,N_18411,N_17038);
and U24659 (N_24659,N_19904,N_16527);
nand U24660 (N_24660,N_15544,N_18181);
nand U24661 (N_24661,N_16924,N_15043);
nand U24662 (N_24662,N_19631,N_18956);
or U24663 (N_24663,N_16197,N_15798);
nand U24664 (N_24664,N_19843,N_19764);
or U24665 (N_24665,N_17526,N_15791);
and U24666 (N_24666,N_17647,N_16126);
nor U24667 (N_24667,N_19213,N_18595);
or U24668 (N_24668,N_16173,N_16091);
or U24669 (N_24669,N_15208,N_17586);
or U24670 (N_24670,N_19608,N_15479);
nand U24671 (N_24671,N_17365,N_16246);
nor U24672 (N_24672,N_19985,N_16919);
and U24673 (N_24673,N_18262,N_17456);
nor U24674 (N_24674,N_18950,N_17868);
or U24675 (N_24675,N_18768,N_17305);
nand U24676 (N_24676,N_16611,N_16739);
nor U24677 (N_24677,N_16593,N_19759);
or U24678 (N_24678,N_18923,N_19003);
nor U24679 (N_24679,N_16352,N_19829);
nor U24680 (N_24680,N_19238,N_15891);
and U24681 (N_24681,N_17853,N_15979);
or U24682 (N_24682,N_15586,N_19844);
xor U24683 (N_24683,N_15274,N_17264);
nor U24684 (N_24684,N_19849,N_15989);
nor U24685 (N_24685,N_17128,N_19621);
or U24686 (N_24686,N_15560,N_16723);
nand U24687 (N_24687,N_16069,N_16432);
nor U24688 (N_24688,N_16276,N_18594);
or U24689 (N_24689,N_19184,N_19085);
or U24690 (N_24690,N_18957,N_17373);
or U24691 (N_24691,N_17358,N_18366);
or U24692 (N_24692,N_16317,N_15956);
nand U24693 (N_24693,N_18350,N_15802);
nand U24694 (N_24694,N_18704,N_18641);
or U24695 (N_24695,N_19376,N_16569);
nand U24696 (N_24696,N_15218,N_16469);
and U24697 (N_24697,N_16642,N_19223);
xor U24698 (N_24698,N_15714,N_17509);
nand U24699 (N_24699,N_18347,N_16485);
and U24700 (N_24700,N_15344,N_19185);
or U24701 (N_24701,N_16219,N_16107);
or U24702 (N_24702,N_17739,N_19989);
and U24703 (N_24703,N_15496,N_19188);
nor U24704 (N_24704,N_19022,N_17120);
or U24705 (N_24705,N_16869,N_18648);
or U24706 (N_24706,N_16747,N_15523);
or U24707 (N_24707,N_16913,N_18060);
and U24708 (N_24708,N_16725,N_15541);
and U24709 (N_24709,N_15816,N_15698);
and U24710 (N_24710,N_16024,N_15532);
nand U24711 (N_24711,N_16609,N_15280);
or U24712 (N_24712,N_19199,N_16515);
nor U24713 (N_24713,N_17945,N_15996);
and U24714 (N_24714,N_17052,N_18722);
or U24715 (N_24715,N_15260,N_18646);
and U24716 (N_24716,N_19117,N_15830);
nand U24717 (N_24717,N_16357,N_16685);
and U24718 (N_24718,N_17962,N_18886);
or U24719 (N_24719,N_15214,N_17669);
nor U24720 (N_24720,N_19470,N_17037);
xnor U24721 (N_24721,N_18251,N_16260);
xnor U24722 (N_24722,N_17301,N_15893);
xor U24723 (N_24723,N_17386,N_15376);
nand U24724 (N_24724,N_18371,N_19572);
xor U24725 (N_24725,N_17755,N_16462);
nor U24726 (N_24726,N_16463,N_19108);
nor U24727 (N_24727,N_19353,N_18273);
xor U24728 (N_24728,N_15625,N_16002);
nand U24729 (N_24729,N_15819,N_18412);
nor U24730 (N_24730,N_15821,N_16376);
or U24731 (N_24731,N_15177,N_18735);
nand U24732 (N_24732,N_17638,N_16046);
nand U24733 (N_24733,N_18649,N_19429);
and U24734 (N_24734,N_16803,N_16550);
nor U24735 (N_24735,N_17210,N_18773);
or U24736 (N_24736,N_16874,N_18605);
or U24737 (N_24737,N_18319,N_16569);
or U24738 (N_24738,N_17183,N_19897);
xnor U24739 (N_24739,N_17767,N_15761);
xor U24740 (N_24740,N_18156,N_19440);
nor U24741 (N_24741,N_18556,N_18654);
nand U24742 (N_24742,N_17453,N_15690);
and U24743 (N_24743,N_18995,N_15452);
xnor U24744 (N_24744,N_17956,N_17998);
nand U24745 (N_24745,N_17610,N_18566);
nand U24746 (N_24746,N_18967,N_18735);
nand U24747 (N_24747,N_18383,N_15084);
and U24748 (N_24748,N_16844,N_15191);
and U24749 (N_24749,N_19888,N_17053);
or U24750 (N_24750,N_18208,N_16374);
or U24751 (N_24751,N_15404,N_19361);
or U24752 (N_24752,N_17358,N_18425);
or U24753 (N_24753,N_15624,N_15879);
nor U24754 (N_24754,N_18773,N_18530);
nor U24755 (N_24755,N_15960,N_18723);
or U24756 (N_24756,N_19410,N_17444);
xor U24757 (N_24757,N_18789,N_16929);
nor U24758 (N_24758,N_18742,N_17518);
and U24759 (N_24759,N_19718,N_15686);
xor U24760 (N_24760,N_19550,N_17511);
or U24761 (N_24761,N_17185,N_18885);
or U24762 (N_24762,N_16732,N_18104);
nor U24763 (N_24763,N_19816,N_18703);
or U24764 (N_24764,N_17741,N_15639);
nor U24765 (N_24765,N_16923,N_19003);
nand U24766 (N_24766,N_15292,N_19834);
nor U24767 (N_24767,N_17728,N_18645);
xor U24768 (N_24768,N_18514,N_15416);
nand U24769 (N_24769,N_15067,N_15066);
nor U24770 (N_24770,N_16295,N_15220);
or U24771 (N_24771,N_19380,N_18879);
nor U24772 (N_24772,N_17574,N_18279);
and U24773 (N_24773,N_18568,N_18353);
nor U24774 (N_24774,N_18541,N_16973);
or U24775 (N_24775,N_17325,N_19413);
and U24776 (N_24776,N_17616,N_17995);
or U24777 (N_24777,N_15329,N_19635);
xor U24778 (N_24778,N_17629,N_15895);
nor U24779 (N_24779,N_17571,N_19562);
nand U24780 (N_24780,N_15994,N_15371);
nand U24781 (N_24781,N_17562,N_17540);
xnor U24782 (N_24782,N_17184,N_19172);
xor U24783 (N_24783,N_18195,N_17469);
nand U24784 (N_24784,N_18162,N_19008);
nand U24785 (N_24785,N_19817,N_15506);
and U24786 (N_24786,N_15793,N_17575);
nor U24787 (N_24787,N_19707,N_16604);
xor U24788 (N_24788,N_18957,N_17328);
nand U24789 (N_24789,N_15055,N_17587);
nand U24790 (N_24790,N_19022,N_19739);
nor U24791 (N_24791,N_15005,N_16883);
or U24792 (N_24792,N_16346,N_15544);
and U24793 (N_24793,N_16188,N_15711);
nor U24794 (N_24794,N_15379,N_18837);
nand U24795 (N_24795,N_17362,N_18367);
and U24796 (N_24796,N_19563,N_16431);
nor U24797 (N_24797,N_15374,N_15249);
nand U24798 (N_24798,N_16599,N_15436);
nor U24799 (N_24799,N_16803,N_18647);
and U24800 (N_24800,N_15113,N_17679);
nand U24801 (N_24801,N_19447,N_15375);
xor U24802 (N_24802,N_15782,N_18520);
nand U24803 (N_24803,N_19103,N_16581);
and U24804 (N_24804,N_18071,N_19972);
xnor U24805 (N_24805,N_16532,N_18779);
xor U24806 (N_24806,N_19213,N_15556);
and U24807 (N_24807,N_16668,N_16126);
or U24808 (N_24808,N_17431,N_18738);
or U24809 (N_24809,N_19577,N_15950);
nor U24810 (N_24810,N_17974,N_16219);
and U24811 (N_24811,N_18289,N_19727);
nand U24812 (N_24812,N_17397,N_15767);
nand U24813 (N_24813,N_15180,N_17443);
and U24814 (N_24814,N_17253,N_18330);
nor U24815 (N_24815,N_17896,N_16537);
nor U24816 (N_24816,N_19517,N_17498);
nor U24817 (N_24817,N_18211,N_16596);
nor U24818 (N_24818,N_15626,N_15653);
nor U24819 (N_24819,N_19694,N_18880);
nor U24820 (N_24820,N_18586,N_17929);
and U24821 (N_24821,N_19250,N_15938);
or U24822 (N_24822,N_19788,N_19727);
xor U24823 (N_24823,N_17711,N_15104);
or U24824 (N_24824,N_15177,N_19216);
and U24825 (N_24825,N_15337,N_18186);
xnor U24826 (N_24826,N_17315,N_15199);
nor U24827 (N_24827,N_15325,N_16147);
nand U24828 (N_24828,N_18169,N_17999);
nand U24829 (N_24829,N_15932,N_18746);
nand U24830 (N_24830,N_19350,N_17656);
nor U24831 (N_24831,N_16985,N_18520);
xnor U24832 (N_24832,N_17312,N_16877);
nor U24833 (N_24833,N_18593,N_16150);
and U24834 (N_24834,N_18023,N_16585);
nor U24835 (N_24835,N_18962,N_16244);
nor U24836 (N_24836,N_16689,N_18193);
or U24837 (N_24837,N_16351,N_18255);
and U24838 (N_24838,N_19792,N_15695);
and U24839 (N_24839,N_15512,N_16245);
nor U24840 (N_24840,N_18770,N_15753);
nand U24841 (N_24841,N_17463,N_17582);
nand U24842 (N_24842,N_17694,N_15633);
nand U24843 (N_24843,N_17909,N_17939);
nor U24844 (N_24844,N_17373,N_19607);
and U24845 (N_24845,N_15742,N_18962);
xnor U24846 (N_24846,N_19537,N_15893);
and U24847 (N_24847,N_18602,N_18448);
xor U24848 (N_24848,N_18106,N_18878);
nand U24849 (N_24849,N_15343,N_19519);
nand U24850 (N_24850,N_16915,N_17644);
nand U24851 (N_24851,N_19052,N_17061);
and U24852 (N_24852,N_15354,N_15248);
nor U24853 (N_24853,N_15504,N_16285);
nor U24854 (N_24854,N_18024,N_17445);
nand U24855 (N_24855,N_18452,N_17349);
nand U24856 (N_24856,N_19823,N_16120);
or U24857 (N_24857,N_15451,N_16795);
nand U24858 (N_24858,N_19124,N_18419);
and U24859 (N_24859,N_19664,N_19948);
xor U24860 (N_24860,N_17844,N_19592);
xor U24861 (N_24861,N_19563,N_15468);
or U24862 (N_24862,N_18385,N_18518);
and U24863 (N_24863,N_17342,N_19123);
xnor U24864 (N_24864,N_18163,N_15269);
and U24865 (N_24865,N_17712,N_17964);
xnor U24866 (N_24866,N_17108,N_19308);
nor U24867 (N_24867,N_16736,N_17073);
nor U24868 (N_24868,N_15963,N_15634);
or U24869 (N_24869,N_19758,N_19222);
nand U24870 (N_24870,N_18369,N_17903);
nor U24871 (N_24871,N_15606,N_17201);
nor U24872 (N_24872,N_18777,N_17160);
or U24873 (N_24873,N_15147,N_18260);
or U24874 (N_24874,N_17908,N_16378);
nor U24875 (N_24875,N_17965,N_16155);
nor U24876 (N_24876,N_16649,N_18200);
and U24877 (N_24877,N_17573,N_15706);
xnor U24878 (N_24878,N_18937,N_17987);
or U24879 (N_24879,N_16731,N_16826);
or U24880 (N_24880,N_19194,N_18611);
and U24881 (N_24881,N_16553,N_17131);
or U24882 (N_24882,N_17625,N_16114);
xnor U24883 (N_24883,N_17656,N_17926);
or U24884 (N_24884,N_19783,N_15858);
and U24885 (N_24885,N_17403,N_16642);
and U24886 (N_24886,N_18015,N_17569);
nand U24887 (N_24887,N_19128,N_17414);
xor U24888 (N_24888,N_17740,N_19447);
and U24889 (N_24889,N_16281,N_18116);
nor U24890 (N_24890,N_19242,N_15300);
nor U24891 (N_24891,N_16232,N_18434);
and U24892 (N_24892,N_16674,N_16554);
nor U24893 (N_24893,N_19842,N_17804);
nand U24894 (N_24894,N_19232,N_15276);
nor U24895 (N_24895,N_16349,N_15993);
nand U24896 (N_24896,N_15760,N_17200);
nor U24897 (N_24897,N_15787,N_15559);
and U24898 (N_24898,N_17642,N_19519);
or U24899 (N_24899,N_19619,N_17899);
xnor U24900 (N_24900,N_18572,N_19194);
nand U24901 (N_24901,N_17890,N_17906);
and U24902 (N_24902,N_19046,N_17460);
nand U24903 (N_24903,N_18062,N_18711);
nand U24904 (N_24904,N_16465,N_16702);
nor U24905 (N_24905,N_19047,N_16626);
or U24906 (N_24906,N_17381,N_18541);
or U24907 (N_24907,N_16938,N_17819);
xnor U24908 (N_24908,N_18735,N_15599);
or U24909 (N_24909,N_16241,N_17979);
or U24910 (N_24910,N_19267,N_17883);
nand U24911 (N_24911,N_16938,N_18740);
or U24912 (N_24912,N_17652,N_16923);
and U24913 (N_24913,N_17947,N_16490);
or U24914 (N_24914,N_18872,N_18657);
and U24915 (N_24915,N_15966,N_17771);
or U24916 (N_24916,N_16759,N_15163);
or U24917 (N_24917,N_19786,N_19332);
nor U24918 (N_24918,N_19095,N_16127);
nand U24919 (N_24919,N_16204,N_18793);
nor U24920 (N_24920,N_15034,N_16511);
or U24921 (N_24921,N_15351,N_17173);
and U24922 (N_24922,N_17977,N_17567);
and U24923 (N_24923,N_15956,N_19922);
nor U24924 (N_24924,N_17504,N_19599);
nand U24925 (N_24925,N_16131,N_16779);
nor U24926 (N_24926,N_16611,N_15482);
nor U24927 (N_24927,N_19970,N_15516);
and U24928 (N_24928,N_18987,N_15275);
or U24929 (N_24929,N_18161,N_17193);
nor U24930 (N_24930,N_16309,N_16086);
xnor U24931 (N_24931,N_17279,N_16902);
and U24932 (N_24932,N_16550,N_16675);
nand U24933 (N_24933,N_17586,N_19381);
nor U24934 (N_24934,N_17435,N_15950);
nand U24935 (N_24935,N_17610,N_16150);
xnor U24936 (N_24936,N_17535,N_19678);
or U24937 (N_24937,N_16798,N_19862);
or U24938 (N_24938,N_15031,N_18223);
nand U24939 (N_24939,N_15146,N_16679);
or U24940 (N_24940,N_16555,N_16812);
and U24941 (N_24941,N_16191,N_19351);
xor U24942 (N_24942,N_15615,N_17735);
and U24943 (N_24943,N_19002,N_17647);
nand U24944 (N_24944,N_15159,N_15248);
and U24945 (N_24945,N_17663,N_18796);
nand U24946 (N_24946,N_17858,N_16395);
nor U24947 (N_24947,N_17803,N_17907);
and U24948 (N_24948,N_16410,N_17293);
or U24949 (N_24949,N_16683,N_18656);
nand U24950 (N_24950,N_18216,N_17874);
or U24951 (N_24951,N_16917,N_19505);
or U24952 (N_24952,N_17912,N_15535);
nor U24953 (N_24953,N_16171,N_19644);
nor U24954 (N_24954,N_15178,N_17476);
nor U24955 (N_24955,N_17565,N_15307);
nand U24956 (N_24956,N_19880,N_18263);
and U24957 (N_24957,N_17688,N_19475);
or U24958 (N_24958,N_17318,N_18908);
and U24959 (N_24959,N_16472,N_15338);
or U24960 (N_24960,N_16003,N_18882);
nand U24961 (N_24961,N_16171,N_19807);
and U24962 (N_24962,N_17201,N_15127);
xnor U24963 (N_24963,N_15091,N_16751);
nand U24964 (N_24964,N_19080,N_16186);
or U24965 (N_24965,N_16296,N_17358);
or U24966 (N_24966,N_18906,N_19674);
nand U24967 (N_24967,N_16510,N_16242);
and U24968 (N_24968,N_16086,N_16060);
or U24969 (N_24969,N_17082,N_18659);
or U24970 (N_24970,N_16117,N_15482);
nand U24971 (N_24971,N_17420,N_18577);
xnor U24972 (N_24972,N_15174,N_15128);
nand U24973 (N_24973,N_19107,N_19040);
or U24974 (N_24974,N_16028,N_18911);
nand U24975 (N_24975,N_17607,N_15762);
nand U24976 (N_24976,N_18650,N_19805);
nor U24977 (N_24977,N_18487,N_16411);
nand U24978 (N_24978,N_18323,N_15693);
nor U24979 (N_24979,N_15836,N_17180);
nor U24980 (N_24980,N_16304,N_15563);
nor U24981 (N_24981,N_15286,N_17667);
and U24982 (N_24982,N_17350,N_16253);
or U24983 (N_24983,N_16076,N_17831);
or U24984 (N_24984,N_15027,N_17147);
and U24985 (N_24985,N_15200,N_19625);
nor U24986 (N_24986,N_16399,N_16159);
nor U24987 (N_24987,N_19358,N_19655);
nor U24988 (N_24988,N_18497,N_17233);
nor U24989 (N_24989,N_15682,N_16635);
xor U24990 (N_24990,N_17559,N_17437);
nand U24991 (N_24991,N_16128,N_19750);
and U24992 (N_24992,N_15179,N_19312);
and U24993 (N_24993,N_15280,N_18519);
and U24994 (N_24994,N_15598,N_15994);
or U24995 (N_24995,N_19951,N_15777);
or U24996 (N_24996,N_18070,N_18600);
nor U24997 (N_24997,N_15541,N_15760);
xor U24998 (N_24998,N_17402,N_15210);
xnor U24999 (N_24999,N_15934,N_16965);
nand UO_0 (O_0,N_20522,N_21483);
nand UO_1 (O_1,N_22627,N_21414);
and UO_2 (O_2,N_21653,N_21530);
nor UO_3 (O_3,N_22560,N_21950);
and UO_4 (O_4,N_24938,N_24781);
nand UO_5 (O_5,N_24968,N_22740);
xnor UO_6 (O_6,N_21843,N_22655);
and UO_7 (O_7,N_20790,N_24143);
nor UO_8 (O_8,N_22205,N_24793);
xnor UO_9 (O_9,N_20145,N_24128);
nor UO_10 (O_10,N_22815,N_20953);
or UO_11 (O_11,N_22487,N_20343);
and UO_12 (O_12,N_23400,N_22499);
and UO_13 (O_13,N_21507,N_21499);
and UO_14 (O_14,N_22300,N_22794);
or UO_15 (O_15,N_23949,N_22165);
or UO_16 (O_16,N_21973,N_23722);
and UO_17 (O_17,N_21013,N_24660);
and UO_18 (O_18,N_24116,N_22647);
nand UO_19 (O_19,N_20869,N_24338);
xnor UO_20 (O_20,N_23300,N_22515);
or UO_21 (O_21,N_24518,N_24697);
and UO_22 (O_22,N_22877,N_24676);
or UO_23 (O_23,N_20765,N_21330);
nand UO_24 (O_24,N_23701,N_24839);
nand UO_25 (O_25,N_22532,N_22833);
or UO_26 (O_26,N_22672,N_24211);
nand UO_27 (O_27,N_20569,N_21787);
nor UO_28 (O_28,N_23755,N_21737);
or UO_29 (O_29,N_24466,N_20695);
and UO_30 (O_30,N_23769,N_24224);
nor UO_31 (O_31,N_22936,N_23839);
and UO_32 (O_32,N_20101,N_23225);
or UO_33 (O_33,N_20546,N_23856);
or UO_34 (O_34,N_22894,N_23972);
or UO_35 (O_35,N_22268,N_24366);
nor UO_36 (O_36,N_23335,N_21022);
nand UO_37 (O_37,N_20148,N_24959);
nor UO_38 (O_38,N_21021,N_20608);
and UO_39 (O_39,N_20453,N_23396);
nor UO_40 (O_40,N_20254,N_24769);
or UO_41 (O_41,N_22652,N_21888);
nand UO_42 (O_42,N_24708,N_23634);
nor UO_43 (O_43,N_24980,N_21529);
nor UO_44 (O_44,N_21638,N_21001);
and UO_45 (O_45,N_22344,N_20019);
and UO_46 (O_46,N_21923,N_20472);
or UO_47 (O_47,N_22198,N_20393);
nand UO_48 (O_48,N_22736,N_23236);
or UO_49 (O_49,N_24017,N_20700);
nor UO_50 (O_50,N_20165,N_21581);
or UO_51 (O_51,N_20055,N_20693);
nand UO_52 (O_52,N_22237,N_24014);
nand UO_53 (O_53,N_20243,N_20473);
and UO_54 (O_54,N_21919,N_20029);
nand UO_55 (O_55,N_23776,N_23840);
or UO_56 (O_56,N_20734,N_20830);
and UO_57 (O_57,N_23510,N_22209);
and UO_58 (O_58,N_20759,N_21434);
or UO_59 (O_59,N_21803,N_22428);
or UO_60 (O_60,N_24249,N_21027);
nand UO_61 (O_61,N_23153,N_21221);
nor UO_62 (O_62,N_23950,N_23518);
nand UO_63 (O_63,N_22839,N_23637);
nor UO_64 (O_64,N_24208,N_20496);
nand UO_65 (O_65,N_21750,N_20806);
and UO_66 (O_66,N_22178,N_21819);
and UO_67 (O_67,N_21298,N_24653);
or UO_68 (O_68,N_20978,N_22531);
xor UO_69 (O_69,N_23617,N_20143);
nor UO_70 (O_70,N_23790,N_24489);
or UO_71 (O_71,N_24301,N_21608);
nor UO_72 (O_72,N_21952,N_23157);
nor UO_73 (O_73,N_20949,N_22097);
and UO_74 (O_74,N_23198,N_23527);
nand UO_75 (O_75,N_22996,N_20838);
or UO_76 (O_76,N_21303,N_24022);
nor UO_77 (O_77,N_23758,N_22854);
nand UO_78 (O_78,N_20528,N_23257);
and UO_79 (O_79,N_20797,N_22153);
nand UO_80 (O_80,N_20282,N_23878);
nor UO_81 (O_81,N_20667,N_22417);
nor UO_82 (O_82,N_22523,N_22761);
and UO_83 (O_83,N_20469,N_23872);
nand UO_84 (O_84,N_24108,N_23679);
or UO_85 (O_85,N_24929,N_22002);
nand UO_86 (O_86,N_20323,N_24855);
xnor UO_87 (O_87,N_20685,N_21484);
and UO_88 (O_88,N_23908,N_21325);
nand UO_89 (O_89,N_20722,N_22992);
or UO_90 (O_90,N_23485,N_21120);
nor UO_91 (O_91,N_24246,N_21830);
and UO_92 (O_92,N_23359,N_24503);
nor UO_93 (O_93,N_22867,N_24065);
and UO_94 (O_94,N_20435,N_20204);
and UO_95 (O_95,N_23708,N_22353);
xor UO_96 (O_96,N_24187,N_24551);
xnor UO_97 (O_97,N_22860,N_24537);
nand UO_98 (O_98,N_23942,N_22910);
or UO_99 (O_99,N_23754,N_24274);
nand UO_100 (O_100,N_24012,N_22974);
or UO_101 (O_101,N_22154,N_20411);
or UO_102 (O_102,N_22017,N_22924);
and UO_103 (O_103,N_24226,N_21450);
or UO_104 (O_104,N_23718,N_20699);
and UO_105 (O_105,N_23853,N_24302);
nor UO_106 (O_106,N_22375,N_23526);
nor UO_107 (O_107,N_20820,N_24740);
and UO_108 (O_108,N_22470,N_24142);
nand UO_109 (O_109,N_22073,N_20286);
nor UO_110 (O_110,N_24252,N_21665);
and UO_111 (O_111,N_21902,N_21311);
and UO_112 (O_112,N_21086,N_20844);
nor UO_113 (O_113,N_22517,N_21616);
nor UO_114 (O_114,N_22873,N_23602);
or UO_115 (O_115,N_24771,N_21805);
nand UO_116 (O_116,N_21575,N_20371);
xnor UO_117 (O_117,N_20552,N_20471);
and UO_118 (O_118,N_23809,N_23166);
and UO_119 (O_119,N_24764,N_20919);
nand UO_120 (O_120,N_21399,N_21542);
nand UO_121 (O_121,N_24655,N_23847);
nor UO_122 (O_122,N_21710,N_21743);
or UO_123 (O_123,N_24276,N_24273);
and UO_124 (O_124,N_23104,N_20913);
nand UO_125 (O_125,N_20764,N_21079);
or UO_126 (O_126,N_24574,N_23158);
and UO_127 (O_127,N_23301,N_23065);
xnor UO_128 (O_128,N_23906,N_22612);
and UO_129 (O_129,N_21730,N_24225);
nor UO_130 (O_130,N_20719,N_22654);
or UO_131 (O_131,N_24088,N_20184);
or UO_132 (O_132,N_23751,N_24385);
or UO_133 (O_133,N_24259,N_22574);
nor UO_134 (O_134,N_21202,N_24178);
xnor UO_135 (O_135,N_20752,N_22305);
or UO_136 (O_136,N_21361,N_22342);
and UO_137 (O_137,N_22835,N_24056);
nor UO_138 (O_138,N_24801,N_21392);
or UO_139 (O_139,N_20175,N_23226);
nand UO_140 (O_140,N_23658,N_24719);
and UO_141 (O_141,N_22535,N_22657);
nor UO_142 (O_142,N_21479,N_21849);
or UO_143 (O_143,N_23688,N_22174);
nand UO_144 (O_144,N_20180,N_24287);
or UO_145 (O_145,N_22335,N_20996);
xor UO_146 (O_146,N_23870,N_23343);
nor UO_147 (O_147,N_20432,N_24707);
xor UO_148 (O_148,N_22730,N_20982);
and UO_149 (O_149,N_22203,N_23959);
nor UO_150 (O_150,N_22128,N_20155);
or UO_151 (O_151,N_24222,N_21807);
xor UO_152 (O_152,N_22516,N_21428);
nor UO_153 (O_153,N_22099,N_23345);
and UO_154 (O_154,N_23793,N_24020);
nor UO_155 (O_155,N_24309,N_23092);
and UO_156 (O_156,N_23168,N_21077);
nand UO_157 (O_157,N_20075,N_22727);
nand UO_158 (O_158,N_21989,N_24910);
nand UO_159 (O_159,N_22893,N_21199);
nor UO_160 (O_160,N_23712,N_21795);
nor UO_161 (O_161,N_20167,N_23183);
nand UO_162 (O_162,N_20004,N_20022);
nand UO_163 (O_163,N_21613,N_20439);
and UO_164 (O_164,N_23001,N_23938);
nand UO_165 (O_165,N_21661,N_22343);
or UO_166 (O_166,N_22226,N_23971);
nand UO_167 (O_167,N_24031,N_24347);
or UO_168 (O_168,N_20348,N_21786);
nor UO_169 (O_169,N_24615,N_24529);
and UO_170 (O_170,N_23741,N_21322);
or UO_171 (O_171,N_21078,N_20142);
xor UO_172 (O_172,N_23072,N_21826);
nand UO_173 (O_173,N_24922,N_24755);
nand UO_174 (O_174,N_24841,N_24444);
nor UO_175 (O_175,N_20925,N_20599);
or UO_176 (O_176,N_22912,N_23902);
nor UO_177 (O_177,N_23451,N_24716);
xnor UO_178 (O_178,N_20841,N_24944);
and UO_179 (O_179,N_23728,N_24344);
nor UO_180 (O_180,N_22699,N_22483);
xnor UO_181 (O_181,N_20385,N_24212);
nand UO_182 (O_182,N_21149,N_22274);
and UO_183 (O_183,N_21211,N_24353);
nand UO_184 (O_184,N_24242,N_23282);
nor UO_185 (O_185,N_24100,N_23952);
and UO_186 (O_186,N_24506,N_20498);
xnor UO_187 (O_187,N_22409,N_23905);
and UO_188 (O_188,N_24358,N_20768);
or UO_189 (O_189,N_20791,N_22434);
and UO_190 (O_190,N_23549,N_22210);
or UO_191 (O_191,N_21157,N_23781);
and UO_192 (O_192,N_24331,N_24836);
and UO_193 (O_193,N_23753,N_21050);
nor UO_194 (O_194,N_24198,N_24731);
or UO_195 (O_195,N_23494,N_24617);
or UO_196 (O_196,N_22648,N_21343);
nand UO_197 (O_197,N_21753,N_22170);
nor UO_198 (O_198,N_24156,N_20523);
nor UO_199 (O_199,N_24355,N_22121);
nor UO_200 (O_200,N_21254,N_21417);
or UO_201 (O_201,N_23401,N_24811);
or UO_202 (O_202,N_21796,N_24673);
or UO_203 (O_203,N_21769,N_21642);
xor UO_204 (O_204,N_24663,N_22631);
nor UO_205 (O_205,N_21775,N_23470);
nand UO_206 (O_206,N_22914,N_23003);
nor UO_207 (O_207,N_20774,N_20587);
and UO_208 (O_208,N_23397,N_23411);
nand UO_209 (O_209,N_20125,N_20349);
nand UO_210 (O_210,N_24153,N_23475);
xnor UO_211 (O_211,N_21538,N_20164);
xor UO_212 (O_212,N_20515,N_21324);
xnor UO_213 (O_213,N_20251,N_22461);
or UO_214 (O_214,N_21827,N_22792);
and UO_215 (O_215,N_23448,N_24329);
or UO_216 (O_216,N_21828,N_24365);
or UO_217 (O_217,N_23019,N_23937);
nor UO_218 (O_218,N_24597,N_21114);
or UO_219 (O_219,N_23509,N_24549);
nand UO_220 (O_220,N_21173,N_20923);
or UO_221 (O_221,N_23006,N_21142);
nand UO_222 (O_222,N_24300,N_24724);
or UO_223 (O_223,N_21407,N_23642);
xnor UO_224 (O_224,N_22668,N_20398);
or UO_225 (O_225,N_20418,N_20556);
nand UO_226 (O_226,N_20316,N_21280);
nand UO_227 (O_227,N_22333,N_20780);
nor UO_228 (O_228,N_20748,N_23573);
or UO_229 (O_229,N_23128,N_24989);
nor UO_230 (O_230,N_21125,N_21720);
or UO_231 (O_231,N_21994,N_24332);
nor UO_232 (O_232,N_24971,N_21461);
and UO_233 (O_233,N_24554,N_20095);
nand UO_234 (O_234,N_20637,N_20186);
nor UO_235 (O_235,N_22413,N_21270);
nor UO_236 (O_236,N_22438,N_21073);
or UO_237 (O_237,N_23187,N_20875);
nor UO_238 (O_238,N_21644,N_24758);
xor UO_239 (O_239,N_21573,N_22323);
or UO_240 (O_240,N_23691,N_20245);
nor UO_241 (O_241,N_20476,N_22718);
nor UO_242 (O_242,N_24447,N_23285);
or UO_243 (O_243,N_22429,N_24970);
nor UO_244 (O_244,N_20220,N_20289);
nand UO_245 (O_245,N_24936,N_21466);
and UO_246 (O_246,N_21901,N_23531);
nand UO_247 (O_247,N_24247,N_21282);
or UO_248 (O_248,N_21204,N_23975);
and UO_249 (O_249,N_22459,N_20969);
and UO_250 (O_250,N_20713,N_22597);
nor UO_251 (O_251,N_21195,N_21393);
and UO_252 (O_252,N_23822,N_22006);
or UO_253 (O_253,N_23421,N_21790);
and UO_254 (O_254,N_23960,N_20156);
nor UO_255 (O_255,N_22920,N_24585);
or UO_256 (O_256,N_23541,N_23650);
and UO_257 (O_257,N_23750,N_21216);
xor UO_258 (O_258,N_22530,N_21314);
nor UO_259 (O_259,N_21135,N_21850);
and UO_260 (O_260,N_21319,N_23934);
nor UO_261 (O_261,N_20708,N_21953);
or UO_262 (O_262,N_22588,N_22250);
nor UO_263 (O_263,N_23638,N_20006);
or UO_264 (O_264,N_20388,N_20117);
or UO_265 (O_265,N_24809,N_20941);
or UO_266 (O_266,N_22288,N_20740);
nand UO_267 (O_267,N_20839,N_24002);
xnor UO_268 (O_268,N_20514,N_23148);
nand UO_269 (O_269,N_21327,N_21855);
nand UO_270 (O_270,N_21728,N_21895);
and UO_271 (O_271,N_23327,N_22537);
nand UO_272 (O_272,N_21081,N_20992);
and UO_273 (O_273,N_24599,N_24481);
nand UO_274 (O_274,N_24851,N_22324);
xnor UO_275 (O_275,N_23779,N_23390);
or UO_276 (O_276,N_23525,N_20187);
nor UO_277 (O_277,N_20808,N_24581);
and UO_278 (O_278,N_23858,N_20848);
nand UO_279 (O_279,N_22137,N_24808);
or UO_280 (O_280,N_22968,N_23592);
nand UO_281 (O_281,N_21731,N_22501);
xnor UO_282 (O_282,N_22230,N_23329);
and UO_283 (O_283,N_23356,N_23309);
or UO_284 (O_284,N_23249,N_24391);
nand UO_285 (O_285,N_22278,N_21345);
or UO_286 (O_286,N_22848,N_24995);
nand UO_287 (O_287,N_20124,N_22639);
or UO_288 (O_288,N_23261,N_21572);
nor UO_289 (O_289,N_20168,N_22377);
and UO_290 (O_290,N_22954,N_21685);
xor UO_291 (O_291,N_20448,N_21054);
and UO_292 (O_292,N_22637,N_21555);
and UO_293 (O_293,N_22927,N_23265);
and UO_294 (O_294,N_23737,N_20690);
xnor UO_295 (O_295,N_24478,N_22649);
and UO_296 (O_296,N_20379,N_24908);
or UO_297 (O_297,N_22598,N_24410);
and UO_298 (O_298,N_23138,N_22905);
nor UO_299 (O_299,N_23556,N_22951);
or UO_300 (O_300,N_23046,N_21570);
or UO_301 (O_301,N_23734,N_20335);
and UO_302 (O_302,N_21656,N_20035);
xor UO_303 (O_303,N_22075,N_21317);
and UO_304 (O_304,N_24702,N_23506);
or UO_305 (O_305,N_21436,N_21401);
or UO_306 (O_306,N_24840,N_22364);
and UO_307 (O_307,N_20802,N_24407);
and UO_308 (O_308,N_22543,N_24798);
nand UO_309 (O_309,N_23612,N_21809);
nor UO_310 (O_310,N_20386,N_23274);
nand UO_311 (O_311,N_22309,N_22796);
xor UO_312 (O_312,N_24881,N_24070);
and UO_313 (O_313,N_24576,N_21365);
and UO_314 (O_314,N_20921,N_23385);
xnor UO_315 (O_315,N_20412,N_24306);
and UO_316 (O_316,N_22626,N_23206);
nand UO_317 (O_317,N_21398,N_21867);
and UO_318 (O_318,N_24281,N_24527);
nor UO_319 (O_319,N_21029,N_21552);
nor UO_320 (O_320,N_20392,N_21341);
nand UO_321 (O_321,N_22492,N_22158);
nor UO_322 (O_322,N_21228,N_22540);
nor UO_323 (O_323,N_21385,N_24861);
nor UO_324 (O_324,N_20895,N_22944);
and UO_325 (O_325,N_20103,N_23048);
nand UO_326 (O_326,N_22525,N_24762);
and UO_327 (O_327,N_24582,N_22732);
xor UO_328 (O_328,N_21637,N_20963);
or UO_329 (O_329,N_20647,N_22619);
nand UO_330 (O_330,N_20937,N_24629);
or UO_331 (O_331,N_22077,N_21060);
nand UO_332 (O_332,N_20593,N_22040);
nand UO_333 (O_333,N_20692,N_22421);
or UO_334 (O_334,N_20359,N_20501);
nand UO_335 (O_335,N_24147,N_24397);
or UO_336 (O_336,N_22180,N_21586);
nor UO_337 (O_337,N_21146,N_21531);
and UO_338 (O_338,N_21203,N_23402);
or UO_339 (O_339,N_22932,N_23632);
and UO_340 (O_340,N_24077,N_22650);
nor UO_341 (O_341,N_23192,N_22798);
nor UO_342 (O_342,N_21147,N_21082);
nand UO_343 (O_343,N_20977,N_21046);
and UO_344 (O_344,N_21210,N_22847);
xor UO_345 (O_345,N_23568,N_21397);
nand UO_346 (O_346,N_24019,N_23234);
xor UO_347 (O_347,N_24803,N_24572);
nor UO_348 (O_348,N_22197,N_23407);
or UO_349 (O_349,N_24982,N_21961);
and UO_350 (O_350,N_24485,N_23266);
nand UO_351 (O_351,N_20108,N_24602);
xor UO_352 (O_352,N_23768,N_22806);
and UO_353 (O_353,N_21909,N_24920);
nor UO_354 (O_354,N_21108,N_24791);
nand UO_355 (O_355,N_21208,N_21512);
and UO_356 (O_356,N_22173,N_21956);
and UO_357 (O_357,N_23994,N_23287);
nor UO_358 (O_358,N_22615,N_22734);
and UO_359 (O_359,N_22832,N_24043);
nor UO_360 (O_360,N_22062,N_21671);
nor UO_361 (O_361,N_20861,N_23852);
or UO_362 (O_362,N_23035,N_21900);
or UO_363 (O_363,N_23667,N_20616);
or UO_364 (O_364,N_24239,N_23672);
or UO_365 (O_365,N_21263,N_20680);
nor UO_366 (O_366,N_23570,N_24440);
nand UO_367 (O_367,N_24364,N_22865);
nor UO_368 (O_368,N_24868,N_22087);
or UO_369 (O_369,N_21235,N_24507);
or UO_370 (O_370,N_24621,N_20660);
nor UO_371 (O_371,N_22478,N_21369);
nor UO_372 (O_372,N_20082,N_22880);
nand UO_373 (O_373,N_20606,N_22320);
nor UO_374 (O_374,N_24446,N_22539);
nand UO_375 (O_375,N_21717,N_24619);
and UO_376 (O_376,N_22143,N_22112);
and UO_377 (O_377,N_23149,N_22861);
nor UO_378 (O_378,N_20783,N_24894);
or UO_379 (O_379,N_22350,N_23094);
xnor UO_380 (O_380,N_24448,N_22952);
xor UO_381 (O_381,N_21893,N_21223);
xor UO_382 (O_382,N_23213,N_21508);
or UO_383 (O_383,N_20486,N_23338);
nand UO_384 (O_384,N_21975,N_20284);
nand UO_385 (O_385,N_24456,N_20850);
and UO_386 (O_386,N_20814,N_24941);
and UO_387 (O_387,N_20018,N_24846);
nor UO_388 (O_388,N_21331,N_22930);
nand UO_389 (O_389,N_22881,N_24169);
and UO_390 (O_390,N_20507,N_22054);
nor UO_391 (O_391,N_21064,N_21792);
and UO_392 (O_392,N_23267,N_24837);
nand UO_393 (O_393,N_23340,N_24490);
nand UO_394 (O_394,N_22890,N_20211);
and UO_395 (O_395,N_24618,N_22347);
nor UO_396 (O_396,N_20898,N_24185);
and UO_397 (O_397,N_22838,N_21139);
nand UO_398 (O_398,N_21691,N_23499);
nor UO_399 (O_399,N_22445,N_21201);
nand UO_400 (O_400,N_21232,N_24172);
xnor UO_401 (O_401,N_23068,N_24500);
and UO_402 (O_402,N_20154,N_24248);
or UO_403 (O_403,N_21601,N_21869);
and UO_404 (O_404,N_22595,N_20907);
nor UO_405 (O_405,N_21025,N_24033);
or UO_406 (O_406,N_22466,N_24742);
nor UO_407 (O_407,N_24806,N_20368);
nor UO_408 (O_408,N_24376,N_20908);
nor UO_409 (O_409,N_22937,N_22363);
nor UO_410 (O_410,N_20743,N_21898);
or UO_411 (O_411,N_23124,N_23074);
nand UO_412 (O_412,N_24165,N_22844);
or UO_413 (O_413,N_21594,N_22050);
or UO_414 (O_414,N_21835,N_21579);
and UO_415 (O_415,N_21265,N_21038);
and UO_416 (O_416,N_22118,N_21926);
nand UO_417 (O_417,N_22127,N_24939);
nand UO_418 (O_418,N_20821,N_20266);
nor UO_419 (O_419,N_20380,N_20857);
and UO_420 (O_420,N_23211,N_23454);
and UO_421 (O_421,N_23252,N_23326);
nand UO_422 (O_422,N_20795,N_21681);
nor UO_423 (O_423,N_24400,N_22680);
and UO_424 (O_424,N_23806,N_21702);
nand UO_425 (O_425,N_22228,N_22829);
and UO_426 (O_426,N_20345,N_21757);
or UO_427 (O_427,N_24879,N_22545);
and UO_428 (O_428,N_24357,N_23077);
or UO_429 (O_429,N_22969,N_22399);
or UO_430 (O_430,N_22509,N_22252);
nand UO_431 (O_431,N_23041,N_23600);
nand UO_432 (O_432,N_20837,N_21376);
nor UO_433 (O_433,N_21186,N_22286);
nor UO_434 (O_434,N_22370,N_24998);
xnor UO_435 (O_435,N_24847,N_20456);
nand UO_436 (O_436,N_21891,N_20793);
nor UO_437 (O_437,N_22706,N_24161);
xnor UO_438 (O_438,N_20120,N_23915);
nand UO_439 (O_439,N_20730,N_21604);
and UO_440 (O_440,N_20571,N_24525);
nand UO_441 (O_441,N_21660,N_22967);
nor UO_442 (O_442,N_23240,N_21597);
and UO_443 (O_443,N_21894,N_22897);
or UO_444 (O_444,N_24046,N_20489);
or UO_445 (O_445,N_22181,N_23389);
nand UO_446 (O_446,N_23880,N_20389);
nand UO_447 (O_447,N_22272,N_24041);
and UO_448 (O_448,N_21964,N_23227);
and UO_449 (O_449,N_21296,N_23312);
nor UO_450 (O_450,N_21630,N_24265);
and UO_451 (O_451,N_21654,N_21104);
nand UO_452 (O_452,N_23384,N_24055);
nor UO_453 (O_453,N_23291,N_24009);
and UO_454 (O_454,N_22217,N_21112);
or UO_455 (O_455,N_23522,N_24199);
nor UO_456 (O_456,N_20011,N_20106);
nand UO_457 (O_457,N_23964,N_22163);
nor UO_458 (O_458,N_22972,N_22804);
nand UO_459 (O_459,N_21733,N_22402);
or UO_460 (O_460,N_20319,N_20465);
or UO_461 (O_461,N_22337,N_20629);
nor UO_462 (O_462,N_24411,N_22613);
nand UO_463 (O_463,N_22600,N_21768);
or UO_464 (O_464,N_23680,N_22818);
nor UO_465 (O_465,N_23540,N_23850);
nand UO_466 (O_466,N_20567,N_22783);
and UO_467 (O_467,N_24728,N_24394);
and UO_468 (O_468,N_23318,N_20596);
or UO_469 (O_469,N_20967,N_23614);
xnor UO_470 (O_470,N_21271,N_23763);
and UO_471 (O_471,N_20718,N_22224);
and UO_472 (O_472,N_23887,N_20994);
nor UO_473 (O_473,N_22430,N_21968);
and UO_474 (O_474,N_20554,N_20689);
nor UO_475 (O_475,N_20427,N_24665);
and UO_476 (O_476,N_22108,N_24349);
nor UO_477 (O_477,N_21017,N_22406);
and UO_478 (O_478,N_21098,N_23843);
or UO_479 (O_479,N_24180,N_21014);
or UO_480 (O_480,N_23391,N_21587);
or UO_481 (O_481,N_23595,N_22923);
nand UO_482 (O_482,N_21914,N_21464);
nand UO_483 (O_483,N_20460,N_23460);
xnor UO_484 (O_484,N_21289,N_24167);
nor UO_485 (O_485,N_24096,N_24215);
nor UO_486 (O_486,N_23030,N_20008);
nor UO_487 (O_487,N_23819,N_23798);
nor UO_488 (O_488,N_24350,N_21215);
nand UO_489 (O_489,N_21993,N_22605);
nand UO_490 (O_490,N_21283,N_22396);
or UO_491 (O_491,N_20051,N_22117);
or UO_492 (O_492,N_23716,N_22467);
nand UO_493 (O_493,N_24218,N_23891);
nor UO_494 (O_494,N_23613,N_24595);
nor UO_495 (O_495,N_22303,N_24759);
nor UO_496 (O_496,N_22970,N_22416);
or UO_497 (O_497,N_22803,N_20846);
xor UO_498 (O_498,N_21287,N_22947);
nand UO_499 (O_499,N_23216,N_24183);
and UO_500 (O_500,N_20649,N_23907);
nor UO_501 (O_501,N_22993,N_23764);
nand UO_502 (O_502,N_21316,N_22172);
nand UO_503 (O_503,N_23997,N_20020);
and UO_504 (O_504,N_20296,N_22213);
nand UO_505 (O_505,N_22622,N_20678);
nor UO_506 (O_506,N_20939,N_21683);
xnor UO_507 (O_507,N_21495,N_24780);
and UO_508 (O_508,N_21514,N_22577);
and UO_509 (O_509,N_24154,N_24689);
and UO_510 (O_510,N_22716,N_24379);
or UO_511 (O_511,N_21825,N_21647);
nor UO_512 (O_512,N_23774,N_24176);
or UO_513 (O_513,N_20840,N_24752);
or UO_514 (O_514,N_20054,N_23830);
xnor UO_515 (O_515,N_23596,N_24557);
and UO_516 (O_516,N_21256,N_23320);
nand UO_517 (O_517,N_23572,N_22559);
nor UO_518 (O_518,N_23917,N_24438);
and UO_519 (O_519,N_22623,N_24393);
nor UO_520 (O_520,N_21118,N_21352);
nand UO_521 (O_521,N_20825,N_21852);
nor UO_522 (O_522,N_20505,N_23709);
and UO_523 (O_523,N_20030,N_21569);
nor UO_524 (O_524,N_23844,N_24661);
nor UO_525 (O_525,N_23517,N_20201);
and UO_526 (O_526,N_21939,N_22264);
and UO_527 (O_527,N_23151,N_22725);
nor UO_528 (O_528,N_24534,N_20260);
or UO_529 (O_529,N_23462,N_22355);
nor UO_530 (O_530,N_21829,N_24144);
and UO_531 (O_531,N_20409,N_20807);
nor UO_532 (O_532,N_20915,N_23876);
and UO_533 (O_533,N_23586,N_23561);
nand UO_534 (O_534,N_24496,N_22119);
nand UO_535 (O_535,N_23428,N_22955);
or UO_536 (O_536,N_20074,N_23496);
or UO_537 (O_537,N_22735,N_20970);
and UO_538 (O_538,N_24788,N_23245);
xnor UO_539 (O_539,N_22057,N_24477);
and UO_540 (O_540,N_23076,N_22677);
and UO_541 (O_541,N_20701,N_23441);
and UO_542 (O_542,N_23109,N_22471);
and UO_543 (O_543,N_21264,N_20829);
nand UO_544 (O_544,N_23859,N_24163);
and UO_545 (O_545,N_24567,N_20543);
nand UO_546 (O_546,N_24395,N_23445);
nand UO_547 (O_547,N_22220,N_24263);
nand UO_548 (O_548,N_20474,N_24918);
or UO_549 (O_549,N_20576,N_21915);
nor UO_550 (O_550,N_22046,N_20219);
xnor UO_551 (O_551,N_24514,N_24262);
and UO_552 (O_552,N_20407,N_24388);
and UO_553 (O_553,N_24897,N_22107);
nand UO_554 (O_554,N_21562,N_20287);
nand UO_555 (O_555,N_23292,N_23083);
nor UO_556 (O_556,N_23665,N_21380);
nand UO_557 (O_557,N_23508,N_24678);
nand UO_558 (O_558,N_20098,N_24497);
or UO_559 (O_559,N_23395,N_20560);
or UO_560 (O_560,N_21501,N_22202);
or UO_561 (O_561,N_21141,N_24885);
nand UO_562 (O_562,N_24679,N_20691);
and UO_563 (O_563,N_24429,N_21856);
nor UO_564 (O_564,N_20045,N_21907);
nand UO_565 (O_565,N_22941,N_20338);
nand UO_566 (O_566,N_23097,N_23368);
or UO_567 (O_567,N_24430,N_22704);
nand UO_568 (O_568,N_22900,N_21680);
nor UO_569 (O_569,N_23246,N_22134);
and UO_570 (O_570,N_22603,N_21641);
or UO_571 (O_571,N_23730,N_21238);
and UO_572 (O_572,N_23720,N_20210);
nor UO_573 (O_573,N_22276,N_23659);
nor UO_574 (O_574,N_22863,N_20529);
nand UO_575 (O_575,N_22875,N_21193);
nor UO_576 (O_576,N_21333,N_21860);
nor UO_577 (O_577,N_21212,N_24351);
and UO_578 (O_578,N_24223,N_21249);
nand UO_579 (O_579,N_21840,N_20372);
and UO_580 (O_580,N_21431,N_22029);
or UO_581 (O_581,N_22225,N_23490);
nor UO_582 (O_582,N_22376,N_23314);
or UO_583 (O_583,N_23467,N_24737);
nor UO_584 (O_584,N_24789,N_21455);
nor UO_585 (O_585,N_21831,N_21375);
or UO_586 (O_586,N_22521,N_21521);
nand UO_587 (O_587,N_22388,N_20509);
or UO_588 (O_588,N_20767,N_21741);
nand UO_589 (O_589,N_22640,N_23201);
nand UO_590 (O_590,N_24699,N_22686);
or UO_591 (O_591,N_21136,N_21711);
or UO_592 (O_592,N_22440,N_22486);
and UO_593 (O_593,N_24069,N_21746);
or UO_594 (O_594,N_24294,N_23476);
or UO_595 (O_595,N_23812,N_23022);
nor UO_596 (O_596,N_21109,N_23064);
and UO_597 (O_597,N_20672,N_22385);
nor UO_598 (O_598,N_21363,N_20086);
nand UO_599 (O_599,N_20889,N_21944);
nand UO_600 (O_600,N_22985,N_24560);
nor UO_601 (O_601,N_24087,N_22386);
and UO_602 (O_602,N_21874,N_24234);
nor UO_603 (O_603,N_23807,N_24021);
nand UO_604 (O_604,N_22221,N_22080);
nand UO_605 (O_605,N_20073,N_22764);
and UO_606 (O_606,N_22381,N_20799);
and UO_607 (O_607,N_22528,N_22997);
xnor UO_608 (O_608,N_20043,N_20406);
and UO_609 (O_609,N_21410,N_22022);
nand UO_610 (O_610,N_24945,N_23824);
nand UO_611 (O_611,N_23648,N_21812);
nand UO_612 (O_612,N_23131,N_20450);
nor UO_613 (O_613,N_22001,N_22182);
nand UO_614 (O_614,N_24862,N_23111);
nand UO_615 (O_615,N_22155,N_20715);
or UO_616 (O_616,N_24786,N_24133);
or UO_617 (O_617,N_23344,N_24591);
xor UO_618 (O_618,N_20169,N_20589);
nor UO_619 (O_619,N_24201,N_20097);
nor UO_620 (O_620,N_23681,N_20487);
nand UO_621 (O_621,N_21603,N_22926);
nor UO_622 (O_622,N_22200,N_21129);
nand UO_623 (O_623,N_22114,N_22047);
and UO_624 (O_624,N_21144,N_20696);
nand UO_625 (O_625,N_22679,N_22518);
or UO_626 (O_626,N_21269,N_23552);
and UO_627 (O_627,N_21297,N_24824);
nand UO_628 (O_628,N_24878,N_24107);
nand UO_629 (O_629,N_24401,N_21838);
and UO_630 (O_630,N_22484,N_22785);
or UO_631 (O_631,N_22751,N_23115);
or UO_632 (O_632,N_21705,N_22265);
or UO_633 (O_633,N_22772,N_22084);
nor UO_634 (O_634,N_23618,N_20614);
nor UO_635 (O_635,N_23782,N_21416);
or UO_636 (O_636,N_22280,N_23136);
xnor UO_637 (O_637,N_21051,N_21183);
and UO_638 (O_638,N_20113,N_22965);
and UO_639 (O_639,N_22722,N_21061);
xnor UO_640 (O_640,N_22762,N_24542);
nand UO_641 (O_641,N_22169,N_24036);
nand UO_642 (O_642,N_23330,N_20763);
and UO_643 (O_643,N_23692,N_24741);
or UO_644 (O_644,N_20458,N_22455);
nand UO_645 (O_645,N_24625,N_21143);
or UO_646 (O_646,N_22036,N_22581);
xnor UO_647 (O_647,N_21445,N_22899);
or UO_648 (O_648,N_23609,N_21596);
or UO_649 (O_649,N_22896,N_20553);
nand UO_650 (O_650,N_21744,N_23127);
nand UO_651 (O_651,N_22692,N_23594);
nand UO_652 (O_652,N_21719,N_23791);
or UO_653 (O_653,N_21004,N_21368);
and UO_654 (O_654,N_22575,N_22670);
or UO_655 (O_655,N_22326,N_24437);
nor UO_656 (O_656,N_23825,N_21688);
xnor UO_657 (O_657,N_21337,N_21154);
and UO_658 (O_658,N_20010,N_21734);
or UO_659 (O_659,N_23551,N_22822);
or UO_660 (O_660,N_23974,N_24405);
nand UO_661 (O_661,N_23542,N_20013);
xnor UO_662 (O_662,N_20962,N_23724);
or UO_663 (O_663,N_23029,N_20463);
or UO_664 (O_664,N_20655,N_24954);
and UO_665 (O_665,N_20943,N_23456);
or UO_666 (O_666,N_20157,N_21617);
nor UO_667 (O_667,N_20137,N_24122);
or UO_668 (O_668,N_21080,N_23723);
nor UO_669 (O_669,N_21067,N_21016);
nand UO_670 (O_670,N_23616,N_24739);
or UO_671 (O_671,N_23874,N_24191);
or UO_672 (O_672,N_24389,N_22256);
nor UO_673 (O_673,N_24607,N_20936);
nor UO_674 (O_674,N_20901,N_23930);
or UO_675 (O_675,N_21706,N_23539);
and UO_676 (O_676,N_24230,N_20877);
or UO_677 (O_677,N_22958,N_23122);
or UO_678 (O_678,N_23788,N_20762);
or UO_679 (O_679,N_20353,N_20468);
or UO_680 (O_680,N_21879,N_23979);
nor UO_681 (O_681,N_24221,N_21076);
or UO_682 (O_682,N_23366,N_24162);
xor UO_683 (O_683,N_24195,N_23185);
nand UO_684 (O_684,N_23520,N_22367);
or UO_685 (O_685,N_23772,N_22194);
xor UO_686 (O_686,N_20646,N_21947);
and UO_687 (O_687,N_24630,N_22380);
nand UO_688 (O_688,N_24726,N_20203);
or UO_689 (O_689,N_21985,N_23674);
and UO_690 (O_690,N_20585,N_21409);
and UO_691 (O_691,N_24896,N_24037);
xnor UO_692 (O_692,N_23511,N_21299);
nand UO_693 (O_693,N_22357,N_23042);
nand UO_694 (O_694,N_22094,N_21599);
nor UO_695 (O_695,N_22738,N_24559);
xnor UO_696 (O_696,N_22115,N_20347);
and UO_697 (O_697,N_21467,N_23748);
or UO_698 (O_698,N_23101,N_21841);
and UO_699 (O_699,N_20749,N_23923);
and UO_700 (O_700,N_24533,N_22673);
xor UO_701 (O_701,N_21367,N_23689);
nor UO_702 (O_702,N_24985,N_20652);
and UO_703 (O_703,N_21580,N_21709);
and UO_704 (O_704,N_22433,N_20663);
nand UO_705 (O_705,N_20484,N_22850);
nor UO_706 (O_706,N_20990,N_24271);
nor UO_707 (O_707,N_20332,N_20738);
nand UO_708 (O_708,N_24664,N_22211);
and UO_709 (O_709,N_22468,N_23683);
or UO_710 (O_710,N_24994,N_21206);
nand UO_711 (O_711,N_21511,N_21934);
nor UO_712 (O_712,N_21725,N_21402);
or UO_713 (O_713,N_21933,N_20182);
and UO_714 (O_714,N_21986,N_23032);
nor UO_715 (O_715,N_21739,N_20153);
or UO_716 (O_716,N_24383,N_24170);
or UO_717 (O_717,N_23842,N_20683);
nand UO_718 (O_718,N_24495,N_22973);
nor UO_719 (O_719,N_23107,N_23598);
or UO_720 (O_720,N_23833,N_24004);
xnor UO_721 (O_721,N_20067,N_23813);
nand UO_722 (O_722,N_23250,N_20924);
nand UO_723 (O_723,N_23834,N_20974);
nor UO_724 (O_724,N_24950,N_24869);
nor UO_725 (O_725,N_24886,N_23450);
and UO_726 (O_726,N_23534,N_23129);
nand UO_727 (O_727,N_22587,N_23284);
and UO_728 (O_728,N_23264,N_21837);
and UO_729 (O_729,N_24193,N_21910);
nor UO_730 (O_730,N_20789,N_20304);
nor UO_731 (O_731,N_22456,N_20413);
and UO_732 (O_732,N_21020,N_23177);
nor UO_733 (O_733,N_21978,N_20865);
and UO_734 (O_734,N_21842,N_20434);
or UO_735 (O_735,N_20613,N_24570);
or UO_736 (O_736,N_23420,N_23130);
and UO_737 (O_737,N_24190,N_22887);
nor UO_738 (O_738,N_22473,N_20321);
nand UO_739 (O_739,N_23981,N_21714);
nor UO_740 (O_740,N_24066,N_22379);
nor UO_741 (O_741,N_21995,N_21472);
nand UO_742 (O_742,N_20504,N_23863);
and UO_743 (O_743,N_21102,N_20061);
nor UO_744 (O_744,N_23239,N_23367);
and UO_745 (O_745,N_21138,N_23879);
nand UO_746 (O_746,N_24860,N_24623);
nor UO_747 (O_747,N_22109,N_22124);
nor UO_748 (O_748,N_23465,N_23233);
nand UO_749 (O_749,N_23283,N_23719);
nand UO_750 (O_750,N_20437,N_23105);
or UO_751 (O_751,N_24072,N_22759);
nand UO_752 (O_752,N_23629,N_23423);
nand UO_753 (O_753,N_20573,N_23615);
nand UO_754 (O_754,N_24307,N_23625);
and UO_755 (O_755,N_22675,N_23966);
or UO_756 (O_756,N_24285,N_20594);
nand UO_757 (O_757,N_23948,N_22548);
nor UO_758 (O_758,N_24698,N_20261);
or UO_759 (O_759,N_24888,N_23660);
or UO_760 (O_760,N_23501,N_23102);
nand UO_761 (O_761,N_22747,N_23702);
or UO_762 (O_762,N_23795,N_24460);
nand UO_763 (O_763,N_21389,N_22267);
and UO_764 (O_764,N_23657,N_21384);
or UO_765 (O_765,N_20714,N_22122);
or UO_766 (O_766,N_24564,N_21788);
nor UO_767 (O_767,N_24799,N_20794);
or UO_768 (O_768,N_20424,N_21442);
and UO_769 (O_769,N_24772,N_20544);
and UO_770 (O_770,N_21836,N_20586);
and UO_771 (O_771,N_23550,N_23463);
xor UO_772 (O_772,N_20997,N_20575);
and UO_773 (O_773,N_24213,N_24253);
or UO_774 (O_774,N_23984,N_23014);
xor UO_775 (O_775,N_23222,N_24593);
or UO_776 (O_776,N_21188,N_23197);
and UO_777 (O_777,N_23328,N_21610);
nand UO_778 (O_778,N_20417,N_21236);
nor UO_779 (O_779,N_21267,N_21941);
xor UO_780 (O_780,N_21639,N_22044);
nor UO_781 (O_781,N_22538,N_20026);
nand UO_782 (O_782,N_23354,N_20656);
or UO_783 (O_783,N_22882,N_21808);
nand UO_784 (O_784,N_20632,N_23875);
nor UO_785 (O_785,N_20138,N_21948);
nor UO_786 (O_786,N_21451,N_24586);
nand UO_787 (O_787,N_23024,N_23276);
nand UO_788 (O_788,N_23978,N_21026);
nand UO_789 (O_789,N_24377,N_21465);
and UO_790 (O_790,N_20263,N_22498);
and UO_791 (O_791,N_23142,N_22551);
nand UO_792 (O_792,N_24765,N_23374);
or UO_793 (O_793,N_23160,N_24119);
nor UO_794 (O_794,N_20374,N_24813);
and UO_795 (O_795,N_21892,N_24552);
nor UO_796 (O_796,N_24796,N_22101);
or UO_797 (O_797,N_23676,N_23376);
and UO_798 (O_798,N_20745,N_22948);
or UO_799 (O_799,N_22495,N_21607);
nor UO_800 (O_800,N_24715,N_24296);
or UO_801 (O_801,N_24168,N_21012);
nand UO_802 (O_802,N_24494,N_24973);
and UO_803 (O_803,N_24427,N_23697);
nand UO_804 (O_804,N_20703,N_24293);
and UO_805 (O_805,N_22711,N_24746);
nor UO_806 (O_806,N_21090,N_20902);
or UO_807 (O_807,N_22586,N_20360);
or UO_808 (O_808,N_21509,N_20516);
and UO_809 (O_809,N_20787,N_24005);
and UO_810 (O_810,N_22823,N_23932);
xor UO_811 (O_811,N_21557,N_23056);
and UO_812 (O_812,N_22604,N_22329);
and UO_813 (O_813,N_24754,N_24370);
nor UO_814 (O_814,N_21689,N_22907);
nor UO_815 (O_815,N_21205,N_22164);
nor UO_816 (O_816,N_22411,N_24384);
and UO_817 (O_817,N_22555,N_20252);
and UO_818 (O_818,N_21904,N_20823);
and UO_819 (O_819,N_20897,N_24268);
nor UO_820 (O_820,N_20502,N_24103);
nor UO_821 (O_821,N_21490,N_21543);
nand UO_822 (O_822,N_20152,N_22405);
nand UO_823 (O_823,N_22443,N_20015);
and UO_824 (O_824,N_20723,N_21563);
and UO_825 (O_825,N_22196,N_20882);
nor UO_826 (O_826,N_23324,N_22257);
and UO_827 (O_827,N_24115,N_20350);
and UO_828 (O_828,N_23547,N_21646);
nor UO_829 (O_829,N_23926,N_23912);
and UO_830 (O_830,N_21658,N_22909);
xnor UO_831 (O_831,N_20358,N_23867);
nor UO_832 (O_832,N_23645,N_21261);
or UO_833 (O_833,N_21473,N_24345);
or UO_834 (O_834,N_20778,N_20114);
nand UO_835 (O_835,N_23849,N_23583);
nand UO_836 (O_836,N_20115,N_24434);
or UO_837 (O_837,N_20188,N_24659);
nand UO_838 (O_838,N_20171,N_24842);
nor UO_839 (O_839,N_24120,N_22013);
nand UO_840 (O_840,N_20123,N_24873);
nand UO_841 (O_841,N_24898,N_21598);
xnor UO_842 (O_842,N_22746,N_23045);
nor UO_843 (O_843,N_20558,N_23317);
nand UO_844 (O_844,N_22500,N_22123);
or UO_845 (O_845,N_20545,N_22031);
or UO_846 (O_846,N_20836,N_24983);
and UO_847 (O_847,N_22005,N_22720);
or UO_848 (O_848,N_20591,N_20785);
nand UO_849 (O_849,N_23529,N_20485);
or UO_850 (O_850,N_22048,N_21101);
nand UO_851 (O_851,N_21084,N_22053);
or UO_852 (O_852,N_22360,N_24756);
nand UO_853 (O_853,N_23965,N_22425);
nand UO_854 (O_854,N_21564,N_24275);
xor UO_855 (O_855,N_22372,N_23695);
and UO_856 (O_856,N_22362,N_24733);
nor UO_857 (O_857,N_22589,N_21672);
or UO_858 (O_858,N_23619,N_23591);
nand UO_859 (O_859,N_23255,N_24590);
or UO_860 (O_860,N_21955,N_24470);
nor UO_861 (O_861,N_21770,N_22830);
and UO_862 (O_862,N_23587,N_22152);
xor UO_863 (O_863,N_24175,N_24472);
nor UO_864 (O_864,N_21833,N_22175);
xnor UO_865 (O_865,N_20267,N_24423);
or UO_866 (O_866,N_21047,N_24895);
xor UO_867 (O_867,N_20750,N_24722);
or UO_868 (O_868,N_20798,N_23350);
nand UO_869 (O_869,N_24508,N_21735);
and UO_870 (O_870,N_23523,N_22207);
and UO_871 (O_871,N_24718,N_21726);
nand UO_872 (O_872,N_21449,N_22665);
nor UO_873 (O_873,N_24232,N_20883);
or UO_874 (O_874,N_20525,N_21732);
and UO_875 (O_875,N_23987,N_20540);
xnor UO_876 (O_876,N_22793,N_23635);
or UO_877 (O_877,N_22065,N_20459);
nand UO_878 (O_878,N_21370,N_23698);
nor UO_879 (O_879,N_23078,N_21533);
or UO_880 (O_880,N_23382,N_20788);
or UO_881 (O_881,N_24797,N_24354);
xor UO_882 (O_882,N_23687,N_22239);
xor UO_883 (O_883,N_22879,N_21659);
nor UO_884 (O_884,N_21541,N_22606);
and UO_885 (O_885,N_23690,N_24324);
and UO_886 (O_886,N_24732,N_24227);
and UO_887 (O_887,N_24382,N_24536);
nor UO_888 (O_888,N_24561,N_23845);
nand UO_889 (O_889,N_24023,N_20199);
nand UO_890 (O_890,N_21851,N_20466);
nor UO_891 (O_891,N_23886,N_20070);
and UO_892 (O_892,N_24749,N_20851);
nand UO_893 (O_893,N_20842,N_21233);
nor UO_894 (O_894,N_22789,N_20920);
and UO_895 (O_895,N_20339,N_20072);
xnor UO_896 (O_896,N_22251,N_22321);
or UO_897 (O_897,N_22302,N_22135);
or UO_898 (O_898,N_20445,N_24937);
nand UO_899 (O_899,N_22024,N_23268);
or UO_900 (O_900,N_20147,N_20547);
or UO_901 (O_901,N_20579,N_21381);
and UO_902 (O_902,N_24272,N_22892);
nor UO_903 (O_903,N_21657,N_21422);
nand UO_904 (O_904,N_22042,N_23593);
and UO_905 (O_905,N_21217,N_24011);
or UO_906 (O_906,N_23200,N_22497);
nand UO_907 (O_907,N_20478,N_24710);
nor UO_908 (O_908,N_23417,N_23098);
nor UO_909 (O_909,N_24942,N_23332);
or UO_910 (O_910,N_22782,N_20891);
nand UO_911 (O_911,N_23785,N_23406);
or UO_912 (O_912,N_24648,N_24126);
xnor UO_913 (O_913,N_20758,N_24203);
nand UO_914 (O_914,N_21359,N_20440);
nand UO_915 (O_915,N_24864,N_24992);
or UO_916 (O_916,N_24068,N_23636);
and UO_917 (O_917,N_21105,N_22479);
and UO_918 (O_918,N_21332,N_23500);
nor UO_919 (O_919,N_23336,N_23585);
nor UO_920 (O_920,N_20675,N_21412);
nand UO_921 (O_921,N_21119,N_24578);
nor UO_922 (O_922,N_22232,N_20513);
and UO_923 (O_923,N_22437,N_24034);
or UO_924 (O_924,N_24424,N_20236);
and UO_925 (O_925,N_22852,N_22325);
and UO_926 (O_926,N_23524,N_21816);
or UO_927 (O_927,N_20709,N_24084);
or UO_928 (O_928,N_23933,N_22404);
and UO_929 (O_929,N_22315,N_21041);
nor UO_930 (O_930,N_20408,N_20081);
or UO_931 (O_931,N_20003,N_22441);
nor UO_932 (O_932,N_22401,N_22033);
nand UO_933 (O_933,N_21364,N_22338);
and UO_934 (O_934,N_23939,N_21595);
nor UO_935 (O_935,N_21075,N_21549);
or UO_936 (O_936,N_24462,N_20611);
and UO_937 (O_937,N_22984,N_22451);
or UO_938 (O_938,N_21391,N_22322);
and UO_939 (O_939,N_23289,N_24912);
or UO_940 (O_940,N_24219,N_22620);
and UO_941 (O_941,N_21127,N_22962);
or UO_942 (O_942,N_24373,N_20669);
nor UO_943 (O_943,N_21505,N_20436);
nand UO_944 (O_944,N_20404,N_20076);
and UO_945 (O_945,N_23305,N_21010);
or UO_946 (O_946,N_21911,N_22964);
nand UO_947 (O_947,N_23590,N_21600);
nor UO_948 (O_948,N_23033,N_21758);
xnor UO_949 (O_949,N_22190,N_24784);
xnor UO_950 (O_950,N_24831,N_24171);
nand UO_951 (O_951,N_20535,N_24932);
or UO_952 (O_952,N_20520,N_23457);
and UO_953 (O_953,N_22279,N_23739);
and UO_954 (O_954,N_21443,N_22966);
nand UO_955 (O_955,N_20892,N_22715);
xnor UO_956 (O_956,N_23706,N_24705);
nand UO_957 (O_957,N_23089,N_23762);
nor UO_958 (O_958,N_22858,N_21662);
and UO_959 (O_959,N_23005,N_22660);
or UO_960 (O_960,N_23993,N_21301);
nor UO_961 (O_961,N_23146,N_21032);
and UO_962 (O_962,N_24957,N_24283);
nand UO_963 (O_963,N_20009,N_22298);
or UO_964 (O_964,N_24935,N_21550);
nor UO_965 (O_965,N_23810,N_20295);
and UO_966 (O_966,N_21366,N_24362);
nand UO_967 (O_967,N_20781,N_23851);
and UO_968 (O_968,N_23455,N_21438);
nor UO_969 (O_969,N_20720,N_22204);
or UO_970 (O_970,N_24029,N_23717);
nand UO_971 (O_971,N_21818,N_24977);
nand UO_972 (O_972,N_23603,N_22933);
nand UO_973 (O_973,N_22840,N_24646);
or UO_974 (O_974,N_22475,N_22100);
and UO_975 (O_975,N_23118,N_24926);
and UO_976 (O_976,N_21406,N_22423);
and UO_977 (O_977,N_20351,N_24336);
nand UO_978 (O_978,N_20623,N_22419);
nor UO_979 (O_979,N_24322,N_24635);
or UO_980 (O_980,N_24280,N_20804);
nor UO_981 (O_981,N_21439,N_22714);
nor UO_982 (O_982,N_21485,N_22602);
nand UO_983 (O_983,N_21545,N_22638);
or UO_984 (O_984,N_20062,N_21518);
and UO_985 (O_985,N_20565,N_23925);
xor UO_986 (O_986,N_23721,N_24102);
and UO_987 (O_987,N_21931,N_21958);
and UO_988 (O_988,N_24965,N_20403);
and UO_989 (O_989,N_24155,N_23155);
and UO_990 (O_990,N_24775,N_24632);
and UO_991 (O_991,N_22231,N_20391);
nand UO_992 (O_992,N_22683,N_20624);
or UO_993 (O_993,N_21626,N_23270);
and UO_994 (O_994,N_24521,N_21920);
and UO_995 (O_995,N_23082,N_24774);
or UO_996 (O_996,N_23571,N_21244);
nand UO_997 (O_997,N_24404,N_22361);
nor UO_998 (O_998,N_21426,N_24848);
nand UO_999 (O_999,N_22868,N_22476);
and UO_1000 (O_1000,N_22240,N_24519);
nand UO_1001 (O_1001,N_24256,N_23888);
nor UO_1002 (O_1002,N_24833,N_24380);
and UO_1003 (O_1003,N_22045,N_22229);
nor UO_1004 (O_1004,N_24008,N_23380);
and UO_1005 (O_1005,N_24966,N_24137);
nor UO_1006 (O_1006,N_24568,N_23188);
and UO_1007 (O_1007,N_24828,N_20442);
or UO_1008 (O_1008,N_24668,N_21000);
and UO_1009 (O_1009,N_23321,N_20577);
and UO_1010 (O_1010,N_22874,N_20390);
nor UO_1011 (O_1011,N_23298,N_20630);
or UO_1012 (O_1012,N_21486,N_24952);
or UO_1013 (O_1013,N_20933,N_21470);
nand UO_1014 (O_1014,N_22780,N_24241);
nor UO_1015 (O_1015,N_21497,N_21151);
and UO_1016 (O_1016,N_22502,N_23472);
nor UO_1017 (O_1017,N_20449,N_22341);
and UO_1018 (O_1018,N_20598,N_23218);
xnor UO_1019 (O_1019,N_24891,N_23208);
xor UO_1020 (O_1020,N_21006,N_23269);
xnor UO_1021 (O_1021,N_24192,N_23004);
or UO_1022 (O_1022,N_22942,N_23043);
nand UO_1023 (O_1023,N_23910,N_22293);
or UO_1024 (O_1024,N_20518,N_23235);
nand UO_1025 (O_1025,N_24596,N_20130);
nand UO_1026 (O_1026,N_21350,N_22176);
and UO_1027 (O_1027,N_22512,N_22553);
and UO_1028 (O_1028,N_20856,N_23182);
nor UO_1029 (O_1029,N_23000,N_21629);
and UO_1030 (O_1030,N_20717,N_22749);
or UO_1031 (O_1031,N_22238,N_20161);
nor UO_1032 (O_1032,N_23099,N_23028);
nor UO_1033 (O_1033,N_21295,N_23904);
and UO_1034 (O_1034,N_21480,N_21675);
nand UO_1035 (O_1035,N_22356,N_21224);
nand UO_1036 (O_1036,N_23700,N_23677);
nor UO_1037 (O_1037,N_21153,N_24098);
nand UO_1038 (O_1038,N_22079,N_20183);
or UO_1039 (O_1039,N_22691,N_21822);
nand UO_1040 (O_1040,N_24339,N_20146);
nor UO_1041 (O_1041,N_21262,N_21166);
nor UO_1042 (O_1042,N_21966,N_23108);
xnor UO_1043 (O_1043,N_22021,N_21791);
nand UO_1044 (O_1044,N_20100,N_23740);
and UO_1045 (O_1045,N_23388,N_20247);
and UO_1046 (O_1046,N_21878,N_20512);
nor UO_1047 (O_1047,N_21106,N_21344);
and UO_1048 (O_1048,N_24250,N_21121);
xnor UO_1049 (O_1049,N_20429,N_21943);
or UO_1050 (O_1050,N_22709,N_22971);
or UO_1051 (O_1051,N_24975,N_24640);
nor UO_1052 (O_1052,N_24964,N_24645);
and UO_1053 (O_1053,N_21930,N_24943);
xnor UO_1054 (O_1054,N_22656,N_23468);
nor UO_1055 (O_1055,N_23566,N_23968);
nor UO_1056 (O_1056,N_21881,N_21057);
nor UO_1057 (O_1057,N_21633,N_24480);
and UO_1058 (O_1058,N_23749,N_21321);
nor UO_1059 (O_1059,N_24834,N_22269);
and UO_1060 (O_1060,N_23103,N_22488);
nand UO_1061 (O_1061,N_22032,N_23178);
nor UO_1062 (O_1062,N_22776,N_22549);
xor UO_1063 (O_1063,N_23582,N_20532);
nand UO_1064 (O_1064,N_22786,N_24818);
or UO_1065 (O_1065,N_22263,N_21674);
nand UO_1066 (O_1066,N_23060,N_20818);
nand UO_1067 (O_1067,N_20601,N_22883);
nor UO_1068 (O_1068,N_21693,N_20396);
nor UO_1069 (O_1069,N_20562,N_20975);
nor UO_1070 (O_1070,N_23020,N_24923);
nand UO_1071 (O_1071,N_22949,N_23883);
nor UO_1072 (O_1072,N_20803,N_22576);
xor UO_1073 (O_1073,N_23331,N_23713);
nand UO_1074 (O_1074,N_22705,N_20341);
nor UO_1075 (O_1075,N_23163,N_24610);
nor UO_1076 (O_1076,N_20177,N_24125);
and UO_1077 (O_1077,N_20344,N_20193);
or UO_1078 (O_1078,N_22208,N_21922);
or UO_1079 (O_1079,N_22807,N_21360);
nand UO_1080 (O_1080,N_21854,N_24018);
and UO_1081 (O_1081,N_23829,N_23554);
nor UO_1082 (O_1082,N_22395,N_22234);
or UO_1083 (O_1083,N_22777,N_21846);
xor UO_1084 (O_1084,N_23601,N_21751);
or UO_1085 (O_1085,N_24875,N_21219);
nand UO_1086 (O_1086,N_20330,N_24064);
and UO_1087 (O_1087,N_20914,N_23147);
nor UO_1088 (O_1088,N_22420,N_20604);
nor UO_1089 (O_1089,N_24081,N_22291);
or UO_1090 (O_1090,N_22105,N_20088);
nor UO_1091 (O_1091,N_23342,N_22125);
or UO_1092 (O_1092,N_23021,N_21115);
nor UO_1093 (O_1093,N_24901,N_23823);
and UO_1094 (O_1094,N_21092,N_20548);
or UO_1095 (O_1095,N_23436,N_20475);
and UO_1096 (O_1096,N_23137,N_21949);
and UO_1097 (O_1097,N_21130,N_22262);
or UO_1098 (O_1098,N_23705,N_22805);
and UO_1099 (O_1099,N_24320,N_22773);
nand UO_1100 (O_1100,N_20775,N_24535);
and UO_1101 (O_1101,N_24160,N_20801);
nor UO_1102 (O_1102,N_22755,N_22721);
nor UO_1103 (O_1103,N_20899,N_22382);
and UO_1104 (O_1104,N_24415,N_22345);
or UO_1105 (O_1105,N_20972,N_22719);
nor UO_1106 (O_1106,N_24024,N_20957);
or UO_1107 (O_1107,N_24101,N_22214);
or UO_1108 (O_1108,N_23039,N_24402);
nor UO_1109 (O_1109,N_22758,N_22931);
nand UO_1110 (O_1110,N_23352,N_20662);
xnor UO_1111 (O_1111,N_24717,N_20862);
nor UO_1112 (O_1112,N_22853,N_23881);
nor UO_1113 (O_1113,N_24650,N_20331);
nand UO_1114 (O_1114,N_22148,N_23914);
or UO_1115 (O_1115,N_24580,N_24874);
nor UO_1116 (O_1116,N_22591,N_24177);
or UO_1117 (O_1117,N_20772,N_20333);
nand UO_1118 (O_1118,N_24736,N_22578);
nor UO_1119 (O_1119,N_22132,N_21970);
nand UO_1120 (O_1120,N_24671,N_20258);
nor UO_1121 (O_1121,N_24483,N_24196);
nor UO_1122 (O_1122,N_20038,N_21458);
or UO_1123 (O_1123,N_20984,N_21334);
nor UO_1124 (O_1124,N_22697,N_23877);
nor UO_1125 (O_1125,N_20226,N_22827);
nand UO_1126 (O_1126,N_23868,N_21342);
nor UO_1127 (O_1127,N_22249,N_21180);
nor UO_1128 (O_1128,N_21513,N_23061);
or UO_1129 (O_1129,N_24512,N_23622);
or UO_1130 (O_1130,N_20716,N_20524);
nor UO_1131 (O_1131,N_23576,N_23821);
nor UO_1132 (O_1132,N_22339,N_22093);
nor UO_1133 (O_1133,N_24880,N_23036);
nand UO_1134 (O_1134,N_23412,N_21942);
and UO_1135 (O_1135,N_21559,N_24063);
or UO_1136 (O_1136,N_24870,N_22596);
or UO_1137 (O_1137,N_21163,N_24667);
xor UO_1138 (O_1138,N_24701,N_23186);
nor UO_1139 (O_1139,N_21890,N_22963);
nand UO_1140 (O_1140,N_21906,N_23399);
nand UO_1141 (O_1141,N_21945,N_22898);
and UO_1142 (O_1142,N_23799,N_23818);
or UO_1143 (O_1143,N_24714,N_22009);
or UO_1144 (O_1144,N_20308,N_23544);
nor UO_1145 (O_1145,N_23624,N_21938);
nor UO_1146 (O_1146,N_24825,N_23956);
xnor UO_1147 (O_1147,N_20405,N_23444);
or UO_1148 (O_1148,N_20207,N_20568);
or UO_1149 (O_1149,N_23015,N_20784);
and UO_1150 (O_1150,N_24649,N_22496);
nand UO_1151 (O_1151,N_21279,N_23663);
nand UO_1152 (O_1152,N_23967,N_20178);
or UO_1153 (O_1153,N_24658,N_24967);
and UO_1154 (O_1154,N_20283,N_20570);
and UO_1155 (O_1155,N_22368,N_24257);
and UO_1156 (O_1156,N_22014,N_22960);
nor UO_1157 (O_1157,N_24086,N_21611);
and UO_1158 (O_1158,N_20159,N_20240);
nand UO_1159 (O_1159,N_22296,N_23062);
xnor UO_1160 (O_1160,N_20044,N_22845);
nor UO_1161 (O_1161,N_20378,N_21834);
nor UO_1162 (O_1162,N_24374,N_20737);
nand UO_1163 (O_1163,N_21088,N_23882);
nor UO_1164 (O_1164,N_23464,N_21859);
xnor UO_1165 (O_1165,N_20834,N_22895);
nor UO_1166 (O_1166,N_21635,N_22254);
or UO_1167 (O_1167,N_20852,N_24600);
nand UO_1168 (O_1168,N_23440,N_24075);
and UO_1169 (O_1169,N_20659,N_22188);
nand UO_1170 (O_1170,N_22206,N_24422);
nand UO_1171 (O_1171,N_21754,N_20250);
and UO_1172 (O_1172,N_20944,N_22255);
nor UO_1173 (O_1173,N_21085,N_20991);
nor UO_1174 (O_1174,N_23732,N_22886);
nor UO_1175 (O_1175,N_24657,N_20307);
and UO_1176 (O_1176,N_23184,N_21845);
xnor UO_1177 (O_1177,N_21404,N_22698);
or UO_1178 (O_1178,N_20265,N_22281);
and UO_1179 (O_1179,N_21433,N_20089);
nor UO_1180 (O_1180,N_24390,N_20771);
xnor UO_1181 (O_1181,N_20916,N_24969);
xnor UO_1182 (O_1182,N_20315,N_20172);
nor UO_1183 (O_1183,N_21239,N_24025);
nand UO_1184 (O_1184,N_22524,N_20227);
and UO_1185 (O_1185,N_24313,N_22744);
or UO_1186 (O_1186,N_20370,N_24455);
xnor UO_1187 (O_1187,N_22359,N_22801);
nand UO_1188 (O_1188,N_22546,N_20482);
nor UO_1189 (O_1189,N_23488,N_24690);
nor UO_1190 (O_1190,N_20235,N_21487);
nand UO_1191 (O_1191,N_24317,N_23302);
and UO_1192 (O_1192,N_23357,N_20224);
nor UO_1193 (O_1193,N_23623,N_20037);
nor UO_1194 (O_1194,N_24688,N_21539);
or UO_1195 (O_1195,N_20786,N_20324);
and UO_1196 (O_1196,N_21155,N_23947);
nor UO_1197 (O_1197,N_23827,N_20668);
nand UO_1198 (O_1198,N_21309,N_23306);
nand UO_1199 (O_1199,N_21053,N_23686);
or UO_1200 (O_1200,N_23360,N_22078);
or UO_1201 (O_1201,N_22244,N_23727);
or UO_1202 (O_1202,N_22739,N_24210);
or UO_1203 (O_1203,N_20060,N_24425);
or UO_1204 (O_1204,N_20542,N_21592);
nor UO_1205 (O_1205,N_22779,N_23631);
xor UO_1206 (O_1206,N_20270,N_21981);
or UO_1207 (O_1207,N_24166,N_20141);
and UO_1208 (O_1208,N_24949,N_22270);
xor UO_1209 (O_1209,N_23620,N_24767);
and UO_1210 (O_1210,N_20230,N_23431);
nand UO_1211 (O_1211,N_22662,N_24787);
or UO_1212 (O_1212,N_24981,N_21290);
nor UO_1213 (O_1213,N_24558,N_20929);
or UO_1214 (O_1214,N_20077,N_20638);
nor UO_1215 (O_1215,N_20200,N_23437);
nand UO_1216 (O_1216,N_22070,N_22159);
nor UO_1217 (O_1217,N_22171,N_21097);
xor UO_1218 (O_1218,N_22572,N_21307);
or UO_1219 (O_1219,N_20563,N_22424);
and UO_1220 (O_1220,N_21326,N_24149);
and UO_1221 (O_1221,N_20704,N_23747);
nand UO_1222 (O_1222,N_21686,N_24372);
and UO_1223 (O_1223,N_22774,N_24795);
and UO_1224 (O_1224,N_22593,N_23398);
or UO_1225 (O_1225,N_24692,N_23126);
xor UO_1226 (O_1226,N_20539,N_20773);
nor UO_1227 (O_1227,N_23223,N_21749);
and UO_1228 (O_1228,N_23513,N_20725);
or UO_1229 (O_1229,N_20564,N_24491);
or UO_1230 (O_1230,N_20111,N_23351);
nand UO_1231 (O_1231,N_20253,N_23425);
and UO_1232 (O_1232,N_20430,N_20402);
nor UO_1233 (O_1233,N_22925,N_21927);
or UO_1234 (O_1234,N_23013,N_23805);
nand UO_1235 (O_1235,N_20215,N_20642);
nor UO_1236 (O_1236,N_20052,N_21037);
and UO_1237 (O_1237,N_24182,N_24547);
or UO_1238 (O_1238,N_24984,N_22177);
nand UO_1239 (O_1239,N_23649,N_23621);
nand UO_1240 (O_1240,N_20966,N_21196);
and UO_1241 (O_1241,N_22599,N_22696);
nor UO_1242 (O_1242,N_21476,N_21553);
and UO_1243 (O_1243,N_22307,N_21260);
nand UO_1244 (O_1244,N_21197,N_20888);
nor UO_1245 (O_1245,N_24924,N_21535);
and UO_1246 (O_1246,N_23848,N_24050);
nand UO_1247 (O_1247,N_21347,N_23815);
nor UO_1248 (O_1248,N_21928,N_23026);
xnor UO_1249 (O_1249,N_22695,N_23931);
or UO_1250 (O_1250,N_21940,N_21698);
xor UO_1251 (O_1251,N_23355,N_20721);
nand UO_1252 (O_1252,N_21150,N_21276);
and UO_1253 (O_1253,N_23735,N_24540);
and UO_1254 (O_1254,N_21971,N_21089);
nor UO_1255 (O_1255,N_22052,N_21039);
nor UO_1256 (O_1256,N_20860,N_24328);
and UO_1257 (O_1257,N_24993,N_21373);
and UO_1258 (O_1258,N_20754,N_22138);
and UO_1259 (O_1259,N_20906,N_24815);
xor UO_1260 (O_1260,N_20813,N_23337);
or UO_1261 (O_1261,N_22651,N_23141);
nor UO_1262 (O_1262,N_23678,N_23970);
and UO_1263 (O_1263,N_22820,N_23736);
and UO_1264 (O_1264,N_24956,N_21070);
xor UO_1265 (O_1265,N_23275,N_23770);
nor UO_1266 (O_1266,N_21625,N_22403);
or UO_1267 (O_1267,N_24927,N_23100);
and UO_1268 (O_1268,N_22071,N_23040);
or UO_1269 (O_1269,N_20705,N_21005);
nor UO_1270 (O_1270,N_24042,N_22219);
or UO_1271 (O_1271,N_21291,N_22090);
or UO_1272 (O_1272,N_24061,N_20357);
and UO_1273 (O_1273,N_24341,N_24035);
and UO_1274 (O_1274,N_23449,N_24082);
nand UO_1275 (O_1275,N_24488,N_24539);
or UO_1276 (O_1276,N_23890,N_21634);
nand UO_1277 (O_1277,N_24778,N_21116);
and UO_1278 (O_1278,N_21977,N_24822);
and UO_1279 (O_1279,N_21980,N_23059);
or UO_1280 (O_1280,N_22407,N_23922);
nor UO_1281 (O_1281,N_21463,N_23466);
or UO_1282 (O_1282,N_21500,N_21008);
nor UO_1283 (O_1283,N_22282,N_23017);
nand UO_1284 (O_1284,N_23086,N_22563);
nand UO_1285 (O_1285,N_21804,N_24999);
xor UO_1286 (O_1286,N_21696,N_21899);
nand UO_1287 (O_1287,N_24934,N_20053);
or UO_1288 (O_1288,N_24651,N_24509);
or UO_1289 (O_1289,N_20248,N_24750);
nor UO_1290 (O_1290,N_20951,N_22816);
or UO_1291 (O_1291,N_21178,N_21182);
nor UO_1292 (O_1292,N_23838,N_22929);
nor UO_1293 (O_1293,N_22485,N_22041);
and UO_1294 (O_1294,N_22480,N_20735);
nand UO_1295 (O_1295,N_23958,N_21503);
or UO_1296 (O_1296,N_23169,N_24109);
and UO_1297 (O_1297,N_21159,N_22454);
nand UO_1298 (O_1298,N_24074,N_21785);
nand UO_1299 (O_1299,N_21493,N_22693);
nor UO_1300 (O_1300,N_24409,N_21234);
xnor UO_1301 (O_1301,N_20521,N_24104);
nor UO_1302 (O_1302,N_24205,N_22737);
or UO_1303 (O_1303,N_22837,N_23521);
nor UO_1304 (O_1304,N_21058,N_21887);
or UO_1305 (O_1305,N_24080,N_24850);
nor UO_1306 (O_1306,N_22913,N_22723);
and UO_1307 (O_1307,N_22458,N_21857);
or UO_1308 (O_1308,N_23288,N_22444);
xnor UO_1309 (O_1309,N_24129,N_24278);
xor UO_1310 (O_1310,N_22465,N_23159);
or UO_1311 (O_1311,N_20085,N_22233);
and UO_1312 (O_1312,N_20880,N_21589);
nor UO_1313 (O_1313,N_20511,N_24158);
and UO_1314 (O_1314,N_22813,N_24314);
and UO_1315 (O_1315,N_23545,N_23383);
or UO_1316 (O_1316,N_20102,N_24335);
nor UO_1317 (O_1317,N_22352,N_24270);
xor UO_1318 (O_1318,N_24220,N_21304);
nand UO_1319 (O_1319,N_22901,N_24251);
or UO_1320 (O_1320,N_23002,N_22049);
and UO_1321 (O_1321,N_22089,N_20728);
and UO_1322 (O_1322,N_22129,N_24807);
and UO_1323 (O_1323,N_23792,N_23560);
and UO_1324 (O_1324,N_24093,N_21474);
nand UO_1325 (O_1325,N_22633,N_23432);
nor UO_1326 (O_1326,N_20947,N_22316);
nor UO_1327 (O_1327,N_23349,N_24356);
or UO_1328 (O_1328,N_24060,N_23505);
nand UO_1329 (O_1329,N_21430,N_23093);
nor UO_1330 (O_1330,N_20300,N_20602);
nor UO_1331 (O_1331,N_24334,N_24666);
and UO_1332 (O_1332,N_20216,N_21128);
or UO_1333 (O_1333,N_20225,N_22435);
nor UO_1334 (O_1334,N_20176,N_22731);
nand UO_1335 (O_1335,N_23871,N_20670);
nor UO_1336 (O_1336,N_21774,N_20241);
nor UO_1337 (O_1337,N_24092,N_21074);
and UO_1338 (O_1338,N_22742,N_21912);
or UO_1339 (O_1339,N_21619,N_23190);
and UO_1340 (O_1340,N_21447,N_20028);
or UO_1341 (O_1341,N_21793,N_24071);
nand UO_1342 (O_1342,N_23416,N_23210);
or UO_1343 (O_1343,N_22116,N_21320);
nor UO_1344 (O_1344,N_20930,N_24289);
and UO_1345 (O_1345,N_24421,N_23909);
and UO_1346 (O_1346,N_20760,N_24588);
xnor UO_1347 (O_1347,N_20531,N_21272);
nor UO_1348 (O_1348,N_22383,N_20612);
xor UO_1349 (O_1349,N_22111,N_21984);
and UO_1350 (O_1350,N_21677,N_23363);
and UO_1351 (O_1351,N_22787,N_21864);
nor UO_1352 (O_1352,N_20968,N_24953);
and UO_1353 (O_1353,N_20561,N_20078);
or UO_1354 (O_1354,N_20158,N_20428);
xor UO_1355 (O_1355,N_21415,N_21832);
nand UO_1356 (O_1356,N_22864,N_21547);
nor UO_1357 (O_1357,N_23202,N_24255);
nand UO_1358 (O_1358,N_22541,N_20517);
xnor UO_1359 (O_1359,N_21903,N_24398);
xnor UO_1360 (O_1360,N_21423,N_20129);
xnor UO_1361 (O_1361,N_22081,N_22621);
nand UO_1362 (O_1362,N_23403,N_21110);
nand UO_1363 (O_1363,N_24814,N_24216);
nand UO_1364 (O_1364,N_23439,N_22630);
nand UO_1365 (O_1365,N_23106,N_23152);
nor UO_1366 (O_1366,N_24261,N_21318);
xor UO_1367 (O_1367,N_21161,N_23079);
xor UO_1368 (O_1368,N_24053,N_21288);
nand UO_1369 (O_1369,N_22086,N_22023);
or UO_1370 (O_1370,N_22906,N_21481);
and UO_1371 (O_1371,N_24420,N_22915);
or UO_1372 (O_1372,N_21606,N_22534);
xnor UO_1373 (O_1373,N_24684,N_21504);
xor UO_1374 (O_1374,N_23209,N_20639);
or UO_1375 (O_1375,N_21551,N_20961);
nand UO_1376 (O_1376,N_23161,N_20237);
or UO_1377 (O_1377,N_20993,N_21353);
and UO_1378 (O_1378,N_23442,N_20866);
and UO_1379 (O_1379,N_21590,N_20259);
or UO_1380 (O_1380,N_24589,N_20399);
nand UO_1381 (O_1381,N_22799,N_22903);
and UO_1382 (O_1382,N_24260,N_24392);
nor UO_1383 (O_1383,N_23532,N_20729);
or UO_1384 (O_1384,N_24996,N_24327);
or UO_1385 (O_1385,N_21437,N_21009);
nand UO_1386 (O_1386,N_22533,N_20779);
or UO_1387 (O_1387,N_21576,N_21226);
nand UO_1388 (O_1388,N_24643,N_24148);
nand UO_1389 (O_1389,N_21967,N_24636);
and UO_1390 (O_1390,N_23901,N_22273);
nand UO_1391 (O_1391,N_24179,N_20603);
or UO_1392 (O_1392,N_24499,N_23862);
and UO_1393 (O_1393,N_24408,N_24804);
nand UO_1394 (O_1394,N_24856,N_21824);
or UO_1395 (O_1395,N_20583,N_20555);
and UO_1396 (O_1396,N_22802,N_23693);
nor UO_1397 (O_1397,N_24573,N_20605);
or UO_1398 (O_1398,N_21925,N_20066);
nor UO_1399 (O_1399,N_20014,N_20687);
and UO_1400 (O_1400,N_20105,N_24819);
and UO_1401 (O_1401,N_24233,N_21087);
nor UO_1402 (O_1402,N_22146,N_21035);
nand UO_1403 (O_1403,N_20057,N_21094);
xor UO_1404 (O_1404,N_22733,N_21678);
and UO_1405 (O_1405,N_20214,N_24859);
nor UO_1406 (O_1406,N_21126,N_24417);
nand UO_1407 (O_1407,N_21124,N_23140);
nor UO_1408 (O_1408,N_21018,N_21960);
nor UO_1409 (O_1409,N_24235,N_22503);
and UO_1410 (O_1410,N_22418,N_20645);
xor UO_1411 (O_1411,N_21335,N_21862);
and UO_1412 (O_1412,N_23310,N_22582);
xor UO_1413 (O_1413,N_21274,N_20238);
nand UO_1414 (O_1414,N_20677,N_20443);
and UO_1415 (O_1415,N_24111,N_23120);
xnor UO_1416 (O_1416,N_20858,N_24760);
nor UO_1417 (O_1417,N_24816,N_22771);
or UO_1418 (O_1418,N_24110,N_21338);
xor UO_1419 (O_1419,N_21621,N_20731);
nor UO_1420 (O_1420,N_23866,N_22389);
xor UO_1421 (O_1421,N_20423,N_22216);
xnor UO_1422 (O_1422,N_20855,N_21740);
and UO_1423 (O_1423,N_24563,N_20099);
or UO_1424 (O_1424,N_22685,N_20935);
xnor UO_1425 (O_1425,N_20311,N_23569);
xor UO_1426 (O_1426,N_20377,N_21670);
or UO_1427 (O_1427,N_21357,N_20025);
nand UO_1428 (O_1428,N_24511,N_21983);
and UO_1429 (O_1429,N_20733,N_22748);
nand UO_1430 (O_1430,N_20096,N_24352);
nor UO_1431 (O_1431,N_24412,N_22140);
nand UO_1432 (O_1432,N_22991,N_23771);
xnor UO_1433 (O_1433,N_24399,N_20776);
nand UO_1434 (O_1434,N_20273,N_20682);
nor UO_1435 (O_1435,N_23646,N_24442);
and UO_1436 (O_1436,N_21250,N_24603);
nor UO_1437 (O_1437,N_20064,N_22678);
nand UO_1438 (O_1438,N_21172,N_20960);
or UO_1439 (O_1439,N_22661,N_21777);
and UO_1440 (O_1440,N_20973,N_24371);
or UO_1441 (O_1441,N_21002,N_22610);
nand UO_1442 (O_1442,N_24613,N_24295);
nand UO_1443 (O_1443,N_24432,N_23181);
nand UO_1444 (O_1444,N_24277,N_22110);
and UO_1445 (O_1445,N_21134,N_23895);
and UO_1446 (O_1446,N_21776,N_22312);
or UO_1447 (O_1447,N_23404,N_23548);
or UO_1448 (O_1448,N_23558,N_21071);
nand UO_1449 (O_1449,N_23608,N_20431);
or UO_1450 (O_1450,N_24316,N_20294);
and UO_1451 (O_1451,N_23405,N_20508);
and UO_1452 (O_1452,N_22285,N_20395);
nor UO_1453 (O_1453,N_21286,N_24186);
or UO_1454 (O_1454,N_21614,N_20640);
nor UO_1455 (O_1455,N_23841,N_20109);
or UO_1456 (O_1456,N_22889,N_24471);
or UO_1457 (O_1457,N_20397,N_24238);
nor UO_1458 (O_1458,N_22935,N_20367);
nor UO_1459 (O_1459,N_20040,N_21524);
or UO_1460 (O_1460,N_24054,N_21916);
or UO_1461 (O_1461,N_20012,N_23976);
xnor UO_1462 (O_1462,N_20648,N_21190);
xor UO_1463 (O_1463,N_23290,N_22921);
and UO_1464 (O_1464,N_20822,N_20694);
nor UO_1465 (O_1465,N_23372,N_22290);
or UO_1466 (O_1466,N_22199,N_21583);
nor UO_1467 (O_1467,N_22253,N_20654);
xor UO_1468 (O_1468,N_24292,N_20277);
nor UO_1469 (O_1469,N_21972,N_23759);
and UO_1470 (O_1470,N_23248,N_20362);
or UO_1471 (O_1471,N_23514,N_20149);
or UO_1472 (O_1472,N_21676,N_20068);
and UO_1473 (O_1473,N_20087,N_24016);
or UO_1474 (O_1474,N_20881,N_22131);
xnor UO_1475 (O_1475,N_23707,N_20526);
nand UO_1476 (O_1476,N_21682,N_21169);
nor UO_1477 (O_1477,N_24931,N_20352);
nand UO_1478 (O_1478,N_24776,N_24450);
and UO_1479 (O_1479,N_21612,N_22330);
and UO_1480 (O_1480,N_23538,N_24955);
or UO_1481 (O_1481,N_21704,N_23864);
nor UO_1482 (O_1482,N_21811,N_24652);
or UO_1483 (O_1483,N_22028,N_22453);
or UO_1484 (O_1484,N_24367,N_20870);
and UO_1485 (O_1485,N_24882,N_20674);
nand UO_1486 (O_1486,N_23203,N_23777);
nand UO_1487 (O_1487,N_21093,N_24204);
nor UO_1488 (O_1488,N_22641,N_24452);
and UO_1489 (O_1489,N_20833,N_23831);
and UO_1490 (O_1490,N_21736,N_22570);
and UO_1491 (O_1491,N_23254,N_23133);
xor UO_1492 (O_1492,N_20107,N_21667);
xnor UO_1493 (O_1493,N_21745,N_21712);
xor UO_1494 (O_1494,N_20420,N_23597);
or UO_1495 (O_1495,N_22505,N_20835);
and UO_1496 (O_1496,N_21453,N_24598);
nor UO_1497 (O_1497,N_23666,N_21976);
nand UO_1498 (O_1498,N_23998,N_20676);
nand UO_1499 (O_1499,N_23095,N_22058);
nor UO_1500 (O_1500,N_24616,N_23639);
and UO_1501 (O_1501,N_24360,N_23165);
nand UO_1502 (O_1502,N_21767,N_24865);
and UO_1503 (O_1503,N_22635,N_21048);
or UO_1504 (O_1504,N_23894,N_23070);
nand UO_1505 (O_1505,N_24032,N_22632);
xor UO_1506 (O_1506,N_21618,N_22756);
nand UO_1507 (O_1507,N_21624,N_22987);
nor UO_1508 (O_1508,N_23662,N_22609);
nand UO_1509 (O_1509,N_20636,N_22261);
nand UO_1510 (O_1510,N_20761,N_24217);
or UO_1511 (O_1511,N_22142,N_22491);
or UO_1512 (O_1512,N_22275,N_20046);
or UO_1513 (O_1513,N_22784,N_23170);
nand UO_1514 (O_1514,N_23796,N_23986);
or UO_1515 (O_1515,N_23773,N_21300);
and UO_1516 (O_1516,N_21242,N_21979);
nand UO_1517 (O_1517,N_23611,N_23945);
nor UO_1518 (O_1518,N_23982,N_24459);
nor UO_1519 (O_1519,N_24501,N_21868);
or UO_1520 (O_1520,N_23219,N_24323);
nand UO_1521 (O_1521,N_22878,N_21305);
nand UO_1522 (O_1522,N_20909,N_23114);
or UO_1523 (O_1523,N_20928,N_23339);
nand UO_1524 (O_1524,N_20625,N_24638);
and UO_1525 (O_1525,N_21266,N_24683);
xor UO_1526 (O_1526,N_20441,N_24662);
nor UO_1527 (O_1527,N_24845,N_21281);
nor UO_1528 (O_1528,N_20479,N_24641);
or UO_1529 (O_1529,N_24644,N_24279);
xor UO_1530 (O_1530,N_20533,N_24887);
or UO_1531 (O_1531,N_22391,N_23651);
nand UO_1532 (O_1532,N_20753,N_21456);
nor UO_1533 (O_1533,N_21729,N_23085);
nand UO_1534 (O_1534,N_21651,N_23121);
xor UO_1535 (O_1535,N_20271,N_20826);
or UO_1536 (O_1536,N_22157,N_24672);
or UO_1537 (O_1537,N_24682,N_24915);
and UO_1538 (O_1538,N_22562,N_20494);
nor UO_1539 (O_1539,N_22939,N_23495);
or UO_1540 (O_1540,N_21241,N_23640);
and UO_1541 (O_1541,N_24948,N_22167);
or UO_1542 (O_1542,N_22959,N_21200);
xnor UO_1543 (O_1543,N_21929,N_23580);
xor UO_1544 (O_1544,N_23069,N_22074);
nand UO_1545 (O_1545,N_23535,N_24835);
nand UO_1546 (O_1546,N_20534,N_22055);
and UO_1547 (O_1547,N_20314,N_21615);
or UO_1548 (O_1548,N_20144,N_20643);
and UO_1549 (O_1549,N_21310,N_20811);
nand UO_1550 (O_1550,N_20864,N_20312);
or UO_1551 (O_1551,N_22091,N_21230);
and UO_1552 (O_1552,N_20426,N_22724);
or UO_1553 (O_1553,N_23641,N_24138);
and UO_1554 (O_1554,N_23066,N_22085);
nor UO_1555 (O_1555,N_23090,N_20162);
and UO_1556 (O_1556,N_23277,N_23491);
nor UO_1557 (O_1557,N_24546,N_20050);
and UO_1558 (O_1558,N_23081,N_20249);
or UO_1559 (O_1559,N_22139,N_20366);
or UO_1560 (O_1560,N_24700,N_20574);
or UO_1561 (O_1561,N_24474,N_24691);
nand UO_1562 (O_1562,N_21772,N_23207);
nand UO_1563 (O_1563,N_24609,N_21873);
nor UO_1564 (O_1564,N_22034,N_23579);
nor UO_1565 (O_1565,N_21478,N_23703);
nor UO_1566 (O_1566,N_24624,N_22195);
and UO_1567 (O_1567,N_20490,N_20519);
or UO_1568 (O_1568,N_24117,N_21935);
nor UO_1569 (O_1569,N_23281,N_21690);
or UO_1570 (O_1570,N_24883,N_20364);
nor UO_1571 (O_1571,N_24045,N_24245);
nor UO_1572 (O_1572,N_22415,N_22393);
or UO_1573 (O_1573,N_24269,N_24141);
and UO_1574 (O_1574,N_20816,N_20635);
or UO_1575 (O_1575,N_24553,N_22550);
or UO_1576 (O_1576,N_23628,N_23238);
nand UO_1577 (O_1577,N_21584,N_20987);
or UO_1578 (O_1578,N_24958,N_22859);
nor UO_1579 (O_1579,N_23921,N_23991);
nand UO_1580 (O_1580,N_20454,N_22754);
nor UO_1581 (O_1581,N_24800,N_21921);
and UO_1582 (O_1582,N_21988,N_23985);
nor UO_1583 (O_1583,N_20192,N_20955);
or UO_1584 (O_1584,N_22979,N_24832);
or UO_1585 (O_1585,N_22398,N_21716);
or UO_1586 (O_1586,N_24057,N_23565);
or UO_1587 (O_1587,N_23473,N_20890);
nand UO_1588 (O_1588,N_23837,N_22728);
and UO_1589 (O_1589,N_21962,N_23567);
nor UO_1590 (O_1590,N_20506,N_24348);
xnor UO_1591 (O_1591,N_22995,N_21561);
nand UO_1592 (O_1592,N_24013,N_20744);
or UO_1593 (O_1593,N_23156,N_21875);
and UO_1594 (O_1594,N_22447,N_23832);
xor UO_1595 (O_1595,N_22507,N_21168);
and UO_1596 (O_1596,N_20470,N_22617);
or UO_1597 (O_1597,N_24493,N_24159);
nand UO_1598 (O_1598,N_24463,N_24555);
and UO_1599 (O_1599,N_23928,N_24106);
nor UO_1600 (O_1600,N_20621,N_20244);
nand UO_1601 (O_1601,N_23644,N_21177);
nor UO_1602 (O_1602,N_21043,N_24051);
xor UO_1603 (O_1603,N_21044,N_21679);
and UO_1604 (O_1604,N_21068,N_21781);
and UO_1605 (O_1605,N_24291,N_24236);
and UO_1606 (O_1606,N_21377,N_24359);
nor UO_1607 (O_1607,N_21042,N_20297);
xnor UO_1608 (O_1608,N_20732,N_20751);
and UO_1609 (O_1609,N_21452,N_21011);
nor UO_1610 (O_1610,N_22150,N_21532);
or UO_1611 (O_1611,N_23049,N_22857);
nand UO_1612 (O_1612,N_20849,N_20878);
and UO_1613 (O_1613,N_21184,N_22810);
or UO_1614 (O_1614,N_24889,N_22592);
nand UO_1615 (O_1615,N_20326,N_23903);
and UO_1616 (O_1616,N_22015,N_20610);
and UO_1617 (O_1617,N_23486,N_20876);
nand UO_1618 (O_1618,N_21396,N_20697);
nor UO_1619 (O_1619,N_22422,N_22439);
nand UO_1620 (O_1620,N_20290,N_23139);
nand UO_1621 (O_1621,N_24785,N_22618);
nor UO_1622 (O_1622,N_20480,N_22082);
nand UO_1623 (O_1623,N_21198,N_23869);
or UO_1624 (O_1624,N_23711,N_20885);
and UO_1625 (O_1625,N_23604,N_22658);
and UO_1626 (O_1626,N_24577,N_20549);
or UO_1627 (O_1627,N_22828,N_20218);
or UO_1628 (O_1628,N_23800,N_20461);
or UO_1629 (O_1629,N_21237,N_20301);
nor UO_1630 (O_1630,N_22585,N_22916);
nand UO_1631 (O_1631,N_24254,N_21225);
and UO_1632 (O_1632,N_22712,N_20007);
xnor UO_1633 (O_1633,N_22808,N_22616);
nor UO_1634 (O_1634,N_22000,N_21386);
nand UO_1635 (O_1635,N_20071,N_20626);
and UO_1636 (O_1636,N_24310,N_23487);
nand UO_1637 (O_1637,N_21444,N_22026);
nand UO_1638 (O_1638,N_23801,N_22856);
nor UO_1639 (O_1639,N_20320,N_21355);
and UO_1640 (O_1640,N_23037,N_24258);
nor UO_1641 (O_1641,N_21605,N_22243);
nand UO_1642 (O_1642,N_22191,N_21817);
xnor UO_1643 (O_1643,N_23710,N_24311);
nor UO_1644 (O_1644,N_23996,N_21527);
and UO_1645 (O_1645,N_23898,N_23144);
xnor UO_1646 (O_1646,N_22527,N_21908);
nor UO_1647 (O_1647,N_24346,N_21482);
and UO_1648 (O_1648,N_20879,N_23010);
nand UO_1649 (O_1649,N_22811,N_20931);
nand UO_1650 (O_1650,N_24622,N_20365);
nor UO_1651 (O_1651,N_23409,N_22051);
or UO_1652 (O_1652,N_22569,N_24396);
nand UO_1653 (O_1653,N_23738,N_24852);
or UO_1654 (O_1654,N_20090,N_20039);
nor UO_1655 (O_1655,N_20644,N_22667);
or UO_1656 (O_1656,N_22869,N_23946);
and UO_1657 (O_1657,N_22374,N_21528);
and UO_1658 (O_1658,N_21419,N_22010);
nand UO_1659 (O_1659,N_23661,N_24049);
nand UO_1660 (O_1660,N_20777,N_20421);
xor UO_1661 (O_1661,N_20002,N_23009);
xnor UO_1662 (O_1662,N_22940,N_23279);
nand UO_1663 (O_1663,N_20828,N_24207);
xnor UO_1664 (O_1664,N_24522,N_21137);
nand UO_1665 (O_1665,N_23325,N_24330);
nor UO_1666 (O_1666,N_20342,N_24974);
nand UO_1667 (O_1667,N_23694,N_22318);
and UO_1668 (O_1668,N_21170,N_22876);
and UO_1669 (O_1669,N_23746,N_24792);
xnor UO_1670 (O_1670,N_20980,N_20658);
or UO_1671 (O_1671,N_23803,N_23258);
nand UO_1672 (O_1672,N_23232,N_24921);
and UO_1673 (O_1673,N_20017,N_22511);
nand UO_1674 (O_1674,N_20770,N_22614);
nand UO_1675 (O_1675,N_20491,N_20530);
or UO_1676 (O_1676,N_23943,N_20264);
nor UO_1677 (O_1677,N_21468,N_24006);
and UO_1678 (O_1678,N_23052,N_23787);
nand UO_1679 (O_1679,N_21328,N_21877);
nor UO_1680 (O_1680,N_22765,N_23999);
or UO_1681 (O_1681,N_23458,N_20191);
and UO_1682 (O_1682,N_23756,N_20727);
nor UO_1683 (O_1683,N_20234,N_21189);
or UO_1684 (O_1684,N_23865,N_23744);
nor UO_1685 (O_1685,N_24286,N_21066);
or UO_1686 (O_1686,N_22095,N_21762);
nand UO_1687 (O_1687,N_22059,N_21773);
nor UO_1688 (O_1688,N_22664,N_23119);
and UO_1689 (O_1689,N_21052,N_22682);
nand UO_1690 (O_1690,N_23297,N_24127);
xor UO_1691 (O_1691,N_21963,N_20934);
nor UO_1692 (O_1692,N_23217,N_23461);
nand UO_1693 (O_1693,N_24112,N_21294);
nor UO_1694 (O_1694,N_22770,N_21578);
nor UO_1695 (O_1695,N_22120,N_22790);
and UO_1696 (O_1696,N_24487,N_20582);
nor UO_1697 (O_1697,N_20698,N_21175);
nor UO_1698 (O_1698,N_21883,N_24768);
nor UO_1699 (O_1699,N_24468,N_22956);
and UO_1700 (O_1700,N_23230,N_24991);
nor UO_1701 (O_1701,N_23627,N_20702);
and UO_1702 (O_1702,N_24548,N_24902);
xor UO_1703 (O_1703,N_23860,N_20387);
or UO_1704 (O_1704,N_23767,N_22030);
nand UO_1705 (O_1705,N_20132,N_24656);
nand UO_1706 (O_1706,N_22819,N_23364);
and UO_1707 (O_1707,N_23055,N_21171);
or UO_1708 (O_1708,N_21424,N_22141);
nand UO_1709 (O_1709,N_23699,N_22726);
nand UO_1710 (O_1710,N_22311,N_21421);
nor UO_1711 (O_1711,N_24810,N_24854);
nor UO_1712 (O_1712,N_22702,N_20580);
and UO_1713 (O_1713,N_22184,N_24730);
xnor UO_1714 (O_1714,N_22653,N_22943);
xnor UO_1715 (O_1715,N_21435,N_22855);
nor UO_1716 (O_1716,N_23962,N_23760);
or UO_1717 (O_1717,N_23504,N_22752);
xnor UO_1718 (O_1718,N_22904,N_22185);
nor UO_1719 (O_1719,N_22663,N_23817);
nor UO_1720 (O_1720,N_22222,N_22160);
nand UO_1721 (O_1721,N_24451,N_23512);
nand UO_1722 (O_1722,N_20940,N_24091);
and UO_1723 (O_1723,N_23145,N_24288);
nor UO_1724 (O_1724,N_23263,N_20293);
or UO_1725 (O_1725,N_20232,N_24904);
or UO_1726 (O_1726,N_21432,N_24140);
xor UO_1727 (O_1727,N_23913,N_22227);
nor UO_1728 (O_1728,N_20617,N_23577);
xnor UO_1729 (O_1729,N_21231,N_22354);
nor UO_1730 (O_1730,N_23319,N_24026);
or UO_1731 (O_1731,N_24520,N_24381);
nand UO_1732 (O_1732,N_23757,N_21713);
or UO_1733 (O_1733,N_20590,N_21936);
nand UO_1734 (O_1734,N_23080,N_21113);
or UO_1735 (O_1735,N_24342,N_23936);
nor UO_1736 (O_1736,N_21759,N_22643);
or UO_1737 (O_1737,N_24118,N_24454);
nor UO_1738 (O_1738,N_24696,N_21164);
and UO_1739 (O_1739,N_24900,N_21167);
nor UO_1740 (O_1740,N_23745,N_21880);
or UO_1741 (O_1741,N_24010,N_23193);
or UO_1742 (O_1742,N_22821,N_20510);
and UO_1743 (O_1743,N_23924,N_23630);
nand UO_1744 (O_1744,N_20213,N_21844);
nand UO_1745 (O_1745,N_23007,N_23194);
or UO_1746 (O_1746,N_23438,N_23134);
and UO_1747 (O_1747,N_21863,N_21526);
nor UO_1748 (O_1748,N_22781,N_20056);
nor UO_1749 (O_1749,N_23944,N_23381);
nor UO_1750 (O_1750,N_21946,N_21133);
or UO_1751 (O_1751,N_20275,N_20042);
or UO_1752 (O_1752,N_24237,N_22775);
nand UO_1753 (O_1753,N_21477,N_21546);
or UO_1754 (O_1754,N_24790,N_22287);
nand UO_1755 (O_1755,N_22308,N_24202);
and UO_1756 (O_1756,N_20938,N_23110);
nand UO_1757 (O_1757,N_24674,N_20871);
xnor UO_1758 (O_1758,N_20031,N_20285);
and UO_1759 (O_1759,N_23025,N_24184);
and UO_1760 (O_1760,N_21782,N_20600);
xor UO_1761 (O_1761,N_21701,N_21220);
or UO_1762 (O_1762,N_21192,N_22460);
nor UO_1763 (O_1763,N_23555,N_22717);
nor UO_1764 (O_1764,N_20292,N_22012);
or UO_1765 (O_1765,N_24214,N_21312);
nor UO_1766 (O_1766,N_21145,N_21162);
nand UO_1767 (O_1767,N_23038,N_20766);
and UO_1768 (O_1768,N_24628,N_22336);
or UO_1769 (O_1769,N_24206,N_22161);
and UO_1770 (O_1770,N_24566,N_21475);
nand UO_1771 (O_1771,N_23954,N_23016);
nand UO_1772 (O_1772,N_24575,N_22814);
nand UO_1773 (O_1773,N_21313,N_22594);
and UO_1774 (O_1774,N_21140,N_20190);
nand UO_1775 (O_1775,N_20979,N_24152);
and UO_1776 (O_1776,N_20000,N_22950);
nand UO_1777 (O_1777,N_21268,N_24777);
or UO_1778 (O_1778,N_20419,N_24962);
or UO_1779 (O_1779,N_20488,N_22812);
or UO_1780 (O_1780,N_23361,N_22558);
or UO_1781 (O_1781,N_21636,N_20209);
nor UO_1782 (O_1782,N_22247,N_21306);
or UO_1783 (O_1783,N_22953,N_20246);
nand UO_1784 (O_1784,N_22849,N_22689);
and UO_1785 (O_1785,N_20948,N_23415);
nand UO_1786 (O_1786,N_23271,N_24634);
and UO_1787 (O_1787,N_24677,N_22982);
and UO_1788 (O_1788,N_21742,N_20059);
xor UO_1789 (O_1789,N_20212,N_22241);
nor UO_1790 (O_1790,N_22628,N_20464);
nand UO_1791 (O_1791,N_24827,N_24562);
xor UO_1792 (O_1792,N_24729,N_22331);
nor UO_1793 (O_1793,N_20150,N_23459);
nor UO_1794 (O_1794,N_22147,N_24467);
nor UO_1795 (O_1795,N_21408,N_24094);
xnor UO_1796 (O_1796,N_21348,N_23018);
xor UO_1797 (O_1797,N_20671,N_23927);
nand UO_1798 (O_1798,N_23215,N_20917);
or UO_1799 (O_1799,N_21566,N_22004);
and UO_1800 (O_1800,N_22245,N_20462);
nand UO_1801 (O_1801,N_21560,N_24753);
nor UO_1802 (O_1802,N_23150,N_23797);
nor UO_1803 (O_1803,N_21246,N_22025);
or UO_1804 (O_1804,N_22870,N_20373);
nor UO_1805 (O_1805,N_24997,N_23626);
and UO_1806 (O_1806,N_22676,N_23562);
or UO_1807 (O_1807,N_20303,N_20894);
or UO_1808 (O_1808,N_24782,N_24579);
or UO_1809 (O_1809,N_24544,N_23780);
nand UO_1810 (O_1810,N_24694,N_22340);
nor UO_1811 (O_1811,N_21760,N_20174);
and UO_1812 (O_1812,N_24594,N_22504);
nand UO_1813 (O_1813,N_22888,N_21349);
or UO_1814 (O_1814,N_23044,N_23530);
xor UO_1815 (O_1815,N_21992,N_22831);
nor UO_1816 (O_1816,N_22133,N_22750);
or UO_1817 (O_1817,N_22063,N_20414);
and UO_1818 (O_1818,N_22037,N_23528);
nand UO_1819 (O_1819,N_21160,N_21631);
nand UO_1820 (O_1820,N_23293,N_22580);
and UO_1821 (O_1821,N_20615,N_21853);
nor UO_1822 (O_1822,N_21905,N_20355);
nor UO_1823 (O_1823,N_21537,N_22235);
nor UO_1824 (O_1824,N_21427,N_21107);
nand UO_1825 (O_1825,N_20618,N_24340);
and UO_1826 (O_1826,N_21411,N_20679);
nand UO_1827 (O_1827,N_21383,N_24465);
and UO_1828 (O_1828,N_24132,N_21885);
nand UO_1829 (O_1829,N_20242,N_23743);
nor UO_1830 (O_1830,N_21258,N_21839);
or UO_1831 (O_1831,N_20945,N_21351);
nor UO_1832 (O_1832,N_22412,N_21388);
and UO_1833 (O_1833,N_20959,N_21031);
or UO_1834 (O_1834,N_22554,N_23112);
and UO_1835 (O_1835,N_21727,N_23682);
nand UO_1836 (O_1836,N_22179,N_20383);
nor UO_1837 (O_1837,N_23873,N_20189);
nand UO_1838 (O_1838,N_22872,N_24626);
xnor UO_1839 (O_1839,N_22192,N_23684);
nor UO_1840 (O_1840,N_24826,N_24893);
xnor UO_1841 (O_1841,N_24090,N_20140);
or UO_1842 (O_1842,N_20724,N_23643);
or UO_1843 (O_1843,N_24872,N_21755);
or UO_1844 (O_1844,N_20988,N_22472);
xor UO_1845 (O_1845,N_22573,N_23091);
or UO_1846 (O_1846,N_20983,N_24003);
and UO_1847 (O_1847,N_22536,N_23418);
nor UO_1848 (O_1848,N_22259,N_21806);
or UO_1849 (O_1849,N_21462,N_24244);
nand UO_1850 (O_1850,N_24458,N_23559);
and UO_1851 (O_1851,N_23237,N_24386);
or UO_1852 (O_1852,N_24308,N_23027);
or UO_1853 (O_1853,N_20255,N_22986);
nand UO_1854 (O_1854,N_23259,N_20971);
or UO_1855 (O_1855,N_20595,N_23322);
xor UO_1856 (O_1856,N_22757,N_23316);
or UO_1857 (O_1857,N_21752,N_22625);
nand UO_1858 (O_1858,N_21765,N_23988);
nand UO_1859 (O_1859,N_23929,N_22064);
or UO_1860 (O_1860,N_24867,N_22008);
or UO_1861 (O_1861,N_21780,N_22666);
nand UO_1862 (O_1862,N_20481,N_23574);
and UO_1863 (O_1863,N_22151,N_21339);
nand UO_1864 (O_1864,N_21425,N_21872);
or UO_1865 (O_1865,N_21998,N_23433);
and UO_1866 (O_1866,N_24475,N_23408);
and UO_1867 (O_1867,N_22365,N_22671);
nor UO_1868 (O_1868,N_20023,N_24531);
nor UO_1869 (O_1869,N_21440,N_21761);
nand UO_1870 (O_1870,N_24687,N_21045);
or UO_1871 (O_1871,N_24378,N_24426);
and UO_1872 (O_1872,N_22506,N_20024);
nor UO_1873 (O_1873,N_20119,N_21028);
or UO_1874 (O_1874,N_22646,N_21593);
xnor UO_1875 (O_1875,N_24369,N_21418);
and UO_1876 (O_1876,N_21820,N_23164);
nor UO_1877 (O_1877,N_23430,N_20995);
nor UO_1878 (O_1878,N_24073,N_22564);
and UO_1879 (O_1879,N_22983,N_23214);
or UO_1880 (O_1880,N_21718,N_24325);
nor UO_1881 (O_1881,N_22126,N_23212);
nand UO_1882 (O_1882,N_24909,N_21491);
nor UO_1883 (O_1883,N_21158,N_21700);
nand UO_1884 (O_1884,N_22745,N_21694);
and UO_1885 (O_1885,N_24526,N_20382);
or UO_1886 (O_1886,N_23446,N_22431);
nand UO_1887 (O_1887,N_23480,N_22457);
nor UO_1888 (O_1888,N_23578,N_23280);
and UO_1889 (O_1889,N_21259,N_22408);
or UO_1890 (O_1890,N_23546,N_22292);
xnor UO_1891 (O_1891,N_24321,N_23731);
or UO_1892 (O_1892,N_23784,N_20887);
and UO_1893 (O_1893,N_23537,N_24858);
nor UO_1894 (O_1894,N_23471,N_23497);
nor UO_1895 (O_1895,N_23174,N_24747);
or UO_1896 (O_1896,N_24343,N_22981);
nor UO_1897 (O_1897,N_23543,N_20661);
nor UO_1898 (O_1898,N_24504,N_20239);
or UO_1899 (O_1899,N_21191,N_24919);
or UO_1900 (O_1900,N_22902,N_23286);
or UO_1901 (O_1901,N_24194,N_23251);
and UO_1902 (O_1902,N_20166,N_20121);
or UO_1903 (O_1903,N_21548,N_20874);
and UO_1904 (O_1904,N_22489,N_21707);
nor UO_1905 (O_1905,N_22306,N_20726);
xnor UO_1906 (O_1906,N_21356,N_22448);
nand UO_1907 (O_1907,N_24326,N_23191);
or UO_1908 (O_1908,N_21132,N_21567);
and UO_1909 (O_1909,N_24188,N_23067);
nand UO_1910 (O_1910,N_24571,N_20394);
and UO_1911 (O_1911,N_22703,N_24757);
or UO_1912 (O_1912,N_24498,N_22334);
and UO_1913 (O_1913,N_21668,N_20650);
and UO_1914 (O_1914,N_21957,N_22908);
xor UO_1915 (O_1915,N_22394,N_23786);
nand UO_1916 (O_1916,N_24502,N_20291);
and UO_1917 (O_1917,N_21209,N_23492);
nor UO_1918 (O_1918,N_21823,N_23347);
nand UO_1919 (O_1919,N_22994,N_24642);
nand UO_1920 (O_1920,N_22246,N_22836);
xnor UO_1921 (O_1921,N_20976,N_23054);
or UO_1922 (O_1922,N_21697,N_20592);
or UO_1923 (O_1923,N_24961,N_22449);
and UO_1924 (O_1924,N_24406,N_23084);
nand UO_1925 (O_1925,N_20588,N_23205);
and UO_1926 (O_1926,N_24976,N_23652);
or UO_1927 (O_1927,N_22707,N_20093);
and UO_1928 (O_1928,N_23323,N_24469);
xnor UO_1929 (O_1929,N_21871,N_20110);
nand UO_1930 (O_1930,N_24987,N_23606);
nor UO_1931 (O_1931,N_24240,N_23180);
nor UO_1932 (O_1932,N_24805,N_20069);
and UO_1933 (O_1933,N_23050,N_21609);
nand UO_1934 (O_1934,N_22687,N_24532);
nand UO_1935 (O_1935,N_23478,N_23664);
and UO_1936 (O_1936,N_24543,N_21448);
xor UO_1937 (O_1937,N_20628,N_20782);
nand UO_1938 (O_1938,N_21185,N_21738);
nor UO_1939 (O_1939,N_22477,N_23447);
and UO_1940 (O_1940,N_22056,N_22561);
xor UO_1941 (O_1941,N_21574,N_22957);
and UO_1942 (O_1942,N_22072,N_22514);
nand UO_1943 (O_1943,N_22980,N_24333);
and UO_1944 (O_1944,N_20800,N_23375);
xor UO_1945 (O_1945,N_20452,N_22096);
and UO_1946 (O_1946,N_24820,N_21810);
nor UO_1947 (O_1947,N_24720,N_23132);
and UO_1948 (O_1948,N_23989,N_22283);
nor UO_1949 (O_1949,N_23977,N_22136);
and UO_1950 (O_1950,N_20033,N_24229);
xnor UO_1951 (O_1951,N_24419,N_21252);
nand UO_1952 (O_1952,N_21990,N_20041);
nand UO_1953 (O_1953,N_22104,N_21403);
nand UO_1954 (O_1954,N_20711,N_21003);
and UO_1955 (O_1955,N_20989,N_21024);
nor UO_1956 (O_1956,N_22346,N_22397);
or UO_1957 (O_1957,N_24947,N_23725);
or UO_1958 (O_1958,N_22871,N_22851);
nand UO_1959 (O_1959,N_21721,N_24829);
xnor UO_1960 (O_1960,N_22464,N_20048);
nor UO_1961 (O_1961,N_23484,N_20609);
nand UO_1962 (O_1962,N_22708,N_23953);
or UO_1963 (O_1963,N_23654,N_24482);
and UO_1964 (O_1964,N_22043,N_23410);
and UO_1965 (O_1965,N_20126,N_24231);
nor UO_1966 (O_1966,N_21794,N_23117);
nor UO_1967 (O_1967,N_24963,N_22566);
or UO_1968 (O_1968,N_21488,N_21207);
xor UO_1969 (O_1969,N_24681,N_20036);
and UO_1970 (O_1970,N_22258,N_24770);
nand UO_1971 (O_1971,N_21766,N_22260);
nor UO_1972 (O_1972,N_24368,N_20309);
nor UO_1973 (O_1973,N_21821,N_21457);
or UO_1974 (O_1974,N_22145,N_21640);
nor UO_1975 (O_1975,N_23892,N_23564);
nand UO_1976 (O_1976,N_23392,N_21645);
nand UO_1977 (O_1977,N_21999,N_20706);
xor UO_1978 (O_1978,N_22436,N_23196);
xnor UO_1979 (O_1979,N_21099,N_23647);
or UO_1980 (O_1980,N_23012,N_21278);
nand UO_1981 (O_1981,N_20805,N_22544);
and UO_1982 (O_1982,N_22189,N_21996);
or UO_1983 (O_1983,N_24761,N_21884);
or UO_1984 (O_1984,N_20354,N_21692);
nand UO_1985 (O_1985,N_23861,N_22611);
or UO_1986 (O_1986,N_23889,N_20021);
and UO_1987 (O_1987,N_24363,N_21387);
nor UO_1988 (O_1988,N_20346,N_20903);
nor UO_1989 (O_1989,N_20196,N_21176);
nand UO_1990 (O_1990,N_20202,N_20181);
xnor UO_1991 (O_1991,N_22977,N_22035);
and UO_1992 (O_1992,N_23884,N_23563);
nand UO_1993 (O_1993,N_24304,N_24433);
nor UO_1994 (O_1994,N_20896,N_22800);
or UO_1995 (O_1995,N_21346,N_21302);
nand UO_1996 (O_1996,N_23778,N_22583);
or UO_1997 (O_1997,N_23893,N_20444);
nand UO_1998 (O_1998,N_22797,N_20541);
nand UO_1999 (O_1999,N_22076,N_22842);
xor UO_2000 (O_2000,N_22607,N_20681);
and UO_2001 (O_2001,N_20792,N_24903);
nand UO_2002 (O_2002,N_24435,N_23696);
or UO_2003 (O_2003,N_20206,N_20001);
nand UO_2004 (O_2004,N_22571,N_20559);
and UO_2005 (O_2005,N_23243,N_22999);
nor UO_2006 (O_2006,N_20080,N_22301);
and UO_2007 (O_2007,N_23726,N_24513);
nor UO_2008 (O_2008,N_21516,N_24928);
nor UO_2009 (O_2009,N_23419,N_22769);
nand UO_2010 (O_2010,N_24685,N_20451);
xnor UO_2011 (O_2011,N_21797,N_20684);
nor UO_2012 (O_2012,N_21072,N_23199);
or UO_2013 (O_2013,N_22215,N_23655);
xnor UO_2014 (O_2014,N_20824,N_24453);
nor UO_2015 (O_2015,N_22809,N_24449);
or UO_2016 (O_2016,N_24838,N_22098);
nand UO_2017 (O_2017,N_23733,N_21932);
xor UO_2018 (O_2018,N_20884,N_23607);
xnor UO_2019 (O_2019,N_22556,N_22557);
and UO_2020 (O_2020,N_20998,N_20756);
and UO_2021 (O_2021,N_20278,N_23087);
or UO_2022 (O_2022,N_22027,N_24113);
and UO_2023 (O_2023,N_20083,N_21801);
nor UO_2024 (O_2024,N_23393,N_21802);
or UO_2025 (O_2025,N_23075,N_23761);
or UO_2026 (O_2026,N_23919,N_20815);
or UO_2027 (O_2027,N_22629,N_22317);
and UO_2028 (O_2028,N_21253,N_21103);
nor UO_2029 (O_2029,N_20268,N_22529);
and UO_2030 (O_2030,N_21784,N_22314);
or UO_2031 (O_2031,N_21814,N_24604);
nand UO_2032 (O_2032,N_24670,N_23669);
nand UO_2033 (O_2033,N_21156,N_24857);
nor UO_2034 (O_2034,N_23294,N_24015);
xnor UO_2035 (O_2035,N_20597,N_24817);
xor UO_2036 (O_2036,N_20999,N_21924);
and UO_2037 (O_2037,N_24123,N_23961);
or UO_2038 (O_2038,N_24584,N_20384);
nor UO_2039 (O_2039,N_23231,N_23123);
nor UO_2040 (O_2040,N_23940,N_24988);
or UO_2041 (O_2041,N_23507,N_21117);
nand UO_2042 (O_2042,N_24095,N_20447);
and UO_2043 (O_2043,N_22061,N_20527);
nand UO_2044 (O_2044,N_20893,N_24916);
nand UO_2045 (O_2045,N_22366,N_21379);
and UO_2046 (O_2046,N_22242,N_23173);
and UO_2047 (O_2047,N_21055,N_21783);
and UO_2048 (O_2048,N_20499,N_23247);
nor UO_2049 (O_2049,N_20135,N_20381);
nand UO_2050 (O_2050,N_22601,N_23957);
or UO_2051 (O_2051,N_22007,N_22020);
nor UO_2052 (O_2052,N_22103,N_22011);
or UO_2053 (O_2053,N_20302,N_23742);
and UO_2054 (O_2054,N_24413,N_20179);
nand UO_2055 (O_2055,N_20127,N_24464);
or UO_2056 (O_2056,N_24299,N_22710);
and UO_2057 (O_2057,N_23346,N_23675);
or UO_2058 (O_2058,N_20336,N_20827);
xor UO_2059 (O_2059,N_20327,N_20281);
xor UO_2060 (O_2060,N_23334,N_22392);
and UO_2061 (O_2061,N_24748,N_23096);
nor UO_2062 (O_2062,N_24062,N_22567);
and UO_2063 (O_2063,N_24763,N_20819);
nand UO_2064 (O_2064,N_23896,N_24007);
xor UO_2065 (O_2065,N_20467,N_23633);
or UO_2066 (O_2066,N_23995,N_22998);
and UO_2067 (O_2067,N_23474,N_22919);
and UO_2068 (O_2068,N_21861,N_24978);
xor UO_2069 (O_2069,N_24315,N_21866);
nor UO_2070 (O_2070,N_24735,N_24139);
xnor UO_2071 (O_2071,N_24849,N_24773);
and UO_2072 (O_2072,N_24606,N_20736);
nand UO_2073 (O_2073,N_20032,N_24627);
xor UO_2074 (O_2074,N_23589,N_24693);
or UO_2075 (O_2075,N_20710,N_22674);
nor UO_2076 (O_2076,N_21227,N_20493);
or UO_2077 (O_2077,N_20755,N_24097);
and UO_2078 (O_2078,N_20433,N_20911);
nor UO_2079 (O_2079,N_21655,N_23424);
nor UO_2080 (O_2080,N_22681,N_20631);
or UO_2081 (O_2081,N_21374,N_23951);
nor UO_2082 (O_2082,N_24297,N_21534);
nand UO_2083 (O_2083,N_20859,N_23304);
and UO_2084 (O_2084,N_20457,N_21652);
or UO_2085 (O_2085,N_23413,N_21620);
nand UO_2086 (O_2086,N_22767,N_24387);
or UO_2087 (O_2087,N_21040,N_24445);
and UO_2088 (O_2088,N_23435,N_22608);
and UO_2089 (O_2089,N_21354,N_21095);
nor UO_2090 (O_2090,N_20900,N_23313);
or UO_2091 (O_2091,N_21308,N_23588);
and UO_2092 (O_2092,N_21152,N_20375);
nand UO_2093 (O_2093,N_24680,N_24783);
xor UO_2094 (O_2094,N_22493,N_22766);
or UO_2095 (O_2095,N_22741,N_22978);
or UO_2096 (O_2096,N_24637,N_20221);
or UO_2097 (O_2097,N_23260,N_24461);
nand UO_2098 (O_2098,N_23154,N_21446);
or UO_2099 (O_2099,N_21100,N_24538);
xnor UO_2100 (O_2100,N_20376,N_20257);
and UO_2101 (O_2101,N_23008,N_23073);
nor UO_2102 (O_2102,N_21602,N_23373);
nor UO_2103 (O_2103,N_24441,N_20369);
nand UO_2104 (O_2104,N_20410,N_23969);
xnor UO_2105 (O_2105,N_24048,N_20810);
or UO_2106 (O_2106,N_20208,N_24713);
or UO_2107 (O_2107,N_20557,N_24228);
nor UO_2108 (O_2108,N_23857,N_24078);
or UO_2109 (O_2109,N_21395,N_20868);
and UO_2110 (O_2110,N_20092,N_21800);
nand UO_2111 (O_2111,N_21965,N_24181);
and UO_2112 (O_2112,N_22327,N_24583);
xnor UO_2113 (O_2113,N_22862,N_23481);
nor UO_2114 (O_2114,N_24079,N_20845);
xor UO_2115 (O_2115,N_21275,N_21429);
nand UO_2116 (O_2116,N_22348,N_23502);
and UO_2117 (O_2117,N_23167,N_24290);
nor UO_2118 (O_2118,N_23489,N_24866);
nand UO_2119 (O_2119,N_21315,N_23244);
nor UO_2120 (O_2120,N_24914,N_21378);
nand UO_2121 (O_2121,N_24135,N_21284);
or UO_2122 (O_2122,N_21664,N_22824);
nand UO_2123 (O_2123,N_22294,N_24913);
and UO_2124 (O_2124,N_23897,N_23242);
nor UO_2125 (O_2125,N_23899,N_20310);
nand UO_2126 (O_2126,N_22186,N_24085);
and UO_2127 (O_2127,N_21779,N_20641);
nand UO_2128 (O_2128,N_24890,N_21240);
nand UO_2129 (O_2129,N_20306,N_21049);
or UO_2130 (O_2130,N_21122,N_21588);
nand UO_2131 (O_2131,N_21069,N_24136);
and UO_2132 (O_2132,N_22156,N_24620);
nand UO_2133 (O_2133,N_22266,N_22520);
nand UO_2134 (O_2134,N_20550,N_20288);
or UO_2135 (O_2135,N_23365,N_23453);
nor UO_2136 (O_2136,N_21502,N_22187);
and UO_2137 (O_2137,N_20356,N_22295);
nor UO_2138 (O_2138,N_23058,N_21019);
or UO_2139 (O_2139,N_23715,N_22713);
nand UO_2140 (O_2140,N_23303,N_22753);
and UO_2141 (O_2141,N_20058,N_23685);
and UO_2142 (O_2142,N_24565,N_24284);
or UO_2143 (O_2143,N_24930,N_24933);
nor UO_2144 (O_2144,N_23047,N_23783);
nand UO_2145 (O_2145,N_21577,N_24925);
and UO_2146 (O_2146,N_22289,N_20538);
and UO_2147 (O_2147,N_20653,N_21650);
nand UO_2148 (O_2148,N_21722,N_21695);
and UO_2149 (O_2149,N_20361,N_21506);
or UO_2150 (O_2150,N_23820,N_20305);
or UO_2151 (O_2151,N_22542,N_22351);
and UO_2152 (O_2152,N_21083,N_21243);
and UO_2153 (O_2153,N_20034,N_22183);
nand UO_2154 (O_2154,N_20809,N_21023);
nor UO_2155 (O_2155,N_21034,N_21063);
and UO_2156 (O_2156,N_22400,N_22144);
or UO_2157 (O_2157,N_20049,N_23854);
nand UO_2158 (O_2158,N_22427,N_21632);
and UO_2159 (O_2159,N_24905,N_23179);
nor UO_2160 (O_2160,N_23802,N_21285);
nand UO_2161 (O_2161,N_22911,N_20318);
nand UO_2162 (O_2162,N_21218,N_21123);
nand UO_2163 (O_2163,N_22088,N_21222);
nor UO_2164 (O_2164,N_21886,N_20269);
nand UO_2165 (O_2165,N_24633,N_24802);
nor UO_2166 (O_2166,N_20664,N_20279);
or UO_2167 (O_2167,N_22645,N_24871);
nand UO_2168 (O_2168,N_21059,N_20222);
nand UO_2169 (O_2169,N_23057,N_23370);
xnor UO_2170 (O_2170,N_21007,N_23610);
and UO_2171 (O_2171,N_22450,N_24569);
and UO_2172 (O_2172,N_20063,N_23088);
nor UO_2173 (O_2173,N_20950,N_21778);
and UO_2174 (O_2174,N_24972,N_24266);
and UO_2175 (O_2175,N_21815,N_21623);
nor UO_2176 (O_2176,N_24173,N_24794);
nand UO_2177 (O_2177,N_21536,N_20942);
nor UO_2178 (O_2178,N_22778,N_24556);
and UO_2179 (O_2179,N_21036,N_21708);
or UO_2180 (O_2180,N_21896,N_24164);
nand UO_2181 (O_2181,N_22946,N_23670);
nand UO_2182 (O_2182,N_22568,N_22313);
and UO_2183 (O_2183,N_24337,N_20500);
nor UO_2184 (O_2184,N_21669,N_20195);
and UO_2185 (O_2185,N_22547,N_22988);
or UO_2186 (O_2186,N_24476,N_23307);
nand UO_2187 (O_2187,N_21213,N_21293);
nor UO_2188 (O_2188,N_20065,N_24124);
nor UO_2189 (O_2189,N_24647,N_21974);
or UO_2190 (O_2190,N_22642,N_20483);
nand UO_2191 (O_2191,N_21460,N_22945);
or UO_2192 (O_2192,N_20131,N_23575);
nand UO_2193 (O_2193,N_21673,N_23516);
and UO_2194 (O_2194,N_21882,N_20886);
nor UO_2195 (O_2195,N_21747,N_20495);
nor UO_2196 (O_2196,N_22371,N_22378);
or UO_2197 (O_2197,N_24114,N_22106);
and UO_2198 (O_2198,N_20272,N_24587);
and UO_2199 (O_2199,N_23353,N_24611);
and UO_2200 (O_2200,N_20578,N_21703);
nor UO_2201 (O_2201,N_21179,N_22490);
or UO_2202 (O_2202,N_20160,N_24030);
and UO_2203 (O_2203,N_21489,N_22843);
nand UO_2204 (O_2204,N_24979,N_22277);
or UO_2205 (O_2205,N_23941,N_23162);
nand UO_2206 (O_2206,N_24990,N_24134);
nor UO_2207 (O_2207,N_21582,N_21684);
and UO_2208 (O_2208,N_23296,N_23483);
nand UO_2209 (O_2209,N_23315,N_23386);
or UO_2210 (O_2210,N_24001,N_20954);
nor UO_2211 (O_2211,N_24038,N_21091);
nor UO_2212 (O_2212,N_21756,N_24473);
nand UO_2213 (O_2213,N_21847,N_23918);
nand UO_2214 (O_2214,N_22432,N_22788);
and UO_2215 (O_2215,N_23533,N_21329);
nand UO_2216 (O_2216,N_23135,N_22522);
or UO_2217 (O_2217,N_24727,N_20116);
and UO_2218 (O_2218,N_24723,N_24743);
nor UO_2219 (O_2219,N_20712,N_23911);
nand UO_2220 (O_2220,N_22579,N_22384);
or UO_2221 (O_2221,N_24303,N_21565);
and UO_2222 (O_2222,N_24039,N_24524);
nand UO_2223 (O_2223,N_23224,N_22426);
or UO_2224 (O_2224,N_24877,N_20854);
nand UO_2225 (O_2225,N_24711,N_20832);
and UO_2226 (O_2226,N_23031,N_24058);
or UO_2227 (O_2227,N_22332,N_24264);
or UO_2228 (O_2228,N_22825,N_23071);
or UO_2229 (O_2229,N_21096,N_22018);
and UO_2230 (O_2230,N_21764,N_21897);
and UO_2231 (O_2231,N_21870,N_23828);
or UO_2232 (O_2232,N_21065,N_23229);
or UO_2233 (O_2233,N_22481,N_20438);
nand UO_2234 (O_2234,N_24844,N_21648);
xor UO_2235 (O_2235,N_24067,N_21649);
nor UO_2236 (O_2236,N_20133,N_22884);
and UO_2237 (O_2237,N_23220,N_24418);
and UO_2238 (O_2238,N_24439,N_23034);
and UO_2239 (O_2239,N_24725,N_23023);
or UO_2240 (O_2240,N_21372,N_20620);
nor UO_2241 (O_2241,N_24282,N_20228);
xor UO_2242 (O_2242,N_24639,N_23752);
or UO_2243 (O_2243,N_20497,N_24911);
nor UO_2244 (O_2244,N_22834,N_22817);
and UO_2245 (O_2245,N_22990,N_23256);
and UO_2246 (O_2246,N_24631,N_23673);
and UO_2247 (O_2247,N_22891,N_23846);
nor UO_2248 (O_2248,N_24121,N_22669);
nand UO_2249 (O_2249,N_20927,N_20047);
and UO_2250 (O_2250,N_22016,N_22414);
or UO_2251 (O_2251,N_20276,N_22743);
nand UO_2252 (O_2252,N_21030,N_22369);
or UO_2253 (O_2253,N_23272,N_22989);
nor UO_2254 (O_2254,N_22462,N_20817);
or UO_2255 (O_2255,N_24027,N_23427);
nor UO_2256 (O_2256,N_22690,N_22223);
or UO_2257 (O_2257,N_20572,N_20280);
xnor UO_2258 (O_2258,N_23414,N_20337);
or UO_2259 (O_2259,N_21858,N_24892);
nor UO_2260 (O_2260,N_21469,N_24960);
and UO_2261 (O_2261,N_21498,N_24361);
xor UO_2262 (O_2262,N_22102,N_22644);
xnor UO_2263 (O_2263,N_21571,N_21510);
nand UO_2264 (O_2264,N_23228,N_24431);
and UO_2265 (O_2265,N_24209,N_20016);
and UO_2266 (O_2266,N_23536,N_22358);
nor UO_2267 (O_2267,N_20746,N_20112);
and UO_2268 (O_2268,N_22846,N_20958);
or UO_2269 (O_2269,N_22928,N_24200);
and UO_2270 (O_2270,N_24189,N_21951);
nand UO_2271 (O_2271,N_24654,N_24145);
xor UO_2272 (O_2272,N_20946,N_24712);
nor UO_2273 (O_2273,N_23308,N_21997);
nand UO_2274 (O_2274,N_23704,N_22271);
xnor UO_2275 (O_2275,N_21798,N_24703);
nand UO_2276 (O_2276,N_21982,N_22885);
and UO_2277 (O_2277,N_23377,N_20118);
nand UO_2278 (O_2278,N_23443,N_24738);
or UO_2279 (O_2279,N_20673,N_23808);
and UO_2280 (O_2280,N_20197,N_23358);
nand UO_2281 (O_2281,N_23935,N_24492);
or UO_2282 (O_2282,N_20005,N_24541);
nand UO_2283 (O_2283,N_20910,N_24695);
or UO_2284 (O_2284,N_24510,N_24305);
xor UO_2285 (O_2285,N_24706,N_20503);
and UO_2286 (O_2286,N_21358,N_22634);
or UO_2287 (O_2287,N_22130,N_24709);
xnor UO_2288 (O_2288,N_20256,N_22003);
nor UO_2289 (O_2289,N_22236,N_22068);
or UO_2290 (O_2290,N_22328,N_21255);
nor UO_2291 (O_2291,N_21148,N_20981);
nand UO_2292 (O_2292,N_21622,N_24044);
and UO_2293 (O_2293,N_20581,N_23836);
nand UO_2294 (O_2294,N_23493,N_21441);
and UO_2295 (O_2295,N_23656,N_20128);
nor UO_2296 (O_2296,N_20627,N_23295);
or UO_2297 (O_2297,N_20747,N_21643);
nand UO_2298 (O_2298,N_22212,N_22526);
nand UO_2299 (O_2299,N_20657,N_22319);
nor UO_2300 (O_2300,N_21517,N_24608);
nor UO_2301 (O_2301,N_21340,N_23371);
nor UO_2302 (O_2302,N_24940,N_20122);
and UO_2303 (O_2303,N_21969,N_21400);
or UO_2304 (O_2304,N_20198,N_23714);
nand UO_2305 (O_2305,N_20298,N_20173);
and UO_2306 (O_2306,N_24734,N_21663);
nand UO_2307 (O_2307,N_20863,N_20084);
nor UO_2308 (O_2308,N_23113,N_24197);
or UO_2309 (O_2309,N_23477,N_21214);
nand UO_2310 (O_2310,N_21918,N_24823);
and UO_2311 (O_2311,N_23379,N_22688);
xnor UO_2312 (O_2312,N_20205,N_24517);
nand UO_2313 (O_2313,N_21273,N_22624);
nor UO_2314 (O_2314,N_22938,N_20918);
nand UO_2315 (O_2315,N_21194,N_22701);
nand UO_2316 (O_2316,N_20537,N_21876);
nand UO_2317 (O_2317,N_23311,N_24669);
or UO_2318 (O_2318,N_22310,N_24047);
xnor UO_2319 (O_2319,N_23387,N_24083);
nor UO_2320 (O_2320,N_24403,N_21522);
and UO_2321 (O_2321,N_21771,N_21724);
xnor UO_2322 (O_2322,N_23816,N_21394);
nor UO_2323 (O_2323,N_20619,N_23299);
nand UO_2324 (O_2324,N_24484,N_23775);
and UO_2325 (O_2325,N_23051,N_24174);
and UO_2326 (O_2326,N_22636,N_20633);
or UO_2327 (O_2327,N_21540,N_22694);
nand UO_2328 (O_2328,N_20027,N_24515);
xnor UO_2329 (O_2329,N_23469,N_21585);
xor UO_2330 (O_2330,N_24812,N_21323);
xor UO_2331 (O_2331,N_20194,N_21277);
or UO_2332 (O_2332,N_20231,N_23189);
or UO_2333 (O_2333,N_21748,N_21131);
nand UO_2334 (O_2334,N_24528,N_24428);
or UO_2335 (O_2335,N_23273,N_22349);
and UO_2336 (O_2336,N_22452,N_20446);
and UO_2337 (O_2337,N_20742,N_21554);
or UO_2338 (O_2338,N_23557,N_24830);
nand UO_2339 (O_2339,N_22866,N_21056);
and UO_2340 (O_2340,N_20686,N_21247);
nor UO_2341 (O_2341,N_22917,N_24267);
nor UO_2342 (O_2342,N_20104,N_24312);
or UO_2343 (O_2343,N_24686,N_24751);
nor UO_2344 (O_2344,N_21515,N_23653);
nor UO_2345 (O_2345,N_20964,N_21181);
nor UO_2346 (O_2346,N_22218,N_24040);
nand UO_2347 (O_2347,N_20873,N_24319);
nand UO_2348 (O_2348,N_23671,N_23503);
and UO_2349 (O_2349,N_22304,N_22067);
and UO_2350 (O_2350,N_21174,N_23980);
and UO_2351 (O_2351,N_23434,N_24414);
or UO_2352 (O_2352,N_20584,N_20229);
nor UO_2353 (O_2353,N_20847,N_22083);
and UO_2354 (O_2354,N_23378,N_23553);
nand UO_2355 (O_2355,N_20170,N_22513);
nor UO_2356 (O_2356,N_24151,N_23333);
and UO_2357 (O_2357,N_20922,N_22918);
nor UO_2358 (O_2358,N_20904,N_20905);
nand UO_2359 (O_2359,N_22193,N_21015);
nor UO_2360 (O_2360,N_24131,N_20163);
nor UO_2361 (O_2361,N_23814,N_24614);
and UO_2362 (O_2362,N_24436,N_22552);
nand UO_2363 (O_2363,N_24416,N_22248);
nor UO_2364 (O_2364,N_21556,N_21913);
and UO_2365 (O_2365,N_23394,N_22795);
and UO_2366 (O_2366,N_24523,N_24946);
or UO_2367 (O_2367,N_20329,N_20094);
nor UO_2368 (O_2368,N_21987,N_20707);
nand UO_2369 (O_2369,N_23175,N_23362);
nor UO_2370 (O_2370,N_20666,N_20965);
nand UO_2371 (O_2371,N_22373,N_23422);
and UO_2372 (O_2372,N_22162,N_21336);
nand UO_2373 (O_2373,N_24375,N_20340);
or UO_2374 (O_2374,N_23429,N_21889);
or UO_2375 (O_2375,N_22469,N_21699);
nor UO_2376 (O_2376,N_21789,N_22039);
nor UO_2377 (O_2377,N_24130,N_24059);
nand UO_2378 (O_2378,N_20151,N_23983);
and UO_2379 (O_2379,N_21591,N_20079);
nor UO_2380 (O_2380,N_20688,N_24744);
nor UO_2381 (O_2381,N_22565,N_21257);
xor UO_2382 (O_2382,N_21033,N_23221);
nor UO_2383 (O_2383,N_20566,N_20769);
xnor UO_2384 (O_2384,N_23766,N_23116);
and UO_2385 (O_2385,N_23053,N_24318);
nor UO_2386 (O_2386,N_21229,N_23668);
nor UO_2387 (O_2387,N_21954,N_20416);
nor UO_2388 (O_2388,N_23171,N_22922);
nor UO_2389 (O_2389,N_23204,N_20317);
and UO_2390 (O_2390,N_23195,N_23992);
nor UO_2391 (O_2391,N_21799,N_21292);
or UO_2392 (O_2392,N_22410,N_21917);
nor UO_2393 (O_2393,N_23581,N_21492);
or UO_2394 (O_2394,N_22826,N_23125);
or UO_2395 (O_2395,N_22390,N_20986);
or UO_2396 (O_2396,N_22284,N_21371);
nand UO_2397 (O_2397,N_21558,N_21813);
and UO_2398 (O_2398,N_22297,N_21666);
nor UO_2399 (O_2399,N_22463,N_22841);
and UO_2400 (O_2400,N_20843,N_21165);
nand UO_2401 (O_2401,N_21248,N_20551);
nor UO_2402 (O_2402,N_21525,N_21519);
or UO_2403 (O_2403,N_23599,N_21111);
or UO_2404 (O_2404,N_20739,N_24675);
and UO_2405 (O_2405,N_20400,N_20322);
or UO_2406 (O_2406,N_20299,N_23973);
nor UO_2407 (O_2407,N_24486,N_21865);
and UO_2408 (O_2408,N_20185,N_23241);
and UO_2409 (O_2409,N_21251,N_22387);
nand UO_2410 (O_2410,N_23482,N_23341);
or UO_2411 (O_2411,N_22494,N_20665);
and UO_2412 (O_2412,N_24052,N_24899);
or UO_2413 (O_2413,N_24853,N_21454);
xnor UO_2414 (O_2414,N_21628,N_24907);
nand UO_2415 (O_2415,N_20853,N_24766);
or UO_2416 (O_2416,N_22299,N_24951);
xor UO_2417 (O_2417,N_21382,N_23855);
xnor UO_2418 (O_2418,N_20757,N_20622);
nand UO_2419 (O_2419,N_20139,N_20313);
nand UO_2420 (O_2420,N_23262,N_20872);
or UO_2421 (O_2421,N_23920,N_23789);
nor UO_2422 (O_2422,N_22684,N_24745);
nand UO_2423 (O_2423,N_24986,N_23498);
and UO_2424 (O_2424,N_23426,N_23990);
and UO_2425 (O_2425,N_23519,N_21937);
or UO_2426 (O_2426,N_22590,N_21544);
nor UO_2427 (O_2427,N_21390,N_20363);
and UO_2428 (O_2428,N_20415,N_20477);
nand UO_2429 (O_2429,N_23765,N_24721);
nand UO_2430 (O_2430,N_23348,N_22019);
or UO_2431 (O_2431,N_20831,N_20536);
and UO_2432 (O_2432,N_22700,N_22060);
or UO_2433 (O_2433,N_22446,N_22584);
xor UO_2434 (O_2434,N_22474,N_23955);
or UO_2435 (O_2435,N_20274,N_24243);
and UO_2436 (O_2436,N_24505,N_22166);
nor UO_2437 (O_2437,N_20812,N_23253);
nor UO_2438 (O_2438,N_23172,N_22149);
nor UO_2439 (O_2439,N_22791,N_24876);
and UO_2440 (O_2440,N_24298,N_20328);
or UO_2441 (O_2441,N_21715,N_24443);
nor UO_2442 (O_2442,N_21420,N_24592);
or UO_2443 (O_2443,N_24457,N_20607);
nor UO_2444 (O_2444,N_24601,N_24843);
xor UO_2445 (O_2445,N_23011,N_20985);
nand UO_2446 (O_2446,N_21959,N_23605);
nand UO_2447 (O_2447,N_20492,N_21848);
nand UO_2448 (O_2448,N_24779,N_20455);
nor UO_2449 (O_2449,N_20425,N_22763);
nand UO_2450 (O_2450,N_24906,N_22442);
or UO_2451 (O_2451,N_22069,N_21471);
nor UO_2452 (O_2452,N_23584,N_21991);
nand UO_2453 (O_2453,N_23885,N_24530);
nor UO_2454 (O_2454,N_24099,N_21413);
or UO_2455 (O_2455,N_21496,N_21723);
and UO_2456 (O_2456,N_20217,N_23515);
or UO_2457 (O_2457,N_24821,N_23916);
nor UO_2458 (O_2458,N_20262,N_22760);
and UO_2459 (O_2459,N_23963,N_21763);
and UO_2460 (O_2460,N_20422,N_22092);
and UO_2461 (O_2461,N_23176,N_21523);
nor UO_2462 (O_2462,N_23063,N_24704);
nand UO_2463 (O_2463,N_22975,N_20134);
and UO_2464 (O_2464,N_22482,N_22768);
nand UO_2465 (O_2465,N_24479,N_23835);
nand UO_2466 (O_2466,N_21459,N_22510);
nand UO_2467 (O_2467,N_23452,N_23826);
nand UO_2468 (O_2468,N_20223,N_20634);
and UO_2469 (O_2469,N_22976,N_22519);
nor UO_2470 (O_2470,N_22168,N_20926);
nor UO_2471 (O_2471,N_21187,N_24917);
and UO_2472 (O_2472,N_20136,N_22961);
and UO_2473 (O_2473,N_22066,N_24028);
xnor UO_2474 (O_2474,N_24545,N_24863);
nand UO_2475 (O_2475,N_20956,N_22201);
xor UO_2476 (O_2476,N_23143,N_20233);
nand UO_2477 (O_2477,N_22659,N_24550);
nand UO_2478 (O_2478,N_20912,N_21494);
nand UO_2479 (O_2479,N_21520,N_24089);
or UO_2480 (O_2480,N_21687,N_22038);
xor UO_2481 (O_2481,N_24884,N_24157);
or UO_2482 (O_2482,N_20952,N_21362);
and UO_2483 (O_2483,N_20334,N_23900);
xor UO_2484 (O_2484,N_21627,N_23369);
or UO_2485 (O_2485,N_22508,N_23794);
xnor UO_2486 (O_2486,N_24605,N_24146);
nor UO_2487 (O_2487,N_24000,N_23729);
nor UO_2488 (O_2488,N_23811,N_24150);
nor UO_2489 (O_2489,N_24076,N_21062);
nand UO_2490 (O_2490,N_20091,N_20796);
and UO_2491 (O_2491,N_24516,N_21405);
nor UO_2492 (O_2492,N_21245,N_20932);
or UO_2493 (O_2493,N_23804,N_20401);
or UO_2494 (O_2494,N_20325,N_23278);
nor UO_2495 (O_2495,N_24105,N_22113);
xor UO_2496 (O_2496,N_20741,N_22729);
or UO_2497 (O_2497,N_24612,N_21568);
xor UO_2498 (O_2498,N_23479,N_20867);
xnor UO_2499 (O_2499,N_20651,N_22934);
nand UO_2500 (O_2500,N_24298,N_23868);
or UO_2501 (O_2501,N_21427,N_23530);
nand UO_2502 (O_2502,N_20076,N_21155);
and UO_2503 (O_2503,N_23309,N_24935);
nor UO_2504 (O_2504,N_20498,N_23672);
nand UO_2505 (O_2505,N_22150,N_24827);
nor UO_2506 (O_2506,N_21472,N_21659);
nor UO_2507 (O_2507,N_24318,N_23960);
nor UO_2508 (O_2508,N_23723,N_23645);
nand UO_2509 (O_2509,N_22284,N_22691);
nand UO_2510 (O_2510,N_24834,N_21677);
nor UO_2511 (O_2511,N_24510,N_20331);
nor UO_2512 (O_2512,N_24206,N_21612);
nand UO_2513 (O_2513,N_24881,N_21767);
nand UO_2514 (O_2514,N_20769,N_20026);
nor UO_2515 (O_2515,N_23688,N_22232);
and UO_2516 (O_2516,N_24147,N_24508);
and UO_2517 (O_2517,N_22797,N_20908);
or UO_2518 (O_2518,N_24613,N_21515);
xor UO_2519 (O_2519,N_22290,N_20833);
or UO_2520 (O_2520,N_23523,N_20091);
or UO_2521 (O_2521,N_21525,N_24749);
and UO_2522 (O_2522,N_23443,N_23708);
xor UO_2523 (O_2523,N_24283,N_23474);
or UO_2524 (O_2524,N_21104,N_24981);
nor UO_2525 (O_2525,N_20587,N_24957);
and UO_2526 (O_2526,N_23784,N_24352);
or UO_2527 (O_2527,N_21872,N_21214);
nand UO_2528 (O_2528,N_20351,N_23209);
xnor UO_2529 (O_2529,N_21704,N_23826);
or UO_2530 (O_2530,N_21379,N_21511);
nand UO_2531 (O_2531,N_24700,N_24971);
nor UO_2532 (O_2532,N_22073,N_23093);
nor UO_2533 (O_2533,N_20347,N_21710);
or UO_2534 (O_2534,N_22666,N_20857);
nand UO_2535 (O_2535,N_20347,N_20375);
xor UO_2536 (O_2536,N_22135,N_23518);
or UO_2537 (O_2537,N_21149,N_24503);
and UO_2538 (O_2538,N_20345,N_21425);
and UO_2539 (O_2539,N_24116,N_23803);
nand UO_2540 (O_2540,N_20356,N_23695);
nand UO_2541 (O_2541,N_20129,N_24412);
or UO_2542 (O_2542,N_22515,N_22238);
or UO_2543 (O_2543,N_24880,N_23942);
xnor UO_2544 (O_2544,N_21260,N_24667);
nand UO_2545 (O_2545,N_20574,N_21677);
or UO_2546 (O_2546,N_21328,N_24633);
and UO_2547 (O_2547,N_20508,N_23795);
nor UO_2548 (O_2548,N_22546,N_22115);
or UO_2549 (O_2549,N_20224,N_21224);
xor UO_2550 (O_2550,N_20074,N_24845);
or UO_2551 (O_2551,N_24496,N_21597);
nand UO_2552 (O_2552,N_22756,N_21365);
and UO_2553 (O_2553,N_21947,N_21053);
nand UO_2554 (O_2554,N_21778,N_22081);
and UO_2555 (O_2555,N_22812,N_22338);
nand UO_2556 (O_2556,N_21736,N_24620);
nor UO_2557 (O_2557,N_20276,N_24326);
xnor UO_2558 (O_2558,N_24054,N_23734);
nor UO_2559 (O_2559,N_23485,N_22186);
or UO_2560 (O_2560,N_22883,N_24573);
nand UO_2561 (O_2561,N_21034,N_24587);
nor UO_2562 (O_2562,N_22513,N_24843);
or UO_2563 (O_2563,N_22300,N_20829);
nand UO_2564 (O_2564,N_23117,N_23558);
nand UO_2565 (O_2565,N_22926,N_23781);
nor UO_2566 (O_2566,N_21842,N_24057);
xor UO_2567 (O_2567,N_23443,N_20794);
xor UO_2568 (O_2568,N_21738,N_24976);
nand UO_2569 (O_2569,N_22730,N_23510);
or UO_2570 (O_2570,N_20909,N_21458);
nand UO_2571 (O_2571,N_21588,N_21235);
xor UO_2572 (O_2572,N_23733,N_24793);
nor UO_2573 (O_2573,N_22611,N_21837);
or UO_2574 (O_2574,N_22315,N_24228);
nand UO_2575 (O_2575,N_22480,N_20527);
nand UO_2576 (O_2576,N_21504,N_24933);
nor UO_2577 (O_2577,N_20481,N_24787);
or UO_2578 (O_2578,N_21037,N_21697);
nor UO_2579 (O_2579,N_22708,N_24119);
nand UO_2580 (O_2580,N_22567,N_20426);
and UO_2581 (O_2581,N_20170,N_23995);
and UO_2582 (O_2582,N_23702,N_21314);
xnor UO_2583 (O_2583,N_21620,N_23435);
nand UO_2584 (O_2584,N_20367,N_22852);
nand UO_2585 (O_2585,N_21605,N_21973);
nor UO_2586 (O_2586,N_24185,N_20212);
xor UO_2587 (O_2587,N_21841,N_20218);
and UO_2588 (O_2588,N_24031,N_23425);
nor UO_2589 (O_2589,N_24004,N_22032);
nand UO_2590 (O_2590,N_20491,N_22809);
or UO_2591 (O_2591,N_23383,N_20870);
nand UO_2592 (O_2592,N_22828,N_21784);
and UO_2593 (O_2593,N_20838,N_22250);
nand UO_2594 (O_2594,N_21850,N_20754);
nand UO_2595 (O_2595,N_22877,N_21535);
nor UO_2596 (O_2596,N_24966,N_21897);
nor UO_2597 (O_2597,N_21561,N_22179);
nor UO_2598 (O_2598,N_20590,N_22089);
and UO_2599 (O_2599,N_20448,N_20959);
and UO_2600 (O_2600,N_24446,N_21843);
and UO_2601 (O_2601,N_21897,N_20708);
xnor UO_2602 (O_2602,N_23327,N_20268);
or UO_2603 (O_2603,N_21344,N_24174);
or UO_2604 (O_2604,N_23402,N_24342);
and UO_2605 (O_2605,N_21963,N_22843);
and UO_2606 (O_2606,N_23610,N_20822);
xnor UO_2607 (O_2607,N_22635,N_20488);
or UO_2608 (O_2608,N_22488,N_23367);
xnor UO_2609 (O_2609,N_20901,N_20453);
nor UO_2610 (O_2610,N_21966,N_21933);
or UO_2611 (O_2611,N_20789,N_20028);
nor UO_2612 (O_2612,N_21530,N_20941);
or UO_2613 (O_2613,N_21373,N_20438);
and UO_2614 (O_2614,N_24715,N_22051);
nand UO_2615 (O_2615,N_23699,N_22437);
nor UO_2616 (O_2616,N_23280,N_23429);
nand UO_2617 (O_2617,N_22012,N_21162);
nor UO_2618 (O_2618,N_23938,N_23235);
or UO_2619 (O_2619,N_21320,N_20697);
nand UO_2620 (O_2620,N_24226,N_20362);
nor UO_2621 (O_2621,N_22974,N_21523);
nor UO_2622 (O_2622,N_22437,N_24589);
and UO_2623 (O_2623,N_23962,N_24395);
nor UO_2624 (O_2624,N_22457,N_20318);
nor UO_2625 (O_2625,N_24491,N_24775);
nand UO_2626 (O_2626,N_21630,N_21611);
nand UO_2627 (O_2627,N_22230,N_21157);
nor UO_2628 (O_2628,N_23564,N_21057);
nor UO_2629 (O_2629,N_23343,N_24262);
nand UO_2630 (O_2630,N_20202,N_24715);
xnor UO_2631 (O_2631,N_24164,N_24233);
and UO_2632 (O_2632,N_24819,N_21927);
nor UO_2633 (O_2633,N_20763,N_21239);
nor UO_2634 (O_2634,N_24764,N_22553);
or UO_2635 (O_2635,N_21662,N_21029);
and UO_2636 (O_2636,N_22308,N_22355);
xnor UO_2637 (O_2637,N_23757,N_23310);
and UO_2638 (O_2638,N_21767,N_20243);
nand UO_2639 (O_2639,N_22671,N_22916);
and UO_2640 (O_2640,N_23621,N_24892);
or UO_2641 (O_2641,N_22126,N_21672);
or UO_2642 (O_2642,N_24974,N_24284);
and UO_2643 (O_2643,N_22542,N_21626);
or UO_2644 (O_2644,N_20542,N_20979);
nand UO_2645 (O_2645,N_24095,N_23901);
and UO_2646 (O_2646,N_21478,N_21695);
and UO_2647 (O_2647,N_24699,N_20687);
nand UO_2648 (O_2648,N_22247,N_21298);
nand UO_2649 (O_2649,N_21419,N_21646);
xor UO_2650 (O_2650,N_20459,N_22227);
or UO_2651 (O_2651,N_20877,N_21577);
nand UO_2652 (O_2652,N_24554,N_20462);
nand UO_2653 (O_2653,N_22361,N_23070);
nand UO_2654 (O_2654,N_20267,N_24918);
nor UO_2655 (O_2655,N_22823,N_24520);
nand UO_2656 (O_2656,N_23275,N_23164);
or UO_2657 (O_2657,N_22237,N_22245);
nand UO_2658 (O_2658,N_23314,N_20333);
and UO_2659 (O_2659,N_22555,N_22986);
or UO_2660 (O_2660,N_20577,N_24624);
nor UO_2661 (O_2661,N_21010,N_24527);
nor UO_2662 (O_2662,N_21275,N_21866);
nand UO_2663 (O_2663,N_21883,N_20942);
or UO_2664 (O_2664,N_24577,N_23794);
and UO_2665 (O_2665,N_21249,N_20072);
or UO_2666 (O_2666,N_21588,N_23273);
nor UO_2667 (O_2667,N_21191,N_22932);
and UO_2668 (O_2668,N_20025,N_24839);
or UO_2669 (O_2669,N_20116,N_20209);
or UO_2670 (O_2670,N_23285,N_22941);
nor UO_2671 (O_2671,N_20485,N_21215);
or UO_2672 (O_2672,N_21556,N_24037);
and UO_2673 (O_2673,N_20603,N_24639);
or UO_2674 (O_2674,N_22085,N_20775);
nand UO_2675 (O_2675,N_22529,N_24660);
xnor UO_2676 (O_2676,N_21856,N_22175);
or UO_2677 (O_2677,N_20890,N_24092);
xnor UO_2678 (O_2678,N_21753,N_20744);
nor UO_2679 (O_2679,N_22813,N_22713);
and UO_2680 (O_2680,N_20991,N_23117);
and UO_2681 (O_2681,N_22810,N_20829);
or UO_2682 (O_2682,N_23506,N_20205);
nor UO_2683 (O_2683,N_24096,N_24972);
nor UO_2684 (O_2684,N_23818,N_23671);
or UO_2685 (O_2685,N_22995,N_20978);
xnor UO_2686 (O_2686,N_22753,N_22462);
xnor UO_2687 (O_2687,N_23510,N_21440);
nor UO_2688 (O_2688,N_24463,N_23727);
and UO_2689 (O_2689,N_20815,N_22634);
or UO_2690 (O_2690,N_23118,N_20523);
and UO_2691 (O_2691,N_22159,N_24264);
nor UO_2692 (O_2692,N_24457,N_22383);
nand UO_2693 (O_2693,N_22109,N_21302);
and UO_2694 (O_2694,N_23240,N_22379);
nand UO_2695 (O_2695,N_22268,N_21158);
xnor UO_2696 (O_2696,N_20308,N_20240);
and UO_2697 (O_2697,N_22864,N_21152);
nand UO_2698 (O_2698,N_20440,N_22083);
nand UO_2699 (O_2699,N_21314,N_20696);
nand UO_2700 (O_2700,N_22829,N_20032);
and UO_2701 (O_2701,N_21872,N_23795);
or UO_2702 (O_2702,N_22774,N_23617);
or UO_2703 (O_2703,N_24355,N_24635);
or UO_2704 (O_2704,N_22145,N_23899);
xnor UO_2705 (O_2705,N_24897,N_23402);
or UO_2706 (O_2706,N_24493,N_23726);
or UO_2707 (O_2707,N_20621,N_21702);
or UO_2708 (O_2708,N_20054,N_22894);
or UO_2709 (O_2709,N_20957,N_21801);
and UO_2710 (O_2710,N_23158,N_23239);
nand UO_2711 (O_2711,N_23467,N_22069);
nand UO_2712 (O_2712,N_21715,N_22940);
xor UO_2713 (O_2713,N_21323,N_22906);
or UO_2714 (O_2714,N_21840,N_21266);
nand UO_2715 (O_2715,N_20274,N_22923);
nand UO_2716 (O_2716,N_20019,N_24305);
nor UO_2717 (O_2717,N_21491,N_21451);
or UO_2718 (O_2718,N_24973,N_22393);
or UO_2719 (O_2719,N_22959,N_20827);
or UO_2720 (O_2720,N_22796,N_22314);
nand UO_2721 (O_2721,N_22971,N_22998);
or UO_2722 (O_2722,N_24360,N_23629);
nand UO_2723 (O_2723,N_24127,N_23098);
nor UO_2724 (O_2724,N_23455,N_24452);
nor UO_2725 (O_2725,N_21888,N_24793);
and UO_2726 (O_2726,N_23955,N_24500);
and UO_2727 (O_2727,N_24947,N_20290);
nand UO_2728 (O_2728,N_21768,N_21248);
xor UO_2729 (O_2729,N_24484,N_22332);
and UO_2730 (O_2730,N_24361,N_20629);
nand UO_2731 (O_2731,N_22927,N_24355);
and UO_2732 (O_2732,N_22792,N_22037);
and UO_2733 (O_2733,N_20313,N_22826);
and UO_2734 (O_2734,N_22041,N_21329);
nand UO_2735 (O_2735,N_23423,N_20235);
xnor UO_2736 (O_2736,N_24713,N_22403);
nand UO_2737 (O_2737,N_23298,N_23439);
nor UO_2738 (O_2738,N_21644,N_21067);
nand UO_2739 (O_2739,N_24436,N_21820);
nor UO_2740 (O_2740,N_22616,N_20737);
and UO_2741 (O_2741,N_21612,N_22448);
or UO_2742 (O_2742,N_22357,N_23629);
nand UO_2743 (O_2743,N_22670,N_23123);
and UO_2744 (O_2744,N_23366,N_23714);
and UO_2745 (O_2745,N_20415,N_22611);
nor UO_2746 (O_2746,N_24935,N_21938);
or UO_2747 (O_2747,N_22080,N_23505);
and UO_2748 (O_2748,N_22430,N_21091);
or UO_2749 (O_2749,N_21855,N_21782);
or UO_2750 (O_2750,N_20504,N_23500);
nor UO_2751 (O_2751,N_20929,N_20015);
or UO_2752 (O_2752,N_24490,N_21546);
and UO_2753 (O_2753,N_24907,N_20714);
nor UO_2754 (O_2754,N_20649,N_23464);
nor UO_2755 (O_2755,N_21032,N_23833);
nor UO_2756 (O_2756,N_23483,N_21973);
nand UO_2757 (O_2757,N_22467,N_23302);
nand UO_2758 (O_2758,N_23463,N_23682);
nor UO_2759 (O_2759,N_22744,N_21695);
and UO_2760 (O_2760,N_20047,N_23990);
or UO_2761 (O_2761,N_21732,N_21577);
and UO_2762 (O_2762,N_21901,N_23960);
nor UO_2763 (O_2763,N_20208,N_23482);
or UO_2764 (O_2764,N_23095,N_22641);
nor UO_2765 (O_2765,N_21284,N_22917);
nand UO_2766 (O_2766,N_20731,N_20814);
xor UO_2767 (O_2767,N_23247,N_21564);
nor UO_2768 (O_2768,N_21404,N_24299);
and UO_2769 (O_2769,N_23018,N_21455);
nor UO_2770 (O_2770,N_20254,N_24256);
nor UO_2771 (O_2771,N_20064,N_24450);
or UO_2772 (O_2772,N_21093,N_21637);
nor UO_2773 (O_2773,N_20622,N_24970);
nand UO_2774 (O_2774,N_22277,N_23164);
nor UO_2775 (O_2775,N_22937,N_23425);
nor UO_2776 (O_2776,N_22600,N_20022);
or UO_2777 (O_2777,N_22096,N_23390);
nand UO_2778 (O_2778,N_24520,N_21959);
nand UO_2779 (O_2779,N_21569,N_24431);
or UO_2780 (O_2780,N_23050,N_21705);
nand UO_2781 (O_2781,N_22214,N_23384);
and UO_2782 (O_2782,N_24747,N_20608);
nand UO_2783 (O_2783,N_21285,N_24087);
or UO_2784 (O_2784,N_23404,N_24551);
nor UO_2785 (O_2785,N_20763,N_22368);
or UO_2786 (O_2786,N_20799,N_24600);
nor UO_2787 (O_2787,N_24314,N_20703);
or UO_2788 (O_2788,N_24603,N_22120);
nand UO_2789 (O_2789,N_22798,N_22860);
nor UO_2790 (O_2790,N_23433,N_20420);
and UO_2791 (O_2791,N_22302,N_20235);
nand UO_2792 (O_2792,N_20952,N_22178);
nand UO_2793 (O_2793,N_21875,N_23237);
nor UO_2794 (O_2794,N_24396,N_21159);
or UO_2795 (O_2795,N_24755,N_22381);
nand UO_2796 (O_2796,N_21952,N_24000);
nor UO_2797 (O_2797,N_22380,N_23757);
or UO_2798 (O_2798,N_21697,N_20308);
nor UO_2799 (O_2799,N_24019,N_20693);
or UO_2800 (O_2800,N_24699,N_22046);
nor UO_2801 (O_2801,N_21724,N_20519);
and UO_2802 (O_2802,N_21939,N_23357);
nor UO_2803 (O_2803,N_24461,N_23375);
nor UO_2804 (O_2804,N_22701,N_23842);
xor UO_2805 (O_2805,N_23229,N_22813);
or UO_2806 (O_2806,N_24872,N_20630);
or UO_2807 (O_2807,N_21332,N_24666);
and UO_2808 (O_2808,N_20330,N_20824);
nor UO_2809 (O_2809,N_20204,N_23536);
or UO_2810 (O_2810,N_23173,N_20381);
nand UO_2811 (O_2811,N_22167,N_24635);
xnor UO_2812 (O_2812,N_24530,N_23856);
or UO_2813 (O_2813,N_22602,N_22119);
xnor UO_2814 (O_2814,N_20532,N_21334);
nor UO_2815 (O_2815,N_21112,N_24097);
and UO_2816 (O_2816,N_23696,N_21114);
nand UO_2817 (O_2817,N_23142,N_23789);
or UO_2818 (O_2818,N_20396,N_24328);
xor UO_2819 (O_2819,N_21822,N_24851);
nand UO_2820 (O_2820,N_24220,N_24973);
or UO_2821 (O_2821,N_20249,N_22740);
nor UO_2822 (O_2822,N_24454,N_22601);
xor UO_2823 (O_2823,N_22011,N_21508);
nand UO_2824 (O_2824,N_20918,N_20343);
nor UO_2825 (O_2825,N_20066,N_22300);
and UO_2826 (O_2826,N_23255,N_22992);
or UO_2827 (O_2827,N_22156,N_20322);
or UO_2828 (O_2828,N_24197,N_22589);
or UO_2829 (O_2829,N_20704,N_22380);
xnor UO_2830 (O_2830,N_23147,N_23178);
xnor UO_2831 (O_2831,N_23377,N_22428);
nor UO_2832 (O_2832,N_24478,N_22905);
nand UO_2833 (O_2833,N_24358,N_22843);
nand UO_2834 (O_2834,N_21749,N_21468);
xor UO_2835 (O_2835,N_23821,N_24174);
nand UO_2836 (O_2836,N_23776,N_23023);
nor UO_2837 (O_2837,N_20008,N_20540);
nand UO_2838 (O_2838,N_20146,N_21829);
or UO_2839 (O_2839,N_22333,N_23738);
or UO_2840 (O_2840,N_23153,N_23266);
and UO_2841 (O_2841,N_23565,N_24082);
or UO_2842 (O_2842,N_22351,N_21359);
and UO_2843 (O_2843,N_24139,N_22618);
and UO_2844 (O_2844,N_20926,N_22189);
nand UO_2845 (O_2845,N_20505,N_21551);
nor UO_2846 (O_2846,N_20169,N_20080);
nor UO_2847 (O_2847,N_20331,N_24686);
nand UO_2848 (O_2848,N_21120,N_20728);
xor UO_2849 (O_2849,N_24547,N_20950);
nor UO_2850 (O_2850,N_22439,N_24809);
xnor UO_2851 (O_2851,N_22811,N_24402);
or UO_2852 (O_2852,N_24534,N_22629);
xor UO_2853 (O_2853,N_23718,N_23073);
and UO_2854 (O_2854,N_24031,N_23220);
or UO_2855 (O_2855,N_22491,N_23644);
nand UO_2856 (O_2856,N_22925,N_20784);
or UO_2857 (O_2857,N_21544,N_23909);
nor UO_2858 (O_2858,N_20308,N_23792);
nand UO_2859 (O_2859,N_22250,N_21147);
nor UO_2860 (O_2860,N_20284,N_20722);
xnor UO_2861 (O_2861,N_22338,N_23971);
xnor UO_2862 (O_2862,N_22380,N_24666);
and UO_2863 (O_2863,N_21803,N_24278);
or UO_2864 (O_2864,N_24091,N_21629);
nand UO_2865 (O_2865,N_22405,N_22608);
or UO_2866 (O_2866,N_20514,N_21525);
or UO_2867 (O_2867,N_20493,N_22973);
or UO_2868 (O_2868,N_24846,N_21479);
or UO_2869 (O_2869,N_23252,N_22953);
xnor UO_2870 (O_2870,N_22577,N_24134);
nor UO_2871 (O_2871,N_23861,N_23743);
and UO_2872 (O_2872,N_24834,N_23314);
nand UO_2873 (O_2873,N_22435,N_22342);
nor UO_2874 (O_2874,N_21911,N_20672);
and UO_2875 (O_2875,N_22831,N_24955);
and UO_2876 (O_2876,N_23262,N_22568);
nor UO_2877 (O_2877,N_20723,N_24150);
or UO_2878 (O_2878,N_21127,N_20288);
nand UO_2879 (O_2879,N_23249,N_24896);
or UO_2880 (O_2880,N_20520,N_22852);
or UO_2881 (O_2881,N_20846,N_23931);
nand UO_2882 (O_2882,N_23151,N_24304);
nand UO_2883 (O_2883,N_20987,N_21958);
xnor UO_2884 (O_2884,N_23403,N_21033);
or UO_2885 (O_2885,N_24599,N_24325);
nand UO_2886 (O_2886,N_23409,N_21903);
and UO_2887 (O_2887,N_24855,N_22196);
nor UO_2888 (O_2888,N_20516,N_21920);
or UO_2889 (O_2889,N_20945,N_23251);
and UO_2890 (O_2890,N_20652,N_23877);
and UO_2891 (O_2891,N_24790,N_22303);
xnor UO_2892 (O_2892,N_21615,N_21346);
and UO_2893 (O_2893,N_20590,N_23168);
nand UO_2894 (O_2894,N_21288,N_22129);
nor UO_2895 (O_2895,N_22716,N_20391);
and UO_2896 (O_2896,N_24426,N_22998);
and UO_2897 (O_2897,N_22845,N_22825);
xor UO_2898 (O_2898,N_20963,N_22794);
xor UO_2899 (O_2899,N_21066,N_21398);
nor UO_2900 (O_2900,N_22741,N_24920);
and UO_2901 (O_2901,N_24093,N_24949);
nor UO_2902 (O_2902,N_24697,N_21260);
nand UO_2903 (O_2903,N_24552,N_24309);
or UO_2904 (O_2904,N_23080,N_21346);
xor UO_2905 (O_2905,N_20076,N_23492);
and UO_2906 (O_2906,N_22905,N_23764);
nor UO_2907 (O_2907,N_23179,N_23937);
nor UO_2908 (O_2908,N_22803,N_21996);
xor UO_2909 (O_2909,N_21519,N_21858);
nand UO_2910 (O_2910,N_24265,N_20716);
nor UO_2911 (O_2911,N_23965,N_20246);
and UO_2912 (O_2912,N_22906,N_24111);
or UO_2913 (O_2913,N_23960,N_21725);
nand UO_2914 (O_2914,N_22301,N_23827);
and UO_2915 (O_2915,N_24996,N_21522);
nand UO_2916 (O_2916,N_23754,N_22129);
xnor UO_2917 (O_2917,N_22297,N_23287);
or UO_2918 (O_2918,N_23325,N_20723);
nand UO_2919 (O_2919,N_22846,N_21802);
or UO_2920 (O_2920,N_21966,N_22775);
nor UO_2921 (O_2921,N_24082,N_22083);
and UO_2922 (O_2922,N_20249,N_22619);
or UO_2923 (O_2923,N_24802,N_21061);
xor UO_2924 (O_2924,N_20653,N_24187);
nor UO_2925 (O_2925,N_23717,N_21331);
nor UO_2926 (O_2926,N_23835,N_22447);
or UO_2927 (O_2927,N_22854,N_20480);
nor UO_2928 (O_2928,N_21265,N_24248);
nor UO_2929 (O_2929,N_23298,N_23793);
or UO_2930 (O_2930,N_24236,N_24858);
nor UO_2931 (O_2931,N_23921,N_21803);
nor UO_2932 (O_2932,N_21611,N_20427);
and UO_2933 (O_2933,N_24474,N_24990);
nor UO_2934 (O_2934,N_20238,N_20274);
xor UO_2935 (O_2935,N_22995,N_22210);
or UO_2936 (O_2936,N_23675,N_21161);
and UO_2937 (O_2937,N_24867,N_22058);
nand UO_2938 (O_2938,N_20107,N_21114);
xnor UO_2939 (O_2939,N_20167,N_22575);
and UO_2940 (O_2940,N_24670,N_23046);
xnor UO_2941 (O_2941,N_23582,N_21478);
and UO_2942 (O_2942,N_23925,N_23090);
and UO_2943 (O_2943,N_24343,N_23726);
nor UO_2944 (O_2944,N_23841,N_23673);
or UO_2945 (O_2945,N_21741,N_24947);
and UO_2946 (O_2946,N_24535,N_24896);
nor UO_2947 (O_2947,N_20815,N_23561);
or UO_2948 (O_2948,N_22654,N_22135);
or UO_2949 (O_2949,N_20743,N_20566);
or UO_2950 (O_2950,N_20009,N_21432);
or UO_2951 (O_2951,N_24427,N_21097);
nand UO_2952 (O_2952,N_23043,N_24695);
and UO_2953 (O_2953,N_23282,N_20157);
nor UO_2954 (O_2954,N_21391,N_21280);
or UO_2955 (O_2955,N_21273,N_20556);
and UO_2956 (O_2956,N_23532,N_22601);
and UO_2957 (O_2957,N_22793,N_21952);
or UO_2958 (O_2958,N_22710,N_20197);
nor UO_2959 (O_2959,N_21891,N_24660);
nand UO_2960 (O_2960,N_24019,N_20288);
nor UO_2961 (O_2961,N_21249,N_22061);
or UO_2962 (O_2962,N_21903,N_23832);
nor UO_2963 (O_2963,N_22788,N_23511);
and UO_2964 (O_2964,N_22430,N_24727);
and UO_2965 (O_2965,N_21727,N_20655);
nor UO_2966 (O_2966,N_22178,N_24683);
and UO_2967 (O_2967,N_23945,N_21149);
nor UO_2968 (O_2968,N_22726,N_21101);
nor UO_2969 (O_2969,N_24953,N_24851);
and UO_2970 (O_2970,N_20722,N_20181);
or UO_2971 (O_2971,N_20738,N_21633);
and UO_2972 (O_2972,N_21448,N_20538);
or UO_2973 (O_2973,N_20909,N_20640);
nand UO_2974 (O_2974,N_21841,N_21369);
and UO_2975 (O_2975,N_20706,N_24795);
or UO_2976 (O_2976,N_23212,N_20992);
or UO_2977 (O_2977,N_24724,N_21145);
and UO_2978 (O_2978,N_24867,N_21277);
nand UO_2979 (O_2979,N_22689,N_24880);
xnor UO_2980 (O_2980,N_20158,N_21992);
and UO_2981 (O_2981,N_22217,N_24476);
nand UO_2982 (O_2982,N_21055,N_23264);
and UO_2983 (O_2983,N_24094,N_23529);
or UO_2984 (O_2984,N_22720,N_22655);
or UO_2985 (O_2985,N_21205,N_21802);
nand UO_2986 (O_2986,N_22673,N_21313);
or UO_2987 (O_2987,N_23714,N_20099);
and UO_2988 (O_2988,N_20990,N_21267);
and UO_2989 (O_2989,N_24571,N_20347);
and UO_2990 (O_2990,N_22608,N_20593);
nor UO_2991 (O_2991,N_22663,N_21649);
nor UO_2992 (O_2992,N_23950,N_23191);
xnor UO_2993 (O_2993,N_20722,N_22959);
or UO_2994 (O_2994,N_23949,N_21038);
nor UO_2995 (O_2995,N_24535,N_21707);
nor UO_2996 (O_2996,N_21456,N_21119);
nand UO_2997 (O_2997,N_21757,N_21203);
nor UO_2998 (O_2998,N_20336,N_22177);
or UO_2999 (O_2999,N_23329,N_22149);
endmodule