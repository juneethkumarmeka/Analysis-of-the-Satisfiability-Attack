module basic_3000_30000_3500_3_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20004,N_20006,N_20007,N_20009,N_20012,N_20013,N_20014,N_20016,N_20017,N_20020,N_20021,N_20024,N_20026,N_20027,N_20031,N_20032,N_20034,N_20035,N_20036,N_20040,N_20041,N_20042,N_20043,N_20044,N_20046,N_20047,N_20048,N_20049,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20066,N_20067,N_20069,N_20071,N_20072,N_20073,N_20074,N_20076,N_20077,N_20079,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20092,N_20093,N_20095,N_20096,N_20097,N_20098,N_20099,N_20101,N_20102,N_20103,N_20104,N_20105,N_20107,N_20108,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20118,N_20119,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20136,N_20137,N_20138,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20161,N_20162,N_20164,N_20165,N_20166,N_20167,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20176,N_20177,N_20178,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20192,N_20194,N_20197,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20210,N_20211,N_20212,N_20216,N_20217,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20230,N_20231,N_20232,N_20233,N_20235,N_20236,N_20237,N_20238,N_20241,N_20242,N_20243,N_20244,N_20246,N_20247,N_20248,N_20250,N_20251,N_20252,N_20253,N_20254,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20263,N_20264,N_20267,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20278,N_20280,N_20282,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20291,N_20292,N_20293,N_20294,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20320,N_20323,N_20325,N_20326,N_20327,N_20328,N_20329,N_20331,N_20332,N_20334,N_20335,N_20337,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20346,N_20347,N_20349,N_20350,N_20351,N_20354,N_20355,N_20356,N_20357,N_20358,N_20360,N_20362,N_20363,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20377,N_20379,N_20380,N_20381,N_20382,N_20384,N_20385,N_20388,N_20390,N_20391,N_20392,N_20393,N_20395,N_20400,N_20403,N_20404,N_20406,N_20407,N_20410,N_20411,N_20413,N_20414,N_20415,N_20417,N_20419,N_20421,N_20422,N_20424,N_20425,N_20426,N_20427,N_20429,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20438,N_20439,N_20440,N_20443,N_20445,N_20446,N_20447,N_20448,N_20450,N_20451,N_20453,N_20454,N_20455,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20466,N_20468,N_20469,N_20470,N_20472,N_20473,N_20474,N_20479,N_20481,N_20482,N_20484,N_20485,N_20487,N_20488,N_20489,N_20491,N_20493,N_20494,N_20497,N_20500,N_20502,N_20503,N_20504,N_20505,N_20507,N_20509,N_20511,N_20513,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20529,N_20531,N_20532,N_20533,N_20534,N_20536,N_20538,N_20539,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20549,N_20550,N_20552,N_20553,N_20555,N_20556,N_20557,N_20558,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20579,N_20580,N_20582,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20604,N_20605,N_20606,N_20608,N_20611,N_20612,N_20619,N_20621,N_20622,N_20623,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20653,N_20655,N_20656,N_20657,N_20658,N_20659,N_20661,N_20662,N_20663,N_20664,N_20666,N_20668,N_20670,N_20672,N_20673,N_20675,N_20676,N_20677,N_20679,N_20680,N_20681,N_20683,N_20684,N_20685,N_20687,N_20688,N_20690,N_20692,N_20693,N_20694,N_20695,N_20697,N_20698,N_20701,N_20702,N_20704,N_20705,N_20706,N_20707,N_20709,N_20712,N_20713,N_20714,N_20716,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20725,N_20726,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20744,N_20746,N_20747,N_20748,N_20749,N_20751,N_20753,N_20755,N_20756,N_20758,N_20760,N_20761,N_20762,N_20763,N_20764,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20786,N_20787,N_20789,N_20790,N_20791,N_20793,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20805,N_20808,N_20809,N_20810,N_20811,N_20812,N_20814,N_20815,N_20817,N_20818,N_20819,N_20821,N_20823,N_20825,N_20826,N_20827,N_20828,N_20830,N_20832,N_20833,N_20836,N_20837,N_20838,N_20839,N_20840,N_20843,N_20844,N_20846,N_20847,N_20848,N_20849,N_20850,N_20852,N_20853,N_20855,N_20857,N_20859,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20874,N_20876,N_20878,N_20880,N_20881,N_20883,N_20885,N_20886,N_20887,N_20888,N_20890,N_20891,N_20892,N_20893,N_20895,N_20896,N_20897,N_20900,N_20902,N_20903,N_20906,N_20908,N_20909,N_20910,N_20911,N_20913,N_20914,N_20916,N_20917,N_20918,N_20920,N_20921,N_20923,N_20924,N_20926,N_20927,N_20928,N_20930,N_20932,N_20933,N_20934,N_20936,N_20937,N_20938,N_20939,N_20941,N_20945,N_20946,N_20947,N_20948,N_20949,N_20951,N_20952,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20964,N_20965,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20976,N_20977,N_20978,N_20980,N_20981,N_20982,N_20983,N_20986,N_20987,N_20988,N_20990,N_20993,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21003,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21034,N_21036,N_21037,N_21038,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21050,N_21051,N_21052,N_21054,N_21057,N_21058,N_21060,N_21061,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21077,N_21078,N_21079,N_21080,N_21082,N_21084,N_21086,N_21087,N_21089,N_21090,N_21091,N_21092,N_21094,N_21095,N_21096,N_21098,N_21099,N_21100,N_21101,N_21103,N_21105,N_21107,N_21109,N_21110,N_21111,N_21114,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21127,N_21128,N_21130,N_21134,N_21135,N_21137,N_21139,N_21140,N_21141,N_21142,N_21143,N_21145,N_21146,N_21147,N_21148,N_21151,N_21152,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21166,N_21167,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21178,N_21182,N_21183,N_21184,N_21186,N_21188,N_21189,N_21190,N_21191,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21205,N_21206,N_21208,N_21209,N_21210,N_21211,N_21212,N_21214,N_21215,N_21216,N_21219,N_21221,N_21222,N_21223,N_21224,N_21225,N_21227,N_21228,N_21229,N_21233,N_21234,N_21235,N_21236,N_21238,N_21239,N_21240,N_21243,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21254,N_21255,N_21258,N_21261,N_21266,N_21268,N_21269,N_21270,N_21271,N_21272,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21286,N_21287,N_21288,N_21289,N_21290,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21299,N_21300,N_21301,N_21302,N_21304,N_21305,N_21307,N_21308,N_21309,N_21311,N_21312,N_21313,N_21315,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21327,N_21328,N_21329,N_21330,N_21333,N_21335,N_21337,N_21338,N_21340,N_21342,N_21343,N_21344,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21359,N_21360,N_21361,N_21362,N_21365,N_21366,N_21367,N_21369,N_21370,N_21373,N_21374,N_21375,N_21376,N_21377,N_21379,N_21380,N_21381,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21416,N_21420,N_21421,N_21422,N_21423,N_21424,N_21426,N_21427,N_21428,N_21429,N_21432,N_21433,N_21434,N_21435,N_21436,N_21438,N_21439,N_21440,N_21442,N_21444,N_21445,N_21446,N_21450,N_21453,N_21454,N_21456,N_21457,N_21459,N_21460,N_21461,N_21462,N_21464,N_21465,N_21468,N_21469,N_21470,N_21471,N_21473,N_21474,N_21475,N_21477,N_21478,N_21479,N_21480,N_21481,N_21484,N_21485,N_21487,N_21488,N_21489,N_21490,N_21492,N_21493,N_21496,N_21497,N_21498,N_21499,N_21501,N_21502,N_21505,N_21507,N_21508,N_21509,N_21511,N_21512,N_21514,N_21516,N_21517,N_21522,N_21524,N_21525,N_21526,N_21527,N_21528,N_21530,N_21531,N_21532,N_21533,N_21536,N_21537,N_21539,N_21540,N_21542,N_21544,N_21545,N_21546,N_21547,N_21549,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21563,N_21564,N_21566,N_21567,N_21569,N_21570,N_21571,N_21574,N_21575,N_21576,N_21578,N_21579,N_21584,N_21585,N_21586,N_21587,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21598,N_21599,N_21601,N_21602,N_21604,N_21605,N_21606,N_21607,N_21608,N_21610,N_21611,N_21612,N_21613,N_21614,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21624,N_21625,N_21626,N_21628,N_21630,N_21631,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21641,N_21642,N_21643,N_21644,N_21647,N_21648,N_21649,N_21650,N_21651,N_21653,N_21655,N_21656,N_21658,N_21660,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21683,N_21684,N_21685,N_21686,N_21687,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21697,N_21698,N_21700,N_21701,N_21703,N_21704,N_21707,N_21709,N_21711,N_21714,N_21715,N_21717,N_21719,N_21720,N_21721,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21731,N_21732,N_21733,N_21734,N_21738,N_21740,N_21741,N_21745,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21758,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21767,N_21768,N_21769,N_21770,N_21772,N_21773,N_21774,N_21775,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21787,N_21788,N_21790,N_21791,N_21793,N_21794,N_21795,N_21797,N_21798,N_21800,N_21802,N_21803,N_21805,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21816,N_21818,N_21819,N_21822,N_21825,N_21828,N_21829,N_21831,N_21832,N_21833,N_21834,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21844,N_21846,N_21849,N_21850,N_21852,N_21856,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21868,N_21869,N_21870,N_21872,N_21873,N_21874,N_21875,N_21876,N_21878,N_21881,N_21885,N_21886,N_21888,N_21889,N_21890,N_21891,N_21892,N_21894,N_21896,N_21898,N_21899,N_21900,N_21901,N_21903,N_21904,N_21905,N_21906,N_21907,N_21909,N_21910,N_21911,N_21913,N_21914,N_21915,N_21917,N_21919,N_21920,N_21921,N_21922,N_21923,N_21926,N_21927,N_21930,N_21931,N_21932,N_21935,N_21936,N_21938,N_21939,N_21941,N_21942,N_21943,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21963,N_21964,N_21965,N_21966,N_21968,N_21970,N_21971,N_21972,N_21975,N_21976,N_21977,N_21980,N_21981,N_21983,N_21985,N_21988,N_21989,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21998,N_22000,N_22001,N_22002,N_22004,N_22005,N_22006,N_22008,N_22009,N_22011,N_22012,N_22013,N_22014,N_22015,N_22017,N_22018,N_22019,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22028,N_22029,N_22030,N_22034,N_22035,N_22037,N_22038,N_22039,N_22041,N_22043,N_22045,N_22046,N_22047,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22059,N_22060,N_22061,N_22063,N_22064,N_22065,N_22068,N_22069,N_22070,N_22074,N_22075,N_22076,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22088,N_22092,N_22093,N_22094,N_22095,N_22096,N_22098,N_22099,N_22100,N_22103,N_22104,N_22107,N_22108,N_22109,N_22110,N_22113,N_22114,N_22115,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22127,N_22128,N_22130,N_22131,N_22132,N_22134,N_22135,N_22136,N_22138,N_22139,N_22140,N_22141,N_22144,N_22145,N_22147,N_22150,N_22151,N_22153,N_22156,N_22158,N_22159,N_22161,N_22163,N_22165,N_22167,N_22169,N_22170,N_22172,N_22174,N_22175,N_22176,N_22177,N_22179,N_22181,N_22182,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22192,N_22193,N_22194,N_22196,N_22197,N_22198,N_22200,N_22203,N_22205,N_22207,N_22208,N_22211,N_22212,N_22213,N_22215,N_22216,N_22217,N_22218,N_22220,N_22222,N_22223,N_22224,N_22225,N_22226,N_22228,N_22229,N_22230,N_22231,N_22233,N_22236,N_22237,N_22238,N_22239,N_22241,N_22242,N_22243,N_22245,N_22246,N_22247,N_22250,N_22251,N_22254,N_22255,N_22256,N_22259,N_22260,N_22261,N_22262,N_22264,N_22265,N_22266,N_22269,N_22272,N_22273,N_22274,N_22276,N_22277,N_22278,N_22281,N_22282,N_22284,N_22285,N_22286,N_22287,N_22289,N_22291,N_22292,N_22295,N_22297,N_22298,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22308,N_22309,N_22311,N_22312,N_22313,N_22314,N_22316,N_22317,N_22320,N_22321,N_22322,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22335,N_22336,N_22338,N_22339,N_22341,N_22342,N_22343,N_22345,N_22346,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22357,N_22358,N_22359,N_22360,N_22364,N_22366,N_22367,N_22368,N_22372,N_22373,N_22375,N_22376,N_22379,N_22384,N_22385,N_22386,N_22387,N_22388,N_22390,N_22392,N_22393,N_22394,N_22396,N_22397,N_22398,N_22399,N_22402,N_22404,N_22405,N_22407,N_22409,N_22410,N_22412,N_22413,N_22416,N_22417,N_22418,N_22420,N_22422,N_22424,N_22426,N_22427,N_22429,N_22430,N_22433,N_22434,N_22436,N_22438,N_22439,N_22440,N_22441,N_22442,N_22444,N_22447,N_22448,N_22451,N_22455,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22483,N_22484,N_22486,N_22487,N_22488,N_22490,N_22492,N_22493,N_22494,N_22496,N_22497,N_22500,N_22502,N_22504,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22520,N_22521,N_22522,N_22523,N_22524,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22539,N_22540,N_22542,N_22545,N_22546,N_22547,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22579,N_22580,N_22581,N_22583,N_22584,N_22585,N_22586,N_22587,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22597,N_22599,N_22600,N_22601,N_22604,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22615,N_22617,N_22620,N_22621,N_22623,N_22624,N_22625,N_22627,N_22629,N_22630,N_22631,N_22632,N_22634,N_22635,N_22636,N_22637,N_22639,N_22641,N_22642,N_22645,N_22646,N_22648,N_22649,N_22650,N_22651,N_22653,N_22656,N_22658,N_22659,N_22661,N_22662,N_22663,N_22665,N_22666,N_22668,N_22669,N_22670,N_22673,N_22675,N_22676,N_22678,N_22679,N_22680,N_22681,N_22683,N_22684,N_22685,N_22688,N_22689,N_22690,N_22692,N_22694,N_22695,N_22697,N_22699,N_22700,N_22704,N_22705,N_22706,N_22707,N_22711,N_22712,N_22713,N_22714,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22723,N_22724,N_22725,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22739,N_22740,N_22741,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22756,N_22757,N_22759,N_22760,N_22762,N_22764,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22774,N_22775,N_22776,N_22778,N_22779,N_22783,N_22784,N_22785,N_22787,N_22788,N_22790,N_22792,N_22793,N_22795,N_22796,N_22797,N_22798,N_22799,N_22801,N_22802,N_22803,N_22805,N_22806,N_22807,N_22808,N_22811,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22820,N_22821,N_22822,N_22823,N_22825,N_22827,N_22828,N_22830,N_22831,N_22832,N_22835,N_22836,N_22837,N_22840,N_22841,N_22844,N_22845,N_22846,N_22847,N_22849,N_22850,N_22851,N_22852,N_22853,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22866,N_22867,N_22869,N_22870,N_22871,N_22874,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22890,N_22891,N_22892,N_22894,N_22895,N_22896,N_22897,N_22900,N_22901,N_22902,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22914,N_22915,N_22917,N_22918,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22929,N_22931,N_22932,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22945,N_22947,N_22949,N_22950,N_22951,N_22952,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22983,N_22984,N_22985,N_22986,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22999,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23010,N_23011,N_23012,N_23016,N_23017,N_23018,N_23020,N_23022,N_23023,N_23024,N_23025,N_23026,N_23029,N_23030,N_23031,N_23033,N_23034,N_23041,N_23042,N_23044,N_23045,N_23047,N_23049,N_23052,N_23053,N_23057,N_23059,N_23060,N_23062,N_23066,N_23067,N_23068,N_23069,N_23070,N_23077,N_23078,N_23081,N_23083,N_23084,N_23087,N_23088,N_23089,N_23090,N_23091,N_23093,N_23094,N_23095,N_23096,N_23097,N_23099,N_23100,N_23103,N_23104,N_23105,N_23106,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23124,N_23125,N_23126,N_23127,N_23128,N_23130,N_23131,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23153,N_23154,N_23156,N_23157,N_23158,N_23159,N_23161,N_23162,N_23165,N_23168,N_23169,N_23171,N_23172,N_23174,N_23175,N_23177,N_23178,N_23179,N_23180,N_23182,N_23183,N_23185,N_23186,N_23187,N_23188,N_23189,N_23191,N_23193,N_23194,N_23196,N_23197,N_23199,N_23200,N_23201,N_23202,N_23204,N_23205,N_23206,N_23208,N_23209,N_23210,N_23211,N_23212,N_23216,N_23217,N_23218,N_23219,N_23220,N_23222,N_23223,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23241,N_23242,N_23244,N_23246,N_23247,N_23248,N_23249,N_23251,N_23252,N_23255,N_23256,N_23258,N_23260,N_23261,N_23262,N_23263,N_23265,N_23266,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23283,N_23284,N_23285,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23297,N_23298,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23311,N_23312,N_23313,N_23314,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23327,N_23331,N_23336,N_23338,N_23342,N_23343,N_23345,N_23347,N_23349,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23361,N_23362,N_23363,N_23364,N_23368,N_23369,N_23371,N_23373,N_23374,N_23376,N_23378,N_23379,N_23380,N_23382,N_23383,N_23386,N_23387,N_23388,N_23389,N_23390,N_23393,N_23394,N_23395,N_23397,N_23398,N_23400,N_23401,N_23403,N_23404,N_23405,N_23407,N_23408,N_23409,N_23411,N_23412,N_23413,N_23414,N_23415,N_23418,N_23419,N_23420,N_23424,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23434,N_23435,N_23438,N_23439,N_23441,N_23442,N_23443,N_23446,N_23448,N_23449,N_23450,N_23451,N_23452,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23470,N_23471,N_23472,N_23473,N_23474,N_23476,N_23477,N_23478,N_23479,N_23481,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23497,N_23498,N_23499,N_23501,N_23503,N_23504,N_23505,N_23508,N_23509,N_23510,N_23511,N_23512,N_23514,N_23516,N_23517,N_23518,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23546,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23557,N_23559,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23568,N_23570,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23579,N_23580,N_23582,N_23583,N_23584,N_23585,N_23587,N_23589,N_23590,N_23591,N_23592,N_23594,N_23595,N_23596,N_23597,N_23598,N_23600,N_23602,N_23604,N_23605,N_23606,N_23607,N_23608,N_23610,N_23613,N_23614,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23624,N_23625,N_23629,N_23630,N_23632,N_23633,N_23636,N_23637,N_23638,N_23639,N_23641,N_23642,N_23644,N_23645,N_23646,N_23647,N_23648,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23658,N_23659,N_23661,N_23662,N_23663,N_23666,N_23667,N_23668,N_23669,N_23672,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23695,N_23698,N_23699,N_23701,N_23702,N_23704,N_23705,N_23707,N_23708,N_23709,N_23710,N_23711,N_23713,N_23715,N_23716,N_23717,N_23719,N_23721,N_23722,N_23723,N_23724,N_23725,N_23727,N_23729,N_23731,N_23732,N_23733,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23744,N_23745,N_23749,N_23750,N_23751,N_23755,N_23756,N_23758,N_23760,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23769,N_23771,N_23772,N_23773,N_23775,N_23776,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23786,N_23787,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23799,N_23801,N_23803,N_23804,N_23806,N_23807,N_23808,N_23814,N_23815,N_23816,N_23817,N_23819,N_23820,N_23821,N_23822,N_23825,N_23826,N_23827,N_23829,N_23830,N_23832,N_23833,N_23835,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23847,N_23850,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23861,N_23862,N_23863,N_23864,N_23865,N_23867,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23896,N_23897,N_23898,N_23899,N_23901,N_23902,N_23903,N_23905,N_23906,N_23907,N_23908,N_23909,N_23911,N_23914,N_23915,N_23916,N_23917,N_23919,N_23921,N_23924,N_23927,N_23928,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23941,N_23942,N_23943,N_23945,N_23946,N_23947,N_23948,N_23951,N_23952,N_23953,N_23955,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23966,N_23967,N_23968,N_23969,N_23970,N_23972,N_23975,N_23976,N_23978,N_23980,N_23981,N_23983,N_23984,N_23985,N_23987,N_23988,N_23990,N_23991,N_23992,N_23994,N_23997,N_24000,N_24001,N_24003,N_24004,N_24007,N_24008,N_24009,N_24010,N_24011,N_24013,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24023,N_24025,N_24027,N_24031,N_24034,N_24035,N_24036,N_24037,N_24038,N_24040,N_24041,N_24043,N_24045,N_24047,N_24048,N_24049,N_24051,N_24052,N_24053,N_24054,N_24055,N_24058,N_24059,N_24060,N_24062,N_24063,N_24064,N_24065,N_24066,N_24068,N_24072,N_24073,N_24074,N_24076,N_24077,N_24081,N_24085,N_24086,N_24088,N_24089,N_24090,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24099,N_24101,N_24102,N_24104,N_24105,N_24107,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24141,N_24143,N_24144,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24159,N_24160,N_24162,N_24163,N_24164,N_24166,N_24167,N_24168,N_24169,N_24170,N_24172,N_24174,N_24177,N_24178,N_24179,N_24180,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24199,N_24200,N_24202,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24227,N_24228,N_24230,N_24231,N_24232,N_24233,N_24235,N_24236,N_24238,N_24239,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24249,N_24250,N_24251,N_24252,N_24254,N_24255,N_24257,N_24258,N_24260,N_24262,N_24263,N_24264,N_24266,N_24267,N_24268,N_24270,N_24273,N_24274,N_24275,N_24276,N_24278,N_24279,N_24280,N_24284,N_24286,N_24288,N_24289,N_24290,N_24292,N_24293,N_24294,N_24295,N_24296,N_24301,N_24303,N_24304,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24318,N_24320,N_24321,N_24322,N_24323,N_24324,N_24327,N_24329,N_24330,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24356,N_24357,N_24359,N_24360,N_24361,N_24363,N_24364,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24383,N_24385,N_24387,N_24388,N_24390,N_24391,N_24392,N_24393,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24404,N_24405,N_24406,N_24407,N_24409,N_24413,N_24414,N_24415,N_24417,N_24419,N_24420,N_24421,N_24422,N_24423,N_24425,N_24427,N_24428,N_24429,N_24430,N_24432,N_24433,N_24434,N_24435,N_24436,N_24438,N_24439,N_24440,N_24442,N_24445,N_24447,N_24449,N_24450,N_24452,N_24454,N_24455,N_24456,N_24458,N_24460,N_24462,N_24463,N_24464,N_24466,N_24467,N_24468,N_24469,N_24473,N_24474,N_24475,N_24476,N_24480,N_24482,N_24483,N_24484,N_24485,N_24487,N_24489,N_24490,N_24492,N_24493,N_24496,N_24497,N_24498,N_24499,N_24501,N_24502,N_24504,N_24506,N_24507,N_24508,N_24509,N_24510,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24520,N_24521,N_24522,N_24523,N_24524,N_24526,N_24527,N_24528,N_24529,N_24530,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24541,N_24542,N_24543,N_24544,N_24545,N_24547,N_24548,N_24551,N_24552,N_24553,N_24555,N_24556,N_24557,N_24558,N_24559,N_24561,N_24562,N_24563,N_24566,N_24567,N_24569,N_24571,N_24572,N_24574,N_24575,N_24576,N_24578,N_24579,N_24580,N_24581,N_24583,N_24584,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24602,N_24603,N_24604,N_24605,N_24608,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24617,N_24618,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24650,N_24652,N_24654,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24665,N_24667,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24684,N_24686,N_24687,N_24689,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24708,N_24709,N_24710,N_24712,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24725,N_24727,N_24731,N_24733,N_24734,N_24737,N_24739,N_24741,N_24742,N_24744,N_24745,N_24746,N_24747,N_24749,N_24750,N_24751,N_24753,N_24755,N_24758,N_24759,N_24760,N_24762,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24773,N_24775,N_24776,N_24777,N_24779,N_24780,N_24781,N_24783,N_24784,N_24785,N_24786,N_24787,N_24790,N_24792,N_24793,N_24795,N_24796,N_24798,N_24799,N_24803,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24838,N_24840,N_24842,N_24843,N_24846,N_24847,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24868,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24880,N_24881,N_24883,N_24884,N_24885,N_24886,N_24889,N_24891,N_24893,N_24894,N_24896,N_24897,N_24898,N_24899,N_24902,N_24904,N_24905,N_24906,N_24907,N_24908,N_24910,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24922,N_24925,N_24926,N_24928,N_24929,N_24930,N_24931,N_24932,N_24934,N_24936,N_24937,N_24938,N_24939,N_24940,N_24942,N_24943,N_24944,N_24947,N_24948,N_24949,N_24951,N_24952,N_24954,N_24956,N_24957,N_24962,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24973,N_24974,N_24975,N_24976,N_24978,N_24979,N_24980,N_24982,N_24983,N_24984,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24994,N_24995,N_24996,N_24997,N_24998,N_25000,N_25001,N_25003,N_25004,N_25005,N_25006,N_25008,N_25010,N_25012,N_25013,N_25014,N_25015,N_25018,N_25019,N_25020,N_25021,N_25022,N_25024,N_25026,N_25027,N_25028,N_25029,N_25032,N_25033,N_25035,N_25036,N_25037,N_25038,N_25039,N_25041,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25054,N_25055,N_25056,N_25058,N_25059,N_25061,N_25062,N_25064,N_25066,N_25067,N_25068,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25081,N_25083,N_25084,N_25085,N_25087,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25097,N_25100,N_25101,N_25102,N_25103,N_25104,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25122,N_25123,N_25125,N_25128,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25138,N_25141,N_25142,N_25144,N_25145,N_25146,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25165,N_25167,N_25168,N_25170,N_25171,N_25173,N_25174,N_25176,N_25177,N_25178,N_25179,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25194,N_25195,N_25196,N_25197,N_25198,N_25202,N_25203,N_25205,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25219,N_25220,N_25222,N_25223,N_25227,N_25232,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25244,N_25245,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25256,N_25258,N_25261,N_25262,N_25265,N_25266,N_25269,N_25270,N_25271,N_25272,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25282,N_25283,N_25285,N_25286,N_25287,N_25288,N_25290,N_25291,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25300,N_25301,N_25304,N_25305,N_25306,N_25307,N_25310,N_25311,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25321,N_25322,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25331,N_25333,N_25335,N_25336,N_25339,N_25340,N_25342,N_25344,N_25345,N_25346,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25359,N_25361,N_25362,N_25363,N_25366,N_25368,N_25369,N_25371,N_25372,N_25374,N_25375,N_25377,N_25379,N_25381,N_25382,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25395,N_25396,N_25397,N_25398,N_25401,N_25402,N_25404,N_25409,N_25411,N_25412,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25435,N_25441,N_25443,N_25445,N_25446,N_25448,N_25449,N_25451,N_25452,N_25453,N_25454,N_25455,N_25457,N_25458,N_25459,N_25461,N_25462,N_25467,N_25468,N_25469,N_25472,N_25473,N_25474,N_25475,N_25476,N_25478,N_25480,N_25481,N_25484,N_25486,N_25487,N_25489,N_25494,N_25495,N_25497,N_25498,N_25499,N_25500,N_25501,N_25503,N_25504,N_25507,N_25508,N_25509,N_25510,N_25511,N_25513,N_25515,N_25519,N_25520,N_25521,N_25522,N_25523,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25537,N_25538,N_25539,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25549,N_25550,N_25551,N_25555,N_25557,N_25558,N_25560,N_25561,N_25562,N_25563,N_25566,N_25567,N_25568,N_25570,N_25572,N_25573,N_25574,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25586,N_25587,N_25588,N_25589,N_25590,N_25594,N_25595,N_25597,N_25598,N_25600,N_25601,N_25603,N_25604,N_25607,N_25608,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25628,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25641,N_25642,N_25643,N_25645,N_25646,N_25648,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25657,N_25658,N_25659,N_25660,N_25662,N_25663,N_25664,N_25666,N_25669,N_25670,N_25672,N_25673,N_25674,N_25675,N_25677,N_25679,N_25681,N_25683,N_25684,N_25685,N_25687,N_25688,N_25690,N_25691,N_25692,N_25693,N_25695,N_25697,N_25698,N_25699,N_25701,N_25703,N_25705,N_25706,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25725,N_25726,N_25727,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25752,N_25753,N_25754,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25769,N_25771,N_25772,N_25774,N_25775,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25796,N_25797,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25807,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25817,N_25819,N_25820,N_25821,N_25822,N_25823,N_25825,N_25826,N_25827,N_25829,N_25832,N_25834,N_25836,N_25837,N_25838,N_25841,N_25842,N_25843,N_25844,N_25847,N_25849,N_25850,N_25851,N_25854,N_25855,N_25856,N_25857,N_25859,N_25860,N_25862,N_25863,N_25865,N_25866,N_25867,N_25869,N_25870,N_25873,N_25874,N_25877,N_25878,N_25879,N_25880,N_25883,N_25884,N_25885,N_25886,N_25887,N_25889,N_25891,N_25893,N_25896,N_25898,N_25899,N_25900,N_25901,N_25907,N_25909,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25921,N_25924,N_25925,N_25927,N_25928,N_25929,N_25930,N_25931,N_25933,N_25934,N_25935,N_25937,N_25939,N_25941,N_25949,N_25950,N_25951,N_25953,N_25954,N_25956,N_25957,N_25959,N_25961,N_25962,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25971,N_25973,N_25975,N_25976,N_25977,N_25979,N_25980,N_25982,N_25986,N_25987,N_25990,N_25991,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_26000,N_26001,N_26002,N_26004,N_26006,N_26008,N_26009,N_26011,N_26012,N_26014,N_26015,N_26017,N_26018,N_26021,N_26022,N_26024,N_26025,N_26026,N_26027,N_26030,N_26031,N_26034,N_26035,N_26036,N_26037,N_26039,N_26040,N_26042,N_26043,N_26044,N_26046,N_26047,N_26049,N_26050,N_26052,N_26055,N_26056,N_26057,N_26059,N_26060,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26072,N_26073,N_26074,N_26078,N_26083,N_26084,N_26085,N_26087,N_26090,N_26092,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26105,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26116,N_26117,N_26118,N_26120,N_26121,N_26123,N_26125,N_26126,N_26127,N_26130,N_26131,N_26132,N_26133,N_26135,N_26138,N_26139,N_26142,N_26143,N_26145,N_26146,N_26147,N_26149,N_26150,N_26152,N_26154,N_26156,N_26159,N_26160,N_26161,N_26163,N_26164,N_26165,N_26166,N_26167,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26186,N_26187,N_26188,N_26189,N_26191,N_26193,N_26195,N_26197,N_26200,N_26201,N_26202,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26216,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26227,N_26230,N_26232,N_26233,N_26234,N_26236,N_26237,N_26238,N_26239,N_26240,N_26243,N_26246,N_26247,N_26251,N_26252,N_26253,N_26255,N_26256,N_26257,N_26259,N_26261,N_26262,N_26264,N_26265,N_26266,N_26267,N_26269,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26281,N_26282,N_26283,N_26284,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26293,N_26296,N_26297,N_26303,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26334,N_26336,N_26337,N_26338,N_26339,N_26341,N_26342,N_26343,N_26344,N_26349,N_26350,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26360,N_26361,N_26362,N_26364,N_26366,N_26367,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26379,N_26380,N_26381,N_26383,N_26385,N_26386,N_26387,N_26389,N_26390,N_26391,N_26392,N_26396,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26423,N_26424,N_26425,N_26426,N_26427,N_26429,N_26430,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26445,N_26446,N_26447,N_26451,N_26454,N_26455,N_26456,N_26458,N_26459,N_26460,N_26461,N_26462,N_26464,N_26467,N_26468,N_26469,N_26471,N_26472,N_26475,N_26477,N_26479,N_26481,N_26482,N_26483,N_26485,N_26486,N_26488,N_26489,N_26490,N_26491,N_26494,N_26495,N_26496,N_26498,N_26500,N_26501,N_26502,N_26506,N_26507,N_26508,N_26509,N_26510,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26519,N_26520,N_26521,N_26522,N_26524,N_26525,N_26526,N_26528,N_26530,N_26531,N_26532,N_26533,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26544,N_26548,N_26549,N_26550,N_26551,N_26552,N_26554,N_26556,N_26557,N_26559,N_26560,N_26561,N_26562,N_26564,N_26566,N_26567,N_26570,N_26571,N_26573,N_26574,N_26577,N_26578,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26593,N_26594,N_26595,N_26596,N_26597,N_26599,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26609,N_26611,N_26612,N_26615,N_26616,N_26619,N_26622,N_26626,N_26627,N_26628,N_26629,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26641,N_26642,N_26643,N_26644,N_26645,N_26647,N_26648,N_26651,N_26652,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26663,N_26665,N_26666,N_26667,N_26670,N_26672,N_26673,N_26674,N_26675,N_26677,N_26678,N_26680,N_26681,N_26683,N_26684,N_26685,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26699,N_26700,N_26701,N_26703,N_26707,N_26708,N_26709,N_26712,N_26713,N_26714,N_26715,N_26717,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26729,N_26731,N_26733,N_26735,N_26736,N_26737,N_26739,N_26740,N_26741,N_26743,N_26744,N_26745,N_26746,N_26748,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26759,N_26760,N_26762,N_26764,N_26765,N_26767,N_26769,N_26770,N_26771,N_26774,N_26775,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26798,N_26799,N_26803,N_26805,N_26806,N_26807,N_26809,N_26811,N_26813,N_26814,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26831,N_26832,N_26835,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26847,N_26848,N_26849,N_26851,N_26852,N_26854,N_26855,N_26856,N_26858,N_26859,N_26860,N_26861,N_26862,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26879,N_26880,N_26881,N_26882,N_26883,N_26885,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26898,N_26900,N_26901,N_26902,N_26904,N_26905,N_26910,N_26912,N_26913,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26941,N_26944,N_26945,N_26946,N_26947,N_26949,N_26950,N_26951,N_26952,N_26953,N_26958,N_26959,N_26960,N_26962,N_26963,N_26964,N_26966,N_26967,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26980,N_26981,N_26983,N_26984,N_26986,N_26987,N_26990,N_26992,N_26993,N_26995,N_26998,N_26999,N_27000,N_27001,N_27002,N_27004,N_27006,N_27007,N_27008,N_27009,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27020,N_27022,N_27023,N_27025,N_27027,N_27029,N_27030,N_27031,N_27032,N_27034,N_27035,N_27036,N_27038,N_27039,N_27040,N_27042,N_27044,N_27045,N_27046,N_27047,N_27048,N_27050,N_27051,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27064,N_27065,N_27067,N_27070,N_27071,N_27072,N_27073,N_27074,N_27077,N_27078,N_27083,N_27086,N_27089,N_27091,N_27092,N_27094,N_27095,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27104,N_27106,N_27107,N_27109,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27119,N_27122,N_27124,N_27125,N_27126,N_27127,N_27132,N_27133,N_27135,N_27137,N_27140,N_27141,N_27142,N_27143,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27159,N_27160,N_27162,N_27165,N_27167,N_27168,N_27169,N_27170,N_27172,N_27175,N_27177,N_27179,N_27181,N_27184,N_27185,N_27187,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27201,N_27202,N_27204,N_27205,N_27208,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27219,N_27221,N_27222,N_27223,N_27226,N_27228,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27241,N_27243,N_27244,N_27245,N_27246,N_27249,N_27250,N_27251,N_27253,N_27254,N_27255,N_27257,N_27258,N_27259,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27271,N_27272,N_27274,N_27275,N_27276,N_27277,N_27278,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27288,N_27289,N_27290,N_27292,N_27296,N_27297,N_27299,N_27300,N_27302,N_27303,N_27304,N_27305,N_27307,N_27309,N_27310,N_27311,N_27312,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27325,N_27326,N_27327,N_27330,N_27331,N_27332,N_27333,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27363,N_27366,N_27367,N_27368,N_27371,N_27372,N_27373,N_27376,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27386,N_27388,N_27389,N_27390,N_27391,N_27394,N_27395,N_27396,N_27397,N_27401,N_27403,N_27404,N_27405,N_27406,N_27408,N_27410,N_27411,N_27413,N_27415,N_27417,N_27418,N_27420,N_27421,N_27422,N_27424,N_27425,N_27426,N_27428,N_27431,N_27432,N_27433,N_27435,N_27436,N_27437,N_27438,N_27440,N_27441,N_27443,N_27444,N_27446,N_27447,N_27449,N_27451,N_27452,N_27453,N_27455,N_27457,N_27458,N_27459,N_27462,N_27464,N_27465,N_27467,N_27468,N_27469,N_27471,N_27472,N_27473,N_27478,N_27482,N_27484,N_27487,N_27489,N_27491,N_27492,N_27493,N_27494,N_27496,N_27498,N_27499,N_27500,N_27501,N_27502,N_27505,N_27506,N_27509,N_27510,N_27512,N_27513,N_27515,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27524,N_27525,N_27526,N_27527,N_27528,N_27530,N_27531,N_27532,N_27533,N_27535,N_27536,N_27539,N_27541,N_27542,N_27545,N_27546,N_27548,N_27549,N_27550,N_27551,N_27554,N_27555,N_27556,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27569,N_27570,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27580,N_27581,N_27584,N_27585,N_27586,N_27587,N_27588,N_27592,N_27593,N_27594,N_27595,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27605,N_27607,N_27609,N_27611,N_27612,N_27613,N_27614,N_27615,N_27617,N_27618,N_27619,N_27621,N_27622,N_27624,N_27625,N_27626,N_27627,N_27630,N_27632,N_27634,N_27635,N_27637,N_27638,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27650,N_27651,N_27652,N_27654,N_27655,N_27656,N_27658,N_27659,N_27661,N_27662,N_27663,N_27665,N_27667,N_27668,N_27670,N_27671,N_27672,N_27674,N_27675,N_27676,N_27679,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27696,N_27697,N_27698,N_27699,N_27700,N_27702,N_27703,N_27705,N_27706,N_27707,N_27708,N_27710,N_27713,N_27716,N_27717,N_27718,N_27719,N_27722,N_27723,N_27725,N_27726,N_27727,N_27729,N_27730,N_27731,N_27733,N_27735,N_27737,N_27739,N_27741,N_27743,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27766,N_27767,N_27768,N_27769,N_27770,N_27772,N_27773,N_27775,N_27776,N_27777,N_27778,N_27779,N_27781,N_27782,N_27784,N_27785,N_27786,N_27788,N_27789,N_27791,N_27792,N_27793,N_27794,N_27795,N_27797,N_27799,N_27801,N_27803,N_27804,N_27805,N_27806,N_27807,N_27813,N_27814,N_27815,N_27817,N_27819,N_27820,N_27821,N_27822,N_27823,N_27825,N_27826,N_27827,N_27829,N_27830,N_27831,N_27833,N_27834,N_27836,N_27837,N_27838,N_27839,N_27842,N_27843,N_27844,N_27845,N_27846,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27857,N_27861,N_27863,N_27864,N_27865,N_27869,N_27870,N_27871,N_27874,N_27875,N_27876,N_27877,N_27878,N_27880,N_27883,N_27884,N_27886,N_27889,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27899,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27909,N_27911,N_27912,N_27913,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27925,N_27929,N_27930,N_27931,N_27932,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27942,N_27943,N_27944,N_27945,N_27947,N_27953,N_27954,N_27956,N_27957,N_27959,N_27960,N_27961,N_27962,N_27965,N_27966,N_27967,N_27969,N_27971,N_27972,N_27974,N_27975,N_27977,N_27981,N_27982,N_27984,N_27985,N_27986,N_27990,N_27991,N_27992,N_27993,N_27994,N_27996,N_27997,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28007,N_28008,N_28009,N_28010,N_28012,N_28015,N_28016,N_28018,N_28020,N_28021,N_28023,N_28024,N_28025,N_28026,N_28027,N_28029,N_28030,N_28031,N_28032,N_28035,N_28037,N_28039,N_28040,N_28042,N_28043,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28054,N_28055,N_28058,N_28059,N_28062,N_28063,N_28064,N_28066,N_28067,N_28069,N_28070,N_28072,N_28073,N_28075,N_28076,N_28077,N_28080,N_28081,N_28082,N_28085,N_28086,N_28087,N_28089,N_28090,N_28091,N_28092,N_28094,N_28096,N_28097,N_28098,N_28101,N_28102,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28143,N_28144,N_28145,N_28146,N_28148,N_28149,N_28152,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28174,N_28175,N_28176,N_28177,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28193,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28227,N_28229,N_28231,N_28233,N_28234,N_28235,N_28238,N_28242,N_28243,N_28245,N_28248,N_28250,N_28251,N_28252,N_28253,N_28255,N_28256,N_28258,N_28259,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28269,N_28270,N_28271,N_28273,N_28274,N_28275,N_28278,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28287,N_28288,N_28289,N_28290,N_28292,N_28293,N_28294,N_28296,N_28297,N_28300,N_28301,N_28302,N_28303,N_28305,N_28306,N_28312,N_28313,N_28315,N_28316,N_28317,N_28320,N_28321,N_28322,N_28324,N_28325,N_28326,N_28328,N_28329,N_28330,N_28331,N_28333,N_28334,N_28335,N_28336,N_28337,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28347,N_28348,N_28350,N_28351,N_28352,N_28355,N_28357,N_28359,N_28360,N_28361,N_28362,N_28363,N_28365,N_28366,N_28367,N_28369,N_28371,N_28374,N_28376,N_28378,N_28379,N_28380,N_28381,N_28383,N_28385,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28395,N_28396,N_28398,N_28399,N_28400,N_28401,N_28404,N_28407,N_28408,N_28410,N_28411,N_28413,N_28416,N_28420,N_28423,N_28424,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28433,N_28434,N_28436,N_28437,N_28439,N_28440,N_28441,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28461,N_28462,N_28466,N_28469,N_28470,N_28471,N_28473,N_28477,N_28478,N_28479,N_28480,N_28482,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28493,N_28494,N_28495,N_28497,N_28498,N_28499,N_28500,N_28501,N_28503,N_28504,N_28508,N_28509,N_28510,N_28512,N_28513,N_28515,N_28516,N_28517,N_28518,N_28519,N_28522,N_28523,N_28525,N_28526,N_28527,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28538,N_28539,N_28543,N_28545,N_28546,N_28548,N_28549,N_28551,N_28553,N_28554,N_28555,N_28556,N_28557,N_28559,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28581,N_28583,N_28585,N_28586,N_28587,N_28588,N_28589,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28599,N_28600,N_28601,N_28604,N_28605,N_28607,N_28608,N_28609,N_28610,N_28612,N_28614,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28627,N_28629,N_28630,N_28631,N_28632,N_28634,N_28635,N_28637,N_28638,N_28639,N_28641,N_28642,N_28643,N_28644,N_28645,N_28647,N_28648,N_28652,N_28653,N_28654,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28689,N_28690,N_28691,N_28695,N_28696,N_28697,N_28698,N_28699,N_28701,N_28702,N_28703,N_28704,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28722,N_28723,N_28725,N_28726,N_28727,N_28728,N_28730,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28749,N_28750,N_28752,N_28753,N_28754,N_28755,N_28756,N_28758,N_28761,N_28762,N_28763,N_28764,N_28765,N_28767,N_28772,N_28773,N_28774,N_28776,N_28777,N_28778,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28802,N_28803,N_28804,N_28806,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28817,N_28819,N_28820,N_28821,N_28822,N_28823,N_28825,N_28826,N_28827,N_28831,N_28832,N_28834,N_28835,N_28837,N_28838,N_28839,N_28840,N_28841,N_28844,N_28846,N_28847,N_28850,N_28851,N_28852,N_28853,N_28855,N_28857,N_28858,N_28859,N_28860,N_28861,N_28863,N_28864,N_28865,N_28866,N_28867,N_28869,N_28870,N_28872,N_28873,N_28874,N_28875,N_28876,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28887,N_28888,N_28891,N_28892,N_28893,N_28895,N_28898,N_28900,N_28901,N_28902,N_28904,N_28906,N_28908,N_28909,N_28911,N_28913,N_28914,N_28916,N_28917,N_28918,N_28921,N_28923,N_28924,N_28925,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28937,N_28938,N_28939,N_28942,N_28943,N_28944,N_28946,N_28947,N_28950,N_28951,N_28953,N_28955,N_28956,N_28957,N_28960,N_28962,N_28964,N_28966,N_28967,N_28968,N_28969,N_28971,N_28973,N_28975,N_28976,N_28977,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28986,N_28987,N_28988,N_28993,N_28994,N_28995,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29010,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29028,N_29029,N_29030,N_29031,N_29032,N_29034,N_29036,N_29037,N_29038,N_29039,N_29040,N_29043,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29052,N_29053,N_29054,N_29058,N_29059,N_29061,N_29062,N_29063,N_29065,N_29067,N_29068,N_29069,N_29070,N_29071,N_29074,N_29076,N_29077,N_29078,N_29081,N_29082,N_29085,N_29087,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29101,N_29102,N_29106,N_29107,N_29109,N_29110,N_29111,N_29112,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29145,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29172,N_29175,N_29176,N_29177,N_29178,N_29180,N_29182,N_29183,N_29184,N_29185,N_29188,N_29189,N_29191,N_29193,N_29194,N_29195,N_29196,N_29197,N_29199,N_29200,N_29201,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29213,N_29214,N_29216,N_29217,N_29218,N_29219,N_29221,N_29223,N_29224,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29234,N_29235,N_29236,N_29238,N_29239,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29249,N_29251,N_29252,N_29254,N_29255,N_29256,N_29259,N_29260,N_29261,N_29264,N_29266,N_29267,N_29268,N_29269,N_29271,N_29272,N_29273,N_29275,N_29277,N_29278,N_29279,N_29280,N_29282,N_29283,N_29284,N_29285,N_29293,N_29294,N_29295,N_29296,N_29298,N_29300,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29314,N_29315,N_29316,N_29317,N_29318,N_29320,N_29321,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29331,N_29332,N_29333,N_29334,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29356,N_29357,N_29358,N_29360,N_29361,N_29363,N_29365,N_29366,N_29368,N_29369,N_29370,N_29371,N_29373,N_29374,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29383,N_29386,N_29388,N_29389,N_29391,N_29393,N_29394,N_29397,N_29398,N_29401,N_29402,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29414,N_29415,N_29416,N_29418,N_29419,N_29420,N_29421,N_29423,N_29424,N_29426,N_29428,N_29430,N_29432,N_29433,N_29436,N_29437,N_29438,N_29439,N_29440,N_29442,N_29443,N_29444,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29456,N_29457,N_29458,N_29460,N_29462,N_29463,N_29464,N_29469,N_29472,N_29473,N_29474,N_29475,N_29477,N_29478,N_29479,N_29480,N_29481,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29491,N_29492,N_29493,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29507,N_29508,N_29509,N_29510,N_29512,N_29513,N_29515,N_29517,N_29518,N_29519,N_29520,N_29523,N_29524,N_29525,N_29528,N_29529,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29541,N_29542,N_29545,N_29548,N_29550,N_29553,N_29554,N_29556,N_29557,N_29558,N_29559,N_29560,N_29562,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29582,N_29585,N_29588,N_29589,N_29590,N_29592,N_29594,N_29595,N_29596,N_29598,N_29599,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29609,N_29610,N_29611,N_29613,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29623,N_29624,N_29626,N_29629,N_29630,N_29631,N_29632,N_29635,N_29636,N_29637,N_29639,N_29640,N_29642,N_29644,N_29645,N_29646,N_29647,N_29649,N_29650,N_29652,N_29653,N_29655,N_29657,N_29658,N_29663,N_29664,N_29666,N_29667,N_29668,N_29670,N_29672,N_29675,N_29676,N_29677,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29688,N_29689,N_29690,N_29692,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29702,N_29703,N_29705,N_29707,N_29709,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29729,N_29730,N_29733,N_29735,N_29736,N_29737,N_29738,N_29739,N_29741,N_29743,N_29746,N_29747,N_29749,N_29750,N_29751,N_29752,N_29755,N_29757,N_29758,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29768,N_29769,N_29771,N_29773,N_29774,N_29775,N_29777,N_29778,N_29780,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29790,N_29791,N_29792,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29801,N_29802,N_29804,N_29807,N_29808,N_29809,N_29810,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29822,N_29824,N_29825,N_29826,N_29827,N_29829,N_29830,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29846,N_29847,N_29848,N_29851,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29864,N_29865,N_29866,N_29867,N_29869,N_29870,N_29871,N_29872,N_29873,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29889,N_29890,N_29891,N_29893,N_29894,N_29895,N_29897,N_29898,N_29899,N_29901,N_29904,N_29905,N_29906,N_29908,N_29909,N_29910,N_29913,N_29915,N_29916,N_29917,N_29918,N_29919,N_29921,N_29922,N_29923,N_29924,N_29925,N_29928,N_29929,N_29931,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29942,N_29943,N_29947,N_29949,N_29950,N_29955,N_29956,N_29957,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29967,N_29968,N_29969,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29984,N_29985,N_29986,N_29987,N_29989,N_29990,N_29991,N_29993,N_29994,N_29996,N_29997,N_29999;
and U0 (N_0,In_733,In_2672);
or U1 (N_1,In_1731,In_266);
or U2 (N_2,In_1038,In_930);
nand U3 (N_3,In_1196,In_1715);
nor U4 (N_4,In_2686,In_2377);
or U5 (N_5,In_256,In_2150);
nor U6 (N_6,In_106,In_2165);
xor U7 (N_7,In_2215,In_2390);
nor U8 (N_8,In_18,In_2486);
nor U9 (N_9,In_767,In_917);
or U10 (N_10,In_471,In_1635);
and U11 (N_11,In_200,In_2476);
nor U12 (N_12,In_1951,In_911);
or U13 (N_13,In_2540,In_275);
and U14 (N_14,In_2644,In_1616);
and U15 (N_15,In_2428,In_257);
nand U16 (N_16,In_722,In_2528);
nand U17 (N_17,In_720,In_2668);
nor U18 (N_18,In_821,In_2512);
or U19 (N_19,In_1321,In_2255);
nand U20 (N_20,In_2507,In_2986);
and U21 (N_21,In_2752,In_2750);
nor U22 (N_22,In_595,In_2396);
nor U23 (N_23,In_186,In_52);
nor U24 (N_24,In_287,In_2744);
nor U25 (N_25,In_831,In_1984);
or U26 (N_26,In_1856,In_2402);
or U27 (N_27,In_2300,In_1424);
nor U28 (N_28,In_1307,In_1587);
or U29 (N_29,In_993,In_482);
nor U30 (N_30,In_2546,In_1278);
nor U31 (N_31,In_128,In_1568);
and U32 (N_32,In_1477,In_2369);
xor U33 (N_33,In_449,In_561);
nand U34 (N_34,In_649,In_127);
nand U35 (N_35,In_2458,In_2501);
or U36 (N_36,In_2778,In_456);
or U37 (N_37,In_1335,In_2849);
nor U38 (N_38,In_2241,In_1252);
or U39 (N_39,In_1834,In_1031);
or U40 (N_40,In_2731,In_1704);
and U41 (N_41,In_73,In_1573);
and U42 (N_42,In_268,In_1146);
nand U43 (N_43,In_1810,In_1860);
and U44 (N_44,In_2292,In_1632);
nor U45 (N_45,In_971,In_963);
nor U46 (N_46,In_204,In_1451);
xor U47 (N_47,In_1903,In_2224);
nand U48 (N_48,In_404,In_1183);
nand U49 (N_49,In_2921,In_1542);
nor U50 (N_50,In_13,In_1311);
and U51 (N_51,In_754,In_2077);
and U52 (N_52,In_786,In_236);
and U53 (N_53,In_1430,In_2149);
or U54 (N_54,In_1833,In_1354);
nor U55 (N_55,In_775,In_473);
nand U56 (N_56,In_2785,In_2814);
xnor U57 (N_57,In_1576,In_771);
nand U58 (N_58,In_1071,In_421);
or U59 (N_59,In_879,In_2757);
or U60 (N_60,In_909,In_2418);
or U61 (N_61,In_2941,In_864);
and U62 (N_62,In_1185,In_2978);
nand U63 (N_63,In_1929,In_1845);
nor U64 (N_64,In_490,In_1709);
or U65 (N_65,In_233,In_1683);
nand U66 (N_66,In_2804,In_2647);
or U67 (N_67,In_1182,In_713);
and U68 (N_68,In_1299,In_1527);
or U69 (N_69,In_1760,In_891);
or U70 (N_70,In_1157,In_232);
nand U71 (N_71,In_847,In_547);
nor U72 (N_72,In_829,In_730);
nand U73 (N_73,In_2837,In_884);
or U74 (N_74,In_1217,In_272);
or U75 (N_75,In_1773,In_472);
nand U76 (N_76,In_701,In_1001);
nand U77 (N_77,In_143,In_1496);
nand U78 (N_78,In_956,In_1256);
nor U79 (N_79,In_1392,In_551);
and U80 (N_80,In_2701,In_860);
nand U81 (N_81,In_298,In_2777);
and U82 (N_82,In_624,In_438);
and U83 (N_83,In_2335,In_1624);
and U84 (N_84,In_1412,In_2243);
or U85 (N_85,In_640,In_528);
nor U86 (N_86,In_1610,In_2200);
xor U87 (N_87,In_2977,In_2805);
nand U88 (N_88,In_850,In_283);
nand U89 (N_89,In_1026,In_2656);
and U90 (N_90,In_2346,In_1420);
or U91 (N_91,In_672,In_586);
or U92 (N_92,In_1047,In_114);
nand U93 (N_93,In_1264,In_182);
nor U94 (N_94,In_832,In_2114);
and U95 (N_95,In_2591,In_2951);
nor U96 (N_96,In_1438,In_2044);
or U97 (N_97,In_1829,In_176);
or U98 (N_98,In_1331,In_80);
or U99 (N_99,In_74,In_407);
nor U100 (N_100,In_2852,In_2787);
nand U101 (N_101,In_147,In_2684);
nor U102 (N_102,In_1896,In_565);
and U103 (N_103,In_2034,In_2705);
or U104 (N_104,In_1965,In_608);
or U105 (N_105,In_377,In_1291);
nor U106 (N_106,In_1763,In_2623);
xnor U107 (N_107,In_218,In_973);
xor U108 (N_108,In_2152,In_2297);
nand U109 (N_109,In_12,In_1663);
nand U110 (N_110,In_1328,In_1265);
nand U111 (N_111,In_727,In_48);
or U112 (N_112,In_1914,In_1705);
nand U113 (N_113,In_1586,In_678);
nand U114 (N_114,In_222,In_2566);
nand U115 (N_115,In_2257,In_1670);
nand U116 (N_116,In_1770,In_873);
and U117 (N_117,In_1140,In_2555);
nand U118 (N_118,In_2557,In_968);
or U119 (N_119,In_88,In_2758);
xnor U120 (N_120,In_862,In_538);
and U121 (N_121,In_2498,In_925);
nor U122 (N_122,In_889,In_1868);
nor U123 (N_123,In_2234,In_2328);
xor U124 (N_124,In_2212,In_782);
nand U125 (N_125,In_295,In_1429);
and U126 (N_126,In_516,In_1764);
xnor U127 (N_127,In_805,In_1161);
and U128 (N_128,In_1651,In_2376);
nor U129 (N_129,In_1563,In_2289);
nand U130 (N_130,In_1675,In_1095);
or U131 (N_131,In_2925,In_812);
or U132 (N_132,In_2975,In_1631);
and U133 (N_133,In_1015,In_2531);
and U134 (N_134,In_2725,In_1032);
nand U135 (N_135,In_1711,In_2992);
nand U136 (N_136,In_282,In_2495);
nand U137 (N_137,In_49,In_2520);
or U138 (N_138,In_2018,In_247);
or U139 (N_139,In_1577,In_2692);
xor U140 (N_140,In_2740,In_1657);
and U141 (N_141,In_2385,In_1019);
and U142 (N_142,In_2947,In_1658);
nor U143 (N_143,In_2043,In_760);
or U144 (N_144,In_1796,In_2188);
and U145 (N_145,In_2201,In_2055);
or U146 (N_146,In_1490,In_843);
nand U147 (N_147,In_1235,In_2131);
and U148 (N_148,In_814,In_818);
nor U149 (N_149,In_1850,In_591);
nor U150 (N_150,In_2301,In_2567);
or U151 (N_151,In_30,In_2197);
or U152 (N_152,In_2859,In_1730);
or U153 (N_153,In_2634,In_387);
or U154 (N_154,In_758,In_2929);
nand U155 (N_155,In_625,In_888);
nor U156 (N_156,In_1339,In_2556);
and U157 (N_157,In_683,In_1021);
nor U158 (N_158,In_2678,In_2467);
nand U159 (N_159,In_681,In_2373);
nand U160 (N_160,In_274,In_2009);
or U161 (N_161,In_1555,In_1945);
nand U162 (N_162,In_1344,In_2545);
nor U163 (N_163,In_2534,In_1963);
xor U164 (N_164,In_2181,In_855);
and U165 (N_165,In_1002,In_2371);
or U166 (N_166,In_2138,In_1158);
nor U167 (N_167,In_2227,In_880);
and U168 (N_168,In_1905,In_1245);
or U169 (N_169,In_2090,In_2135);
nor U170 (N_170,In_588,In_944);
or U171 (N_171,In_2040,In_63);
xor U172 (N_172,In_2105,In_597);
nor U173 (N_173,In_2329,In_2683);
and U174 (N_174,In_2931,In_334);
nand U175 (N_175,In_1213,In_43);
or U176 (N_176,In_2326,In_265);
and U177 (N_177,In_2544,In_2961);
nand U178 (N_178,In_2351,In_1150);
nor U179 (N_179,In_1584,In_281);
and U180 (N_180,In_599,In_2356);
and U181 (N_181,In_2422,In_2988);
nor U182 (N_182,In_221,In_2437);
nand U183 (N_183,In_484,In_2155);
nor U184 (N_184,In_60,In_1493);
nand U185 (N_185,In_19,In_2824);
nor U186 (N_186,In_2287,In_1838);
or U187 (N_187,In_81,In_2115);
or U188 (N_188,In_2828,In_1063);
or U189 (N_189,In_1706,In_373);
nor U190 (N_190,In_1911,In_89);
nor U191 (N_191,In_662,In_2509);
or U192 (N_192,In_842,In_1491);
and U193 (N_193,In_2271,In_153);
and U194 (N_194,In_2160,In_2596);
and U195 (N_195,In_1014,In_724);
and U196 (N_196,In_1585,In_1590);
or U197 (N_197,In_305,In_2399);
nor U198 (N_198,In_1457,In_187);
nor U199 (N_199,In_1877,In_2801);
or U200 (N_200,In_406,In_2885);
or U201 (N_201,In_2882,In_803);
nand U202 (N_202,In_2915,In_2734);
nand U203 (N_203,In_2378,In_2167);
nor U204 (N_204,In_393,In_2020);
nor U205 (N_205,In_1289,In_2096);
xnor U206 (N_206,In_2216,In_653);
or U207 (N_207,In_255,In_251);
nor U208 (N_208,In_2876,In_2345);
nor U209 (N_209,In_1687,In_11);
nor U210 (N_210,In_2997,In_1572);
or U211 (N_211,In_1201,In_2424);
or U212 (N_212,In_2614,In_2480);
or U213 (N_213,In_2677,In_2796);
and U214 (N_214,In_780,In_1093);
nand U215 (N_215,In_1895,In_1506);
nand U216 (N_216,In_2370,In_427);
xor U217 (N_217,In_2946,In_1839);
or U218 (N_218,In_1094,In_619);
nand U219 (N_219,In_1756,In_1788);
nand U220 (N_220,In_1292,In_962);
and U221 (N_221,In_2884,In_871);
and U222 (N_222,In_371,In_1917);
xnor U223 (N_223,In_2184,In_1154);
and U224 (N_224,In_1613,In_1888);
and U225 (N_225,In_523,In_2802);
or U226 (N_226,In_712,In_8);
and U227 (N_227,In_964,In_2963);
and U228 (N_228,In_2795,In_2967);
or U229 (N_229,In_1503,In_788);
nor U230 (N_230,In_1907,In_1);
or U231 (N_231,In_1197,In_1598);
and U232 (N_232,In_1776,In_447);
and U233 (N_233,In_1743,In_337);
and U234 (N_234,In_2117,In_1969);
nor U235 (N_235,In_249,In_2879);
nor U236 (N_236,In_1611,In_1575);
nand U237 (N_237,In_195,In_2918);
or U238 (N_238,In_576,In_857);
and U239 (N_239,In_1456,In_2854);
and U240 (N_240,In_1302,In_2039);
nand U241 (N_241,In_254,In_1761);
and U242 (N_242,In_2790,In_458);
nor U243 (N_243,In_1667,In_940);
nand U244 (N_244,In_777,In_2367);
and U245 (N_245,In_2898,In_673);
and U246 (N_246,In_2139,In_297);
or U247 (N_247,In_1008,In_2912);
nand U248 (N_248,In_526,In_1044);
nor U249 (N_249,In_1700,In_3);
nor U250 (N_250,In_69,In_2283);
or U251 (N_251,In_119,In_2343);
nor U252 (N_252,In_2330,In_1507);
nand U253 (N_253,In_1600,In_1099);
nand U254 (N_254,In_1558,In_1027);
and U255 (N_255,In_2006,In_2553);
nand U256 (N_256,In_2010,In_2170);
or U257 (N_257,In_1097,In_2514);
xor U258 (N_258,In_1475,In_1733);
nand U259 (N_259,In_2219,In_248);
xnor U260 (N_260,In_316,In_2927);
nor U261 (N_261,In_480,In_1740);
or U262 (N_262,In_1474,In_212);
or U263 (N_263,In_359,In_1554);
and U264 (N_264,In_338,In_1592);
and U265 (N_265,In_1938,In_2938);
nor U266 (N_266,In_2336,In_2896);
and U267 (N_267,In_2353,In_2078);
nand U268 (N_268,In_1380,In_379);
nand U269 (N_269,In_910,In_1842);
nand U270 (N_270,In_2934,In_1612);
and U271 (N_271,In_2982,In_188);
or U272 (N_272,In_2249,In_949);
nor U273 (N_273,In_2535,In_1665);
nor U274 (N_274,In_1222,In_2471);
nor U275 (N_275,In_429,In_2084);
nor U276 (N_276,In_1083,In_35);
or U277 (N_277,In_2771,In_2542);
and U278 (N_278,In_1853,In_726);
and U279 (N_279,In_6,In_2788);
and U280 (N_280,In_1241,In_1151);
and U281 (N_281,In_2917,In_654);
xnor U282 (N_282,In_318,In_1793);
or U283 (N_283,In_96,In_2881);
and U284 (N_284,In_762,In_1797);
or U285 (N_285,In_1696,In_1594);
nor U286 (N_286,In_2107,In_2615);
nor U287 (N_287,In_870,In_1803);
and U288 (N_288,In_1249,In_2488);
or U289 (N_289,In_518,In_415);
nand U290 (N_290,In_428,In_2570);
and U291 (N_291,In_1862,In_1061);
and U292 (N_292,In_2667,In_702);
nor U293 (N_293,In_2209,In_2945);
or U294 (N_294,In_423,In_23);
and U295 (N_295,In_1142,In_2087);
or U296 (N_296,In_736,In_1463);
and U297 (N_297,In_900,In_1359);
or U298 (N_298,In_2291,In_1734);
or U299 (N_299,In_1989,In_2483);
or U300 (N_300,In_1618,In_2459);
xor U301 (N_301,In_2416,In_2940);
nand U302 (N_302,In_2064,In_2060);
nor U303 (N_303,In_1040,In_354);
nor U304 (N_304,In_149,In_848);
nor U305 (N_305,In_1341,In_320);
and U306 (N_306,In_2826,In_1255);
nor U307 (N_307,In_2479,In_1268);
or U308 (N_308,In_2425,In_1408);
nor U309 (N_309,In_2832,In_1821);
or U310 (N_310,In_1997,In_977);
or U311 (N_311,In_2245,In_723);
or U312 (N_312,In_2720,In_2156);
and U313 (N_313,In_446,In_2900);
xor U314 (N_314,In_1648,In_979);
and U315 (N_315,In_238,In_987);
or U316 (N_316,In_704,In_93);
nor U317 (N_317,In_477,In_2264);
nand U318 (N_318,In_659,In_955);
and U319 (N_319,In_1208,In_2054);
nand U320 (N_320,In_1275,In_2955);
nor U321 (N_321,In_922,In_975);
and U322 (N_322,In_2624,In_2104);
nand U323 (N_323,In_2993,In_1781);
nand U324 (N_324,In_1262,In_2022);
xor U325 (N_325,In_972,In_300);
and U326 (N_326,In_2529,In_1692);
nor U327 (N_327,In_2908,In_953);
nor U328 (N_328,In_1221,In_2061);
nor U329 (N_329,In_2724,In_36);
nand U330 (N_330,In_905,In_196);
nor U331 (N_331,In_445,In_2387);
xnor U332 (N_332,In_2751,In_312);
nor U333 (N_333,In_54,In_1155);
nor U334 (N_334,In_1902,In_2630);
xor U335 (N_335,In_542,In_2470);
nor U336 (N_336,In_2485,In_1237);
nor U337 (N_337,In_1187,In_2350);
or U338 (N_338,In_982,In_2123);
nor U339 (N_339,In_1464,In_1104);
and U340 (N_340,In_345,In_172);
nor U341 (N_341,In_1534,In_580);
or U342 (N_342,In_622,In_705);
and U343 (N_343,In_809,In_742);
and U344 (N_344,In_711,In_693);
or U345 (N_345,In_1317,In_2284);
nand U346 (N_346,In_1045,In_1415);
nor U347 (N_347,In_2738,In_457);
or U348 (N_348,In_1090,In_985);
or U349 (N_349,In_2404,In_2338);
nor U350 (N_350,In_258,In_264);
xor U351 (N_351,In_2062,In_2780);
nand U352 (N_352,In_839,In_496);
nand U353 (N_353,In_462,In_1520);
nor U354 (N_354,In_1224,In_79);
and U355 (N_355,In_2013,In_1831);
nor U356 (N_356,In_1133,In_546);
nand U357 (N_357,In_2238,In_2847);
or U358 (N_358,In_1702,In_1349);
nand U359 (N_359,In_2456,In_2874);
nand U360 (N_360,In_1041,In_273);
nand U361 (N_361,In_2666,In_1096);
nand U362 (N_362,In_2413,In_331);
and U363 (N_363,In_1580,In_409);
nor U364 (N_364,In_1024,In_1596);
or U365 (N_365,In_2503,In_2932);
and U366 (N_366,In_2059,In_868);
nand U367 (N_367,In_2990,In_867);
xor U368 (N_368,In_921,In_1921);
or U369 (N_369,In_118,In_1976);
or U370 (N_370,In_1165,In_1004);
nand U371 (N_371,In_2268,In_1108);
nor U372 (N_372,In_2579,In_2916);
and U373 (N_373,In_1633,In_1425);
and U374 (N_374,In_1285,In_443);
and U375 (N_375,In_2178,In_303);
xnor U376 (N_376,In_1772,In_159);
or U377 (N_377,In_845,In_638);
xor U378 (N_378,In_460,In_686);
nand U379 (N_379,In_2072,In_1070);
nor U380 (N_380,In_1413,In_519);
xor U381 (N_381,In_2251,In_2333);
and U382 (N_382,In_2920,In_2973);
nor U383 (N_383,In_833,In_2682);
nand U384 (N_384,In_2058,In_1578);
nor U385 (N_385,In_2162,In_629);
and U386 (N_386,In_947,In_637);
and U387 (N_387,In_941,In_17);
and U388 (N_388,In_437,In_557);
or U389 (N_389,In_413,In_1199);
or U390 (N_390,In_541,In_28);
or U391 (N_391,In_2194,In_1202);
nand U392 (N_392,In_1295,In_2440);
nand U393 (N_393,In_1020,In_1878);
nor U394 (N_394,In_2708,In_2173);
or U395 (N_395,In_1214,In_1149);
nor U396 (N_396,In_2491,In_2718);
xor U397 (N_397,In_2368,In_2549);
or U398 (N_398,In_1362,In_567);
nand U399 (N_399,In_202,In_1684);
and U400 (N_400,In_358,In_826);
nor U401 (N_401,In_1977,In_1012);
nand U402 (N_402,In_494,In_2619);
and U403 (N_403,In_1057,In_1721);
xnor U404 (N_404,In_1866,In_1009);
nand U405 (N_405,In_1712,In_1739);
and U406 (N_406,In_590,In_641);
nor U407 (N_407,In_698,In_615);
nand U408 (N_408,In_1274,In_548);
and U409 (N_409,In_1968,In_2384);
or U410 (N_410,In_1472,In_592);
and U411 (N_411,In_1680,In_2609);
and U412 (N_412,In_746,In_1771);
or U413 (N_413,In_1322,In_1276);
nor U414 (N_414,In_2517,In_2959);
or U415 (N_415,In_2122,In_1982);
nand U416 (N_416,In_1912,In_863);
nand U417 (N_417,In_898,In_852);
nand U418 (N_418,In_790,In_2462);
and U419 (N_419,In_569,In_721);
nor U420 (N_420,In_1053,In_2056);
and U421 (N_421,In_244,In_1869);
xor U422 (N_422,In_205,In_2019);
or U423 (N_423,In_1942,In_2585);
and U424 (N_424,In_1243,In_2391);
xor U425 (N_425,In_568,In_2575);
nand U426 (N_426,In_1735,In_2365);
and U427 (N_427,In_1082,In_1267);
nand U428 (N_428,In_278,In_1055);
or U429 (N_429,In_1210,In_1356);
nand U430 (N_430,In_162,In_2032);
nor U431 (N_431,In_927,In_2948);
nor U432 (N_432,In_1498,In_1792);
nand U433 (N_433,In_448,In_574);
nor U434 (N_434,In_2833,In_1310);
and U435 (N_435,In_1173,In_601);
and U436 (N_436,In_2168,In_2163);
or U437 (N_437,In_1003,In_2258);
xor U438 (N_438,In_1767,In_2957);
or U439 (N_439,In_908,In_866);
and U440 (N_440,In_2547,In_743);
or U441 (N_441,In_2956,In_1660);
or U442 (N_442,In_2712,In_161);
nor U443 (N_443,In_418,In_1930);
nor U444 (N_444,In_1674,In_2527);
nand U445 (N_445,In_2492,In_1323);
and U446 (N_446,In_1784,In_1402);
and U447 (N_447,In_2379,In_225);
nor U448 (N_448,In_509,In_2204);
and U449 (N_449,In_1646,In_124);
and U450 (N_450,In_1634,In_1148);
and U451 (N_451,In_112,In_1067);
or U452 (N_452,In_224,In_1435);
nand U453 (N_453,In_2976,In_1107);
and U454 (N_454,In_651,In_1483);
or U455 (N_455,In_416,In_806);
and U456 (N_456,In_1282,In_1549);
and U457 (N_457,In_1143,In_1901);
nand U458 (N_458,In_2341,In_131);
nand U459 (N_459,In_1987,In_2095);
nand U460 (N_460,In_2980,In_306);
nor U461 (N_461,In_1179,In_328);
nand U462 (N_462,In_1085,In_2202);
nand U463 (N_463,In_2302,In_308);
or U464 (N_464,In_134,In_639);
nand U465 (N_465,In_2521,In_532);
or U466 (N_466,In_2831,In_1485);
nand U467 (N_467,In_2484,In_677);
and U468 (N_468,In_2433,In_825);
nor U469 (N_469,In_1076,In_483);
nor U470 (N_470,In_148,In_960);
or U471 (N_471,In_1433,In_375);
or U472 (N_472,In_699,In_2049);
nor U473 (N_473,In_342,In_2588);
or U474 (N_474,In_1897,In_1172);
nor U475 (N_475,In_2574,In_2237);
and U476 (N_476,In_133,In_2690);
nor U477 (N_477,In_1664,In_1326);
or U478 (N_478,In_797,In_419);
and U479 (N_479,In_2183,In_2092);
and U480 (N_480,In_353,In_29);
and U481 (N_481,In_2664,In_1092);
or U482 (N_482,In_998,In_1159);
nand U483 (N_483,In_1944,In_327);
nand U484 (N_484,In_410,In_2449);
nand U485 (N_485,In_1927,In_2893);
nand U486 (N_486,In_658,In_1988);
or U487 (N_487,In_1537,In_2776);
nand U488 (N_488,In_151,In_1419);
nor U489 (N_489,In_2323,In_2821);
and U490 (N_490,In_111,In_902);
or U491 (N_491,In_543,In_14);
nand U492 (N_492,In_1832,In_2560);
or U493 (N_493,In_103,In_364);
nor U494 (N_494,In_2016,In_2126);
and U495 (N_495,In_2628,In_1488);
nand U496 (N_496,In_1231,In_2595);
nor U497 (N_497,In_136,In_564);
nor U498 (N_498,In_2745,In_2887);
nor U499 (N_499,In_2841,In_1511);
nor U500 (N_500,In_1673,In_219);
and U501 (N_501,In_1778,In_2767);
xor U502 (N_502,In_1049,In_1909);
and U503 (N_503,In_2648,In_84);
or U504 (N_504,In_578,In_1974);
nor U505 (N_505,In_2172,In_2372);
nand U506 (N_506,In_1867,In_2144);
nor U507 (N_507,In_1703,In_664);
or U508 (N_508,In_367,In_1487);
or U509 (N_509,In_123,In_1765);
or U510 (N_510,In_1314,In_1894);
or U511 (N_511,In_1417,In_2774);
nor U512 (N_512,In_1844,In_1309);
nand U513 (N_513,In_2157,In_2511);
nor U514 (N_514,In_58,In_2746);
or U515 (N_515,In_2743,In_381);
xnor U516 (N_516,In_1259,In_1959);
xor U517 (N_517,In_2696,In_1431);
nor U518 (N_518,In_648,In_1943);
and U519 (N_519,In_2454,In_2923);
nor U520 (N_520,In_675,In_2526);
nand U521 (N_521,In_2532,In_2226);
xor U522 (N_522,In_1186,In_798);
xnor U523 (N_523,In_2050,In_2082);
nand U524 (N_524,In_1389,In_53);
nand U525 (N_525,In_1641,In_1736);
nand U526 (N_526,In_2282,In_1180);
nand U527 (N_527,In_1716,In_2400);
nor U528 (N_528,In_2792,In_2401);
nand U529 (N_529,In_102,In_226);
and U530 (N_530,In_1919,In_770);
nand U531 (N_531,In_2186,In_1913);
nand U532 (N_532,In_178,In_374);
nand U533 (N_533,In_2063,In_104);
nor U534 (N_534,In_1134,In_2862);
nand U535 (N_535,In_1661,In_294);
nand U536 (N_536,In_135,In_1975);
and U537 (N_537,In_2913,In_2116);
or U538 (N_538,In_2048,In_109);
and U539 (N_539,In_2334,In_2844);
or U540 (N_540,In_1553,In_2136);
or U541 (N_541,In_1622,In_2419);
or U542 (N_542,In_2823,In_1995);
nand U543 (N_543,In_464,In_2551);
nor U544 (N_544,In_1524,In_976);
or U545 (N_545,In_1290,In_370);
nand U546 (N_546,In_2374,In_2671);
or U547 (N_547,In_1080,In_799);
xor U548 (N_548,In_34,In_1468);
nand U549 (N_549,In_2706,In_1497);
xnor U550 (N_550,In_555,In_525);
nand U551 (N_551,In_1513,In_1540);
and U552 (N_552,In_1297,In_0);
and U553 (N_553,In_2093,In_1353);
nor U554 (N_554,In_372,In_1294);
nand U555 (N_555,In_878,In_2606);
and U556 (N_556,In_2891,In_970);
or U557 (N_557,In_2290,In_2661);
and U558 (N_558,In_2794,In_1672);
nor U559 (N_559,In_2576,In_2129);
and U560 (N_560,In_1998,In_1247);
or U561 (N_561,In_2618,In_534);
and U562 (N_562,In_2298,In_1861);
nand U563 (N_563,In_2930,In_378);
or U564 (N_564,In_2177,In_1205);
nor U565 (N_565,In_807,In_2926);
nand U566 (N_566,In_185,In_2244);
and U567 (N_567,In_1113,In_1355);
nand U568 (N_568,In_2352,In_150);
nor U569 (N_569,In_173,In_1873);
xnor U570 (N_570,In_887,In_269);
or U571 (N_571,In_2733,In_984);
nand U572 (N_572,In_2278,In_465);
and U573 (N_573,In_1599,In_861);
nor U574 (N_574,In_734,In_958);
or U575 (N_575,In_434,In_2229);
or U576 (N_576,In_671,In_1985);
or U577 (N_577,In_1029,In_2789);
xnor U578 (N_578,In_2295,In_2246);
or U579 (N_579,In_2147,In_967);
and U580 (N_580,In_243,In_572);
and U581 (N_581,In_392,In_1368);
xor U582 (N_582,In_1226,In_787);
or U583 (N_583,In_2808,In_90);
and U584 (N_584,In_718,In_1961);
and U585 (N_585,In_2046,In_1601);
or U586 (N_586,In_1644,In_1242);
xnor U587 (N_587,In_2119,In_912);
or U588 (N_588,In_2863,In_2616);
and U589 (N_589,In_2303,In_1177);
and U590 (N_590,In_459,In_2361);
nor U591 (N_591,In_933,In_1386);
nand U592 (N_592,In_1482,In_2636);
or U593 (N_593,In_1167,In_1372);
or U594 (N_594,In_796,In_1439);
nor U595 (N_595,In_1659,In_774);
nand U596 (N_596,In_630,In_503);
nand U597 (N_597,In_319,In_1970);
nor U598 (N_598,In_486,In_660);
or U599 (N_599,In_420,In_1526);
xor U600 (N_600,In_1738,In_1865);
or U601 (N_601,In_468,In_51);
nor U602 (N_602,In_750,In_737);
nand U603 (N_603,In_1212,In_2439);
and U604 (N_604,In_179,In_22);
nor U605 (N_605,In_2504,In_1544);
or U606 (N_606,In_1629,In_2652);
or U607 (N_607,In_405,In_1169);
or U608 (N_608,In_1522,In_800);
and U609 (N_609,In_655,In_2109);
and U610 (N_610,In_2014,In_1752);
and U611 (N_611,In_2490,In_2002);
xor U612 (N_612,In_2094,In_1397);
and U613 (N_613,In_2053,In_802);
or U614 (N_614,In_1614,In_533);
nand U615 (N_615,In_2468,In_1744);
nor U616 (N_616,In_2897,In_1694);
nor U617 (N_617,In_2651,In_2137);
nor U618 (N_618,In_2603,In_1676);
xnor U619 (N_619,In_335,In_913);
nand U620 (N_620,In_2590,In_563);
nor U621 (N_621,In_1343,In_1514);
nand U622 (N_622,In_2220,In_2175);
nor U623 (N_623,In_1636,In_2421);
nand U624 (N_624,In_1218,In_680);
nor U625 (N_625,In_141,In_1394);
and U626 (N_626,In_2159,In_2877);
and U627 (N_627,In_2765,In_2427);
and U628 (N_628,In_2154,In_1418);
nand U629 (N_629,In_293,In_1348);
nand U630 (N_630,In_1375,In_980);
or U631 (N_631,In_152,In_1382);
xnor U632 (N_632,In_764,In_94);
nor U633 (N_633,In_98,In_1164);
or U634 (N_634,In_1649,In_2592);
nand U635 (N_635,In_2513,In_652);
nor U636 (N_636,In_587,In_974);
and U637 (N_637,In_697,In_2442);
nand U638 (N_638,In_1645,In_1062);
or U639 (N_639,In_117,In_1195);
nand U640 (N_640,In_2602,In_2420);
or U641 (N_641,In_2791,In_313);
xor U642 (N_642,In_1955,In_1774);
xnor U643 (N_643,In_535,In_332);
and U644 (N_644,In_1434,In_56);
or U645 (N_645,In_936,In_1500);
nand U646 (N_646,In_349,In_1971);
nor U647 (N_647,In_1495,In_1209);
or U648 (N_648,In_2455,In_361);
and U649 (N_649,In_1830,In_2723);
and U650 (N_650,In_50,In_2627);
nand U651 (N_651,In_926,In_355);
nand U652 (N_652,In_1211,In_621);
xnor U653 (N_653,In_2487,In_602);
or U654 (N_654,In_1678,In_2607);
nand U655 (N_655,In_2180,In_137);
and U656 (N_656,In_2066,In_1129);
nand U657 (N_657,In_2306,In_2571);
nand U658 (N_658,In_695,In_1017);
xnor U659 (N_659,In_1854,In_57);
nand U660 (N_660,In_2313,In_1250);
xor U661 (N_661,In_433,In_2075);
nor U662 (N_662,In_614,In_1697);
and U663 (N_663,In_1013,In_2561);
and U664 (N_664,In_1075,In_424);
nand U665 (N_665,In_2469,In_2052);
or U666 (N_666,In_336,In_2228);
nor U667 (N_667,In_97,In_999);
and U668 (N_668,In_2415,In_347);
and U669 (N_669,In_1455,In_1579);
nor U670 (N_670,In_1652,In_1627);
or U671 (N_671,In_2537,In_2388);
and U672 (N_672,In_1777,In_981);
or U673 (N_673,In_2029,In_830);
nand U674 (N_674,In_1145,In_2809);
and U675 (N_675,In_2360,In_1808);
nand U676 (N_676,In_366,In_194);
nor U677 (N_677,In_539,In_2450);
nand U678 (N_678,In_550,In_1918);
and U679 (N_679,In_575,In_235);
and U680 (N_680,In_531,In_795);
xnor U681 (N_681,In_2953,In_1036);
nand U682 (N_682,In_2263,In_263);
nor U683 (N_683,In_1746,In_2024);
nand U684 (N_684,In_2981,In_605);
nor U685 (N_685,In_1621,In_2827);
xor U686 (N_686,In_1583,In_380);
and U687 (N_687,In_107,In_500);
and U688 (N_688,In_2629,In_573);
or U689 (N_689,In_1701,In_1690);
and U690 (N_690,In_2754,In_4);
nand U691 (N_691,In_2461,In_2968);
nand U692 (N_692,In_1422,In_267);
nand U693 (N_693,In_1864,In_290);
and U694 (N_694,In_759,In_1364);
nor U695 (N_695,In_475,In_1550);
nand U696 (N_696,In_1118,In_16);
or U697 (N_697,In_280,In_752);
and U698 (N_698,In_2856,In_356);
or U699 (N_699,In_383,In_1682);
nand U700 (N_700,In_166,In_192);
or U701 (N_701,In_2151,In_1440);
or U702 (N_702,In_1589,In_1445);
nor U703 (N_703,In_270,In_1361);
or U704 (N_704,In_2375,In_277);
and U705 (N_705,In_1991,In_2153);
nand U706 (N_706,In_344,In_2314);
nor U707 (N_707,In_2125,In_64);
and U708 (N_708,In_1597,In_2681);
or U709 (N_709,In_781,In_552);
nor U710 (N_710,In_2713,In_1940);
or U711 (N_711,In_1462,In_923);
nand U712 (N_712,In_1898,In_2023);
and U713 (N_713,In_1227,In_2867);
nand U714 (N_714,In_1393,In_2822);
or U715 (N_715,In_2552,In_1405);
nand U716 (N_716,In_674,In_1908);
or U717 (N_717,In_928,In_2405);
nand U718 (N_718,In_417,In_1804);
nand U719 (N_719,In_1699,In_1395);
nor U720 (N_720,In_1416,In_1531);
and U721 (N_721,In_1841,In_1301);
nand U722 (N_722,In_1593,In_2568);
and U723 (N_723,In_2460,In_1688);
or U724 (N_724,In_986,In_499);
and U725 (N_725,In_772,In_1766);
nand U726 (N_726,In_1691,In_1028);
and U727 (N_727,In_307,In_1204);
or U728 (N_728,In_2834,In_616);
and U729 (N_729,In_2099,In_2031);
or U730 (N_730,In_333,In_745);
and U731 (N_731,In_1720,In_2779);
or U732 (N_732,In_512,In_401);
nor U733 (N_733,In_382,In_1303);
or U734 (N_734,In_1139,In_2525);
nand U735 (N_735,In_1135,In_2403);
nor U736 (N_736,In_2407,In_2098);
nor U737 (N_737,In_1119,In_369);
or U738 (N_738,In_755,In_491);
nor U739 (N_739,In_1306,In_2730);
nor U740 (N_740,In_156,In_1184);
and U741 (N_741,In_2482,In_2543);
and U742 (N_742,In_2047,In_571);
and U743 (N_743,In_2729,In_804);
nand U744 (N_744,In_2079,In_2317);
nand U745 (N_745,In_2905,In_690);
nand U746 (N_746,In_945,In_1280);
nor U747 (N_747,In_476,In_1899);
nor U748 (N_748,In_1442,In_1484);
and U749 (N_749,In_2320,In_85);
nand U750 (N_750,In_1234,In_1427);
and U751 (N_751,In_856,In_2033);
and U752 (N_752,In_2645,In_506);
and U753 (N_753,In_1390,In_2861);
nor U754 (N_754,In_689,In_2937);
and U755 (N_755,In_2318,In_560);
or U756 (N_756,In_1751,In_644);
or U757 (N_757,In_1327,In_1820);
nor U758 (N_758,In_766,In_78);
nor U759 (N_759,In_59,In_647);
or U760 (N_760,In_931,In_2145);
or U761 (N_761,In_2739,In_2728);
nor U762 (N_762,In_2673,In_2106);
xor U763 (N_763,In_1748,In_1073);
nand U764 (N_764,In_1742,In_1480);
and U765 (N_765,In_190,In_1443);
or U766 (N_766,In_2233,In_1874);
or U767 (N_767,In_2924,In_1758);
nor U768 (N_768,In_2803,In_2389);
or U769 (N_769,In_2355,In_1952);
nand U770 (N_770,In_2735,In_2563);
nor U771 (N_771,In_451,In_1993);
nor U772 (N_772,In_1383,In_2689);
nor U773 (N_773,In_784,In_311);
and U774 (N_774,In_776,In_1823);
nor U775 (N_775,In_2816,In_174);
xor U776 (N_776,In_2208,In_1728);
nand U777 (N_777,In_1994,In_1602);
and U778 (N_778,In_2569,In_1088);
nand U779 (N_779,In_2662,In_1545);
xor U780 (N_780,In_505,In_47);
xor U781 (N_781,In_2481,In_846);
xnor U782 (N_782,In_2453,In_2536);
nand U783 (N_783,In_992,In_1043);
nor U784 (N_784,In_1710,In_481);
and U785 (N_785,In_2310,In_2296);
and U786 (N_786,In_2252,In_2001);
nand U787 (N_787,In_1452,In_1023);
nand U788 (N_788,In_1347,In_1926);
nor U789 (N_789,In_1072,In_2236);
nor U790 (N_790,In_2475,In_632);
nor U791 (N_791,In_322,In_83);
or U792 (N_792,In_2688,In_1465);
nand U793 (N_793,In_1608,In_389);
nand U794 (N_794,In_827,In_841);
nor U795 (N_795,In_634,In_1388);
or U796 (N_796,In_2472,In_2017);
nand U797 (N_797,In_517,In_1138);
nor U798 (N_798,In_2565,In_1011);
nor U799 (N_799,In_1656,In_1479);
and U800 (N_800,In_55,In_1203);
nand U801 (N_801,In_1852,In_2633);
xnor U802 (N_802,In_2904,In_2559);
nor U803 (N_803,In_2191,In_304);
nor U804 (N_804,In_1337,In_2722);
or U805 (N_805,In_1399,In_2889);
or U806 (N_806,In_2755,In_907);
and U807 (N_807,In_385,In_1381);
and U808 (N_808,In_1857,In_1225);
nor U809 (N_809,In_2658,In_2176);
and U810 (N_810,In_679,In_1713);
and U811 (N_811,In_2362,In_988);
nor U812 (N_812,In_2477,In_2441);
and U813 (N_813,In_160,In_1263);
xnor U814 (N_814,In_2842,In_291);
or U815 (N_815,In_317,In_515);
nand U816 (N_816,In_213,In_1588);
or U817 (N_817,In_1625,In_2665);
or U818 (N_818,In_2068,In_789);
xor U819 (N_819,In_487,In_139);
nor U820 (N_820,In_2192,In_400);
nor U821 (N_821,In_2112,In_2431);
or U822 (N_822,In_489,In_2190);
and U823 (N_823,In_1152,In_1876);
xnor U824 (N_824,In_2259,In_2280);
nor U825 (N_825,In_1787,In_2270);
nand U826 (N_826,In_763,In_2581);
xnor U827 (N_827,In_556,In_1846);
or U828 (N_828,In_628,In_688);
nand U829 (N_829,In_1607,In_1050);
and U830 (N_830,In_411,In_1979);
nor U831 (N_831,In_2496,In_2025);
xor U832 (N_832,In_2818,In_2587);
nor U833 (N_833,In_1768,In_2584);
nor U834 (N_834,In_1741,In_216);
or U835 (N_835,In_966,In_2749);
and U836 (N_836,In_1471,In_1446);
nand U837 (N_837,In_2901,In_2562);
nand U838 (N_838,In_2996,In_2782);
nand U839 (N_839,In_2817,In_76);
nor U840 (N_840,In_2349,In_1565);
and U841 (N_841,In_2711,In_1192);
nor U842 (N_842,In_2036,In_1745);
nor U843 (N_843,In_2174,In_271);
and U844 (N_844,In_100,In_1996);
or U845 (N_845,In_633,In_2770);
and U846 (N_846,In_2108,In_1007);
nand U847 (N_847,In_368,In_946);
nor U848 (N_848,In_1160,In_2214);
or U849 (N_849,In_2083,In_1283);
and U850 (N_850,In_1098,In_2637);
and U851 (N_851,In_2702,In_1035);
nand U852 (N_852,In_2866,In_1737);
xnor U853 (N_853,In_2102,In_302);
and U854 (N_854,In_2593,In_991);
nor U855 (N_855,In_566,In_215);
xor U856 (N_856,In_2691,In_1469);
nand U857 (N_857,In_504,In_2985);
or U858 (N_858,In_2873,In_1603);
or U859 (N_859,In_1329,In_1609);
nor U860 (N_860,In_579,In_2118);
nor U861 (N_861,In_1461,In_2435);
or U862 (N_862,In_1230,In_20);
and U863 (N_863,In_386,In_125);
or U864 (N_864,In_2970,In_1654);
and U865 (N_865,In_2262,In_663);
nand U866 (N_866,In_2275,In_877);
and U867 (N_867,In_2417,In_2895);
xor U868 (N_868,In_2693,In_1374);
nor U869 (N_869,In_885,In_892);
and U870 (N_870,In_1123,In_2143);
xor U871 (N_871,In_163,In_2641);
nand U872 (N_872,In_875,In_2218);
or U873 (N_873,In_1937,In_2276);
nor U874 (N_874,In_2196,In_1366);
nor U875 (N_875,In_1960,In_260);
and U876 (N_876,In_508,In_292);
nor U877 (N_877,In_1859,In_1387);
nor U878 (N_878,In_513,In_2070);
or U879 (N_879,In_259,In_2443);
nor U880 (N_880,In_1200,In_1883);
nand U881 (N_881,In_2065,In_768);
or U882 (N_882,In_1966,In_1109);
and U883 (N_883,In_1707,In_906);
xor U884 (N_884,In_365,In_399);
nand U885 (N_885,In_514,In_1817);
nand U886 (N_886,In_1144,In_2182);
and U887 (N_887,In_692,In_142);
nand U888 (N_888,In_1087,In_620);
and U889 (N_889,In_1566,In_1855);
nand U890 (N_890,In_1714,In_2983);
nor U891 (N_891,In_2363,In_1539);
xor U892 (N_892,In_1115,In_1884);
or U893 (N_893,In_310,In_2952);
nand U894 (N_894,In_1316,In_2660);
or U895 (N_895,In_1947,In_2621);
nand U896 (N_896,In_2960,In_2747);
nand U897 (N_897,In_2383,In_1924);
or U898 (N_898,In_1279,In_2021);
nand U899 (N_899,In_2638,In_2337);
nand U900 (N_900,In_537,In_2538);
or U901 (N_901,In_2928,In_2872);
xnor U902 (N_902,In_607,In_180);
nand U903 (N_903,In_2653,In_2674);
or U904 (N_904,In_738,In_529);
nor U905 (N_905,In_1369,In_1269);
and U906 (N_906,In_2342,In_2254);
or U907 (N_907,In_2510,In_25);
or U908 (N_908,In_488,In_808);
and U909 (N_909,In_2494,In_470);
and U910 (N_910,In_1671,In_1174);
nor U911 (N_911,In_783,In_116);
nand U912 (N_912,In_1801,In_728);
and U913 (N_913,In_1130,In_1964);
or U914 (N_914,In_2393,In_1515);
nor U915 (N_915,In_2203,In_2784);
and U916 (N_916,In_983,In_321);
or U917 (N_917,In_865,In_1941);
or U918 (N_918,In_2843,In_914);
or U919 (N_919,In_2121,In_2865);
nand U920 (N_920,In_2768,In_2580);
or U921 (N_921,In_2829,In_903);
nand U922 (N_922,In_2669,In_2111);
or U923 (N_923,In_1708,In_1885);
nand U924 (N_924,In_408,In_357);
nand U925 (N_925,In_1421,In_323);
nor U926 (N_926,In_598,In_2299);
nand U927 (N_927,In_1653,In_1207);
or U928 (N_928,In_2432,In_2643);
nor U929 (N_929,In_242,In_191);
xnor U930 (N_930,In_444,In_2366);
nor U931 (N_931,In_894,In_2447);
nor U932 (N_932,In_2715,In_2497);
nor U933 (N_933,In_969,In_2502);
and U934 (N_934,In_391,In_2466);
and U935 (N_935,In_2995,In_1619);
nand U936 (N_936,In_1560,In_793);
and U937 (N_937,In_932,In_450);
xor U938 (N_938,In_1643,In_1816);
nand U939 (N_939,In_2650,In_1727);
nand U940 (N_940,In_2835,In_2211);
xnor U941 (N_941,In_77,In_2260);
and U942 (N_942,In_1889,In_2799);
nand U943 (N_943,In_1582,In_978);
xor U944 (N_944,In_1562,In_122);
xnor U945 (N_945,In_2583,In_2444);
and U946 (N_946,In_1103,In_2463);
nand U947 (N_947,In_2719,In_1147);
nor U948 (N_948,In_1437,In_1837);
or U949 (N_949,In_1571,In_603);
nand U950 (N_950,In_230,In_140);
or U951 (N_951,In_2103,In_2076);
and U952 (N_952,In_326,In_432);
nor U953 (N_953,In_1176,In_1018);
nand U954 (N_954,In_2008,In_2969);
or U955 (N_955,In_1567,In_1460);
nand U956 (N_956,In_1978,In_618);
or U957 (N_957,In_1426,In_2737);
and U958 (N_958,In_2892,In_2586);
and U959 (N_959,In_1385,In_2836);
nor U960 (N_960,In_2830,In_1220);
xnor U961 (N_961,In_703,In_261);
xnor U962 (N_962,In_177,In_2085);
nand U963 (N_963,In_1640,In_1872);
and U964 (N_964,In_1287,In_1835);
xnor U965 (N_965,In_1882,In_325);
nor U966 (N_966,In_2000,In_1783);
nand U967 (N_967,In_1548,In_1517);
or U968 (N_968,In_45,In_1825);
and U969 (N_969,In_1042,In_581);
and U970 (N_970,In_1064,In_1893);
nand U971 (N_971,In_2838,In_2030);
and U972 (N_972,In_2707,In_2169);
nor U973 (N_973,In_1755,In_1116);
or U974 (N_974,In_1033,In_2193);
nor U975 (N_975,In_895,In_1216);
nand U976 (N_976,In_558,In_340);
and U977 (N_977,In_396,In_1121);
xnor U978 (N_978,In_1750,In_2281);
nor U979 (N_979,In_2906,In_2594);
nand U980 (N_980,In_2038,In_208);
nor U981 (N_981,In_62,In_42);
nand U982 (N_982,In_794,In_522);
nor U983 (N_983,In_296,In_1194);
or U984 (N_984,In_1934,In_276);
and U985 (N_985,In_1338,In_1060);
nor U986 (N_986,In_740,In_719);
and U987 (N_987,In_2519,In_67);
nand U988 (N_988,In_611,In_1037);
nor U989 (N_989,In_1376,In_2411);
nor U990 (N_990,In_1510,In_1084);
or U991 (N_991,In_1384,In_2132);
and U992 (N_992,In_1906,In_1407);
and U993 (N_993,In_360,In_2331);
or U994 (N_994,In_1128,In_2239);
and U995 (N_995,In_199,In_1595);
nor U996 (N_996,In_553,In_757);
nor U997 (N_997,In_1749,In_1698);
nor U998 (N_998,In_2741,In_376);
nand U999 (N_999,In_1819,In_2886);
nand U1000 (N_1000,In_584,In_1669);
and U1001 (N_1001,In_2426,In_498);
nor U1002 (N_1002,In_1473,In_694);
nor U1003 (N_1003,In_2949,In_2775);
nand U1004 (N_1004,In_785,In_1059);
and U1005 (N_1005,In_1305,In_2312);
or U1006 (N_1006,In_2922,In_2057);
nor U1007 (N_1007,In_549,In_2091);
nor U1008 (N_1008,In_2769,In_479);
or U1009 (N_1009,In_1920,In_495);
and U1010 (N_1010,In_709,In_924);
and U1011 (N_1011,In_1849,In_72);
and U1012 (N_1012,In_1127,In_2726);
nor U1013 (N_1013,In_2878,In_2625);
xnor U1014 (N_1014,In_1525,In_635);
or U1015 (N_1015,In_1170,In_612);
nand U1016 (N_1016,In_1298,In_2759);
or U1017 (N_1017,In_2958,In_1112);
nand U1018 (N_1018,In_1246,In_1812);
and U1019 (N_1019,In_1818,In_731);
nand U1020 (N_1020,In_2558,In_700);
or U1021 (N_1021,In_2304,In_1851);
or U1022 (N_1022,In_1377,In_1779);
and U1023 (N_1023,In_2950,In_1536);
nor U1024 (N_1024,In_2875,In_1193);
or U1025 (N_1025,In_223,In_2309);
xnor U1026 (N_1026,In_474,In_837);
nor U1027 (N_1027,In_1546,In_1863);
xnor U1028 (N_1028,In_570,In_1681);
and U1029 (N_1029,In_2230,In_1824);
and U1030 (N_1030,In_1805,In_2680);
xnor U1031 (N_1031,In_1523,In_2522);
and U1032 (N_1032,In_285,In_2635);
and U1033 (N_1033,In_2248,In_2699);
xnor U1034 (N_1034,In_1048,In_237);
xor U1035 (N_1035,In_1628,In_1564);
nor U1036 (N_1036,In_881,In_2324);
and U1037 (N_1037,In_1324,In_610);
nor U1038 (N_1038,In_657,In_1077);
nand U1039 (N_1039,In_617,In_165);
and U1040 (N_1040,In_915,In_1494);
and U1041 (N_1041,In_2398,In_1642);
nor U1042 (N_1042,In_1248,In_1686);
or U1043 (N_1043,In_430,In_2819);
and U1044 (N_1044,In_1051,In_2714);
nand U1045 (N_1045,In_901,In_2256);
nor U1046 (N_1046,In_1910,In_853);
or U1047 (N_1047,In_2185,In_2071);
nor U1048 (N_1048,In_442,In_497);
nand U1049 (N_1049,In_1620,In_39);
or U1050 (N_1050,In_1695,In_1521);
nand U1051 (N_1051,In_1258,In_2319);
nor U1052 (N_1052,In_2727,In_1504);
xor U1053 (N_1053,In_1171,In_2269);
or U1054 (N_1054,In_2423,In_1724);
nand U1055 (N_1055,In_1189,In_989);
nor U1056 (N_1056,In_732,In_2516);
nand U1057 (N_1057,In_2316,In_286);
nor U1058 (N_1058,In_1935,In_2850);
nand U1059 (N_1059,In_715,In_1378);
nand U1060 (N_1060,In_751,In_1005);
and U1061 (N_1061,In_2539,In_193);
or U1062 (N_1062,In_2195,In_66);
or U1063 (N_1063,In_250,In_1126);
nor U1064 (N_1064,In_2773,In_1351);
nand U1065 (N_1065,In_1718,In_710);
and U1066 (N_1066,In_1105,In_939);
nor U1067 (N_1067,In_2919,In_2134);
nor U1068 (N_1068,In_2676,In_527);
or U1069 (N_1069,In_1436,In_1458);
nand U1070 (N_1070,In_1637,In_113);
nor U1071 (N_1071,In_9,In_1892);
nand U1072 (N_1072,In_2894,In_1840);
xnor U1073 (N_1073,In_2798,In_934);
nand U1074 (N_1074,In_82,In_1191);
nor U1075 (N_1075,In_1371,In_454);
nand U1076 (N_1076,In_2572,In_228);
or U1077 (N_1077,In_1647,In_1958);
or U1078 (N_1078,In_1552,In_478);
or U1079 (N_1079,In_1342,In_1124);
nand U1080 (N_1080,In_26,In_2240);
nor U1081 (N_1081,In_2840,In_1962);
or U1082 (N_1082,In_1272,In_2073);
and U1083 (N_1083,In_2045,In_1775);
and U1084 (N_1084,In_2089,In_1254);
nor U1085 (N_1085,In_1459,In_2124);
or U1086 (N_1086,In_1450,In_951);
and U1087 (N_1087,In_2612,In_33);
and U1088 (N_1088,In_646,In_893);
and U1089 (N_1089,In_2753,In_1313);
nand U1090 (N_1090,In_2308,In_1693);
xor U1091 (N_1091,In_41,In_314);
nor U1092 (N_1092,In_1953,In_1277);
nand U1093 (N_1093,In_897,In_2703);
xor U1094 (N_1094,In_1626,In_469);
nor U1095 (N_1095,In_1219,In_1228);
nand U1096 (N_1096,In_171,In_24);
and U1097 (N_1097,In_2820,In_1065);
nor U1098 (N_1098,In_1125,In_1722);
and U1099 (N_1099,In_904,In_1373);
nor U1100 (N_1100,In_1685,In_1813);
nor U1101 (N_1101,In_362,In_899);
nand U1102 (N_1102,In_2911,In_684);
nand U1103 (N_1103,In_2902,In_279);
or U1104 (N_1104,In_2253,In_2382);
xor U1105 (N_1105,In_245,In_2074);
and U1106 (N_1106,In_1106,In_1300);
or U1107 (N_1107,In_2294,In_348);
nand U1108 (N_1108,In_1318,In_2035);
nor U1109 (N_1109,In_1650,In_2935);
or U1110 (N_1110,In_2984,In_38);
nor U1111 (N_1111,In_1444,In_1615);
nand U1112 (N_1112,In_341,In_2452);
xnor U1113 (N_1113,In_1604,In_289);
nor U1114 (N_1114,In_1244,In_883);
and U1115 (N_1115,In_2864,In_1928);
and U1116 (N_1116,In_1875,In_744);
nor U1117 (N_1117,In_1486,In_2266);
xnor U1118 (N_1118,In_339,In_203);
or U1119 (N_1119,In_2438,In_2434);
nor U1120 (N_1120,In_1478,In_2293);
nor U1121 (N_1121,In_1163,In_1581);
nor U1122 (N_1122,In_1925,In_2599);
and U1123 (N_1123,In_741,In_2080);
nor U1124 (N_1124,In_1312,In_1370);
or U1125 (N_1125,In_351,In_2042);
nand U1126 (N_1126,In_144,In_390);
nor U1127 (N_1127,In_435,In_2392);
and U1128 (N_1128,In_2395,In_183);
nand U1129 (N_1129,In_40,In_201);
nand U1130 (N_1130,In_1827,In_2120);
or U1131 (N_1131,In_492,In_1365);
nand U1132 (N_1132,In_1114,In_2041);
and U1133 (N_1133,In_1518,In_1078);
xor U1134 (N_1134,In_2793,In_2910);
nand U1135 (N_1135,In_2464,In_2764);
nand U1136 (N_1136,In_536,In_2364);
or U1137 (N_1137,In_582,In_1509);
and U1138 (N_1138,In_2011,In_1058);
nand U1139 (N_1139,In_2550,In_2409);
or U1140 (N_1140,In_824,In_414);
or U1141 (N_1141,In_2171,In_2564);
and U1142 (N_1142,In_2573,In_2142);
xor U1143 (N_1143,In_65,In_1723);
nand U1144 (N_1144,In_1717,In_1815);
and U1145 (N_1145,In_252,In_1320);
or U1146 (N_1146,In_1785,In_849);
nand U1147 (N_1147,In_1453,In_2971);
xor U1148 (N_1148,In_1802,In_402);
and U1149 (N_1149,In_1541,In_2386);
and U1150 (N_1150,In_656,In_120);
nand U1151 (N_1151,In_2474,In_1340);
nor U1152 (N_1152,In_1870,In_613);
and U1153 (N_1153,In_1454,In_1253);
nor U1154 (N_1154,In_1181,In_2999);
nor U1155 (N_1155,In_214,In_110);
xnor U1156 (N_1156,In_2626,In_761);
nor U1157 (N_1157,In_1530,In_1466);
nand U1158 (N_1158,In_583,In_2307);
nor U1159 (N_1159,In_2140,In_70);
or U1160 (N_1160,In_685,In_2631);
and U1161 (N_1161,In_1136,In_1843);
and U1162 (N_1162,In_858,In_2851);
xor U1163 (N_1163,In_2846,In_2860);
nand U1164 (N_1164,In_2436,In_669);
or U1165 (N_1165,In_1570,In_189);
nor U1166 (N_1166,In_859,In_1367);
nand U1167 (N_1167,In_1946,In_2670);
nand U1168 (N_1168,In_869,In_1950);
nor U1169 (N_1169,In_2272,In_2274);
or U1170 (N_1170,In_1346,In_2210);
or U1171 (N_1171,In_2286,In_1789);
and U1172 (N_1172,In_2265,In_129);
xor U1173 (N_1173,In_559,In_747);
xnor U1174 (N_1174,In_1284,In_1639);
nand U1175 (N_1175,In_994,In_288);
or U1176 (N_1176,In_2189,In_2786);
or U1177 (N_1177,In_714,In_2848);
xor U1178 (N_1178,In_2148,In_2914);
nor U1179 (N_1179,In_890,In_596);
xor U1180 (N_1180,In_1357,In_2797);
or U1181 (N_1181,In_2505,In_2261);
nand U1182 (N_1182,In_1296,In_2101);
nand U1183 (N_1183,In_708,In_2242);
or U1184 (N_1184,In_1822,In_301);
or U1185 (N_1185,In_1557,In_485);
or U1186 (N_1186,In_1847,In_1132);
nand U1187 (N_1187,In_1010,In_1508);
and U1188 (N_1188,In_1363,In_2998);
or U1189 (N_1189,In_1215,In_2883);
nand U1190 (N_1190,In_844,In_636);
nand U1191 (N_1191,In_716,In_1336);
and U1192 (N_1192,In_1198,In_2989);
nand U1193 (N_1193,In_2515,In_1273);
nand U1194 (N_1194,In_2756,In_461);
nand U1195 (N_1195,In_950,In_916);
or U1196 (N_1196,In_2357,In_170);
nor U1197 (N_1197,In_241,In_363);
nand U1198 (N_1198,In_431,In_197);
or U1199 (N_1199,In_2600,In_1532);
or U1200 (N_1200,In_31,In_155);
and U1201 (N_1201,In_2340,In_2871);
nor U1202 (N_1202,In_2709,In_1512);
nand U1203 (N_1203,In_811,In_2321);
nor U1204 (N_1204,In_1786,In_511);
nand U1205 (N_1205,In_2807,In_466);
nor U1206 (N_1206,In_227,In_2868);
nor U1207 (N_1207,In_1795,In_1501);
nand U1208 (N_1208,In_2523,In_2530);
xor U1209 (N_1209,In_819,In_682);
and U1210 (N_1210,In_2250,In_388);
nor U1211 (N_1211,In_791,In_820);
and U1212 (N_1212,In_75,In_2974);
nor U1213 (N_1213,In_1806,In_2994);
and U1214 (N_1214,In_1923,In_2133);
nand U1215 (N_1215,In_2857,In_2327);
or U1216 (N_1216,In_2870,In_1949);
nor U1217 (N_1217,In_2810,In_1986);
or U1218 (N_1218,In_562,In_1166);
nor U1219 (N_1219,In_769,In_1345);
and U1220 (N_1220,In_239,In_1190);
and U1221 (N_1221,In_1729,In_965);
and U1222 (N_1222,In_1074,In_2005);
xnor U1223 (N_1223,In_2687,In_240);
and U1224 (N_1224,In_2344,In_2598);
and U1225 (N_1225,In_1677,In_2166);
and U1226 (N_1226,In_2772,In_2548);
nor U1227 (N_1227,In_1992,In_439);
and U1228 (N_1228,In_1288,In_1753);
nor U1229 (N_1229,In_2610,In_778);
nor U1230 (N_1230,In_2554,In_1502);
nor U1231 (N_1231,In_2332,In_2742);
or U1232 (N_1232,In_593,In_2);
and U1233 (N_1233,In_1811,In_748);
nand U1234 (N_1234,In_2508,In_2222);
nand U1235 (N_1235,In_1025,In_835);
nor U1236 (N_1236,In_1826,In_851);
and U1237 (N_1237,In_2979,In_138);
nor U1238 (N_1238,In_2642,In_1308);
and U1239 (N_1239,In_2223,In_154);
nor U1240 (N_1240,In_957,In_2880);
nor U1241 (N_1241,In_1936,In_1529);
or U1242 (N_1242,In_2815,In_1409);
nand U1243 (N_1243,In_1569,In_544);
or U1244 (N_1244,In_1890,In_1315);
xnor U1245 (N_1245,In_1623,In_108);
nor U1246 (N_1246,In_1261,In_874);
nor U1247 (N_1247,In_687,In_1726);
xor U1248 (N_1248,In_1240,In_1257);
xor U1249 (N_1249,In_896,In_2657);
nor U1250 (N_1250,In_7,In_667);
or U1251 (N_1251,In_577,In_2339);
xor U1252 (N_1252,In_1319,In_2622);
and U1253 (N_1253,In_2578,In_1360);
and U1254 (N_1254,In_2943,In_2760);
or U1255 (N_1255,In_1967,In_2158);
and U1256 (N_1256,In_1206,In_2617);
nand U1257 (N_1257,In_2448,In_1794);
nor U1258 (N_1258,In_937,In_175);
or U1259 (N_1259,In_1973,In_1886);
and U1260 (N_1260,In_105,In_2097);
or U1261 (N_1261,In_600,In_1120);
or U1262 (N_1262,In_997,In_2012);
nand U1263 (N_1263,In_2698,In_2311);
nand U1264 (N_1264,In_2736,In_1481);
or U1265 (N_1265,In_817,In_350);
nand U1266 (N_1266,In_2027,In_1499);
nand U1267 (N_1267,In_792,In_521);
nor U1268 (N_1268,In_1535,In_2907);
and U1269 (N_1269,In_1239,In_1401);
or U1270 (N_1270,In_1880,In_210);
nand U1271 (N_1271,In_2199,In_1398);
or U1272 (N_1272,In_206,In_1079);
and U1273 (N_1273,In_37,In_467);
nand U1274 (N_1274,In_756,In_1931);
and U1275 (N_1275,In_61,In_2589);
and U1276 (N_1276,In_1091,In_207);
nand U1277 (N_1277,In_1957,In_1800);
or U1278 (N_1278,In_2654,In_540);
nor U1279 (N_1279,In_220,In_661);
or U1280 (N_1280,In_229,In_2207);
nor U1281 (N_1281,In_1039,In_520);
and U1282 (N_1282,In_2605,In_836);
nand U1283 (N_1283,In_2763,In_1330);
nor U1284 (N_1284,In_1561,In_1406);
and U1285 (N_1285,In_840,In_706);
and U1286 (N_1286,In_1836,In_717);
or U1287 (N_1287,In_1881,In_1848);
nand U1288 (N_1288,In_1334,In_2141);
or U1289 (N_1289,In_1551,In_1543);
xnor U1290 (N_1290,In_1238,In_1476);
and U1291 (N_1291,In_929,In_554);
nor U1292 (N_1292,In_920,In_1679);
and U1293 (N_1293,In_2081,In_749);
xor U1294 (N_1294,In_10,In_1100);
nor U1295 (N_1295,In_1980,In_1188);
nand U1296 (N_1296,In_2430,In_2965);
nor U1297 (N_1297,In_609,In_1655);
or U1298 (N_1298,In_2231,In_2806);
nor U1299 (N_1299,In_209,In_1762);
and U1300 (N_1300,In_2899,In_384);
or U1301 (N_1301,In_234,In_2903);
nor U1302 (N_1302,In_463,In_284);
xnor U1303 (N_1303,In_2933,In_666);
nor U1304 (N_1304,In_2655,In_246);
and U1305 (N_1305,In_815,In_2716);
or U1306 (N_1306,In_2322,In_2088);
xnor U1307 (N_1307,In_1662,In_606);
nor U1308 (N_1308,In_1956,In_2408);
and U1309 (N_1309,In_645,In_2206);
and U1310 (N_1310,In_2451,In_1232);
nand U1311 (N_1311,In_2853,In_2987);
nor U1312 (N_1312,In_2113,In_1606);
nand U1313 (N_1313,In_952,In_918);
and U1314 (N_1314,In_2028,In_1251);
xor U1315 (N_1315,In_1666,In_2936);
xor U1316 (N_1316,In_2939,In_886);
nand U1317 (N_1317,In_2499,In_2695);
and U1318 (N_1318,In_838,In_510);
or U1319 (N_1319,In_2414,In_1759);
nor U1320 (N_1320,In_2608,In_665);
nor U1321 (N_1321,In_954,In_440);
or U1322 (N_1322,In_854,In_2679);
nand U1323 (N_1323,In_262,In_1719);
nand U1324 (N_1324,In_343,In_68);
and U1325 (N_1325,In_739,In_828);
nor U1326 (N_1326,In_1533,In_1547);
nor U1327 (N_1327,In_493,In_959);
or U1328 (N_1328,In_2473,In_1891);
nand U1329 (N_1329,In_2100,In_422);
and U1330 (N_1330,In_453,In_643);
and U1331 (N_1331,In_2288,In_1052);
nand U1332 (N_1332,In_2279,In_44);
or U1333 (N_1333,In_2845,In_441);
xor U1334 (N_1334,In_2348,In_1111);
nor U1335 (N_1335,In_436,In_604);
nor U1336 (N_1336,In_1948,In_990);
nand U1337 (N_1337,In_1069,In_146);
and U1338 (N_1338,In_1809,In_2762);
nor U1339 (N_1339,In_1379,In_2675);
and U1340 (N_1340,In_1538,In_1270);
nand U1341 (N_1341,In_725,In_2954);
and U1342 (N_1342,In_2710,In_2858);
and U1343 (N_1343,In_2397,In_1617);
nand U1344 (N_1344,In_2942,In_2051);
nor U1345 (N_1345,In_211,In_2429);
xor U1346 (N_1346,In_1391,In_1141);
nand U1347 (N_1347,In_1086,In_2410);
or U1348 (N_1348,In_309,In_2541);
and U1349 (N_1349,In_164,In_872);
nand U1350 (N_1350,In_1754,In_2748);
and U1351 (N_1351,In_1266,In_2697);
nor U1352 (N_1352,In_810,In_834);
nor U1353 (N_1353,In_1519,In_1447);
and U1354 (N_1354,In_2213,In_1725);
xor U1355 (N_1355,In_2235,In_507);
nand U1356 (N_1356,In_2315,In_452);
nor U1357 (N_1357,In_2962,In_2620);
and U1358 (N_1358,In_1006,In_502);
or U1359 (N_1359,In_1689,In_1887);
or U1360 (N_1360,In_2305,In_2381);
nand U1361 (N_1361,In_299,In_2110);
or U1362 (N_1362,In_352,In_2717);
xor U1363 (N_1363,In_642,In_2267);
nor U1364 (N_1364,In_2015,In_623);
or U1365 (N_1365,In_2406,In_1352);
or U1366 (N_1366,In_121,In_2394);
nor U1367 (N_1367,In_1556,In_130);
and U1368 (N_1368,In_145,In_2685);
or U1369 (N_1369,In_1999,In_2067);
xnor U1370 (N_1370,In_1858,In_2026);
xnor U1371 (N_1371,In_2524,In_1414);
and U1372 (N_1372,In_2966,In_1922);
xor U1373 (N_1373,In_1223,In_2632);
and U1374 (N_1374,In_1871,In_1467);
nand U1375 (N_1375,In_1358,In_455);
nor U1376 (N_1376,In_1137,In_753);
or U1377 (N_1377,In_2506,In_2007);
or U1378 (N_1378,In_1175,In_1782);
and U1379 (N_1379,In_1131,In_2869);
or U1380 (N_1380,In_1428,In_1162);
nand U1381 (N_1381,In_943,In_330);
and U1382 (N_1382,In_876,In_1732);
nor U1383 (N_1383,In_2465,In_1790);
and U1384 (N_1384,In_115,In_995);
nor U1385 (N_1385,In_1757,In_1981);
and U1386 (N_1386,In_2783,In_816);
nor U1387 (N_1387,In_2813,In_2478);
nor U1388 (N_1388,In_1423,In_1304);
and U1389 (N_1389,In_1798,In_2358);
or U1390 (N_1390,In_1769,In_2721);
nand U1391 (N_1391,In_2964,In_2161);
nor U1392 (N_1392,In_86,In_1022);
nand U1393 (N_1393,In_2533,In_2972);
and U1394 (N_1394,In_315,In_1574);
xor U1395 (N_1395,In_1528,In_2700);
nand U1396 (N_1396,In_168,In_1168);
nor U1397 (N_1397,In_2359,In_2130);
nand U1398 (N_1398,In_696,In_91);
and U1399 (N_1399,In_1030,In_585);
and U1400 (N_1400,In_765,In_2446);
or U1401 (N_1401,In_2825,In_1747);
and U1402 (N_1402,In_2146,In_2855);
nand U1403 (N_1403,In_2277,In_813);
or U1404 (N_1404,In_2811,In_1271);
or U1405 (N_1405,In_1605,In_426);
and U1406 (N_1406,In_2649,In_1229);
nand U1407 (N_1407,In_403,In_2991);
nand U1408 (N_1408,In_2217,In_1591);
nor U1409 (N_1409,In_1916,In_2704);
xnor U1410 (N_1410,In_21,In_1056);
nand U1411 (N_1411,In_2582,In_2812);
and U1412 (N_1412,In_92,In_2247);
nand U1413 (N_1413,In_397,In_126);
and U1414 (N_1414,In_707,In_1046);
xnor U1415 (N_1415,In_1396,In_2613);
nor U1416 (N_1416,In_729,In_691);
and U1417 (N_1417,In_2597,In_329);
nor U1418 (N_1418,In_2347,In_2944);
and U1419 (N_1419,In_2086,In_2187);
nor U1420 (N_1420,In_1668,In_1791);
or U1421 (N_1421,In_2198,In_1799);
nand U1422 (N_1422,In_1448,In_801);
or U1423 (N_1423,In_1638,In_919);
nor U1424 (N_1424,In_394,In_95);
nand U1425 (N_1425,In_2489,In_2412);
xnor U1426 (N_1426,In_324,In_1236);
or U1427 (N_1427,In_501,In_1489);
or U1428 (N_1428,In_1122,In_99);
nor U1429 (N_1429,In_779,In_2380);
nand U1430 (N_1430,In_524,In_882);
nand U1431 (N_1431,In_1470,In_676);
xnor U1432 (N_1432,In_1505,In_2285);
xor U1433 (N_1433,In_2518,In_2890);
nand U1434 (N_1434,In_1054,In_1101);
nand U1435 (N_1435,In_1900,In_1000);
nand U1436 (N_1436,In_1932,In_530);
nor U1437 (N_1437,In_942,In_15);
xor U1438 (N_1438,In_1153,In_1983);
xor U1439 (N_1439,In_169,In_1403);
and U1440 (N_1440,In_346,In_948);
nand U1441 (N_1441,In_1260,In_735);
nor U1442 (N_1442,In_181,In_1933);
and U1443 (N_1443,In_2888,In_2640);
nand U1444 (N_1444,In_71,In_1990);
nand U1445 (N_1445,In_1156,In_2639);
nor U1446 (N_1446,In_1066,In_412);
nand U1447 (N_1447,In_425,In_2761);
and U1448 (N_1448,In_2004,In_46);
or U1449 (N_1449,In_2909,In_1404);
nand U1450 (N_1450,In_1432,In_589);
xor U1451 (N_1451,In_668,In_1441);
or U1452 (N_1452,In_2445,In_1089);
and U1453 (N_1453,In_2577,In_961);
xnor U1454 (N_1454,In_2232,In_1449);
and U1455 (N_1455,In_1178,In_2732);
and U1456 (N_1456,In_2493,In_650);
and U1457 (N_1457,In_2646,In_1286);
and U1458 (N_1458,In_2037,In_1915);
nand U1459 (N_1459,In_822,In_627);
nand U1460 (N_1460,In_1780,In_1293);
and U1461 (N_1461,In_132,In_2221);
nand U1462 (N_1462,In_1117,In_2663);
nand U1463 (N_1463,In_1332,In_1828);
xnor U1464 (N_1464,In_1411,In_2069);
or U1465 (N_1465,In_2694,In_2611);
nand U1466 (N_1466,In_2127,In_1233);
nand U1467 (N_1467,In_217,In_1879);
xnor U1468 (N_1468,In_2273,In_231);
xnor U1469 (N_1469,In_27,In_670);
or U1470 (N_1470,In_87,In_1400);
nand U1471 (N_1471,In_1034,In_2457);
xnor U1472 (N_1472,In_1939,In_184);
or U1473 (N_1473,In_1559,In_996);
nand U1474 (N_1474,In_1630,In_1904);
nand U1475 (N_1475,In_2800,In_2205);
xnor U1476 (N_1476,In_1516,In_1492);
or U1477 (N_1477,In_1110,In_2128);
nand U1478 (N_1478,In_32,In_935);
nor U1479 (N_1479,In_1350,In_1410);
and U1480 (N_1480,In_2003,In_2164);
xnor U1481 (N_1481,In_2325,In_2659);
and U1482 (N_1482,In_2839,In_1807);
nand U1483 (N_1483,In_2354,In_938);
and U1484 (N_1484,In_158,In_1068);
and U1485 (N_1485,In_1102,In_398);
nand U1486 (N_1486,In_167,In_395);
nand U1487 (N_1487,In_1972,In_2781);
nand U1488 (N_1488,In_1081,In_101);
nor U1489 (N_1489,In_545,In_1814);
nor U1490 (N_1490,In_594,In_2225);
nor U1491 (N_1491,In_626,In_198);
and U1492 (N_1492,In_1016,In_5);
and U1493 (N_1493,In_2766,In_1325);
or U1494 (N_1494,In_1333,In_157);
and U1495 (N_1495,In_2500,In_631);
nor U1496 (N_1496,In_2179,In_2604);
nand U1497 (N_1497,In_773,In_2601);
nand U1498 (N_1498,In_823,In_253);
nor U1499 (N_1499,In_1281,In_1954);
xor U1500 (N_1500,In_39,In_1871);
and U1501 (N_1501,In_1548,In_2498);
nor U1502 (N_1502,In_2481,In_1331);
nor U1503 (N_1503,In_2632,In_1969);
or U1504 (N_1504,In_1244,In_2029);
or U1505 (N_1505,In_474,In_2227);
and U1506 (N_1506,In_2036,In_2874);
nor U1507 (N_1507,In_2474,In_600);
and U1508 (N_1508,In_942,In_2495);
nor U1509 (N_1509,In_2194,In_1715);
and U1510 (N_1510,In_1364,In_2091);
or U1511 (N_1511,In_2363,In_636);
and U1512 (N_1512,In_2970,In_2780);
or U1513 (N_1513,In_993,In_2620);
xnor U1514 (N_1514,In_770,In_2045);
nor U1515 (N_1515,In_159,In_760);
nand U1516 (N_1516,In_415,In_1711);
and U1517 (N_1517,In_385,In_834);
nand U1518 (N_1518,In_2055,In_2790);
nand U1519 (N_1519,In_272,In_1635);
and U1520 (N_1520,In_1327,In_840);
nor U1521 (N_1521,In_294,In_426);
or U1522 (N_1522,In_1644,In_263);
or U1523 (N_1523,In_712,In_224);
or U1524 (N_1524,In_1400,In_2837);
nand U1525 (N_1525,In_2493,In_2562);
and U1526 (N_1526,In_2385,In_2706);
nor U1527 (N_1527,In_96,In_2497);
nand U1528 (N_1528,In_2218,In_2443);
or U1529 (N_1529,In_672,In_443);
xnor U1530 (N_1530,In_1413,In_2648);
nand U1531 (N_1531,In_1973,In_443);
nand U1532 (N_1532,In_1138,In_889);
nor U1533 (N_1533,In_570,In_2845);
nand U1534 (N_1534,In_1949,In_1455);
and U1535 (N_1535,In_2113,In_937);
nand U1536 (N_1536,In_1645,In_458);
xor U1537 (N_1537,In_1420,In_1734);
nand U1538 (N_1538,In_1224,In_1099);
nor U1539 (N_1539,In_1950,In_1238);
xnor U1540 (N_1540,In_2176,In_2148);
and U1541 (N_1541,In_590,In_2874);
nor U1542 (N_1542,In_1800,In_1784);
or U1543 (N_1543,In_2150,In_1841);
or U1544 (N_1544,In_788,In_1809);
xor U1545 (N_1545,In_614,In_925);
nand U1546 (N_1546,In_2212,In_2263);
nand U1547 (N_1547,In_586,In_2662);
nor U1548 (N_1548,In_715,In_2042);
or U1549 (N_1549,In_726,In_364);
nand U1550 (N_1550,In_1707,In_2147);
or U1551 (N_1551,In_729,In_1394);
nor U1552 (N_1552,In_787,In_2451);
or U1553 (N_1553,In_231,In_1546);
and U1554 (N_1554,In_2614,In_2942);
or U1555 (N_1555,In_2680,In_285);
or U1556 (N_1556,In_1549,In_2181);
nor U1557 (N_1557,In_2364,In_2206);
xnor U1558 (N_1558,In_2623,In_916);
nor U1559 (N_1559,In_1712,In_2235);
nor U1560 (N_1560,In_1419,In_1200);
and U1561 (N_1561,In_672,In_568);
nor U1562 (N_1562,In_526,In_2345);
and U1563 (N_1563,In_222,In_292);
nor U1564 (N_1564,In_2000,In_158);
and U1565 (N_1565,In_311,In_962);
nor U1566 (N_1566,In_2252,In_2078);
and U1567 (N_1567,In_293,In_353);
nor U1568 (N_1568,In_2312,In_496);
nor U1569 (N_1569,In_2234,In_389);
nand U1570 (N_1570,In_1617,In_2024);
xor U1571 (N_1571,In_2059,In_1301);
and U1572 (N_1572,In_671,In_2751);
nand U1573 (N_1573,In_864,In_1782);
nor U1574 (N_1574,In_754,In_843);
or U1575 (N_1575,In_2304,In_741);
or U1576 (N_1576,In_747,In_1983);
nand U1577 (N_1577,In_247,In_1690);
nand U1578 (N_1578,In_2654,In_1203);
or U1579 (N_1579,In_2555,In_2977);
or U1580 (N_1580,In_659,In_938);
nor U1581 (N_1581,In_1165,In_1513);
nand U1582 (N_1582,In_1587,In_1698);
nand U1583 (N_1583,In_673,In_1532);
nor U1584 (N_1584,In_1891,In_443);
and U1585 (N_1585,In_2476,In_2482);
and U1586 (N_1586,In_907,In_1657);
xor U1587 (N_1587,In_2306,In_2586);
and U1588 (N_1588,In_192,In_1467);
and U1589 (N_1589,In_132,In_2478);
or U1590 (N_1590,In_2567,In_100);
nor U1591 (N_1591,In_2133,In_562);
and U1592 (N_1592,In_510,In_1397);
or U1593 (N_1593,In_652,In_614);
nor U1594 (N_1594,In_1974,In_59);
nor U1595 (N_1595,In_389,In_2356);
and U1596 (N_1596,In_1096,In_516);
or U1597 (N_1597,In_2258,In_2388);
and U1598 (N_1598,In_2316,In_1028);
xor U1599 (N_1599,In_2166,In_1057);
nor U1600 (N_1600,In_165,In_1559);
nor U1601 (N_1601,In_547,In_241);
or U1602 (N_1602,In_2516,In_904);
xor U1603 (N_1603,In_1476,In_789);
nand U1604 (N_1604,In_1665,In_74);
nor U1605 (N_1605,In_1806,In_1399);
nor U1606 (N_1606,In_2967,In_53);
or U1607 (N_1607,In_149,In_1498);
or U1608 (N_1608,In_1949,In_1634);
nand U1609 (N_1609,In_1914,In_813);
or U1610 (N_1610,In_2198,In_1756);
nor U1611 (N_1611,In_988,In_1069);
and U1612 (N_1612,In_470,In_893);
or U1613 (N_1613,In_2716,In_1067);
nand U1614 (N_1614,In_2005,In_1348);
and U1615 (N_1615,In_1522,In_2691);
nor U1616 (N_1616,In_1773,In_226);
nand U1617 (N_1617,In_874,In_152);
and U1618 (N_1618,In_1972,In_909);
or U1619 (N_1619,In_141,In_506);
xor U1620 (N_1620,In_1196,In_1114);
nand U1621 (N_1621,In_1921,In_1525);
or U1622 (N_1622,In_2600,In_1666);
nor U1623 (N_1623,In_730,In_726);
or U1624 (N_1624,In_1718,In_995);
and U1625 (N_1625,In_2071,In_2999);
nand U1626 (N_1626,In_2374,In_2557);
nor U1627 (N_1627,In_730,In_2485);
nor U1628 (N_1628,In_374,In_1898);
xor U1629 (N_1629,In_2744,In_2025);
or U1630 (N_1630,In_671,In_1409);
and U1631 (N_1631,In_166,In_507);
nand U1632 (N_1632,In_2417,In_1074);
nand U1633 (N_1633,In_56,In_652);
nand U1634 (N_1634,In_1179,In_2978);
and U1635 (N_1635,In_2250,In_1326);
nand U1636 (N_1636,In_2647,In_1420);
nor U1637 (N_1637,In_751,In_2319);
nand U1638 (N_1638,In_747,In_1248);
nor U1639 (N_1639,In_1789,In_653);
and U1640 (N_1640,In_706,In_2873);
and U1641 (N_1641,In_499,In_1409);
or U1642 (N_1642,In_1632,In_1102);
nor U1643 (N_1643,In_928,In_2408);
nor U1644 (N_1644,In_2635,In_800);
nand U1645 (N_1645,In_558,In_1696);
nor U1646 (N_1646,In_285,In_1151);
or U1647 (N_1647,In_1211,In_2152);
and U1648 (N_1648,In_2092,In_1958);
nor U1649 (N_1649,In_1686,In_2546);
nor U1650 (N_1650,In_2744,In_1535);
or U1651 (N_1651,In_2896,In_69);
nand U1652 (N_1652,In_720,In_2688);
or U1653 (N_1653,In_2604,In_1137);
nor U1654 (N_1654,In_2182,In_355);
or U1655 (N_1655,In_2554,In_1322);
or U1656 (N_1656,In_244,In_2695);
or U1657 (N_1657,In_1542,In_1449);
nand U1658 (N_1658,In_457,In_1984);
nor U1659 (N_1659,In_2880,In_318);
and U1660 (N_1660,In_1202,In_2682);
nor U1661 (N_1661,In_993,In_647);
nand U1662 (N_1662,In_242,In_1948);
or U1663 (N_1663,In_2043,In_1257);
nand U1664 (N_1664,In_2164,In_1218);
or U1665 (N_1665,In_1227,In_1981);
xor U1666 (N_1666,In_1947,In_262);
nor U1667 (N_1667,In_528,In_1403);
nand U1668 (N_1668,In_1501,In_309);
nand U1669 (N_1669,In_2775,In_2410);
or U1670 (N_1670,In_1273,In_714);
nand U1671 (N_1671,In_899,In_842);
and U1672 (N_1672,In_2315,In_2025);
and U1673 (N_1673,In_1358,In_2580);
or U1674 (N_1674,In_1807,In_2031);
and U1675 (N_1675,In_484,In_2886);
nand U1676 (N_1676,In_1799,In_156);
nor U1677 (N_1677,In_1274,In_2433);
and U1678 (N_1678,In_597,In_448);
nor U1679 (N_1679,In_1115,In_2962);
or U1680 (N_1680,In_2309,In_2252);
or U1681 (N_1681,In_2746,In_2008);
nor U1682 (N_1682,In_586,In_1656);
and U1683 (N_1683,In_1809,In_2808);
and U1684 (N_1684,In_963,In_797);
nand U1685 (N_1685,In_50,In_2617);
nand U1686 (N_1686,In_1575,In_2539);
nor U1687 (N_1687,In_2333,In_2271);
and U1688 (N_1688,In_2345,In_2287);
and U1689 (N_1689,In_564,In_2753);
and U1690 (N_1690,In_2247,In_2010);
or U1691 (N_1691,In_138,In_1367);
and U1692 (N_1692,In_1781,In_1831);
or U1693 (N_1693,In_2880,In_1283);
xnor U1694 (N_1694,In_2055,In_2742);
nor U1695 (N_1695,In_9,In_1498);
xor U1696 (N_1696,In_253,In_942);
and U1697 (N_1697,In_1717,In_1933);
and U1698 (N_1698,In_2292,In_1527);
and U1699 (N_1699,In_2312,In_1443);
xor U1700 (N_1700,In_1427,In_2329);
and U1701 (N_1701,In_2255,In_1524);
and U1702 (N_1702,In_2139,In_1409);
and U1703 (N_1703,In_1102,In_2749);
or U1704 (N_1704,In_1631,In_2586);
xnor U1705 (N_1705,In_2935,In_617);
nor U1706 (N_1706,In_90,In_2237);
nor U1707 (N_1707,In_1882,In_190);
nand U1708 (N_1708,In_2316,In_2968);
nor U1709 (N_1709,In_1923,In_396);
nand U1710 (N_1710,In_2534,In_2744);
and U1711 (N_1711,In_2929,In_531);
nand U1712 (N_1712,In_2085,In_1937);
and U1713 (N_1713,In_1743,In_1777);
or U1714 (N_1714,In_610,In_1218);
or U1715 (N_1715,In_2838,In_1092);
and U1716 (N_1716,In_1044,In_1475);
nor U1717 (N_1717,In_722,In_1471);
and U1718 (N_1718,In_2173,In_1657);
nand U1719 (N_1719,In_625,In_2244);
and U1720 (N_1720,In_2494,In_267);
or U1721 (N_1721,In_781,In_1208);
nand U1722 (N_1722,In_998,In_1558);
nor U1723 (N_1723,In_1500,In_1842);
or U1724 (N_1724,In_1707,In_591);
xnor U1725 (N_1725,In_1085,In_1535);
nand U1726 (N_1726,In_1142,In_382);
nor U1727 (N_1727,In_783,In_1394);
or U1728 (N_1728,In_1859,In_13);
and U1729 (N_1729,In_1153,In_2222);
xor U1730 (N_1730,In_591,In_454);
nor U1731 (N_1731,In_1582,In_866);
xnor U1732 (N_1732,In_1876,In_1235);
and U1733 (N_1733,In_1337,In_102);
and U1734 (N_1734,In_2117,In_2345);
nand U1735 (N_1735,In_2053,In_1679);
xnor U1736 (N_1736,In_958,In_622);
or U1737 (N_1737,In_1845,In_1894);
nor U1738 (N_1738,In_1258,In_2823);
nand U1739 (N_1739,In_1464,In_655);
nor U1740 (N_1740,In_762,In_1751);
nand U1741 (N_1741,In_2370,In_797);
and U1742 (N_1742,In_1951,In_601);
nand U1743 (N_1743,In_262,In_2273);
and U1744 (N_1744,In_2223,In_2577);
and U1745 (N_1745,In_2545,In_1615);
nor U1746 (N_1746,In_440,In_1209);
or U1747 (N_1747,In_1727,In_319);
and U1748 (N_1748,In_540,In_2503);
nor U1749 (N_1749,In_1678,In_615);
nor U1750 (N_1750,In_1994,In_181);
or U1751 (N_1751,In_2818,In_76);
or U1752 (N_1752,In_2478,In_1110);
xor U1753 (N_1753,In_868,In_1228);
nand U1754 (N_1754,In_1763,In_981);
nor U1755 (N_1755,In_1598,In_1419);
or U1756 (N_1756,In_2392,In_1401);
and U1757 (N_1757,In_2298,In_2156);
nor U1758 (N_1758,In_1215,In_2418);
or U1759 (N_1759,In_1147,In_2654);
or U1760 (N_1760,In_2531,In_1486);
nor U1761 (N_1761,In_651,In_504);
nand U1762 (N_1762,In_373,In_2514);
xnor U1763 (N_1763,In_2290,In_2728);
and U1764 (N_1764,In_1246,In_929);
nand U1765 (N_1765,In_2635,In_1970);
or U1766 (N_1766,In_1640,In_2840);
nor U1767 (N_1767,In_2149,In_352);
and U1768 (N_1768,In_1215,In_2022);
or U1769 (N_1769,In_1809,In_1727);
nand U1770 (N_1770,In_1004,In_568);
nand U1771 (N_1771,In_566,In_610);
nor U1772 (N_1772,In_1251,In_1379);
nor U1773 (N_1773,In_715,In_92);
and U1774 (N_1774,In_60,In_1860);
nand U1775 (N_1775,In_808,In_2192);
nand U1776 (N_1776,In_1589,In_2220);
or U1777 (N_1777,In_729,In_2700);
and U1778 (N_1778,In_2180,In_2760);
nor U1779 (N_1779,In_1228,In_1169);
or U1780 (N_1780,In_1762,In_1146);
xor U1781 (N_1781,In_2827,In_1305);
nand U1782 (N_1782,In_2897,In_773);
nand U1783 (N_1783,In_1936,In_472);
xnor U1784 (N_1784,In_672,In_1694);
and U1785 (N_1785,In_158,In_2733);
nand U1786 (N_1786,In_2591,In_879);
nand U1787 (N_1787,In_2414,In_2291);
or U1788 (N_1788,In_1655,In_873);
and U1789 (N_1789,In_1256,In_1912);
nor U1790 (N_1790,In_2532,In_644);
xnor U1791 (N_1791,In_1238,In_1873);
nor U1792 (N_1792,In_2054,In_1031);
and U1793 (N_1793,In_2832,In_255);
nand U1794 (N_1794,In_2630,In_2410);
nand U1795 (N_1795,In_1194,In_1568);
or U1796 (N_1796,In_835,In_1985);
or U1797 (N_1797,In_1044,In_2777);
nand U1798 (N_1798,In_2604,In_643);
nor U1799 (N_1799,In_1571,In_2347);
nand U1800 (N_1800,In_875,In_1597);
xor U1801 (N_1801,In_2278,In_1034);
nand U1802 (N_1802,In_1806,In_825);
nor U1803 (N_1803,In_1770,In_1276);
nand U1804 (N_1804,In_395,In_781);
nor U1805 (N_1805,In_1882,In_1339);
nand U1806 (N_1806,In_274,In_2515);
or U1807 (N_1807,In_2513,In_2231);
xor U1808 (N_1808,In_1270,In_1909);
and U1809 (N_1809,In_1610,In_2212);
or U1810 (N_1810,In_2603,In_374);
nand U1811 (N_1811,In_1172,In_2114);
nor U1812 (N_1812,In_2753,In_265);
or U1813 (N_1813,In_2124,In_1102);
nor U1814 (N_1814,In_157,In_2777);
nor U1815 (N_1815,In_589,In_1721);
nand U1816 (N_1816,In_1958,In_1149);
nor U1817 (N_1817,In_2012,In_1334);
nand U1818 (N_1818,In_479,In_2360);
or U1819 (N_1819,In_1157,In_324);
and U1820 (N_1820,In_1520,In_2728);
and U1821 (N_1821,In_2671,In_1489);
or U1822 (N_1822,In_2886,In_469);
or U1823 (N_1823,In_1960,In_767);
or U1824 (N_1824,In_123,In_1422);
nor U1825 (N_1825,In_2975,In_2687);
nand U1826 (N_1826,In_1235,In_830);
nand U1827 (N_1827,In_764,In_1847);
or U1828 (N_1828,In_1556,In_1528);
nor U1829 (N_1829,In_1799,In_1062);
nand U1830 (N_1830,In_171,In_2334);
and U1831 (N_1831,In_1919,In_1479);
or U1832 (N_1832,In_1594,In_2518);
nor U1833 (N_1833,In_1722,In_1868);
nor U1834 (N_1834,In_1218,In_312);
and U1835 (N_1835,In_1289,In_981);
nor U1836 (N_1836,In_658,In_2916);
and U1837 (N_1837,In_2030,In_1598);
xnor U1838 (N_1838,In_1080,In_2282);
and U1839 (N_1839,In_594,In_623);
nand U1840 (N_1840,In_2138,In_859);
nor U1841 (N_1841,In_177,In_22);
and U1842 (N_1842,In_1781,In_1105);
or U1843 (N_1843,In_2968,In_1579);
nor U1844 (N_1844,In_2159,In_1518);
nor U1845 (N_1845,In_791,In_1837);
nor U1846 (N_1846,In_776,In_542);
xor U1847 (N_1847,In_876,In_1003);
and U1848 (N_1848,In_199,In_657);
or U1849 (N_1849,In_1819,In_1356);
nand U1850 (N_1850,In_2034,In_2739);
nor U1851 (N_1851,In_1475,In_807);
nand U1852 (N_1852,In_1840,In_363);
xor U1853 (N_1853,In_598,In_2712);
or U1854 (N_1854,In_772,In_1157);
nand U1855 (N_1855,In_1942,In_2125);
xnor U1856 (N_1856,In_938,In_2803);
or U1857 (N_1857,In_1748,In_1182);
and U1858 (N_1858,In_140,In_1747);
nand U1859 (N_1859,In_1205,In_1469);
nor U1860 (N_1860,In_88,In_539);
or U1861 (N_1861,In_77,In_178);
nand U1862 (N_1862,In_1798,In_2577);
nor U1863 (N_1863,In_2863,In_1010);
nand U1864 (N_1864,In_1633,In_1374);
xnor U1865 (N_1865,In_401,In_302);
nand U1866 (N_1866,In_2763,In_1574);
nor U1867 (N_1867,In_1222,In_2048);
and U1868 (N_1868,In_2982,In_936);
xnor U1869 (N_1869,In_321,In_252);
xor U1870 (N_1870,In_791,In_288);
nand U1871 (N_1871,In_444,In_1456);
nand U1872 (N_1872,In_2537,In_1792);
or U1873 (N_1873,In_2486,In_2361);
and U1874 (N_1874,In_362,In_236);
and U1875 (N_1875,In_1594,In_1039);
nand U1876 (N_1876,In_1709,In_852);
nand U1877 (N_1877,In_2688,In_1693);
and U1878 (N_1878,In_1729,In_1826);
or U1879 (N_1879,In_2791,In_928);
or U1880 (N_1880,In_2813,In_1258);
or U1881 (N_1881,In_38,In_1421);
or U1882 (N_1882,In_1761,In_2303);
and U1883 (N_1883,In_1048,In_1885);
or U1884 (N_1884,In_845,In_348);
or U1885 (N_1885,In_1057,In_1616);
or U1886 (N_1886,In_1268,In_27);
xor U1887 (N_1887,In_2232,In_2145);
xnor U1888 (N_1888,In_2079,In_439);
or U1889 (N_1889,In_1879,In_1063);
and U1890 (N_1890,In_2886,In_1156);
nand U1891 (N_1891,In_2031,In_1959);
nor U1892 (N_1892,In_2289,In_1671);
or U1893 (N_1893,In_649,In_2098);
and U1894 (N_1894,In_1544,In_2082);
nor U1895 (N_1895,In_2367,In_35);
nand U1896 (N_1896,In_1331,In_52);
and U1897 (N_1897,In_1528,In_1905);
or U1898 (N_1898,In_2114,In_1007);
and U1899 (N_1899,In_1911,In_1443);
or U1900 (N_1900,In_1414,In_750);
nor U1901 (N_1901,In_2346,In_1051);
nand U1902 (N_1902,In_708,In_63);
nor U1903 (N_1903,In_177,In_1813);
nand U1904 (N_1904,In_1021,In_2666);
or U1905 (N_1905,In_24,In_1584);
nand U1906 (N_1906,In_671,In_1602);
nand U1907 (N_1907,In_2736,In_7);
or U1908 (N_1908,In_2363,In_831);
nand U1909 (N_1909,In_0,In_1623);
nand U1910 (N_1910,In_1136,In_220);
nand U1911 (N_1911,In_1504,In_861);
nand U1912 (N_1912,In_895,In_2716);
or U1913 (N_1913,In_1785,In_650);
or U1914 (N_1914,In_1629,In_1034);
xor U1915 (N_1915,In_1947,In_1815);
or U1916 (N_1916,In_1645,In_597);
nor U1917 (N_1917,In_1858,In_1912);
and U1918 (N_1918,In_427,In_2351);
nand U1919 (N_1919,In_2350,In_381);
nand U1920 (N_1920,In_294,In_937);
or U1921 (N_1921,In_1143,In_1490);
xor U1922 (N_1922,In_1724,In_1344);
and U1923 (N_1923,In_2959,In_638);
and U1924 (N_1924,In_1755,In_360);
nor U1925 (N_1925,In_905,In_172);
or U1926 (N_1926,In_1171,In_1345);
or U1927 (N_1927,In_2868,In_2186);
nand U1928 (N_1928,In_628,In_841);
or U1929 (N_1929,In_772,In_1134);
and U1930 (N_1930,In_921,In_9);
or U1931 (N_1931,In_765,In_2376);
nand U1932 (N_1932,In_2658,In_594);
nand U1933 (N_1933,In_1102,In_2496);
nor U1934 (N_1934,In_2359,In_2352);
nand U1935 (N_1935,In_2203,In_316);
nor U1936 (N_1936,In_509,In_2812);
and U1937 (N_1937,In_2396,In_317);
and U1938 (N_1938,In_2972,In_2380);
nor U1939 (N_1939,In_1409,In_634);
xnor U1940 (N_1940,In_2880,In_1138);
nor U1941 (N_1941,In_1287,In_2388);
nor U1942 (N_1942,In_2496,In_1974);
nor U1943 (N_1943,In_1170,In_829);
nor U1944 (N_1944,In_893,In_2108);
nor U1945 (N_1945,In_2739,In_513);
and U1946 (N_1946,In_2779,In_2410);
or U1947 (N_1947,In_1555,In_1528);
xor U1948 (N_1948,In_257,In_537);
and U1949 (N_1949,In_636,In_283);
nor U1950 (N_1950,In_2258,In_2819);
nand U1951 (N_1951,In_2853,In_558);
xor U1952 (N_1952,In_27,In_1041);
xnor U1953 (N_1953,In_1904,In_1810);
or U1954 (N_1954,In_2266,In_1811);
and U1955 (N_1955,In_1688,In_1198);
or U1956 (N_1956,In_418,In_2045);
nand U1957 (N_1957,In_1835,In_761);
or U1958 (N_1958,In_1317,In_2712);
nor U1959 (N_1959,In_596,In_180);
xor U1960 (N_1960,In_554,In_2468);
and U1961 (N_1961,In_478,In_2520);
or U1962 (N_1962,In_302,In_2529);
nand U1963 (N_1963,In_2539,In_1021);
xor U1964 (N_1964,In_2498,In_1641);
nand U1965 (N_1965,In_1652,In_1425);
xor U1966 (N_1966,In_319,In_723);
nor U1967 (N_1967,In_2388,In_1594);
nor U1968 (N_1968,In_1549,In_383);
xor U1969 (N_1969,In_255,In_536);
or U1970 (N_1970,In_733,In_332);
and U1971 (N_1971,In_1404,In_2194);
nor U1972 (N_1972,In_2153,In_1474);
and U1973 (N_1973,In_553,In_2879);
nor U1974 (N_1974,In_2259,In_740);
or U1975 (N_1975,In_1677,In_2774);
nor U1976 (N_1976,In_812,In_1036);
xor U1977 (N_1977,In_2387,In_2433);
nor U1978 (N_1978,In_804,In_1201);
or U1979 (N_1979,In_821,In_349);
nand U1980 (N_1980,In_1806,In_155);
nor U1981 (N_1981,In_1075,In_602);
nand U1982 (N_1982,In_226,In_504);
or U1983 (N_1983,In_2582,In_962);
nand U1984 (N_1984,In_2206,In_1992);
nor U1985 (N_1985,In_1281,In_1043);
and U1986 (N_1986,In_1086,In_217);
nand U1987 (N_1987,In_167,In_705);
nor U1988 (N_1988,In_2616,In_1301);
nor U1989 (N_1989,In_1915,In_323);
or U1990 (N_1990,In_622,In_1947);
and U1991 (N_1991,In_2278,In_2206);
and U1992 (N_1992,In_1611,In_395);
and U1993 (N_1993,In_2262,In_2531);
nand U1994 (N_1994,In_1794,In_969);
or U1995 (N_1995,In_885,In_2256);
nand U1996 (N_1996,In_2776,In_2817);
nand U1997 (N_1997,In_1723,In_1901);
nand U1998 (N_1998,In_1633,In_2271);
and U1999 (N_1999,In_2838,In_2740);
or U2000 (N_2000,In_235,In_2262);
and U2001 (N_2001,In_517,In_2391);
xnor U2002 (N_2002,In_2022,In_1904);
or U2003 (N_2003,In_217,In_1717);
or U2004 (N_2004,In_917,In_601);
nand U2005 (N_2005,In_2033,In_810);
nand U2006 (N_2006,In_2031,In_649);
nor U2007 (N_2007,In_34,In_415);
and U2008 (N_2008,In_365,In_2556);
nor U2009 (N_2009,In_1644,In_498);
or U2010 (N_2010,In_2317,In_740);
or U2011 (N_2011,In_2432,In_2031);
and U2012 (N_2012,In_2963,In_745);
or U2013 (N_2013,In_443,In_151);
or U2014 (N_2014,In_937,In_1129);
nand U2015 (N_2015,In_2615,In_307);
nand U2016 (N_2016,In_25,In_277);
nor U2017 (N_2017,In_2351,In_511);
and U2018 (N_2018,In_88,In_716);
and U2019 (N_2019,In_2375,In_2936);
or U2020 (N_2020,In_284,In_25);
or U2021 (N_2021,In_558,In_2216);
or U2022 (N_2022,In_2382,In_713);
nor U2023 (N_2023,In_2120,In_2815);
or U2024 (N_2024,In_22,In_2347);
xor U2025 (N_2025,In_1461,In_1609);
or U2026 (N_2026,In_1609,In_2172);
nor U2027 (N_2027,In_310,In_1912);
nand U2028 (N_2028,In_2320,In_2801);
nand U2029 (N_2029,In_2384,In_2151);
and U2030 (N_2030,In_1802,In_72);
nor U2031 (N_2031,In_2902,In_536);
and U2032 (N_2032,In_1715,In_1544);
nor U2033 (N_2033,In_1312,In_1106);
or U2034 (N_2034,In_1952,In_2816);
nand U2035 (N_2035,In_2997,In_199);
or U2036 (N_2036,In_628,In_843);
or U2037 (N_2037,In_1088,In_1937);
nand U2038 (N_2038,In_999,In_941);
or U2039 (N_2039,In_2048,In_1890);
nor U2040 (N_2040,In_314,In_361);
and U2041 (N_2041,In_2902,In_1945);
nor U2042 (N_2042,In_2427,In_1677);
or U2043 (N_2043,In_2730,In_1227);
nor U2044 (N_2044,In_2897,In_1125);
or U2045 (N_2045,In_581,In_2140);
nand U2046 (N_2046,In_1388,In_2777);
and U2047 (N_2047,In_1041,In_1463);
or U2048 (N_2048,In_1374,In_1240);
and U2049 (N_2049,In_2629,In_1049);
nand U2050 (N_2050,In_264,In_1888);
nand U2051 (N_2051,In_422,In_1680);
nand U2052 (N_2052,In_2619,In_2648);
nand U2053 (N_2053,In_2095,In_2661);
or U2054 (N_2054,In_714,In_2112);
and U2055 (N_2055,In_314,In_1404);
nand U2056 (N_2056,In_1177,In_482);
nand U2057 (N_2057,In_2744,In_450);
nor U2058 (N_2058,In_1742,In_2682);
nor U2059 (N_2059,In_2843,In_2033);
or U2060 (N_2060,In_2953,In_366);
and U2061 (N_2061,In_2996,In_833);
and U2062 (N_2062,In_2734,In_2248);
nor U2063 (N_2063,In_1812,In_758);
nand U2064 (N_2064,In_1926,In_2886);
or U2065 (N_2065,In_1557,In_2581);
nor U2066 (N_2066,In_859,In_860);
xnor U2067 (N_2067,In_1805,In_1004);
or U2068 (N_2068,In_2967,In_36);
or U2069 (N_2069,In_588,In_380);
xor U2070 (N_2070,In_1478,In_8);
or U2071 (N_2071,In_2392,In_2806);
nand U2072 (N_2072,In_1008,In_1040);
or U2073 (N_2073,In_2348,In_1306);
or U2074 (N_2074,In_641,In_1100);
nor U2075 (N_2075,In_2009,In_2107);
nand U2076 (N_2076,In_443,In_411);
or U2077 (N_2077,In_888,In_2133);
or U2078 (N_2078,In_2647,In_865);
xor U2079 (N_2079,In_2726,In_2552);
xnor U2080 (N_2080,In_1339,In_2441);
nand U2081 (N_2081,In_518,In_1517);
nor U2082 (N_2082,In_2684,In_1652);
nand U2083 (N_2083,In_533,In_289);
nand U2084 (N_2084,In_1214,In_1331);
or U2085 (N_2085,In_2200,In_1083);
nand U2086 (N_2086,In_2101,In_2119);
nor U2087 (N_2087,In_481,In_1439);
nand U2088 (N_2088,In_819,In_2025);
and U2089 (N_2089,In_2028,In_1098);
nand U2090 (N_2090,In_1789,In_929);
nor U2091 (N_2091,In_2817,In_2016);
nor U2092 (N_2092,In_1456,In_907);
nor U2093 (N_2093,In_1478,In_794);
or U2094 (N_2094,In_2718,In_258);
or U2095 (N_2095,In_59,In_637);
nand U2096 (N_2096,In_252,In_2216);
xor U2097 (N_2097,In_265,In_726);
nand U2098 (N_2098,In_2906,In_528);
nor U2099 (N_2099,In_656,In_833);
nor U2100 (N_2100,In_1382,In_2271);
nor U2101 (N_2101,In_1796,In_1424);
nor U2102 (N_2102,In_2117,In_354);
and U2103 (N_2103,In_54,In_2831);
and U2104 (N_2104,In_2978,In_522);
or U2105 (N_2105,In_2524,In_841);
nor U2106 (N_2106,In_2837,In_2211);
or U2107 (N_2107,In_2843,In_2533);
nand U2108 (N_2108,In_1090,In_1967);
nor U2109 (N_2109,In_1039,In_1786);
or U2110 (N_2110,In_1030,In_2121);
xor U2111 (N_2111,In_2315,In_2687);
nand U2112 (N_2112,In_2977,In_43);
nand U2113 (N_2113,In_2926,In_648);
or U2114 (N_2114,In_1737,In_2226);
xnor U2115 (N_2115,In_1072,In_2531);
nor U2116 (N_2116,In_2011,In_1607);
nor U2117 (N_2117,In_725,In_1548);
nor U2118 (N_2118,In_2658,In_1437);
or U2119 (N_2119,In_640,In_1942);
or U2120 (N_2120,In_183,In_2493);
nand U2121 (N_2121,In_1709,In_1012);
and U2122 (N_2122,In_2352,In_671);
nor U2123 (N_2123,In_475,In_2727);
nand U2124 (N_2124,In_2549,In_2761);
or U2125 (N_2125,In_901,In_1308);
or U2126 (N_2126,In_1239,In_1820);
nor U2127 (N_2127,In_2442,In_64);
nor U2128 (N_2128,In_1535,In_1287);
nand U2129 (N_2129,In_904,In_858);
or U2130 (N_2130,In_1976,In_2340);
nor U2131 (N_2131,In_1249,In_1919);
xor U2132 (N_2132,In_2021,In_2018);
nor U2133 (N_2133,In_151,In_1336);
or U2134 (N_2134,In_1812,In_1592);
and U2135 (N_2135,In_1452,In_2444);
and U2136 (N_2136,In_236,In_1232);
nor U2137 (N_2137,In_1146,In_283);
nand U2138 (N_2138,In_686,In_1552);
and U2139 (N_2139,In_169,In_1667);
nand U2140 (N_2140,In_367,In_2490);
and U2141 (N_2141,In_1383,In_682);
or U2142 (N_2142,In_342,In_131);
or U2143 (N_2143,In_2418,In_2873);
and U2144 (N_2144,In_1103,In_1658);
nor U2145 (N_2145,In_216,In_25);
or U2146 (N_2146,In_1312,In_686);
or U2147 (N_2147,In_1305,In_2002);
or U2148 (N_2148,In_2397,In_2615);
and U2149 (N_2149,In_1498,In_759);
nand U2150 (N_2150,In_1554,In_2629);
and U2151 (N_2151,In_2636,In_2792);
and U2152 (N_2152,In_350,In_264);
or U2153 (N_2153,In_1453,In_2218);
or U2154 (N_2154,In_192,In_2244);
or U2155 (N_2155,In_682,In_2462);
nor U2156 (N_2156,In_2413,In_1010);
and U2157 (N_2157,In_1536,In_1375);
or U2158 (N_2158,In_553,In_2065);
nand U2159 (N_2159,In_276,In_1317);
and U2160 (N_2160,In_146,In_2934);
or U2161 (N_2161,In_2993,In_2222);
and U2162 (N_2162,In_2857,In_2874);
or U2163 (N_2163,In_770,In_886);
or U2164 (N_2164,In_305,In_186);
nor U2165 (N_2165,In_969,In_2530);
xnor U2166 (N_2166,In_255,In_2732);
nand U2167 (N_2167,In_2332,In_2746);
nor U2168 (N_2168,In_308,In_1287);
nor U2169 (N_2169,In_1845,In_1031);
nand U2170 (N_2170,In_1379,In_1802);
or U2171 (N_2171,In_1051,In_490);
and U2172 (N_2172,In_1681,In_2730);
and U2173 (N_2173,In_2760,In_2866);
and U2174 (N_2174,In_2055,In_604);
or U2175 (N_2175,In_584,In_634);
and U2176 (N_2176,In_2160,In_1765);
xor U2177 (N_2177,In_1127,In_630);
xnor U2178 (N_2178,In_32,In_1031);
and U2179 (N_2179,In_1335,In_1112);
or U2180 (N_2180,In_2724,In_772);
or U2181 (N_2181,In_109,In_2263);
nor U2182 (N_2182,In_1759,In_2409);
or U2183 (N_2183,In_1189,In_2546);
or U2184 (N_2184,In_2024,In_371);
or U2185 (N_2185,In_88,In_2084);
or U2186 (N_2186,In_1137,In_931);
xnor U2187 (N_2187,In_2102,In_1229);
nor U2188 (N_2188,In_770,In_1592);
xnor U2189 (N_2189,In_411,In_2191);
nor U2190 (N_2190,In_444,In_1778);
or U2191 (N_2191,In_1289,In_1543);
or U2192 (N_2192,In_2793,In_2736);
or U2193 (N_2193,In_582,In_350);
nor U2194 (N_2194,In_138,In_2584);
and U2195 (N_2195,In_2031,In_2215);
nor U2196 (N_2196,In_737,In_2247);
nor U2197 (N_2197,In_904,In_39);
or U2198 (N_2198,In_515,In_2125);
nor U2199 (N_2199,In_2829,In_314);
nand U2200 (N_2200,In_2790,In_2487);
and U2201 (N_2201,In_1360,In_736);
nand U2202 (N_2202,In_1783,In_2440);
nor U2203 (N_2203,In_1239,In_2081);
xnor U2204 (N_2204,In_1261,In_1451);
nor U2205 (N_2205,In_2718,In_704);
and U2206 (N_2206,In_2047,In_2966);
or U2207 (N_2207,In_2457,In_2944);
and U2208 (N_2208,In_1362,In_1160);
and U2209 (N_2209,In_642,In_102);
nor U2210 (N_2210,In_1552,In_999);
nor U2211 (N_2211,In_1682,In_2880);
and U2212 (N_2212,In_2863,In_1247);
nor U2213 (N_2213,In_549,In_53);
or U2214 (N_2214,In_2794,In_2927);
and U2215 (N_2215,In_718,In_2615);
or U2216 (N_2216,In_1509,In_2948);
and U2217 (N_2217,In_2910,In_2619);
and U2218 (N_2218,In_409,In_281);
nor U2219 (N_2219,In_2268,In_603);
nand U2220 (N_2220,In_2532,In_1044);
and U2221 (N_2221,In_1016,In_1655);
nor U2222 (N_2222,In_2557,In_1511);
nor U2223 (N_2223,In_938,In_2344);
nor U2224 (N_2224,In_2595,In_825);
or U2225 (N_2225,In_1955,In_2290);
xnor U2226 (N_2226,In_2594,In_1274);
nand U2227 (N_2227,In_1710,In_452);
or U2228 (N_2228,In_1315,In_2677);
nand U2229 (N_2229,In_1574,In_1938);
and U2230 (N_2230,In_2827,In_2637);
and U2231 (N_2231,In_2849,In_975);
nand U2232 (N_2232,In_1419,In_896);
nor U2233 (N_2233,In_2651,In_1970);
nand U2234 (N_2234,In_630,In_1738);
and U2235 (N_2235,In_2488,In_938);
nand U2236 (N_2236,In_1742,In_2094);
or U2237 (N_2237,In_1703,In_779);
and U2238 (N_2238,In_826,In_2231);
nor U2239 (N_2239,In_1693,In_2646);
or U2240 (N_2240,In_2030,In_2355);
nor U2241 (N_2241,In_2605,In_2919);
nand U2242 (N_2242,In_216,In_2572);
and U2243 (N_2243,In_2614,In_1989);
nor U2244 (N_2244,In_2052,In_700);
or U2245 (N_2245,In_1586,In_951);
nor U2246 (N_2246,In_2648,In_2401);
or U2247 (N_2247,In_2689,In_1822);
nor U2248 (N_2248,In_1949,In_835);
and U2249 (N_2249,In_802,In_1003);
and U2250 (N_2250,In_387,In_1597);
or U2251 (N_2251,In_2871,In_919);
and U2252 (N_2252,In_1536,In_2488);
and U2253 (N_2253,In_2752,In_2873);
nor U2254 (N_2254,In_371,In_6);
and U2255 (N_2255,In_742,In_60);
nor U2256 (N_2256,In_2644,In_891);
nand U2257 (N_2257,In_2328,In_1589);
nand U2258 (N_2258,In_2824,In_441);
and U2259 (N_2259,In_2357,In_1030);
or U2260 (N_2260,In_2293,In_446);
or U2261 (N_2261,In_1337,In_2380);
nand U2262 (N_2262,In_2174,In_755);
and U2263 (N_2263,In_1240,In_287);
or U2264 (N_2264,In_2847,In_1190);
or U2265 (N_2265,In_450,In_1406);
nor U2266 (N_2266,In_2401,In_2785);
nand U2267 (N_2267,In_1841,In_2104);
nor U2268 (N_2268,In_2921,In_2077);
nor U2269 (N_2269,In_2634,In_2251);
nand U2270 (N_2270,In_2525,In_2391);
nor U2271 (N_2271,In_408,In_1174);
nor U2272 (N_2272,In_846,In_1204);
nand U2273 (N_2273,In_182,In_2087);
nand U2274 (N_2274,In_247,In_1268);
or U2275 (N_2275,In_1086,In_1231);
or U2276 (N_2276,In_429,In_1260);
and U2277 (N_2277,In_2810,In_728);
or U2278 (N_2278,In_2692,In_231);
nand U2279 (N_2279,In_1954,In_2953);
and U2280 (N_2280,In_524,In_1996);
nand U2281 (N_2281,In_430,In_2010);
nor U2282 (N_2282,In_800,In_2753);
nor U2283 (N_2283,In_1257,In_680);
or U2284 (N_2284,In_319,In_1089);
or U2285 (N_2285,In_1594,In_1835);
or U2286 (N_2286,In_1443,In_1696);
nor U2287 (N_2287,In_1336,In_348);
nor U2288 (N_2288,In_2719,In_2947);
nand U2289 (N_2289,In_2451,In_2933);
nor U2290 (N_2290,In_1388,In_490);
and U2291 (N_2291,In_790,In_1243);
nor U2292 (N_2292,In_1656,In_740);
nand U2293 (N_2293,In_2955,In_2775);
nor U2294 (N_2294,In_1945,In_705);
and U2295 (N_2295,In_386,In_1351);
or U2296 (N_2296,In_118,In_861);
and U2297 (N_2297,In_2132,In_1107);
nand U2298 (N_2298,In_1878,In_900);
nor U2299 (N_2299,In_31,In_1063);
xor U2300 (N_2300,In_1966,In_1799);
and U2301 (N_2301,In_850,In_1831);
xor U2302 (N_2302,In_2832,In_1999);
xor U2303 (N_2303,In_2173,In_2631);
nor U2304 (N_2304,In_622,In_2568);
nor U2305 (N_2305,In_2684,In_2162);
nand U2306 (N_2306,In_2982,In_2326);
nor U2307 (N_2307,In_2121,In_2788);
and U2308 (N_2308,In_226,In_2701);
nor U2309 (N_2309,In_951,In_1423);
or U2310 (N_2310,In_1981,In_1215);
or U2311 (N_2311,In_730,In_2378);
nor U2312 (N_2312,In_2631,In_2262);
nor U2313 (N_2313,In_2137,In_1687);
nor U2314 (N_2314,In_553,In_2036);
nand U2315 (N_2315,In_2306,In_363);
nand U2316 (N_2316,In_2495,In_1629);
nand U2317 (N_2317,In_1102,In_2540);
and U2318 (N_2318,In_931,In_142);
or U2319 (N_2319,In_829,In_1846);
and U2320 (N_2320,In_690,In_1142);
xnor U2321 (N_2321,In_6,In_488);
and U2322 (N_2322,In_2894,In_1101);
nor U2323 (N_2323,In_1722,In_1786);
nand U2324 (N_2324,In_2182,In_2108);
nand U2325 (N_2325,In_826,In_797);
xnor U2326 (N_2326,In_2248,In_26);
nor U2327 (N_2327,In_326,In_2844);
nand U2328 (N_2328,In_1404,In_1214);
nor U2329 (N_2329,In_228,In_1423);
nand U2330 (N_2330,In_2048,In_1437);
and U2331 (N_2331,In_2980,In_580);
nor U2332 (N_2332,In_624,In_2927);
or U2333 (N_2333,In_2939,In_1819);
and U2334 (N_2334,In_158,In_2508);
nor U2335 (N_2335,In_1491,In_1581);
nor U2336 (N_2336,In_1444,In_1812);
and U2337 (N_2337,In_2054,In_600);
xor U2338 (N_2338,In_1409,In_389);
or U2339 (N_2339,In_2973,In_1542);
and U2340 (N_2340,In_1694,In_349);
and U2341 (N_2341,In_1000,In_2789);
and U2342 (N_2342,In_1813,In_2163);
nand U2343 (N_2343,In_2482,In_1922);
or U2344 (N_2344,In_1873,In_479);
or U2345 (N_2345,In_1731,In_117);
or U2346 (N_2346,In_530,In_1856);
or U2347 (N_2347,In_1204,In_720);
nand U2348 (N_2348,In_2687,In_1886);
nor U2349 (N_2349,In_105,In_1040);
nor U2350 (N_2350,In_1125,In_1376);
or U2351 (N_2351,In_1287,In_517);
and U2352 (N_2352,In_188,In_2629);
or U2353 (N_2353,In_2386,In_2018);
nor U2354 (N_2354,In_2809,In_1250);
xor U2355 (N_2355,In_1964,In_2932);
nand U2356 (N_2356,In_493,In_1780);
nor U2357 (N_2357,In_213,In_145);
or U2358 (N_2358,In_2447,In_1405);
nand U2359 (N_2359,In_768,In_2027);
xor U2360 (N_2360,In_1259,In_1444);
nand U2361 (N_2361,In_2971,In_1698);
nand U2362 (N_2362,In_5,In_970);
or U2363 (N_2363,In_1190,In_2842);
and U2364 (N_2364,In_1705,In_2197);
xor U2365 (N_2365,In_836,In_1972);
and U2366 (N_2366,In_99,In_1106);
and U2367 (N_2367,In_2307,In_716);
nor U2368 (N_2368,In_2546,In_1850);
nor U2369 (N_2369,In_1230,In_1036);
or U2370 (N_2370,In_2665,In_1569);
nor U2371 (N_2371,In_1365,In_407);
or U2372 (N_2372,In_2435,In_1710);
nor U2373 (N_2373,In_1076,In_1937);
and U2374 (N_2374,In_872,In_272);
or U2375 (N_2375,In_1644,In_747);
or U2376 (N_2376,In_740,In_511);
and U2377 (N_2377,In_1822,In_262);
xnor U2378 (N_2378,In_1049,In_111);
nor U2379 (N_2379,In_2258,In_1649);
or U2380 (N_2380,In_390,In_367);
and U2381 (N_2381,In_2279,In_2680);
nand U2382 (N_2382,In_1915,In_683);
xnor U2383 (N_2383,In_1630,In_371);
or U2384 (N_2384,In_1153,In_350);
nor U2385 (N_2385,In_2124,In_192);
nand U2386 (N_2386,In_2343,In_1065);
or U2387 (N_2387,In_1605,In_835);
xor U2388 (N_2388,In_727,In_2536);
nor U2389 (N_2389,In_2536,In_974);
nor U2390 (N_2390,In_2123,In_2071);
or U2391 (N_2391,In_315,In_2634);
nand U2392 (N_2392,In_47,In_703);
xor U2393 (N_2393,In_2776,In_1333);
nor U2394 (N_2394,In_28,In_675);
or U2395 (N_2395,In_2264,In_440);
or U2396 (N_2396,In_2483,In_2984);
or U2397 (N_2397,In_2655,In_1682);
and U2398 (N_2398,In_1327,In_64);
nand U2399 (N_2399,In_2242,In_144);
nor U2400 (N_2400,In_2792,In_2756);
nor U2401 (N_2401,In_1525,In_325);
nor U2402 (N_2402,In_2862,In_1933);
and U2403 (N_2403,In_2751,In_2939);
nand U2404 (N_2404,In_1624,In_1464);
nand U2405 (N_2405,In_2093,In_946);
or U2406 (N_2406,In_289,In_1789);
nor U2407 (N_2407,In_1313,In_1959);
nor U2408 (N_2408,In_1087,In_1994);
nor U2409 (N_2409,In_2935,In_356);
and U2410 (N_2410,In_1424,In_1252);
xnor U2411 (N_2411,In_1605,In_479);
nor U2412 (N_2412,In_881,In_949);
or U2413 (N_2413,In_1694,In_2612);
nor U2414 (N_2414,In_122,In_756);
nand U2415 (N_2415,In_2846,In_2292);
nor U2416 (N_2416,In_1379,In_1187);
nand U2417 (N_2417,In_242,In_1967);
and U2418 (N_2418,In_877,In_463);
and U2419 (N_2419,In_1051,In_2059);
or U2420 (N_2420,In_1840,In_2186);
xnor U2421 (N_2421,In_27,In_733);
and U2422 (N_2422,In_2430,In_2304);
or U2423 (N_2423,In_2142,In_1270);
nand U2424 (N_2424,In_2741,In_1358);
nand U2425 (N_2425,In_2501,In_1802);
xnor U2426 (N_2426,In_1849,In_2300);
or U2427 (N_2427,In_2369,In_2418);
or U2428 (N_2428,In_849,In_2571);
or U2429 (N_2429,In_1909,In_221);
nor U2430 (N_2430,In_746,In_214);
and U2431 (N_2431,In_947,In_2403);
nor U2432 (N_2432,In_2619,In_207);
nand U2433 (N_2433,In_1553,In_156);
nand U2434 (N_2434,In_1849,In_2416);
or U2435 (N_2435,In_1284,In_2313);
xor U2436 (N_2436,In_1088,In_2524);
nor U2437 (N_2437,In_905,In_1051);
and U2438 (N_2438,In_1265,In_2953);
nand U2439 (N_2439,In_2135,In_1188);
nor U2440 (N_2440,In_705,In_1435);
xnor U2441 (N_2441,In_776,In_1103);
nand U2442 (N_2442,In_235,In_1155);
nor U2443 (N_2443,In_1432,In_2549);
or U2444 (N_2444,In_441,In_2215);
nor U2445 (N_2445,In_1951,In_1712);
nand U2446 (N_2446,In_1917,In_563);
xnor U2447 (N_2447,In_2796,In_906);
and U2448 (N_2448,In_407,In_2889);
and U2449 (N_2449,In_666,In_308);
xnor U2450 (N_2450,In_266,In_1210);
or U2451 (N_2451,In_26,In_2342);
nor U2452 (N_2452,In_2137,In_2105);
or U2453 (N_2453,In_2254,In_890);
nor U2454 (N_2454,In_1294,In_2649);
nand U2455 (N_2455,In_2869,In_2824);
nor U2456 (N_2456,In_505,In_1434);
and U2457 (N_2457,In_766,In_2859);
or U2458 (N_2458,In_358,In_2699);
nand U2459 (N_2459,In_1313,In_2007);
xor U2460 (N_2460,In_1517,In_805);
nor U2461 (N_2461,In_2488,In_298);
nor U2462 (N_2462,In_2942,In_232);
nand U2463 (N_2463,In_1220,In_825);
and U2464 (N_2464,In_2697,In_833);
xor U2465 (N_2465,In_894,In_1590);
nor U2466 (N_2466,In_1664,In_1645);
and U2467 (N_2467,In_1227,In_1660);
xnor U2468 (N_2468,In_624,In_1774);
and U2469 (N_2469,In_1411,In_647);
xnor U2470 (N_2470,In_1666,In_989);
nand U2471 (N_2471,In_255,In_1246);
nand U2472 (N_2472,In_1482,In_2578);
nand U2473 (N_2473,In_1786,In_701);
nand U2474 (N_2474,In_168,In_2242);
xor U2475 (N_2475,In_1693,In_2407);
or U2476 (N_2476,In_75,In_1380);
nand U2477 (N_2477,In_104,In_1134);
or U2478 (N_2478,In_2015,In_2029);
nand U2479 (N_2479,In_2580,In_64);
and U2480 (N_2480,In_2486,In_362);
nor U2481 (N_2481,In_1259,In_458);
and U2482 (N_2482,In_936,In_1048);
nand U2483 (N_2483,In_635,In_2250);
nor U2484 (N_2484,In_2144,In_1597);
and U2485 (N_2485,In_2632,In_473);
and U2486 (N_2486,In_485,In_391);
xnor U2487 (N_2487,In_1777,In_1460);
nor U2488 (N_2488,In_2436,In_1978);
nor U2489 (N_2489,In_1313,In_2563);
or U2490 (N_2490,In_1241,In_2314);
xor U2491 (N_2491,In_557,In_2070);
nor U2492 (N_2492,In_580,In_2341);
and U2493 (N_2493,In_1994,In_2443);
nand U2494 (N_2494,In_1239,In_456);
nand U2495 (N_2495,In_1399,In_1786);
and U2496 (N_2496,In_2943,In_1696);
and U2497 (N_2497,In_1134,In_1874);
and U2498 (N_2498,In_2089,In_2406);
or U2499 (N_2499,In_1074,In_1539);
or U2500 (N_2500,In_1979,In_537);
nand U2501 (N_2501,In_1772,In_1696);
or U2502 (N_2502,In_527,In_1559);
nand U2503 (N_2503,In_2760,In_1217);
and U2504 (N_2504,In_1132,In_348);
nand U2505 (N_2505,In_2467,In_2416);
and U2506 (N_2506,In_1013,In_1572);
or U2507 (N_2507,In_2379,In_386);
nor U2508 (N_2508,In_1963,In_988);
nor U2509 (N_2509,In_39,In_1521);
and U2510 (N_2510,In_1997,In_693);
nor U2511 (N_2511,In_1846,In_583);
nor U2512 (N_2512,In_1017,In_1666);
and U2513 (N_2513,In_1362,In_772);
xnor U2514 (N_2514,In_408,In_681);
and U2515 (N_2515,In_2924,In_1895);
and U2516 (N_2516,In_2264,In_2289);
or U2517 (N_2517,In_312,In_1470);
or U2518 (N_2518,In_1079,In_36);
and U2519 (N_2519,In_1722,In_277);
nand U2520 (N_2520,In_900,In_2995);
xor U2521 (N_2521,In_1906,In_2042);
nand U2522 (N_2522,In_1991,In_1405);
xor U2523 (N_2523,In_2030,In_2282);
and U2524 (N_2524,In_255,In_1474);
and U2525 (N_2525,In_1694,In_110);
xor U2526 (N_2526,In_2174,In_2683);
and U2527 (N_2527,In_1905,In_2198);
nor U2528 (N_2528,In_1690,In_27);
and U2529 (N_2529,In_1699,In_406);
nand U2530 (N_2530,In_2625,In_693);
or U2531 (N_2531,In_465,In_2543);
nand U2532 (N_2532,In_2309,In_1998);
nor U2533 (N_2533,In_1964,In_1040);
nor U2534 (N_2534,In_2112,In_2267);
nand U2535 (N_2535,In_1578,In_755);
nor U2536 (N_2536,In_2487,In_1311);
nand U2537 (N_2537,In_2053,In_2677);
or U2538 (N_2538,In_534,In_2473);
nand U2539 (N_2539,In_2990,In_953);
or U2540 (N_2540,In_2179,In_2801);
nand U2541 (N_2541,In_2130,In_359);
nor U2542 (N_2542,In_378,In_2947);
nand U2543 (N_2543,In_730,In_197);
and U2544 (N_2544,In_2078,In_2917);
nand U2545 (N_2545,In_504,In_1841);
and U2546 (N_2546,In_1010,In_2071);
and U2547 (N_2547,In_888,In_1970);
nor U2548 (N_2548,In_1654,In_1697);
or U2549 (N_2549,In_1793,In_726);
and U2550 (N_2550,In_1036,In_416);
nand U2551 (N_2551,In_681,In_0);
nand U2552 (N_2552,In_935,In_444);
xnor U2553 (N_2553,In_674,In_333);
and U2554 (N_2554,In_2458,In_2978);
and U2555 (N_2555,In_920,In_1080);
or U2556 (N_2556,In_2590,In_321);
nor U2557 (N_2557,In_2566,In_2968);
and U2558 (N_2558,In_1815,In_2236);
xnor U2559 (N_2559,In_2605,In_2810);
xor U2560 (N_2560,In_97,In_2695);
nor U2561 (N_2561,In_2470,In_1235);
or U2562 (N_2562,In_1843,In_1050);
or U2563 (N_2563,In_2491,In_462);
and U2564 (N_2564,In_964,In_782);
and U2565 (N_2565,In_903,In_349);
or U2566 (N_2566,In_593,In_1221);
nor U2567 (N_2567,In_2272,In_1814);
nand U2568 (N_2568,In_2565,In_2414);
and U2569 (N_2569,In_287,In_1736);
nand U2570 (N_2570,In_2387,In_1287);
nor U2571 (N_2571,In_2037,In_2452);
nand U2572 (N_2572,In_712,In_1623);
or U2573 (N_2573,In_1281,In_2512);
xnor U2574 (N_2574,In_2087,In_649);
or U2575 (N_2575,In_1324,In_1315);
nand U2576 (N_2576,In_926,In_2747);
nor U2577 (N_2577,In_388,In_1443);
xnor U2578 (N_2578,In_1409,In_1955);
and U2579 (N_2579,In_281,In_1598);
or U2580 (N_2580,In_1496,In_2166);
nand U2581 (N_2581,In_1158,In_1420);
nand U2582 (N_2582,In_1238,In_2973);
nor U2583 (N_2583,In_606,In_734);
nand U2584 (N_2584,In_2600,In_1681);
nor U2585 (N_2585,In_2107,In_1455);
and U2586 (N_2586,In_2707,In_469);
nand U2587 (N_2587,In_974,In_282);
xor U2588 (N_2588,In_2184,In_1974);
nor U2589 (N_2589,In_1519,In_1579);
xor U2590 (N_2590,In_219,In_853);
nand U2591 (N_2591,In_2559,In_1292);
nor U2592 (N_2592,In_1445,In_2792);
or U2593 (N_2593,In_1366,In_2682);
and U2594 (N_2594,In_2087,In_2751);
or U2595 (N_2595,In_1361,In_277);
nand U2596 (N_2596,In_2565,In_986);
nor U2597 (N_2597,In_97,In_1175);
and U2598 (N_2598,In_2541,In_9);
or U2599 (N_2599,In_2588,In_2430);
xor U2600 (N_2600,In_2011,In_2030);
nand U2601 (N_2601,In_1539,In_2800);
and U2602 (N_2602,In_2257,In_1899);
nand U2603 (N_2603,In_313,In_205);
nor U2604 (N_2604,In_2162,In_1678);
nand U2605 (N_2605,In_1068,In_2863);
nand U2606 (N_2606,In_2598,In_377);
and U2607 (N_2607,In_806,In_406);
nand U2608 (N_2608,In_2051,In_482);
xor U2609 (N_2609,In_102,In_2759);
nor U2610 (N_2610,In_2865,In_1147);
or U2611 (N_2611,In_664,In_2411);
nor U2612 (N_2612,In_2062,In_2009);
or U2613 (N_2613,In_2538,In_194);
nand U2614 (N_2614,In_1226,In_1842);
nor U2615 (N_2615,In_502,In_2799);
or U2616 (N_2616,In_2627,In_2066);
nor U2617 (N_2617,In_2260,In_2778);
and U2618 (N_2618,In_2646,In_1558);
nand U2619 (N_2619,In_1997,In_1399);
and U2620 (N_2620,In_2319,In_2521);
and U2621 (N_2621,In_1668,In_2625);
or U2622 (N_2622,In_1529,In_2283);
and U2623 (N_2623,In_1934,In_2970);
xor U2624 (N_2624,In_930,In_148);
and U2625 (N_2625,In_2553,In_1809);
or U2626 (N_2626,In_1382,In_2173);
nor U2627 (N_2627,In_1944,In_1377);
nand U2628 (N_2628,In_211,In_2484);
nor U2629 (N_2629,In_1811,In_546);
nor U2630 (N_2630,In_1994,In_991);
nand U2631 (N_2631,In_613,In_1685);
xnor U2632 (N_2632,In_1369,In_467);
nand U2633 (N_2633,In_192,In_1617);
nand U2634 (N_2634,In_2292,In_2929);
nor U2635 (N_2635,In_2941,In_880);
nand U2636 (N_2636,In_265,In_2047);
nand U2637 (N_2637,In_271,In_1860);
nand U2638 (N_2638,In_2207,In_958);
nand U2639 (N_2639,In_2561,In_1370);
nand U2640 (N_2640,In_594,In_778);
and U2641 (N_2641,In_527,In_2265);
or U2642 (N_2642,In_2292,In_1912);
or U2643 (N_2643,In_2755,In_2058);
and U2644 (N_2644,In_2140,In_180);
and U2645 (N_2645,In_606,In_2508);
nand U2646 (N_2646,In_2846,In_1233);
nor U2647 (N_2647,In_2915,In_814);
or U2648 (N_2648,In_2429,In_1190);
and U2649 (N_2649,In_240,In_42);
nor U2650 (N_2650,In_2473,In_823);
xor U2651 (N_2651,In_1674,In_2691);
and U2652 (N_2652,In_2919,In_2365);
nand U2653 (N_2653,In_90,In_2158);
or U2654 (N_2654,In_331,In_1659);
nand U2655 (N_2655,In_2238,In_8);
nand U2656 (N_2656,In_387,In_1761);
or U2657 (N_2657,In_521,In_2981);
xnor U2658 (N_2658,In_462,In_2512);
and U2659 (N_2659,In_1667,In_1805);
nor U2660 (N_2660,In_1458,In_1370);
or U2661 (N_2661,In_74,In_466);
or U2662 (N_2662,In_1720,In_208);
or U2663 (N_2663,In_51,In_498);
or U2664 (N_2664,In_2431,In_2047);
xor U2665 (N_2665,In_623,In_1614);
nand U2666 (N_2666,In_1080,In_1567);
xor U2667 (N_2667,In_905,In_942);
nor U2668 (N_2668,In_975,In_2291);
or U2669 (N_2669,In_482,In_2524);
nor U2670 (N_2670,In_1990,In_2417);
or U2671 (N_2671,In_527,In_697);
or U2672 (N_2672,In_619,In_1067);
or U2673 (N_2673,In_2722,In_742);
and U2674 (N_2674,In_2683,In_403);
nand U2675 (N_2675,In_393,In_2221);
xnor U2676 (N_2676,In_2870,In_2680);
and U2677 (N_2677,In_26,In_333);
nand U2678 (N_2678,In_1174,In_309);
and U2679 (N_2679,In_61,In_2112);
nor U2680 (N_2680,In_1532,In_466);
nand U2681 (N_2681,In_1783,In_1541);
nand U2682 (N_2682,In_1018,In_973);
nor U2683 (N_2683,In_58,In_1465);
nor U2684 (N_2684,In_17,In_1481);
or U2685 (N_2685,In_1355,In_810);
and U2686 (N_2686,In_2623,In_2480);
nor U2687 (N_2687,In_1701,In_2634);
nand U2688 (N_2688,In_2385,In_1381);
nor U2689 (N_2689,In_1369,In_2796);
and U2690 (N_2690,In_77,In_2674);
or U2691 (N_2691,In_2698,In_2167);
nand U2692 (N_2692,In_124,In_256);
and U2693 (N_2693,In_1693,In_806);
xnor U2694 (N_2694,In_1252,In_437);
and U2695 (N_2695,In_1800,In_588);
and U2696 (N_2696,In_1842,In_2506);
and U2697 (N_2697,In_1669,In_315);
and U2698 (N_2698,In_2495,In_721);
nor U2699 (N_2699,In_2326,In_1084);
or U2700 (N_2700,In_2111,In_2086);
nand U2701 (N_2701,In_1580,In_1425);
nand U2702 (N_2702,In_2721,In_2663);
nand U2703 (N_2703,In_1914,In_503);
and U2704 (N_2704,In_534,In_2917);
xor U2705 (N_2705,In_2291,In_1498);
and U2706 (N_2706,In_469,In_622);
xnor U2707 (N_2707,In_2831,In_329);
or U2708 (N_2708,In_68,In_864);
and U2709 (N_2709,In_1880,In_1001);
or U2710 (N_2710,In_2608,In_1917);
xnor U2711 (N_2711,In_2198,In_2623);
or U2712 (N_2712,In_538,In_1289);
nor U2713 (N_2713,In_539,In_2583);
nand U2714 (N_2714,In_176,In_417);
nor U2715 (N_2715,In_1398,In_1601);
or U2716 (N_2716,In_1173,In_2769);
nand U2717 (N_2717,In_2367,In_1796);
nor U2718 (N_2718,In_54,In_873);
or U2719 (N_2719,In_2078,In_483);
nor U2720 (N_2720,In_1292,In_1022);
or U2721 (N_2721,In_2065,In_802);
and U2722 (N_2722,In_2442,In_2695);
and U2723 (N_2723,In_180,In_729);
nand U2724 (N_2724,In_1204,In_2903);
nor U2725 (N_2725,In_2298,In_551);
or U2726 (N_2726,In_2818,In_1497);
and U2727 (N_2727,In_1343,In_1980);
or U2728 (N_2728,In_1173,In_2002);
nor U2729 (N_2729,In_2365,In_1332);
or U2730 (N_2730,In_735,In_2913);
or U2731 (N_2731,In_2069,In_808);
or U2732 (N_2732,In_2376,In_66);
and U2733 (N_2733,In_2303,In_2147);
nor U2734 (N_2734,In_2913,In_1558);
nor U2735 (N_2735,In_483,In_1613);
nor U2736 (N_2736,In_1025,In_2689);
nand U2737 (N_2737,In_1570,In_1021);
nor U2738 (N_2738,In_946,In_933);
and U2739 (N_2739,In_1341,In_2321);
or U2740 (N_2740,In_1059,In_2438);
and U2741 (N_2741,In_2167,In_1307);
and U2742 (N_2742,In_2604,In_2083);
or U2743 (N_2743,In_1250,In_2573);
nand U2744 (N_2744,In_1603,In_2914);
nand U2745 (N_2745,In_1334,In_340);
and U2746 (N_2746,In_445,In_2089);
nand U2747 (N_2747,In_1053,In_1076);
nor U2748 (N_2748,In_1693,In_2760);
nand U2749 (N_2749,In_424,In_2879);
xor U2750 (N_2750,In_2297,In_1186);
nand U2751 (N_2751,In_1928,In_629);
nand U2752 (N_2752,In_2779,In_2858);
or U2753 (N_2753,In_1102,In_21);
nand U2754 (N_2754,In_666,In_683);
nand U2755 (N_2755,In_1205,In_298);
or U2756 (N_2756,In_2720,In_1892);
nor U2757 (N_2757,In_1379,In_341);
or U2758 (N_2758,In_2609,In_2447);
and U2759 (N_2759,In_1895,In_2299);
and U2760 (N_2760,In_1133,In_354);
nor U2761 (N_2761,In_2759,In_1041);
and U2762 (N_2762,In_368,In_1340);
xor U2763 (N_2763,In_1340,In_861);
xor U2764 (N_2764,In_1679,In_2869);
nand U2765 (N_2765,In_1318,In_1979);
or U2766 (N_2766,In_119,In_2750);
nor U2767 (N_2767,In_2575,In_2185);
or U2768 (N_2768,In_1059,In_2423);
nand U2769 (N_2769,In_2648,In_116);
nand U2770 (N_2770,In_1543,In_195);
or U2771 (N_2771,In_1051,In_2062);
and U2772 (N_2772,In_1913,In_578);
and U2773 (N_2773,In_2481,In_58);
nor U2774 (N_2774,In_695,In_737);
nor U2775 (N_2775,In_979,In_537);
nand U2776 (N_2776,In_410,In_2735);
or U2777 (N_2777,In_954,In_2100);
and U2778 (N_2778,In_1998,In_1352);
or U2779 (N_2779,In_2847,In_178);
nand U2780 (N_2780,In_2120,In_2796);
nor U2781 (N_2781,In_936,In_686);
nor U2782 (N_2782,In_730,In_2871);
and U2783 (N_2783,In_625,In_2203);
or U2784 (N_2784,In_1206,In_2901);
or U2785 (N_2785,In_1517,In_440);
nor U2786 (N_2786,In_132,In_516);
or U2787 (N_2787,In_867,In_2257);
nand U2788 (N_2788,In_1400,In_1260);
or U2789 (N_2789,In_795,In_598);
nor U2790 (N_2790,In_615,In_2482);
or U2791 (N_2791,In_2025,In_2408);
or U2792 (N_2792,In_219,In_1176);
nand U2793 (N_2793,In_1547,In_2566);
or U2794 (N_2794,In_1574,In_320);
nand U2795 (N_2795,In_673,In_96);
or U2796 (N_2796,In_1757,In_2137);
and U2797 (N_2797,In_1683,In_498);
xnor U2798 (N_2798,In_1273,In_2472);
nor U2799 (N_2799,In_2748,In_1156);
nor U2800 (N_2800,In_2110,In_1090);
nor U2801 (N_2801,In_2464,In_2314);
nand U2802 (N_2802,In_2770,In_2614);
nand U2803 (N_2803,In_513,In_2941);
nand U2804 (N_2804,In_1807,In_1815);
or U2805 (N_2805,In_2979,In_1533);
or U2806 (N_2806,In_280,In_1376);
xnor U2807 (N_2807,In_896,In_1923);
or U2808 (N_2808,In_2332,In_1937);
and U2809 (N_2809,In_2062,In_1976);
nor U2810 (N_2810,In_112,In_1394);
nor U2811 (N_2811,In_607,In_2813);
and U2812 (N_2812,In_1752,In_1570);
nand U2813 (N_2813,In_68,In_1917);
or U2814 (N_2814,In_2074,In_310);
and U2815 (N_2815,In_905,In_2477);
nand U2816 (N_2816,In_2512,In_2774);
nor U2817 (N_2817,In_434,In_2696);
nand U2818 (N_2818,In_2873,In_1933);
or U2819 (N_2819,In_2537,In_2913);
or U2820 (N_2820,In_975,In_1861);
and U2821 (N_2821,In_872,In_1228);
and U2822 (N_2822,In_1936,In_556);
and U2823 (N_2823,In_2791,In_2573);
nor U2824 (N_2824,In_1388,In_59);
nor U2825 (N_2825,In_691,In_975);
or U2826 (N_2826,In_2128,In_1326);
nor U2827 (N_2827,In_1950,In_1483);
nor U2828 (N_2828,In_1129,In_2172);
and U2829 (N_2829,In_1984,In_1448);
nand U2830 (N_2830,In_2847,In_983);
or U2831 (N_2831,In_2143,In_1004);
and U2832 (N_2832,In_1089,In_1150);
nor U2833 (N_2833,In_2069,In_981);
nor U2834 (N_2834,In_1067,In_2457);
nor U2835 (N_2835,In_745,In_1240);
and U2836 (N_2836,In_672,In_1315);
nand U2837 (N_2837,In_2062,In_1878);
or U2838 (N_2838,In_758,In_570);
and U2839 (N_2839,In_573,In_162);
nand U2840 (N_2840,In_1903,In_2367);
or U2841 (N_2841,In_400,In_741);
or U2842 (N_2842,In_1836,In_2054);
nor U2843 (N_2843,In_1558,In_2503);
and U2844 (N_2844,In_1620,In_1029);
nor U2845 (N_2845,In_2653,In_2918);
nor U2846 (N_2846,In_851,In_2836);
nor U2847 (N_2847,In_2601,In_423);
nand U2848 (N_2848,In_201,In_90);
and U2849 (N_2849,In_491,In_69);
or U2850 (N_2850,In_2690,In_2033);
xor U2851 (N_2851,In_442,In_1813);
or U2852 (N_2852,In_424,In_1814);
or U2853 (N_2853,In_821,In_1410);
nor U2854 (N_2854,In_1407,In_2451);
nor U2855 (N_2855,In_808,In_2254);
or U2856 (N_2856,In_1627,In_2221);
or U2857 (N_2857,In_1820,In_423);
nand U2858 (N_2858,In_821,In_1631);
xor U2859 (N_2859,In_2787,In_768);
or U2860 (N_2860,In_2423,In_737);
or U2861 (N_2861,In_2282,In_2496);
and U2862 (N_2862,In_1678,In_1827);
nor U2863 (N_2863,In_1120,In_634);
and U2864 (N_2864,In_32,In_2870);
nor U2865 (N_2865,In_2225,In_2027);
nor U2866 (N_2866,In_1732,In_1921);
and U2867 (N_2867,In_1123,In_372);
xnor U2868 (N_2868,In_265,In_1982);
and U2869 (N_2869,In_1641,In_946);
nand U2870 (N_2870,In_2486,In_2436);
xnor U2871 (N_2871,In_1714,In_1863);
nor U2872 (N_2872,In_2479,In_2453);
and U2873 (N_2873,In_1724,In_2454);
or U2874 (N_2874,In_393,In_761);
nor U2875 (N_2875,In_303,In_1417);
and U2876 (N_2876,In_430,In_1107);
and U2877 (N_2877,In_1700,In_862);
nor U2878 (N_2878,In_846,In_269);
nand U2879 (N_2879,In_2387,In_32);
nand U2880 (N_2880,In_2305,In_251);
and U2881 (N_2881,In_2896,In_230);
nand U2882 (N_2882,In_361,In_920);
or U2883 (N_2883,In_1527,In_291);
and U2884 (N_2884,In_1636,In_1527);
and U2885 (N_2885,In_155,In_1535);
nor U2886 (N_2886,In_106,In_2547);
nand U2887 (N_2887,In_1618,In_984);
or U2888 (N_2888,In_237,In_2328);
xor U2889 (N_2889,In_2752,In_1746);
nor U2890 (N_2890,In_356,In_601);
and U2891 (N_2891,In_227,In_833);
and U2892 (N_2892,In_713,In_471);
and U2893 (N_2893,In_364,In_2588);
xnor U2894 (N_2894,In_431,In_2776);
and U2895 (N_2895,In_1263,In_186);
nor U2896 (N_2896,In_2542,In_2518);
and U2897 (N_2897,In_128,In_2050);
nor U2898 (N_2898,In_322,In_2901);
nor U2899 (N_2899,In_1355,In_1675);
nand U2900 (N_2900,In_992,In_578);
or U2901 (N_2901,In_2258,In_1448);
and U2902 (N_2902,In_1356,In_974);
xor U2903 (N_2903,In_1976,In_2808);
nor U2904 (N_2904,In_1271,In_2370);
nor U2905 (N_2905,In_537,In_2315);
or U2906 (N_2906,In_2633,In_1096);
nor U2907 (N_2907,In_2821,In_113);
and U2908 (N_2908,In_1291,In_1659);
nor U2909 (N_2909,In_904,In_284);
and U2910 (N_2910,In_1995,In_932);
and U2911 (N_2911,In_139,In_160);
nand U2912 (N_2912,In_2118,In_2600);
nand U2913 (N_2913,In_1509,In_2122);
and U2914 (N_2914,In_534,In_2022);
and U2915 (N_2915,In_2724,In_189);
xor U2916 (N_2916,In_2214,In_2867);
xor U2917 (N_2917,In_793,In_1214);
nor U2918 (N_2918,In_2553,In_407);
and U2919 (N_2919,In_786,In_790);
nor U2920 (N_2920,In_1128,In_520);
and U2921 (N_2921,In_1422,In_210);
nand U2922 (N_2922,In_2267,In_2303);
and U2923 (N_2923,In_2126,In_979);
nand U2924 (N_2924,In_2376,In_724);
and U2925 (N_2925,In_2052,In_1664);
or U2926 (N_2926,In_567,In_997);
nor U2927 (N_2927,In_659,In_2062);
xnor U2928 (N_2928,In_1131,In_2416);
nor U2929 (N_2929,In_1925,In_879);
or U2930 (N_2930,In_2652,In_1153);
xor U2931 (N_2931,In_529,In_280);
or U2932 (N_2932,In_1940,In_287);
and U2933 (N_2933,In_2567,In_107);
and U2934 (N_2934,In_1016,In_1534);
and U2935 (N_2935,In_2568,In_604);
nand U2936 (N_2936,In_2608,In_1063);
nor U2937 (N_2937,In_1081,In_1789);
xnor U2938 (N_2938,In_1615,In_2145);
and U2939 (N_2939,In_1347,In_2372);
nor U2940 (N_2940,In_1906,In_2386);
xnor U2941 (N_2941,In_2484,In_864);
and U2942 (N_2942,In_436,In_321);
and U2943 (N_2943,In_216,In_717);
and U2944 (N_2944,In_2720,In_1723);
nand U2945 (N_2945,In_2103,In_614);
or U2946 (N_2946,In_367,In_2775);
and U2947 (N_2947,In_201,In_1654);
nor U2948 (N_2948,In_1989,In_2473);
and U2949 (N_2949,In_2986,In_1598);
nand U2950 (N_2950,In_2795,In_1650);
or U2951 (N_2951,In_515,In_146);
xnor U2952 (N_2952,In_2336,In_2212);
and U2953 (N_2953,In_2363,In_2959);
nor U2954 (N_2954,In_40,In_1347);
nand U2955 (N_2955,In_2507,In_1651);
and U2956 (N_2956,In_13,In_2667);
and U2957 (N_2957,In_2525,In_1002);
xor U2958 (N_2958,In_1085,In_311);
and U2959 (N_2959,In_1635,In_1923);
nand U2960 (N_2960,In_2828,In_2401);
and U2961 (N_2961,In_1801,In_2472);
xnor U2962 (N_2962,In_2241,In_2526);
and U2963 (N_2963,In_1377,In_1724);
nand U2964 (N_2964,In_2450,In_1602);
and U2965 (N_2965,In_361,In_1760);
or U2966 (N_2966,In_1804,In_852);
nor U2967 (N_2967,In_2672,In_951);
nand U2968 (N_2968,In_1551,In_1653);
nand U2969 (N_2969,In_1365,In_2814);
nor U2970 (N_2970,In_1609,In_1154);
nand U2971 (N_2971,In_1810,In_2732);
or U2972 (N_2972,In_2826,In_1094);
nand U2973 (N_2973,In_1293,In_734);
or U2974 (N_2974,In_2738,In_801);
nor U2975 (N_2975,In_1186,In_2616);
xnor U2976 (N_2976,In_84,In_22);
nand U2977 (N_2977,In_2825,In_2617);
nor U2978 (N_2978,In_2188,In_830);
xnor U2979 (N_2979,In_288,In_1988);
nand U2980 (N_2980,In_937,In_2553);
nor U2981 (N_2981,In_1312,In_1502);
nand U2982 (N_2982,In_2151,In_1432);
nand U2983 (N_2983,In_2236,In_1309);
or U2984 (N_2984,In_72,In_585);
and U2985 (N_2985,In_2282,In_2036);
nand U2986 (N_2986,In_2545,In_1427);
or U2987 (N_2987,In_2428,In_1594);
or U2988 (N_2988,In_2675,In_2831);
and U2989 (N_2989,In_583,In_162);
or U2990 (N_2990,In_893,In_340);
or U2991 (N_2991,In_1502,In_1906);
nor U2992 (N_2992,In_1798,In_2869);
or U2993 (N_2993,In_833,In_18);
xor U2994 (N_2994,In_2091,In_247);
nand U2995 (N_2995,In_2239,In_2817);
and U2996 (N_2996,In_92,In_24);
nor U2997 (N_2997,In_282,In_2424);
nor U2998 (N_2998,In_2996,In_156);
nor U2999 (N_2999,In_1378,In_455);
and U3000 (N_3000,In_164,In_2023);
nand U3001 (N_3001,In_386,In_140);
or U3002 (N_3002,In_894,In_1338);
nand U3003 (N_3003,In_2621,In_154);
nand U3004 (N_3004,In_1378,In_1368);
and U3005 (N_3005,In_2676,In_2684);
and U3006 (N_3006,In_1884,In_157);
nor U3007 (N_3007,In_2096,In_2158);
or U3008 (N_3008,In_1298,In_928);
xnor U3009 (N_3009,In_1807,In_2785);
nand U3010 (N_3010,In_1895,In_682);
nor U3011 (N_3011,In_190,In_536);
or U3012 (N_3012,In_628,In_2162);
and U3013 (N_3013,In_896,In_1677);
or U3014 (N_3014,In_173,In_2888);
nand U3015 (N_3015,In_2226,In_273);
and U3016 (N_3016,In_2061,In_1467);
nand U3017 (N_3017,In_685,In_1467);
nand U3018 (N_3018,In_930,In_657);
and U3019 (N_3019,In_1537,In_1944);
and U3020 (N_3020,In_746,In_591);
nor U3021 (N_3021,In_2507,In_682);
nor U3022 (N_3022,In_2918,In_1233);
nand U3023 (N_3023,In_121,In_728);
nand U3024 (N_3024,In_809,In_349);
nand U3025 (N_3025,In_2170,In_2686);
nand U3026 (N_3026,In_1765,In_2181);
nor U3027 (N_3027,In_287,In_793);
or U3028 (N_3028,In_2296,In_2605);
or U3029 (N_3029,In_2781,In_785);
or U3030 (N_3030,In_2760,In_1204);
and U3031 (N_3031,In_1395,In_210);
nor U3032 (N_3032,In_1818,In_1043);
nand U3033 (N_3033,In_1072,In_873);
nor U3034 (N_3034,In_86,In_1707);
and U3035 (N_3035,In_2599,In_2092);
nand U3036 (N_3036,In_2685,In_1434);
nand U3037 (N_3037,In_2152,In_1191);
and U3038 (N_3038,In_471,In_2884);
nor U3039 (N_3039,In_902,In_1232);
or U3040 (N_3040,In_1292,In_926);
and U3041 (N_3041,In_64,In_637);
nor U3042 (N_3042,In_2129,In_2152);
nor U3043 (N_3043,In_338,In_2081);
nand U3044 (N_3044,In_1550,In_1195);
and U3045 (N_3045,In_2594,In_2075);
nor U3046 (N_3046,In_2057,In_1291);
nand U3047 (N_3047,In_1299,In_2001);
and U3048 (N_3048,In_217,In_1931);
nor U3049 (N_3049,In_864,In_127);
nor U3050 (N_3050,In_1519,In_1552);
xor U3051 (N_3051,In_739,In_2440);
nand U3052 (N_3052,In_1958,In_1748);
and U3053 (N_3053,In_722,In_597);
or U3054 (N_3054,In_1257,In_2849);
xor U3055 (N_3055,In_201,In_650);
nand U3056 (N_3056,In_1113,In_548);
and U3057 (N_3057,In_638,In_1200);
or U3058 (N_3058,In_2984,In_420);
nand U3059 (N_3059,In_1179,In_2887);
and U3060 (N_3060,In_2925,In_2128);
and U3061 (N_3061,In_1933,In_896);
and U3062 (N_3062,In_1496,In_2590);
xnor U3063 (N_3063,In_1433,In_2412);
or U3064 (N_3064,In_2217,In_837);
or U3065 (N_3065,In_2240,In_1131);
and U3066 (N_3066,In_92,In_2331);
nor U3067 (N_3067,In_2888,In_604);
nor U3068 (N_3068,In_216,In_922);
xnor U3069 (N_3069,In_633,In_899);
or U3070 (N_3070,In_2219,In_468);
and U3071 (N_3071,In_514,In_2861);
and U3072 (N_3072,In_907,In_1390);
or U3073 (N_3073,In_2895,In_2273);
nand U3074 (N_3074,In_440,In_2653);
or U3075 (N_3075,In_967,In_743);
nor U3076 (N_3076,In_760,In_2289);
and U3077 (N_3077,In_761,In_1679);
and U3078 (N_3078,In_1196,In_1241);
xor U3079 (N_3079,In_1584,In_280);
and U3080 (N_3080,In_765,In_64);
xor U3081 (N_3081,In_1754,In_2789);
nand U3082 (N_3082,In_1720,In_969);
and U3083 (N_3083,In_411,In_1375);
nor U3084 (N_3084,In_2091,In_1898);
nor U3085 (N_3085,In_1873,In_19);
or U3086 (N_3086,In_394,In_692);
and U3087 (N_3087,In_349,In_570);
nor U3088 (N_3088,In_2787,In_1026);
and U3089 (N_3089,In_2209,In_620);
nand U3090 (N_3090,In_427,In_1059);
nor U3091 (N_3091,In_2081,In_2656);
or U3092 (N_3092,In_2793,In_103);
and U3093 (N_3093,In_1393,In_1004);
xnor U3094 (N_3094,In_2411,In_1567);
nor U3095 (N_3095,In_2999,In_453);
nand U3096 (N_3096,In_728,In_2380);
and U3097 (N_3097,In_2193,In_2327);
xor U3098 (N_3098,In_415,In_1740);
and U3099 (N_3099,In_743,In_1532);
nand U3100 (N_3100,In_2180,In_1121);
and U3101 (N_3101,In_2858,In_1232);
nor U3102 (N_3102,In_2824,In_2008);
xor U3103 (N_3103,In_1282,In_476);
nand U3104 (N_3104,In_2138,In_1452);
or U3105 (N_3105,In_2985,In_1917);
or U3106 (N_3106,In_1093,In_1277);
or U3107 (N_3107,In_1171,In_2196);
nand U3108 (N_3108,In_1944,In_2737);
and U3109 (N_3109,In_1379,In_398);
or U3110 (N_3110,In_1558,In_1973);
xnor U3111 (N_3111,In_1936,In_1285);
or U3112 (N_3112,In_2171,In_1187);
nand U3113 (N_3113,In_352,In_1673);
nor U3114 (N_3114,In_720,In_2976);
and U3115 (N_3115,In_657,In_979);
and U3116 (N_3116,In_1844,In_2440);
and U3117 (N_3117,In_1903,In_453);
or U3118 (N_3118,In_1323,In_1584);
nor U3119 (N_3119,In_1443,In_343);
and U3120 (N_3120,In_471,In_197);
and U3121 (N_3121,In_199,In_1851);
xnor U3122 (N_3122,In_2345,In_2930);
nand U3123 (N_3123,In_1181,In_646);
and U3124 (N_3124,In_1293,In_1807);
nor U3125 (N_3125,In_1907,In_1299);
nand U3126 (N_3126,In_506,In_607);
or U3127 (N_3127,In_387,In_49);
nor U3128 (N_3128,In_247,In_922);
or U3129 (N_3129,In_810,In_1153);
and U3130 (N_3130,In_150,In_2307);
nor U3131 (N_3131,In_56,In_876);
xnor U3132 (N_3132,In_2186,In_1772);
nand U3133 (N_3133,In_785,In_885);
nor U3134 (N_3134,In_1805,In_1185);
nor U3135 (N_3135,In_1548,In_2037);
or U3136 (N_3136,In_1715,In_2115);
nor U3137 (N_3137,In_1406,In_1901);
and U3138 (N_3138,In_306,In_2947);
nor U3139 (N_3139,In_2909,In_814);
or U3140 (N_3140,In_1436,In_1712);
or U3141 (N_3141,In_58,In_947);
or U3142 (N_3142,In_366,In_2574);
nor U3143 (N_3143,In_1302,In_1413);
or U3144 (N_3144,In_832,In_2732);
nor U3145 (N_3145,In_2874,In_1576);
or U3146 (N_3146,In_1698,In_1302);
nor U3147 (N_3147,In_567,In_1156);
and U3148 (N_3148,In_1788,In_204);
nand U3149 (N_3149,In_2518,In_2828);
nor U3150 (N_3150,In_2827,In_2308);
nand U3151 (N_3151,In_1290,In_2984);
xnor U3152 (N_3152,In_1460,In_2529);
xor U3153 (N_3153,In_1617,In_699);
nor U3154 (N_3154,In_2790,In_1104);
and U3155 (N_3155,In_679,In_2704);
or U3156 (N_3156,In_669,In_129);
nand U3157 (N_3157,In_1172,In_1029);
and U3158 (N_3158,In_851,In_2327);
and U3159 (N_3159,In_1772,In_1149);
nor U3160 (N_3160,In_982,In_2676);
nand U3161 (N_3161,In_2693,In_198);
and U3162 (N_3162,In_2605,In_938);
and U3163 (N_3163,In_2309,In_349);
or U3164 (N_3164,In_1564,In_2713);
and U3165 (N_3165,In_926,In_2714);
nor U3166 (N_3166,In_555,In_47);
nand U3167 (N_3167,In_1346,In_96);
nand U3168 (N_3168,In_2335,In_841);
or U3169 (N_3169,In_409,In_2528);
and U3170 (N_3170,In_210,In_2791);
nor U3171 (N_3171,In_1799,In_2059);
nand U3172 (N_3172,In_1383,In_1788);
or U3173 (N_3173,In_2467,In_1448);
xor U3174 (N_3174,In_6,In_300);
xor U3175 (N_3175,In_1133,In_1912);
or U3176 (N_3176,In_2105,In_2648);
nand U3177 (N_3177,In_598,In_1970);
nor U3178 (N_3178,In_763,In_936);
xor U3179 (N_3179,In_1357,In_2619);
nand U3180 (N_3180,In_2211,In_262);
nand U3181 (N_3181,In_1911,In_2742);
or U3182 (N_3182,In_1193,In_1600);
nand U3183 (N_3183,In_1085,In_2378);
nand U3184 (N_3184,In_2145,In_249);
nor U3185 (N_3185,In_1611,In_2769);
nor U3186 (N_3186,In_2941,In_2965);
nand U3187 (N_3187,In_1677,In_44);
xor U3188 (N_3188,In_1065,In_1206);
nand U3189 (N_3189,In_2503,In_2350);
or U3190 (N_3190,In_2023,In_656);
or U3191 (N_3191,In_668,In_1351);
or U3192 (N_3192,In_1692,In_958);
and U3193 (N_3193,In_2217,In_757);
and U3194 (N_3194,In_1349,In_2597);
nand U3195 (N_3195,In_1814,In_2013);
nand U3196 (N_3196,In_1912,In_1766);
or U3197 (N_3197,In_1361,In_393);
nand U3198 (N_3198,In_1597,In_2076);
nand U3199 (N_3199,In_2043,In_1388);
and U3200 (N_3200,In_880,In_193);
nor U3201 (N_3201,In_845,In_336);
or U3202 (N_3202,In_859,In_2527);
nand U3203 (N_3203,In_139,In_731);
nor U3204 (N_3204,In_1390,In_2428);
nand U3205 (N_3205,In_1136,In_2758);
or U3206 (N_3206,In_1596,In_2094);
nor U3207 (N_3207,In_1976,In_1581);
xor U3208 (N_3208,In_790,In_1244);
nand U3209 (N_3209,In_142,In_1718);
or U3210 (N_3210,In_544,In_2071);
or U3211 (N_3211,In_247,In_1288);
nand U3212 (N_3212,In_2658,In_1050);
and U3213 (N_3213,In_1824,In_1825);
and U3214 (N_3214,In_2688,In_2634);
nand U3215 (N_3215,In_2666,In_2436);
nor U3216 (N_3216,In_1146,In_779);
and U3217 (N_3217,In_2546,In_2718);
and U3218 (N_3218,In_49,In_1773);
nand U3219 (N_3219,In_2164,In_2805);
nand U3220 (N_3220,In_2228,In_1692);
or U3221 (N_3221,In_1694,In_2149);
nand U3222 (N_3222,In_1058,In_1928);
or U3223 (N_3223,In_326,In_2117);
xor U3224 (N_3224,In_1912,In_334);
nand U3225 (N_3225,In_1807,In_245);
nand U3226 (N_3226,In_1770,In_771);
nand U3227 (N_3227,In_644,In_2212);
nor U3228 (N_3228,In_1889,In_770);
and U3229 (N_3229,In_2637,In_1405);
nand U3230 (N_3230,In_1806,In_2811);
nor U3231 (N_3231,In_2619,In_906);
nand U3232 (N_3232,In_2925,In_1039);
and U3233 (N_3233,In_890,In_1021);
nand U3234 (N_3234,In_1627,In_2324);
nand U3235 (N_3235,In_1617,In_1630);
xor U3236 (N_3236,In_991,In_2881);
nor U3237 (N_3237,In_763,In_2795);
xnor U3238 (N_3238,In_2710,In_890);
or U3239 (N_3239,In_763,In_2324);
nor U3240 (N_3240,In_869,In_804);
nor U3241 (N_3241,In_2744,In_2570);
nand U3242 (N_3242,In_1735,In_2939);
and U3243 (N_3243,In_2702,In_2097);
and U3244 (N_3244,In_2393,In_2976);
or U3245 (N_3245,In_1009,In_1200);
nor U3246 (N_3246,In_1429,In_1);
or U3247 (N_3247,In_2146,In_2026);
or U3248 (N_3248,In_153,In_1525);
nand U3249 (N_3249,In_1071,In_906);
nand U3250 (N_3250,In_353,In_639);
and U3251 (N_3251,In_415,In_2335);
and U3252 (N_3252,In_2963,In_1917);
xor U3253 (N_3253,In_2128,In_746);
nand U3254 (N_3254,In_934,In_2674);
nand U3255 (N_3255,In_2059,In_2711);
or U3256 (N_3256,In_2481,In_2100);
nor U3257 (N_3257,In_657,In_1249);
nor U3258 (N_3258,In_2765,In_1108);
nand U3259 (N_3259,In_779,In_1288);
nand U3260 (N_3260,In_1452,In_1728);
and U3261 (N_3261,In_886,In_1428);
and U3262 (N_3262,In_1646,In_2754);
nand U3263 (N_3263,In_168,In_2939);
xnor U3264 (N_3264,In_2468,In_868);
nand U3265 (N_3265,In_1857,In_1727);
nor U3266 (N_3266,In_19,In_2462);
nand U3267 (N_3267,In_637,In_820);
nand U3268 (N_3268,In_2839,In_2904);
nor U3269 (N_3269,In_1656,In_2622);
and U3270 (N_3270,In_621,In_480);
or U3271 (N_3271,In_948,In_406);
nand U3272 (N_3272,In_2581,In_1128);
nand U3273 (N_3273,In_397,In_2733);
and U3274 (N_3274,In_1999,In_324);
xnor U3275 (N_3275,In_2658,In_2972);
nand U3276 (N_3276,In_1697,In_2049);
nor U3277 (N_3277,In_2235,In_178);
xnor U3278 (N_3278,In_1543,In_4);
and U3279 (N_3279,In_92,In_2657);
xnor U3280 (N_3280,In_1516,In_529);
and U3281 (N_3281,In_1950,In_2495);
or U3282 (N_3282,In_2467,In_1817);
nor U3283 (N_3283,In_1082,In_146);
xnor U3284 (N_3284,In_1099,In_1429);
nor U3285 (N_3285,In_1572,In_2349);
and U3286 (N_3286,In_202,In_2675);
and U3287 (N_3287,In_2507,In_672);
nand U3288 (N_3288,In_2342,In_1058);
xnor U3289 (N_3289,In_436,In_2669);
and U3290 (N_3290,In_2453,In_1604);
xnor U3291 (N_3291,In_2202,In_2847);
nor U3292 (N_3292,In_700,In_733);
nor U3293 (N_3293,In_1631,In_2307);
or U3294 (N_3294,In_2875,In_702);
nor U3295 (N_3295,In_1993,In_168);
or U3296 (N_3296,In_1371,In_160);
or U3297 (N_3297,In_1444,In_1357);
nor U3298 (N_3298,In_1495,In_1596);
nand U3299 (N_3299,In_1402,In_159);
or U3300 (N_3300,In_1908,In_955);
nand U3301 (N_3301,In_823,In_35);
nor U3302 (N_3302,In_245,In_2124);
and U3303 (N_3303,In_1509,In_1261);
nor U3304 (N_3304,In_2475,In_1626);
nor U3305 (N_3305,In_2724,In_176);
and U3306 (N_3306,In_1027,In_2172);
nor U3307 (N_3307,In_145,In_1879);
xor U3308 (N_3308,In_2963,In_2123);
nor U3309 (N_3309,In_200,In_194);
or U3310 (N_3310,In_1685,In_463);
nand U3311 (N_3311,In_1645,In_1684);
nand U3312 (N_3312,In_677,In_2726);
or U3313 (N_3313,In_2012,In_2439);
nand U3314 (N_3314,In_2117,In_2492);
or U3315 (N_3315,In_2984,In_1569);
nand U3316 (N_3316,In_825,In_879);
nor U3317 (N_3317,In_501,In_420);
and U3318 (N_3318,In_2887,In_70);
and U3319 (N_3319,In_930,In_2450);
nand U3320 (N_3320,In_2796,In_2933);
nand U3321 (N_3321,In_119,In_943);
and U3322 (N_3322,In_2122,In_518);
nand U3323 (N_3323,In_2013,In_1703);
and U3324 (N_3324,In_296,In_1763);
xor U3325 (N_3325,In_936,In_1589);
and U3326 (N_3326,In_1824,In_387);
nand U3327 (N_3327,In_52,In_178);
or U3328 (N_3328,In_537,In_2008);
nand U3329 (N_3329,In_1255,In_2160);
and U3330 (N_3330,In_2040,In_2495);
or U3331 (N_3331,In_2572,In_2058);
nor U3332 (N_3332,In_114,In_769);
and U3333 (N_3333,In_1243,In_2620);
xor U3334 (N_3334,In_2790,In_36);
nand U3335 (N_3335,In_2392,In_349);
or U3336 (N_3336,In_2652,In_2514);
nor U3337 (N_3337,In_539,In_2212);
nand U3338 (N_3338,In_2478,In_1633);
xnor U3339 (N_3339,In_1249,In_967);
nand U3340 (N_3340,In_2504,In_2787);
nand U3341 (N_3341,In_2989,In_879);
xnor U3342 (N_3342,In_2576,In_2257);
nor U3343 (N_3343,In_905,In_49);
or U3344 (N_3344,In_120,In_1710);
nor U3345 (N_3345,In_191,In_2919);
nor U3346 (N_3346,In_1615,In_2404);
or U3347 (N_3347,In_2657,In_1388);
nor U3348 (N_3348,In_674,In_959);
nor U3349 (N_3349,In_1244,In_730);
nor U3350 (N_3350,In_2528,In_820);
and U3351 (N_3351,In_1677,In_1047);
nand U3352 (N_3352,In_315,In_2401);
or U3353 (N_3353,In_2731,In_727);
or U3354 (N_3354,In_2228,In_927);
and U3355 (N_3355,In_101,In_1454);
xor U3356 (N_3356,In_2872,In_1889);
xor U3357 (N_3357,In_605,In_504);
or U3358 (N_3358,In_2770,In_1161);
nand U3359 (N_3359,In_2038,In_2990);
nand U3360 (N_3360,In_2063,In_1099);
and U3361 (N_3361,In_840,In_1118);
or U3362 (N_3362,In_1366,In_1598);
and U3363 (N_3363,In_605,In_1682);
and U3364 (N_3364,In_954,In_2429);
or U3365 (N_3365,In_2265,In_31);
and U3366 (N_3366,In_918,In_132);
and U3367 (N_3367,In_1548,In_1164);
nand U3368 (N_3368,In_485,In_2061);
nor U3369 (N_3369,In_1015,In_2339);
nor U3370 (N_3370,In_1482,In_738);
nand U3371 (N_3371,In_39,In_455);
nand U3372 (N_3372,In_2450,In_1209);
and U3373 (N_3373,In_2753,In_2572);
nor U3374 (N_3374,In_1422,In_2032);
and U3375 (N_3375,In_2886,In_909);
nand U3376 (N_3376,In_2103,In_158);
and U3377 (N_3377,In_2059,In_2629);
nor U3378 (N_3378,In_2912,In_267);
or U3379 (N_3379,In_1241,In_1824);
nand U3380 (N_3380,In_1826,In_1142);
and U3381 (N_3381,In_1387,In_623);
nand U3382 (N_3382,In_157,In_2017);
nand U3383 (N_3383,In_859,In_77);
or U3384 (N_3384,In_2582,In_1005);
and U3385 (N_3385,In_2818,In_2632);
nor U3386 (N_3386,In_1549,In_465);
nand U3387 (N_3387,In_203,In_34);
or U3388 (N_3388,In_2772,In_2351);
xnor U3389 (N_3389,In_2260,In_2380);
or U3390 (N_3390,In_2497,In_1409);
nand U3391 (N_3391,In_1352,In_1743);
xnor U3392 (N_3392,In_1801,In_2079);
nand U3393 (N_3393,In_1304,In_1060);
nor U3394 (N_3394,In_1658,In_132);
nand U3395 (N_3395,In_2365,In_421);
nand U3396 (N_3396,In_992,In_1239);
nor U3397 (N_3397,In_698,In_1651);
and U3398 (N_3398,In_1407,In_1543);
nand U3399 (N_3399,In_2290,In_2447);
and U3400 (N_3400,In_1065,In_1727);
nor U3401 (N_3401,In_2898,In_1340);
nand U3402 (N_3402,In_1523,In_861);
nor U3403 (N_3403,In_611,In_771);
nand U3404 (N_3404,In_572,In_2283);
nand U3405 (N_3405,In_2836,In_2566);
nand U3406 (N_3406,In_736,In_1427);
nand U3407 (N_3407,In_2227,In_101);
and U3408 (N_3408,In_1100,In_2633);
xor U3409 (N_3409,In_782,In_1543);
or U3410 (N_3410,In_2788,In_105);
nor U3411 (N_3411,In_2284,In_926);
or U3412 (N_3412,In_2506,In_847);
xnor U3413 (N_3413,In_373,In_1922);
and U3414 (N_3414,In_1838,In_2148);
or U3415 (N_3415,In_1014,In_1114);
nand U3416 (N_3416,In_2366,In_441);
nor U3417 (N_3417,In_501,In_2810);
or U3418 (N_3418,In_49,In_103);
nand U3419 (N_3419,In_943,In_1404);
nand U3420 (N_3420,In_1848,In_1579);
or U3421 (N_3421,In_1047,In_2181);
nand U3422 (N_3422,In_1568,In_1638);
and U3423 (N_3423,In_12,In_1515);
nand U3424 (N_3424,In_2773,In_2133);
or U3425 (N_3425,In_2907,In_1492);
nor U3426 (N_3426,In_2983,In_290);
nor U3427 (N_3427,In_1063,In_92);
or U3428 (N_3428,In_627,In_1472);
nor U3429 (N_3429,In_322,In_1133);
nor U3430 (N_3430,In_1409,In_1252);
or U3431 (N_3431,In_2572,In_2450);
or U3432 (N_3432,In_2490,In_519);
nor U3433 (N_3433,In_2943,In_859);
nand U3434 (N_3434,In_2245,In_478);
nand U3435 (N_3435,In_920,In_1492);
nand U3436 (N_3436,In_783,In_1538);
and U3437 (N_3437,In_1628,In_2563);
nor U3438 (N_3438,In_724,In_1434);
nand U3439 (N_3439,In_1768,In_1901);
and U3440 (N_3440,In_2634,In_2627);
nor U3441 (N_3441,In_1598,In_1721);
nand U3442 (N_3442,In_2405,In_53);
nand U3443 (N_3443,In_2986,In_2983);
or U3444 (N_3444,In_1824,In_430);
xnor U3445 (N_3445,In_2416,In_1536);
or U3446 (N_3446,In_1315,In_705);
nand U3447 (N_3447,In_675,In_2137);
nand U3448 (N_3448,In_1333,In_2896);
or U3449 (N_3449,In_1724,In_114);
or U3450 (N_3450,In_676,In_728);
nor U3451 (N_3451,In_2139,In_329);
nor U3452 (N_3452,In_746,In_2379);
nor U3453 (N_3453,In_318,In_517);
or U3454 (N_3454,In_2917,In_2299);
and U3455 (N_3455,In_1373,In_2722);
nand U3456 (N_3456,In_1645,In_2185);
nor U3457 (N_3457,In_1400,In_2692);
and U3458 (N_3458,In_125,In_511);
xor U3459 (N_3459,In_2143,In_2100);
or U3460 (N_3460,In_2351,In_1753);
nor U3461 (N_3461,In_2662,In_2284);
and U3462 (N_3462,In_2785,In_963);
nand U3463 (N_3463,In_886,In_611);
or U3464 (N_3464,In_1569,In_326);
nand U3465 (N_3465,In_1413,In_266);
nor U3466 (N_3466,In_358,In_1034);
nand U3467 (N_3467,In_2530,In_1897);
nand U3468 (N_3468,In_1933,In_2201);
or U3469 (N_3469,In_1863,In_0);
nand U3470 (N_3470,In_171,In_2765);
nand U3471 (N_3471,In_1873,In_688);
and U3472 (N_3472,In_1172,In_2770);
nand U3473 (N_3473,In_1203,In_1963);
nand U3474 (N_3474,In_2163,In_1795);
nor U3475 (N_3475,In_1265,In_118);
and U3476 (N_3476,In_1996,In_887);
nand U3477 (N_3477,In_768,In_789);
nand U3478 (N_3478,In_202,In_1510);
or U3479 (N_3479,In_2213,In_2407);
or U3480 (N_3480,In_744,In_1197);
nand U3481 (N_3481,In_313,In_1914);
or U3482 (N_3482,In_255,In_844);
nand U3483 (N_3483,In_2020,In_1009);
and U3484 (N_3484,In_2430,In_2249);
nor U3485 (N_3485,In_2073,In_212);
nor U3486 (N_3486,In_2513,In_1880);
and U3487 (N_3487,In_2086,In_709);
nor U3488 (N_3488,In_216,In_2265);
nand U3489 (N_3489,In_529,In_2597);
nand U3490 (N_3490,In_635,In_1005);
nor U3491 (N_3491,In_1799,In_2658);
and U3492 (N_3492,In_2612,In_1589);
and U3493 (N_3493,In_350,In_9);
xnor U3494 (N_3494,In_2754,In_1806);
or U3495 (N_3495,In_389,In_24);
nor U3496 (N_3496,In_1813,In_531);
or U3497 (N_3497,In_1566,In_691);
nand U3498 (N_3498,In_790,In_1092);
or U3499 (N_3499,In_330,In_64);
and U3500 (N_3500,In_70,In_360);
nand U3501 (N_3501,In_2812,In_1809);
nor U3502 (N_3502,In_1048,In_2209);
nand U3503 (N_3503,In_1846,In_1951);
and U3504 (N_3504,In_494,In_1768);
xnor U3505 (N_3505,In_2587,In_692);
nor U3506 (N_3506,In_1676,In_2273);
xor U3507 (N_3507,In_784,In_1399);
xor U3508 (N_3508,In_2209,In_2832);
nand U3509 (N_3509,In_1113,In_1466);
or U3510 (N_3510,In_1916,In_982);
or U3511 (N_3511,In_1026,In_306);
nor U3512 (N_3512,In_295,In_21);
xor U3513 (N_3513,In_1199,In_437);
nand U3514 (N_3514,In_2641,In_1940);
or U3515 (N_3515,In_312,In_151);
and U3516 (N_3516,In_488,In_2524);
or U3517 (N_3517,In_2474,In_412);
and U3518 (N_3518,In_448,In_461);
nor U3519 (N_3519,In_1045,In_2955);
and U3520 (N_3520,In_184,In_2453);
nand U3521 (N_3521,In_375,In_1343);
and U3522 (N_3522,In_509,In_245);
nand U3523 (N_3523,In_1993,In_1479);
xnor U3524 (N_3524,In_1481,In_383);
xnor U3525 (N_3525,In_633,In_644);
nor U3526 (N_3526,In_408,In_1794);
and U3527 (N_3527,In_922,In_2223);
and U3528 (N_3528,In_1057,In_1160);
nand U3529 (N_3529,In_2005,In_966);
xnor U3530 (N_3530,In_2645,In_350);
nand U3531 (N_3531,In_130,In_2030);
nand U3532 (N_3532,In_2759,In_181);
nand U3533 (N_3533,In_1079,In_949);
or U3534 (N_3534,In_1406,In_2159);
and U3535 (N_3535,In_2831,In_2625);
nand U3536 (N_3536,In_746,In_1340);
or U3537 (N_3537,In_2202,In_747);
or U3538 (N_3538,In_1366,In_2194);
or U3539 (N_3539,In_511,In_2281);
or U3540 (N_3540,In_1735,In_2101);
nand U3541 (N_3541,In_2141,In_2485);
nand U3542 (N_3542,In_879,In_2984);
nand U3543 (N_3543,In_2526,In_600);
or U3544 (N_3544,In_1492,In_2259);
nand U3545 (N_3545,In_655,In_2007);
xnor U3546 (N_3546,In_1403,In_1444);
nor U3547 (N_3547,In_1422,In_195);
nand U3548 (N_3548,In_185,In_478);
nand U3549 (N_3549,In_923,In_1181);
or U3550 (N_3550,In_620,In_1015);
nand U3551 (N_3551,In_1745,In_1312);
nand U3552 (N_3552,In_242,In_1712);
or U3553 (N_3553,In_1812,In_2862);
and U3554 (N_3554,In_987,In_217);
nor U3555 (N_3555,In_662,In_2023);
or U3556 (N_3556,In_2774,In_2960);
nand U3557 (N_3557,In_2146,In_1458);
and U3558 (N_3558,In_1306,In_347);
or U3559 (N_3559,In_2407,In_2002);
or U3560 (N_3560,In_1516,In_386);
or U3561 (N_3561,In_2782,In_715);
nor U3562 (N_3562,In_2277,In_2506);
or U3563 (N_3563,In_1208,In_2712);
nor U3564 (N_3564,In_1167,In_817);
or U3565 (N_3565,In_2060,In_827);
or U3566 (N_3566,In_2409,In_2278);
and U3567 (N_3567,In_2813,In_630);
and U3568 (N_3568,In_1170,In_673);
nor U3569 (N_3569,In_1861,In_646);
or U3570 (N_3570,In_2736,In_752);
nand U3571 (N_3571,In_86,In_1905);
nand U3572 (N_3572,In_933,In_760);
nand U3573 (N_3573,In_533,In_1391);
and U3574 (N_3574,In_2059,In_1056);
xnor U3575 (N_3575,In_1749,In_823);
or U3576 (N_3576,In_614,In_2981);
and U3577 (N_3577,In_2124,In_521);
and U3578 (N_3578,In_35,In_1391);
and U3579 (N_3579,In_2242,In_2917);
or U3580 (N_3580,In_2478,In_2840);
or U3581 (N_3581,In_2932,In_1172);
nor U3582 (N_3582,In_1949,In_397);
or U3583 (N_3583,In_130,In_2340);
and U3584 (N_3584,In_687,In_297);
nand U3585 (N_3585,In_641,In_1556);
nor U3586 (N_3586,In_2611,In_2725);
and U3587 (N_3587,In_220,In_1541);
or U3588 (N_3588,In_406,In_1464);
nand U3589 (N_3589,In_120,In_2278);
nand U3590 (N_3590,In_2422,In_2450);
and U3591 (N_3591,In_2990,In_251);
or U3592 (N_3592,In_1759,In_1493);
nor U3593 (N_3593,In_2393,In_2376);
nand U3594 (N_3594,In_2965,In_1275);
nor U3595 (N_3595,In_1243,In_809);
and U3596 (N_3596,In_1601,In_1547);
or U3597 (N_3597,In_1453,In_2831);
nor U3598 (N_3598,In_2954,In_343);
and U3599 (N_3599,In_1532,In_263);
nand U3600 (N_3600,In_662,In_2927);
nand U3601 (N_3601,In_2575,In_1783);
xnor U3602 (N_3602,In_1028,In_1359);
and U3603 (N_3603,In_2726,In_1484);
nand U3604 (N_3604,In_270,In_2191);
nor U3605 (N_3605,In_1136,In_2422);
nor U3606 (N_3606,In_982,In_13);
or U3607 (N_3607,In_2863,In_1280);
or U3608 (N_3608,In_21,In_2136);
and U3609 (N_3609,In_1530,In_1273);
nand U3610 (N_3610,In_2044,In_2711);
and U3611 (N_3611,In_2768,In_2865);
or U3612 (N_3612,In_314,In_1237);
or U3613 (N_3613,In_2476,In_588);
nand U3614 (N_3614,In_629,In_805);
and U3615 (N_3615,In_2471,In_2521);
nor U3616 (N_3616,In_1761,In_1019);
nor U3617 (N_3617,In_2081,In_1732);
nand U3618 (N_3618,In_1620,In_1743);
or U3619 (N_3619,In_2632,In_563);
and U3620 (N_3620,In_2120,In_1834);
nand U3621 (N_3621,In_1023,In_2593);
and U3622 (N_3622,In_1225,In_2417);
nand U3623 (N_3623,In_2268,In_930);
nor U3624 (N_3624,In_1868,In_2810);
nand U3625 (N_3625,In_1324,In_517);
and U3626 (N_3626,In_569,In_2652);
or U3627 (N_3627,In_2709,In_2670);
and U3628 (N_3628,In_971,In_547);
and U3629 (N_3629,In_965,In_621);
and U3630 (N_3630,In_766,In_2604);
or U3631 (N_3631,In_1209,In_1819);
and U3632 (N_3632,In_361,In_2932);
or U3633 (N_3633,In_2840,In_248);
or U3634 (N_3634,In_1618,In_670);
xor U3635 (N_3635,In_1070,In_2581);
nand U3636 (N_3636,In_193,In_1200);
nor U3637 (N_3637,In_1653,In_2638);
nor U3638 (N_3638,In_385,In_1894);
nor U3639 (N_3639,In_1632,In_726);
or U3640 (N_3640,In_987,In_944);
xnor U3641 (N_3641,In_1694,In_757);
nor U3642 (N_3642,In_462,In_299);
nand U3643 (N_3643,In_668,In_2372);
nand U3644 (N_3644,In_1048,In_1992);
nand U3645 (N_3645,In_1136,In_852);
nor U3646 (N_3646,In_2711,In_2772);
nor U3647 (N_3647,In_2602,In_1509);
or U3648 (N_3648,In_415,In_1688);
or U3649 (N_3649,In_2662,In_1984);
xor U3650 (N_3650,In_413,In_2238);
and U3651 (N_3651,In_2749,In_2678);
xnor U3652 (N_3652,In_1430,In_1807);
and U3653 (N_3653,In_260,In_420);
nor U3654 (N_3654,In_2174,In_1163);
or U3655 (N_3655,In_320,In_1729);
or U3656 (N_3656,In_1827,In_772);
and U3657 (N_3657,In_2615,In_1507);
nand U3658 (N_3658,In_513,In_2062);
and U3659 (N_3659,In_2425,In_1500);
nand U3660 (N_3660,In_1905,In_1912);
xor U3661 (N_3661,In_2414,In_1395);
and U3662 (N_3662,In_2873,In_614);
nor U3663 (N_3663,In_2804,In_2807);
and U3664 (N_3664,In_1129,In_1594);
xnor U3665 (N_3665,In_2937,In_316);
nor U3666 (N_3666,In_610,In_337);
and U3667 (N_3667,In_1347,In_336);
nand U3668 (N_3668,In_2454,In_1054);
nand U3669 (N_3669,In_903,In_1684);
and U3670 (N_3670,In_412,In_1266);
or U3671 (N_3671,In_2768,In_110);
and U3672 (N_3672,In_1935,In_2619);
nor U3673 (N_3673,In_792,In_419);
nand U3674 (N_3674,In_2149,In_1383);
xnor U3675 (N_3675,In_668,In_1435);
nor U3676 (N_3676,In_2387,In_1698);
nand U3677 (N_3677,In_104,In_2634);
and U3678 (N_3678,In_846,In_1551);
and U3679 (N_3679,In_1679,In_1797);
or U3680 (N_3680,In_1019,In_2185);
and U3681 (N_3681,In_2791,In_2288);
or U3682 (N_3682,In_1128,In_849);
nand U3683 (N_3683,In_1416,In_625);
nand U3684 (N_3684,In_1314,In_2805);
and U3685 (N_3685,In_1818,In_1993);
nor U3686 (N_3686,In_277,In_1475);
or U3687 (N_3687,In_2133,In_692);
and U3688 (N_3688,In_1218,In_2166);
and U3689 (N_3689,In_2722,In_92);
or U3690 (N_3690,In_2193,In_2491);
nor U3691 (N_3691,In_268,In_2461);
nor U3692 (N_3692,In_1382,In_1766);
nor U3693 (N_3693,In_1548,In_937);
and U3694 (N_3694,In_2172,In_2463);
and U3695 (N_3695,In_881,In_211);
nand U3696 (N_3696,In_2346,In_1517);
and U3697 (N_3697,In_1705,In_1524);
nand U3698 (N_3698,In_178,In_2525);
and U3699 (N_3699,In_1811,In_765);
or U3700 (N_3700,In_425,In_1666);
or U3701 (N_3701,In_2189,In_1592);
nor U3702 (N_3702,In_2799,In_1227);
nor U3703 (N_3703,In_2338,In_324);
nand U3704 (N_3704,In_1650,In_2802);
and U3705 (N_3705,In_520,In_465);
nor U3706 (N_3706,In_1117,In_235);
or U3707 (N_3707,In_224,In_2790);
nor U3708 (N_3708,In_616,In_389);
and U3709 (N_3709,In_1733,In_794);
nand U3710 (N_3710,In_517,In_1698);
nor U3711 (N_3711,In_1933,In_1673);
nor U3712 (N_3712,In_2693,In_825);
nand U3713 (N_3713,In_1925,In_1027);
nand U3714 (N_3714,In_2045,In_1807);
xor U3715 (N_3715,In_2664,In_762);
nand U3716 (N_3716,In_1365,In_1691);
and U3717 (N_3717,In_2028,In_2923);
or U3718 (N_3718,In_2994,In_1956);
nor U3719 (N_3719,In_1206,In_652);
nand U3720 (N_3720,In_1099,In_2454);
and U3721 (N_3721,In_2169,In_2455);
nand U3722 (N_3722,In_2638,In_2679);
nand U3723 (N_3723,In_2219,In_1191);
nor U3724 (N_3724,In_1263,In_69);
or U3725 (N_3725,In_7,In_566);
xor U3726 (N_3726,In_2114,In_1495);
nand U3727 (N_3727,In_2054,In_2806);
and U3728 (N_3728,In_1415,In_1755);
nand U3729 (N_3729,In_876,In_1342);
or U3730 (N_3730,In_860,In_1682);
nor U3731 (N_3731,In_332,In_866);
or U3732 (N_3732,In_459,In_1643);
and U3733 (N_3733,In_1532,In_368);
and U3734 (N_3734,In_1294,In_573);
xnor U3735 (N_3735,In_2433,In_896);
xor U3736 (N_3736,In_1530,In_67);
or U3737 (N_3737,In_2225,In_1809);
and U3738 (N_3738,In_1356,In_2759);
nand U3739 (N_3739,In_2475,In_1408);
and U3740 (N_3740,In_2644,In_1547);
and U3741 (N_3741,In_1017,In_2812);
nor U3742 (N_3742,In_1029,In_2664);
nor U3743 (N_3743,In_2617,In_921);
or U3744 (N_3744,In_369,In_1067);
or U3745 (N_3745,In_1005,In_267);
nor U3746 (N_3746,In_0,In_1772);
nand U3747 (N_3747,In_305,In_233);
xnor U3748 (N_3748,In_2057,In_204);
and U3749 (N_3749,In_2595,In_1235);
nand U3750 (N_3750,In_828,In_395);
nand U3751 (N_3751,In_2736,In_152);
and U3752 (N_3752,In_2126,In_1911);
nand U3753 (N_3753,In_907,In_1111);
nor U3754 (N_3754,In_2108,In_1281);
nor U3755 (N_3755,In_1446,In_449);
or U3756 (N_3756,In_2866,In_2793);
xor U3757 (N_3757,In_445,In_819);
or U3758 (N_3758,In_1999,In_679);
nand U3759 (N_3759,In_44,In_495);
nor U3760 (N_3760,In_184,In_1160);
nand U3761 (N_3761,In_1477,In_169);
and U3762 (N_3762,In_2831,In_2936);
nand U3763 (N_3763,In_1792,In_1689);
or U3764 (N_3764,In_1894,In_171);
nand U3765 (N_3765,In_2664,In_2);
and U3766 (N_3766,In_913,In_1373);
nor U3767 (N_3767,In_2290,In_824);
and U3768 (N_3768,In_2811,In_1075);
nand U3769 (N_3769,In_2965,In_337);
and U3770 (N_3770,In_2911,In_1870);
nor U3771 (N_3771,In_1902,In_1463);
nor U3772 (N_3772,In_1329,In_1630);
and U3773 (N_3773,In_2620,In_1958);
nor U3774 (N_3774,In_1699,In_1019);
nor U3775 (N_3775,In_24,In_121);
or U3776 (N_3776,In_1221,In_1261);
nor U3777 (N_3777,In_21,In_458);
nor U3778 (N_3778,In_2879,In_2308);
nor U3779 (N_3779,In_1462,In_2852);
or U3780 (N_3780,In_1145,In_1554);
xor U3781 (N_3781,In_43,In_643);
or U3782 (N_3782,In_375,In_2497);
nand U3783 (N_3783,In_98,In_296);
or U3784 (N_3784,In_2901,In_480);
nand U3785 (N_3785,In_2186,In_56);
or U3786 (N_3786,In_437,In_2935);
or U3787 (N_3787,In_830,In_2176);
or U3788 (N_3788,In_1629,In_204);
and U3789 (N_3789,In_407,In_79);
nor U3790 (N_3790,In_2908,In_2145);
nor U3791 (N_3791,In_2426,In_2064);
and U3792 (N_3792,In_1255,In_96);
nand U3793 (N_3793,In_1093,In_2324);
nor U3794 (N_3794,In_438,In_1190);
or U3795 (N_3795,In_51,In_514);
nand U3796 (N_3796,In_2491,In_625);
nor U3797 (N_3797,In_1809,In_1726);
or U3798 (N_3798,In_2122,In_1262);
xnor U3799 (N_3799,In_291,In_2387);
and U3800 (N_3800,In_1981,In_2597);
or U3801 (N_3801,In_22,In_1144);
or U3802 (N_3802,In_1224,In_1802);
xor U3803 (N_3803,In_2147,In_466);
nand U3804 (N_3804,In_94,In_515);
and U3805 (N_3805,In_723,In_675);
nand U3806 (N_3806,In_2463,In_815);
or U3807 (N_3807,In_611,In_55);
or U3808 (N_3808,In_495,In_2003);
nor U3809 (N_3809,In_548,In_81);
and U3810 (N_3810,In_307,In_219);
nand U3811 (N_3811,In_991,In_224);
and U3812 (N_3812,In_2507,In_2353);
or U3813 (N_3813,In_587,In_1684);
and U3814 (N_3814,In_350,In_2778);
nor U3815 (N_3815,In_903,In_2097);
or U3816 (N_3816,In_1260,In_1506);
nand U3817 (N_3817,In_2520,In_628);
or U3818 (N_3818,In_861,In_1460);
and U3819 (N_3819,In_144,In_222);
nor U3820 (N_3820,In_1647,In_2107);
nor U3821 (N_3821,In_2042,In_144);
nor U3822 (N_3822,In_2571,In_1177);
or U3823 (N_3823,In_2471,In_1176);
or U3824 (N_3824,In_1710,In_2583);
nand U3825 (N_3825,In_645,In_1704);
nand U3826 (N_3826,In_2905,In_754);
or U3827 (N_3827,In_2631,In_36);
nand U3828 (N_3828,In_1826,In_1331);
xor U3829 (N_3829,In_703,In_994);
and U3830 (N_3830,In_962,In_2231);
nor U3831 (N_3831,In_109,In_110);
nor U3832 (N_3832,In_2192,In_1571);
and U3833 (N_3833,In_2365,In_2160);
or U3834 (N_3834,In_1841,In_2941);
or U3835 (N_3835,In_2203,In_915);
and U3836 (N_3836,In_1329,In_718);
or U3837 (N_3837,In_370,In_695);
and U3838 (N_3838,In_2868,In_1854);
or U3839 (N_3839,In_1163,In_466);
nand U3840 (N_3840,In_1017,In_2856);
and U3841 (N_3841,In_2228,In_2565);
and U3842 (N_3842,In_1270,In_2214);
nor U3843 (N_3843,In_1138,In_873);
nor U3844 (N_3844,In_744,In_2593);
and U3845 (N_3845,In_104,In_1282);
and U3846 (N_3846,In_2275,In_1636);
and U3847 (N_3847,In_2151,In_841);
or U3848 (N_3848,In_727,In_2094);
or U3849 (N_3849,In_1558,In_2505);
nor U3850 (N_3850,In_236,In_2988);
nand U3851 (N_3851,In_2565,In_2066);
nor U3852 (N_3852,In_1151,In_2240);
or U3853 (N_3853,In_2456,In_408);
and U3854 (N_3854,In_930,In_1022);
or U3855 (N_3855,In_345,In_92);
nand U3856 (N_3856,In_2111,In_2241);
nand U3857 (N_3857,In_1664,In_1857);
and U3858 (N_3858,In_1948,In_1072);
nor U3859 (N_3859,In_2085,In_1512);
nand U3860 (N_3860,In_1099,In_2287);
nand U3861 (N_3861,In_1248,In_2250);
and U3862 (N_3862,In_267,In_946);
and U3863 (N_3863,In_2582,In_2049);
or U3864 (N_3864,In_1985,In_831);
and U3865 (N_3865,In_1299,In_891);
nor U3866 (N_3866,In_2234,In_2895);
nand U3867 (N_3867,In_2693,In_44);
nor U3868 (N_3868,In_540,In_2867);
or U3869 (N_3869,In_2178,In_1461);
nor U3870 (N_3870,In_2844,In_2178);
nand U3871 (N_3871,In_2192,In_1541);
nor U3872 (N_3872,In_1832,In_2334);
nand U3873 (N_3873,In_2980,In_1775);
nor U3874 (N_3874,In_2504,In_1555);
and U3875 (N_3875,In_2543,In_1562);
or U3876 (N_3876,In_1490,In_7);
and U3877 (N_3877,In_1391,In_2065);
nand U3878 (N_3878,In_867,In_1342);
nor U3879 (N_3879,In_1435,In_2674);
or U3880 (N_3880,In_531,In_660);
nor U3881 (N_3881,In_244,In_1049);
nand U3882 (N_3882,In_2972,In_1207);
nand U3883 (N_3883,In_1194,In_372);
and U3884 (N_3884,In_1232,In_102);
and U3885 (N_3885,In_2694,In_2463);
and U3886 (N_3886,In_2855,In_2851);
nand U3887 (N_3887,In_559,In_1287);
nor U3888 (N_3888,In_1621,In_651);
nand U3889 (N_3889,In_2996,In_2838);
or U3890 (N_3890,In_2652,In_1953);
or U3891 (N_3891,In_66,In_1619);
nand U3892 (N_3892,In_2381,In_981);
and U3893 (N_3893,In_1582,In_1722);
and U3894 (N_3894,In_2037,In_2817);
and U3895 (N_3895,In_800,In_1370);
and U3896 (N_3896,In_2417,In_31);
and U3897 (N_3897,In_222,In_1817);
nor U3898 (N_3898,In_1555,In_1917);
or U3899 (N_3899,In_2375,In_151);
xor U3900 (N_3900,In_2890,In_1052);
nand U3901 (N_3901,In_1422,In_834);
or U3902 (N_3902,In_1764,In_660);
and U3903 (N_3903,In_658,In_985);
or U3904 (N_3904,In_1608,In_2963);
xnor U3905 (N_3905,In_2267,In_2840);
nor U3906 (N_3906,In_1658,In_377);
nand U3907 (N_3907,In_2463,In_1530);
and U3908 (N_3908,In_343,In_2770);
nor U3909 (N_3909,In_500,In_0);
nand U3910 (N_3910,In_1816,In_573);
or U3911 (N_3911,In_765,In_1830);
nand U3912 (N_3912,In_2582,In_1046);
nor U3913 (N_3913,In_242,In_2719);
nor U3914 (N_3914,In_487,In_1039);
xnor U3915 (N_3915,In_1158,In_2262);
nor U3916 (N_3916,In_2743,In_1232);
nand U3917 (N_3917,In_568,In_1077);
nand U3918 (N_3918,In_203,In_576);
or U3919 (N_3919,In_430,In_150);
and U3920 (N_3920,In_1810,In_2341);
nor U3921 (N_3921,In_2474,In_2043);
and U3922 (N_3922,In_1944,In_811);
and U3923 (N_3923,In_541,In_2139);
nand U3924 (N_3924,In_1526,In_1706);
nor U3925 (N_3925,In_1439,In_2751);
and U3926 (N_3926,In_2821,In_1104);
nor U3927 (N_3927,In_2860,In_2916);
nand U3928 (N_3928,In_1210,In_289);
nand U3929 (N_3929,In_2938,In_1304);
nor U3930 (N_3930,In_1244,In_1969);
nand U3931 (N_3931,In_2886,In_2567);
nor U3932 (N_3932,In_2154,In_2256);
or U3933 (N_3933,In_437,In_1046);
nand U3934 (N_3934,In_426,In_1512);
xnor U3935 (N_3935,In_1810,In_2935);
or U3936 (N_3936,In_744,In_2029);
and U3937 (N_3937,In_85,In_1318);
xnor U3938 (N_3938,In_1456,In_1186);
or U3939 (N_3939,In_2813,In_893);
or U3940 (N_3940,In_678,In_1077);
and U3941 (N_3941,In_1793,In_1755);
nand U3942 (N_3942,In_2758,In_1347);
nor U3943 (N_3943,In_1239,In_2733);
xnor U3944 (N_3944,In_452,In_1403);
or U3945 (N_3945,In_2942,In_1921);
nand U3946 (N_3946,In_586,In_1083);
xnor U3947 (N_3947,In_769,In_1051);
nand U3948 (N_3948,In_221,In_2879);
nand U3949 (N_3949,In_2737,In_371);
xnor U3950 (N_3950,In_532,In_258);
and U3951 (N_3951,In_281,In_1034);
and U3952 (N_3952,In_1425,In_2494);
or U3953 (N_3953,In_1616,In_2637);
or U3954 (N_3954,In_2351,In_2259);
nand U3955 (N_3955,In_134,In_1410);
or U3956 (N_3956,In_2572,In_1133);
nor U3957 (N_3957,In_1604,In_1086);
or U3958 (N_3958,In_882,In_232);
or U3959 (N_3959,In_96,In_2259);
and U3960 (N_3960,In_266,In_571);
and U3961 (N_3961,In_2035,In_2146);
nor U3962 (N_3962,In_1751,In_1626);
or U3963 (N_3963,In_2768,In_162);
nand U3964 (N_3964,In_932,In_2090);
or U3965 (N_3965,In_1502,In_1307);
nor U3966 (N_3966,In_566,In_1035);
or U3967 (N_3967,In_2785,In_1283);
and U3968 (N_3968,In_2775,In_582);
nor U3969 (N_3969,In_1810,In_1963);
nor U3970 (N_3970,In_2400,In_2462);
or U3971 (N_3971,In_1723,In_1079);
and U3972 (N_3972,In_131,In_2687);
or U3973 (N_3973,In_2656,In_912);
xor U3974 (N_3974,In_1068,In_1090);
and U3975 (N_3975,In_2644,In_2820);
nand U3976 (N_3976,In_2391,In_1216);
and U3977 (N_3977,In_1970,In_1040);
or U3978 (N_3978,In_47,In_62);
xnor U3979 (N_3979,In_1843,In_2862);
and U3980 (N_3980,In_1802,In_1116);
nand U3981 (N_3981,In_822,In_1899);
nand U3982 (N_3982,In_1448,In_1411);
nand U3983 (N_3983,In_991,In_1958);
nand U3984 (N_3984,In_1320,In_70);
or U3985 (N_3985,In_2737,In_2618);
nand U3986 (N_3986,In_1442,In_2187);
or U3987 (N_3987,In_2229,In_1974);
nor U3988 (N_3988,In_2976,In_213);
nand U3989 (N_3989,In_1297,In_1254);
and U3990 (N_3990,In_2594,In_2660);
xnor U3991 (N_3991,In_1500,In_876);
or U3992 (N_3992,In_1764,In_1414);
or U3993 (N_3993,In_64,In_2209);
nor U3994 (N_3994,In_1758,In_2608);
xor U3995 (N_3995,In_1834,In_1998);
nor U3996 (N_3996,In_460,In_791);
nand U3997 (N_3997,In_679,In_1132);
nor U3998 (N_3998,In_2759,In_2932);
and U3999 (N_3999,In_230,In_1662);
nand U4000 (N_4000,In_1671,In_1336);
nand U4001 (N_4001,In_1399,In_1472);
or U4002 (N_4002,In_82,In_1784);
nand U4003 (N_4003,In_132,In_257);
or U4004 (N_4004,In_324,In_2476);
nand U4005 (N_4005,In_1234,In_401);
or U4006 (N_4006,In_2169,In_389);
or U4007 (N_4007,In_877,In_1632);
or U4008 (N_4008,In_2236,In_2768);
and U4009 (N_4009,In_1488,In_1900);
or U4010 (N_4010,In_1695,In_2584);
or U4011 (N_4011,In_1553,In_2776);
xor U4012 (N_4012,In_297,In_2561);
nor U4013 (N_4013,In_2067,In_904);
or U4014 (N_4014,In_44,In_157);
xor U4015 (N_4015,In_2449,In_1735);
or U4016 (N_4016,In_2378,In_2333);
nand U4017 (N_4017,In_2149,In_1332);
nor U4018 (N_4018,In_2977,In_1399);
nand U4019 (N_4019,In_1726,In_1131);
and U4020 (N_4020,In_1835,In_1428);
xor U4021 (N_4021,In_792,In_1569);
xnor U4022 (N_4022,In_2060,In_123);
nand U4023 (N_4023,In_580,In_509);
or U4024 (N_4024,In_1505,In_1004);
nor U4025 (N_4025,In_1069,In_2890);
nand U4026 (N_4026,In_1351,In_2454);
and U4027 (N_4027,In_1109,In_2328);
nor U4028 (N_4028,In_2908,In_1450);
or U4029 (N_4029,In_804,In_79);
and U4030 (N_4030,In_840,In_2646);
nand U4031 (N_4031,In_2798,In_906);
and U4032 (N_4032,In_41,In_221);
or U4033 (N_4033,In_1138,In_1725);
and U4034 (N_4034,In_542,In_2901);
and U4035 (N_4035,In_1358,In_2532);
nor U4036 (N_4036,In_2451,In_1063);
and U4037 (N_4037,In_447,In_2154);
nor U4038 (N_4038,In_2691,In_836);
and U4039 (N_4039,In_171,In_2862);
nand U4040 (N_4040,In_2205,In_1464);
and U4041 (N_4041,In_2745,In_603);
nand U4042 (N_4042,In_1279,In_1745);
or U4043 (N_4043,In_1037,In_144);
nand U4044 (N_4044,In_491,In_1678);
nor U4045 (N_4045,In_794,In_2700);
and U4046 (N_4046,In_90,In_2579);
nor U4047 (N_4047,In_488,In_2167);
nand U4048 (N_4048,In_119,In_2455);
and U4049 (N_4049,In_1341,In_2029);
or U4050 (N_4050,In_1463,In_1546);
and U4051 (N_4051,In_2848,In_364);
xor U4052 (N_4052,In_1558,In_2525);
nand U4053 (N_4053,In_1840,In_280);
or U4054 (N_4054,In_1907,In_2379);
and U4055 (N_4055,In_2944,In_2441);
nand U4056 (N_4056,In_2804,In_735);
xor U4057 (N_4057,In_3,In_1528);
nand U4058 (N_4058,In_1110,In_1796);
and U4059 (N_4059,In_1341,In_1698);
and U4060 (N_4060,In_1185,In_1787);
or U4061 (N_4061,In_2381,In_140);
or U4062 (N_4062,In_1108,In_589);
nand U4063 (N_4063,In_983,In_1388);
nand U4064 (N_4064,In_2143,In_1124);
nand U4065 (N_4065,In_680,In_259);
and U4066 (N_4066,In_1980,In_1000);
or U4067 (N_4067,In_846,In_663);
and U4068 (N_4068,In_1508,In_2960);
or U4069 (N_4069,In_1507,In_1672);
xor U4070 (N_4070,In_2780,In_1834);
nand U4071 (N_4071,In_980,In_1559);
and U4072 (N_4072,In_967,In_1311);
nor U4073 (N_4073,In_1479,In_1593);
nor U4074 (N_4074,In_1458,In_875);
or U4075 (N_4075,In_2443,In_1226);
nor U4076 (N_4076,In_574,In_690);
or U4077 (N_4077,In_1180,In_790);
nor U4078 (N_4078,In_1105,In_716);
nand U4079 (N_4079,In_1565,In_2546);
xor U4080 (N_4080,In_2211,In_648);
nand U4081 (N_4081,In_418,In_847);
nand U4082 (N_4082,In_536,In_1402);
or U4083 (N_4083,In_80,In_2675);
and U4084 (N_4084,In_1570,In_14);
nor U4085 (N_4085,In_667,In_2768);
nand U4086 (N_4086,In_51,In_1153);
nor U4087 (N_4087,In_643,In_1817);
nand U4088 (N_4088,In_2333,In_2678);
or U4089 (N_4089,In_2,In_2114);
nand U4090 (N_4090,In_2333,In_842);
nand U4091 (N_4091,In_1745,In_632);
nor U4092 (N_4092,In_1510,In_2935);
nand U4093 (N_4093,In_2310,In_2813);
nor U4094 (N_4094,In_161,In_703);
or U4095 (N_4095,In_1758,In_1764);
or U4096 (N_4096,In_563,In_96);
nor U4097 (N_4097,In_1424,In_432);
or U4098 (N_4098,In_88,In_551);
and U4099 (N_4099,In_1006,In_1833);
nand U4100 (N_4100,In_1350,In_2);
nand U4101 (N_4101,In_1230,In_1793);
nand U4102 (N_4102,In_2994,In_2378);
and U4103 (N_4103,In_1135,In_2709);
and U4104 (N_4104,In_373,In_1059);
xor U4105 (N_4105,In_815,In_1385);
and U4106 (N_4106,In_909,In_1888);
xor U4107 (N_4107,In_329,In_857);
and U4108 (N_4108,In_1587,In_2374);
nand U4109 (N_4109,In_960,In_1133);
xor U4110 (N_4110,In_262,In_533);
xor U4111 (N_4111,In_2487,In_1188);
and U4112 (N_4112,In_769,In_1408);
nand U4113 (N_4113,In_1395,In_2009);
or U4114 (N_4114,In_1532,In_110);
nand U4115 (N_4115,In_2821,In_2947);
or U4116 (N_4116,In_1983,In_1494);
xor U4117 (N_4117,In_2686,In_2465);
and U4118 (N_4118,In_2171,In_1081);
and U4119 (N_4119,In_1760,In_2461);
nor U4120 (N_4120,In_1221,In_779);
xnor U4121 (N_4121,In_2922,In_134);
xnor U4122 (N_4122,In_1836,In_2612);
nor U4123 (N_4123,In_1486,In_815);
nor U4124 (N_4124,In_1314,In_1530);
nand U4125 (N_4125,In_2496,In_1632);
xnor U4126 (N_4126,In_2485,In_1363);
nand U4127 (N_4127,In_2559,In_2902);
nand U4128 (N_4128,In_171,In_2236);
and U4129 (N_4129,In_1064,In_873);
or U4130 (N_4130,In_2911,In_1081);
or U4131 (N_4131,In_1870,In_1852);
and U4132 (N_4132,In_1021,In_167);
or U4133 (N_4133,In_30,In_890);
nor U4134 (N_4134,In_1456,In_2738);
nand U4135 (N_4135,In_353,In_855);
or U4136 (N_4136,In_1905,In_2002);
nor U4137 (N_4137,In_967,In_0);
or U4138 (N_4138,In_2894,In_2114);
nand U4139 (N_4139,In_491,In_1412);
nor U4140 (N_4140,In_1894,In_2540);
and U4141 (N_4141,In_138,In_1027);
nor U4142 (N_4142,In_1855,In_44);
nor U4143 (N_4143,In_630,In_2585);
nor U4144 (N_4144,In_617,In_946);
nor U4145 (N_4145,In_1567,In_1028);
and U4146 (N_4146,In_2291,In_800);
or U4147 (N_4147,In_1651,In_446);
and U4148 (N_4148,In_642,In_251);
xnor U4149 (N_4149,In_1886,In_2322);
and U4150 (N_4150,In_1855,In_466);
nor U4151 (N_4151,In_2682,In_2404);
and U4152 (N_4152,In_53,In_796);
or U4153 (N_4153,In_1421,In_1536);
and U4154 (N_4154,In_2455,In_1820);
nor U4155 (N_4155,In_119,In_7);
nand U4156 (N_4156,In_2026,In_1887);
or U4157 (N_4157,In_1750,In_2609);
and U4158 (N_4158,In_94,In_96);
nor U4159 (N_4159,In_1504,In_2671);
and U4160 (N_4160,In_2728,In_1936);
nand U4161 (N_4161,In_681,In_304);
and U4162 (N_4162,In_2873,In_2869);
nand U4163 (N_4163,In_1166,In_876);
nor U4164 (N_4164,In_2103,In_676);
nand U4165 (N_4165,In_1688,In_932);
and U4166 (N_4166,In_1980,In_290);
or U4167 (N_4167,In_719,In_120);
nand U4168 (N_4168,In_170,In_2345);
and U4169 (N_4169,In_1252,In_138);
nand U4170 (N_4170,In_824,In_281);
or U4171 (N_4171,In_1226,In_4);
nor U4172 (N_4172,In_597,In_2682);
nor U4173 (N_4173,In_269,In_465);
nor U4174 (N_4174,In_1634,In_1335);
nand U4175 (N_4175,In_2958,In_1219);
or U4176 (N_4176,In_1555,In_379);
nand U4177 (N_4177,In_2180,In_2241);
and U4178 (N_4178,In_2020,In_642);
nand U4179 (N_4179,In_900,In_1333);
and U4180 (N_4180,In_626,In_1823);
nand U4181 (N_4181,In_952,In_2541);
and U4182 (N_4182,In_2978,In_2193);
and U4183 (N_4183,In_319,In_553);
nor U4184 (N_4184,In_1244,In_1054);
nor U4185 (N_4185,In_904,In_1700);
nand U4186 (N_4186,In_1090,In_1789);
nor U4187 (N_4187,In_1394,In_304);
or U4188 (N_4188,In_2326,In_1445);
nor U4189 (N_4189,In_2118,In_649);
or U4190 (N_4190,In_1298,In_1282);
and U4191 (N_4191,In_1251,In_2975);
nor U4192 (N_4192,In_2004,In_821);
nor U4193 (N_4193,In_1691,In_170);
nor U4194 (N_4194,In_1502,In_1967);
xor U4195 (N_4195,In_25,In_442);
and U4196 (N_4196,In_1263,In_1930);
xnor U4197 (N_4197,In_1559,In_2589);
or U4198 (N_4198,In_1894,In_2988);
nand U4199 (N_4199,In_759,In_2797);
nor U4200 (N_4200,In_2734,In_517);
nor U4201 (N_4201,In_434,In_1788);
and U4202 (N_4202,In_430,In_2696);
or U4203 (N_4203,In_2709,In_2658);
nand U4204 (N_4204,In_1385,In_2232);
nand U4205 (N_4205,In_547,In_1145);
or U4206 (N_4206,In_27,In_2454);
and U4207 (N_4207,In_31,In_1881);
and U4208 (N_4208,In_948,In_2768);
or U4209 (N_4209,In_1293,In_1432);
nor U4210 (N_4210,In_1806,In_226);
and U4211 (N_4211,In_685,In_1673);
and U4212 (N_4212,In_180,In_404);
and U4213 (N_4213,In_1253,In_2446);
xor U4214 (N_4214,In_2769,In_2937);
and U4215 (N_4215,In_2060,In_1536);
and U4216 (N_4216,In_84,In_621);
and U4217 (N_4217,In_2147,In_1146);
or U4218 (N_4218,In_397,In_939);
or U4219 (N_4219,In_971,In_2453);
or U4220 (N_4220,In_2387,In_1814);
or U4221 (N_4221,In_2770,In_1392);
nor U4222 (N_4222,In_1544,In_840);
or U4223 (N_4223,In_2249,In_1639);
and U4224 (N_4224,In_2564,In_1748);
nor U4225 (N_4225,In_2058,In_2559);
nand U4226 (N_4226,In_1833,In_330);
nand U4227 (N_4227,In_666,In_1456);
nor U4228 (N_4228,In_812,In_1173);
nor U4229 (N_4229,In_713,In_937);
or U4230 (N_4230,In_2110,In_1078);
nor U4231 (N_4231,In_1362,In_2633);
nand U4232 (N_4232,In_442,In_2453);
or U4233 (N_4233,In_2596,In_2745);
and U4234 (N_4234,In_867,In_870);
or U4235 (N_4235,In_2384,In_1623);
nor U4236 (N_4236,In_1122,In_1166);
and U4237 (N_4237,In_925,In_1045);
nand U4238 (N_4238,In_2977,In_2202);
nand U4239 (N_4239,In_376,In_1818);
nand U4240 (N_4240,In_1708,In_1536);
nand U4241 (N_4241,In_2562,In_450);
and U4242 (N_4242,In_1291,In_1751);
nand U4243 (N_4243,In_1739,In_2773);
and U4244 (N_4244,In_1339,In_1601);
or U4245 (N_4245,In_1948,In_2451);
or U4246 (N_4246,In_2869,In_2726);
nand U4247 (N_4247,In_2006,In_1063);
nor U4248 (N_4248,In_792,In_141);
and U4249 (N_4249,In_2338,In_1560);
and U4250 (N_4250,In_179,In_1881);
or U4251 (N_4251,In_1386,In_79);
and U4252 (N_4252,In_94,In_2275);
or U4253 (N_4253,In_2823,In_2568);
or U4254 (N_4254,In_1111,In_2937);
nor U4255 (N_4255,In_246,In_1748);
nor U4256 (N_4256,In_763,In_1887);
nand U4257 (N_4257,In_2474,In_1467);
nor U4258 (N_4258,In_2421,In_695);
or U4259 (N_4259,In_451,In_657);
xor U4260 (N_4260,In_2742,In_741);
and U4261 (N_4261,In_657,In_918);
nor U4262 (N_4262,In_1701,In_2566);
nor U4263 (N_4263,In_420,In_1648);
xor U4264 (N_4264,In_905,In_2221);
nor U4265 (N_4265,In_2897,In_2195);
nor U4266 (N_4266,In_1629,In_2466);
nor U4267 (N_4267,In_548,In_39);
nor U4268 (N_4268,In_376,In_815);
xnor U4269 (N_4269,In_1697,In_2282);
nor U4270 (N_4270,In_2098,In_1499);
and U4271 (N_4271,In_1609,In_1234);
or U4272 (N_4272,In_621,In_108);
and U4273 (N_4273,In_2566,In_1668);
nand U4274 (N_4274,In_1874,In_303);
or U4275 (N_4275,In_1887,In_52);
and U4276 (N_4276,In_192,In_2547);
nand U4277 (N_4277,In_337,In_952);
and U4278 (N_4278,In_1141,In_738);
nand U4279 (N_4279,In_2667,In_2618);
nor U4280 (N_4280,In_2528,In_2382);
nor U4281 (N_4281,In_276,In_1198);
nor U4282 (N_4282,In_1394,In_2088);
or U4283 (N_4283,In_264,In_2062);
nand U4284 (N_4284,In_398,In_421);
and U4285 (N_4285,In_1084,In_1196);
nor U4286 (N_4286,In_2597,In_1532);
nand U4287 (N_4287,In_1916,In_2436);
nor U4288 (N_4288,In_1587,In_2484);
nor U4289 (N_4289,In_64,In_1444);
nand U4290 (N_4290,In_993,In_1689);
nand U4291 (N_4291,In_1136,In_336);
nand U4292 (N_4292,In_1352,In_1090);
nor U4293 (N_4293,In_1133,In_1867);
and U4294 (N_4294,In_1831,In_2682);
or U4295 (N_4295,In_567,In_2749);
or U4296 (N_4296,In_2843,In_1054);
and U4297 (N_4297,In_2184,In_315);
nor U4298 (N_4298,In_947,In_1194);
nand U4299 (N_4299,In_277,In_507);
nand U4300 (N_4300,In_734,In_1351);
and U4301 (N_4301,In_1082,In_2582);
or U4302 (N_4302,In_1262,In_50);
nand U4303 (N_4303,In_2585,In_2360);
nor U4304 (N_4304,In_2972,In_2903);
or U4305 (N_4305,In_2043,In_911);
and U4306 (N_4306,In_2387,In_114);
or U4307 (N_4307,In_2099,In_757);
or U4308 (N_4308,In_2712,In_1249);
or U4309 (N_4309,In_1413,In_734);
and U4310 (N_4310,In_1056,In_1188);
and U4311 (N_4311,In_434,In_949);
nand U4312 (N_4312,In_640,In_2475);
nor U4313 (N_4313,In_1603,In_2561);
or U4314 (N_4314,In_2783,In_1100);
and U4315 (N_4315,In_2849,In_866);
and U4316 (N_4316,In_111,In_1615);
and U4317 (N_4317,In_1154,In_1771);
nor U4318 (N_4318,In_2105,In_2630);
nor U4319 (N_4319,In_2540,In_1831);
nor U4320 (N_4320,In_1648,In_2261);
and U4321 (N_4321,In_2580,In_2714);
xor U4322 (N_4322,In_839,In_935);
nand U4323 (N_4323,In_2659,In_852);
or U4324 (N_4324,In_4,In_1865);
and U4325 (N_4325,In_468,In_2000);
nor U4326 (N_4326,In_2675,In_455);
or U4327 (N_4327,In_2008,In_732);
nand U4328 (N_4328,In_241,In_1514);
and U4329 (N_4329,In_1907,In_2859);
and U4330 (N_4330,In_936,In_237);
xor U4331 (N_4331,In_882,In_1465);
nor U4332 (N_4332,In_1450,In_823);
or U4333 (N_4333,In_2661,In_2178);
xnor U4334 (N_4334,In_387,In_201);
nand U4335 (N_4335,In_1504,In_727);
nand U4336 (N_4336,In_48,In_107);
nor U4337 (N_4337,In_715,In_1744);
nor U4338 (N_4338,In_217,In_708);
or U4339 (N_4339,In_1366,In_2586);
and U4340 (N_4340,In_2392,In_2999);
and U4341 (N_4341,In_1203,In_203);
nand U4342 (N_4342,In_1089,In_1262);
nor U4343 (N_4343,In_1134,In_2025);
and U4344 (N_4344,In_2327,In_2877);
nand U4345 (N_4345,In_1010,In_62);
xor U4346 (N_4346,In_2167,In_244);
or U4347 (N_4347,In_2784,In_1857);
and U4348 (N_4348,In_1492,In_1463);
nand U4349 (N_4349,In_749,In_1132);
xnor U4350 (N_4350,In_747,In_314);
or U4351 (N_4351,In_464,In_17);
xor U4352 (N_4352,In_2304,In_2327);
nand U4353 (N_4353,In_70,In_2596);
or U4354 (N_4354,In_528,In_1031);
nand U4355 (N_4355,In_1134,In_1336);
nor U4356 (N_4356,In_272,In_1546);
or U4357 (N_4357,In_337,In_1707);
or U4358 (N_4358,In_2798,In_1983);
and U4359 (N_4359,In_1061,In_841);
nor U4360 (N_4360,In_1874,In_834);
xor U4361 (N_4361,In_64,In_958);
and U4362 (N_4362,In_438,In_85);
and U4363 (N_4363,In_1935,In_2621);
xor U4364 (N_4364,In_171,In_2181);
nor U4365 (N_4365,In_1241,In_443);
nand U4366 (N_4366,In_1943,In_1808);
and U4367 (N_4367,In_2194,In_2787);
or U4368 (N_4368,In_51,In_1269);
xnor U4369 (N_4369,In_1849,In_2147);
nor U4370 (N_4370,In_976,In_1847);
nor U4371 (N_4371,In_12,In_758);
and U4372 (N_4372,In_937,In_2394);
nor U4373 (N_4373,In_2022,In_1337);
nor U4374 (N_4374,In_956,In_49);
nand U4375 (N_4375,In_1462,In_816);
nand U4376 (N_4376,In_1996,In_1020);
nand U4377 (N_4377,In_2977,In_1964);
nor U4378 (N_4378,In_589,In_1976);
nor U4379 (N_4379,In_1045,In_193);
and U4380 (N_4380,In_2290,In_2121);
and U4381 (N_4381,In_2883,In_2892);
and U4382 (N_4382,In_1999,In_2114);
nor U4383 (N_4383,In_1792,In_2663);
nor U4384 (N_4384,In_1761,In_207);
nand U4385 (N_4385,In_1620,In_1034);
xnor U4386 (N_4386,In_1988,In_2820);
nand U4387 (N_4387,In_2425,In_2137);
nand U4388 (N_4388,In_742,In_2538);
and U4389 (N_4389,In_950,In_1313);
or U4390 (N_4390,In_1445,In_2898);
nor U4391 (N_4391,In_747,In_2186);
nor U4392 (N_4392,In_1873,In_1998);
nand U4393 (N_4393,In_2240,In_346);
nor U4394 (N_4394,In_530,In_1079);
nand U4395 (N_4395,In_902,In_2802);
and U4396 (N_4396,In_2195,In_1349);
or U4397 (N_4397,In_2895,In_2988);
nand U4398 (N_4398,In_2371,In_2395);
nand U4399 (N_4399,In_413,In_2050);
nand U4400 (N_4400,In_2154,In_1480);
nand U4401 (N_4401,In_1011,In_1809);
or U4402 (N_4402,In_1617,In_2504);
nand U4403 (N_4403,In_2887,In_1144);
nor U4404 (N_4404,In_1446,In_858);
or U4405 (N_4405,In_2759,In_339);
and U4406 (N_4406,In_1288,In_1985);
nor U4407 (N_4407,In_2521,In_1027);
and U4408 (N_4408,In_314,In_2492);
or U4409 (N_4409,In_827,In_879);
and U4410 (N_4410,In_2248,In_1980);
and U4411 (N_4411,In_2417,In_1757);
or U4412 (N_4412,In_989,In_1462);
and U4413 (N_4413,In_342,In_436);
nor U4414 (N_4414,In_1780,In_936);
or U4415 (N_4415,In_2969,In_1594);
and U4416 (N_4416,In_2629,In_1675);
nand U4417 (N_4417,In_1290,In_61);
nand U4418 (N_4418,In_2425,In_342);
xnor U4419 (N_4419,In_988,In_2198);
nor U4420 (N_4420,In_1763,In_2154);
nor U4421 (N_4421,In_1715,In_1893);
or U4422 (N_4422,In_1154,In_1167);
or U4423 (N_4423,In_2230,In_1614);
or U4424 (N_4424,In_1500,In_2750);
nor U4425 (N_4425,In_817,In_1396);
xnor U4426 (N_4426,In_1736,In_2729);
xor U4427 (N_4427,In_2248,In_2685);
xor U4428 (N_4428,In_2415,In_2570);
nand U4429 (N_4429,In_517,In_1805);
nor U4430 (N_4430,In_994,In_2774);
and U4431 (N_4431,In_930,In_1676);
nor U4432 (N_4432,In_1512,In_2798);
nor U4433 (N_4433,In_2390,In_934);
or U4434 (N_4434,In_2457,In_1922);
nand U4435 (N_4435,In_796,In_1841);
xor U4436 (N_4436,In_2915,In_1386);
nand U4437 (N_4437,In_13,In_1923);
or U4438 (N_4438,In_1973,In_302);
nand U4439 (N_4439,In_2754,In_1472);
nand U4440 (N_4440,In_812,In_296);
nand U4441 (N_4441,In_2913,In_1588);
and U4442 (N_4442,In_1010,In_2428);
nor U4443 (N_4443,In_901,In_480);
nor U4444 (N_4444,In_2482,In_2797);
and U4445 (N_4445,In_992,In_1464);
nor U4446 (N_4446,In_1812,In_1922);
or U4447 (N_4447,In_858,In_1735);
nor U4448 (N_4448,In_171,In_1230);
nor U4449 (N_4449,In_2883,In_1577);
nand U4450 (N_4450,In_1115,In_915);
nand U4451 (N_4451,In_1046,In_1701);
nor U4452 (N_4452,In_1352,In_2010);
and U4453 (N_4453,In_2209,In_2046);
nor U4454 (N_4454,In_1220,In_1400);
or U4455 (N_4455,In_2228,In_1007);
nand U4456 (N_4456,In_2532,In_2593);
or U4457 (N_4457,In_1807,In_649);
nand U4458 (N_4458,In_125,In_1036);
or U4459 (N_4459,In_1852,In_955);
and U4460 (N_4460,In_1824,In_2721);
nor U4461 (N_4461,In_874,In_2678);
nand U4462 (N_4462,In_390,In_1454);
nand U4463 (N_4463,In_1650,In_1633);
nand U4464 (N_4464,In_2442,In_1015);
or U4465 (N_4465,In_2370,In_1929);
or U4466 (N_4466,In_1882,In_2456);
or U4467 (N_4467,In_2552,In_1884);
or U4468 (N_4468,In_2987,In_2036);
xnor U4469 (N_4469,In_2435,In_1104);
nor U4470 (N_4470,In_476,In_1860);
or U4471 (N_4471,In_1697,In_103);
or U4472 (N_4472,In_1352,In_328);
or U4473 (N_4473,In_1055,In_387);
nand U4474 (N_4474,In_2978,In_914);
nor U4475 (N_4475,In_2782,In_571);
and U4476 (N_4476,In_1441,In_288);
nand U4477 (N_4477,In_2887,In_1884);
or U4478 (N_4478,In_959,In_2440);
xor U4479 (N_4479,In_2269,In_2581);
nand U4480 (N_4480,In_2890,In_1803);
nand U4481 (N_4481,In_2228,In_2542);
or U4482 (N_4482,In_187,In_2050);
nand U4483 (N_4483,In_1763,In_802);
xnor U4484 (N_4484,In_670,In_475);
nand U4485 (N_4485,In_1388,In_2357);
and U4486 (N_4486,In_1367,In_2508);
or U4487 (N_4487,In_1448,In_2139);
nand U4488 (N_4488,In_121,In_2315);
nor U4489 (N_4489,In_2540,In_1388);
xnor U4490 (N_4490,In_2126,In_1980);
and U4491 (N_4491,In_1298,In_2714);
and U4492 (N_4492,In_617,In_2691);
or U4493 (N_4493,In_1106,In_2480);
and U4494 (N_4494,In_419,In_1859);
nand U4495 (N_4495,In_2103,In_1601);
or U4496 (N_4496,In_1337,In_413);
nor U4497 (N_4497,In_2302,In_415);
nand U4498 (N_4498,In_2935,In_1569);
and U4499 (N_4499,In_789,In_2651);
or U4500 (N_4500,In_317,In_697);
and U4501 (N_4501,In_109,In_1607);
or U4502 (N_4502,In_238,In_548);
nand U4503 (N_4503,In_2338,In_2108);
nor U4504 (N_4504,In_648,In_2026);
or U4505 (N_4505,In_1211,In_2751);
or U4506 (N_4506,In_158,In_2725);
nor U4507 (N_4507,In_2318,In_2649);
or U4508 (N_4508,In_2342,In_917);
and U4509 (N_4509,In_1918,In_2757);
and U4510 (N_4510,In_2399,In_2212);
nand U4511 (N_4511,In_1473,In_10);
nand U4512 (N_4512,In_1737,In_2048);
nor U4513 (N_4513,In_1343,In_492);
and U4514 (N_4514,In_1650,In_2186);
nand U4515 (N_4515,In_2097,In_1156);
nand U4516 (N_4516,In_288,In_1326);
nor U4517 (N_4517,In_18,In_1382);
and U4518 (N_4518,In_2116,In_2258);
nor U4519 (N_4519,In_1847,In_2695);
or U4520 (N_4520,In_1666,In_1296);
nand U4521 (N_4521,In_1044,In_2470);
nor U4522 (N_4522,In_1465,In_1401);
nor U4523 (N_4523,In_2225,In_1461);
or U4524 (N_4524,In_2912,In_1727);
xnor U4525 (N_4525,In_632,In_1715);
nand U4526 (N_4526,In_1271,In_2516);
or U4527 (N_4527,In_780,In_347);
or U4528 (N_4528,In_589,In_2775);
or U4529 (N_4529,In_1351,In_4);
xor U4530 (N_4530,In_2526,In_456);
nand U4531 (N_4531,In_728,In_1001);
nor U4532 (N_4532,In_1868,In_2349);
nand U4533 (N_4533,In_2323,In_1122);
nor U4534 (N_4534,In_1545,In_2837);
nand U4535 (N_4535,In_2000,In_2523);
nor U4536 (N_4536,In_2463,In_1082);
nor U4537 (N_4537,In_311,In_1504);
nor U4538 (N_4538,In_988,In_372);
xor U4539 (N_4539,In_923,In_2832);
xnor U4540 (N_4540,In_2526,In_2911);
or U4541 (N_4541,In_544,In_2437);
or U4542 (N_4542,In_1497,In_2455);
xor U4543 (N_4543,In_2561,In_1189);
and U4544 (N_4544,In_1511,In_2566);
nor U4545 (N_4545,In_541,In_2786);
nand U4546 (N_4546,In_1593,In_2142);
and U4547 (N_4547,In_1353,In_134);
nor U4548 (N_4548,In_1607,In_439);
or U4549 (N_4549,In_2939,In_1519);
and U4550 (N_4550,In_1984,In_119);
nand U4551 (N_4551,In_258,In_1789);
nor U4552 (N_4552,In_1611,In_241);
nand U4553 (N_4553,In_87,In_428);
nand U4554 (N_4554,In_1417,In_858);
nand U4555 (N_4555,In_619,In_896);
nand U4556 (N_4556,In_2078,In_1351);
and U4557 (N_4557,In_2639,In_2203);
nor U4558 (N_4558,In_1899,In_2136);
and U4559 (N_4559,In_2583,In_2946);
and U4560 (N_4560,In_2794,In_2346);
and U4561 (N_4561,In_1849,In_1635);
or U4562 (N_4562,In_2969,In_507);
nand U4563 (N_4563,In_2525,In_690);
nor U4564 (N_4564,In_1745,In_1604);
xor U4565 (N_4565,In_2103,In_2423);
and U4566 (N_4566,In_2304,In_2975);
or U4567 (N_4567,In_2834,In_2962);
nand U4568 (N_4568,In_777,In_241);
and U4569 (N_4569,In_2791,In_282);
nand U4570 (N_4570,In_1665,In_200);
and U4571 (N_4571,In_2857,In_1434);
or U4572 (N_4572,In_2203,In_2783);
nor U4573 (N_4573,In_135,In_546);
or U4574 (N_4574,In_1858,In_1197);
xor U4575 (N_4575,In_319,In_2641);
nor U4576 (N_4576,In_2660,In_2773);
xnor U4577 (N_4577,In_2468,In_2760);
nor U4578 (N_4578,In_2628,In_208);
xnor U4579 (N_4579,In_1300,In_727);
nand U4580 (N_4580,In_1818,In_821);
or U4581 (N_4581,In_292,In_1534);
xor U4582 (N_4582,In_1190,In_2609);
and U4583 (N_4583,In_2100,In_664);
nand U4584 (N_4584,In_2118,In_233);
nand U4585 (N_4585,In_2865,In_1216);
and U4586 (N_4586,In_2750,In_710);
xnor U4587 (N_4587,In_655,In_1360);
xor U4588 (N_4588,In_2357,In_2795);
and U4589 (N_4589,In_1333,In_1095);
nand U4590 (N_4590,In_1217,In_1773);
nand U4591 (N_4591,In_1673,In_1649);
nand U4592 (N_4592,In_2731,In_368);
and U4593 (N_4593,In_1102,In_2184);
nor U4594 (N_4594,In_752,In_953);
and U4595 (N_4595,In_1519,In_2991);
nand U4596 (N_4596,In_1427,In_869);
and U4597 (N_4597,In_1746,In_959);
or U4598 (N_4598,In_2207,In_2479);
or U4599 (N_4599,In_2586,In_2649);
and U4600 (N_4600,In_2063,In_2410);
and U4601 (N_4601,In_1870,In_1903);
and U4602 (N_4602,In_271,In_2980);
and U4603 (N_4603,In_2596,In_251);
nand U4604 (N_4604,In_888,In_228);
and U4605 (N_4605,In_930,In_2132);
xnor U4606 (N_4606,In_1990,In_1390);
and U4607 (N_4607,In_2614,In_1439);
or U4608 (N_4608,In_1364,In_222);
nor U4609 (N_4609,In_2274,In_80);
or U4610 (N_4610,In_682,In_1810);
nand U4611 (N_4611,In_774,In_887);
or U4612 (N_4612,In_2985,In_2147);
and U4613 (N_4613,In_1870,In_2662);
xnor U4614 (N_4614,In_1521,In_1402);
and U4615 (N_4615,In_2766,In_1905);
or U4616 (N_4616,In_1728,In_1983);
nand U4617 (N_4617,In_1538,In_2588);
and U4618 (N_4618,In_2217,In_1636);
or U4619 (N_4619,In_2321,In_598);
nor U4620 (N_4620,In_2427,In_2475);
and U4621 (N_4621,In_1427,In_1606);
nor U4622 (N_4622,In_55,In_622);
nand U4623 (N_4623,In_2973,In_1480);
nand U4624 (N_4624,In_354,In_420);
and U4625 (N_4625,In_2839,In_1841);
or U4626 (N_4626,In_1543,In_119);
nor U4627 (N_4627,In_1459,In_1198);
nand U4628 (N_4628,In_1145,In_1906);
nand U4629 (N_4629,In_1048,In_1691);
nor U4630 (N_4630,In_2998,In_1663);
or U4631 (N_4631,In_392,In_1784);
and U4632 (N_4632,In_2734,In_2818);
or U4633 (N_4633,In_1251,In_398);
and U4634 (N_4634,In_1763,In_1374);
nand U4635 (N_4635,In_1992,In_1143);
or U4636 (N_4636,In_11,In_1586);
nand U4637 (N_4637,In_2184,In_1197);
nand U4638 (N_4638,In_1432,In_1987);
nand U4639 (N_4639,In_1701,In_2945);
or U4640 (N_4640,In_1695,In_165);
and U4641 (N_4641,In_955,In_1264);
or U4642 (N_4642,In_246,In_374);
xnor U4643 (N_4643,In_560,In_1960);
nor U4644 (N_4644,In_2294,In_620);
nor U4645 (N_4645,In_2425,In_2055);
or U4646 (N_4646,In_1851,In_764);
or U4647 (N_4647,In_1695,In_421);
or U4648 (N_4648,In_1359,In_2492);
nor U4649 (N_4649,In_632,In_304);
or U4650 (N_4650,In_1234,In_2706);
and U4651 (N_4651,In_988,In_2335);
nor U4652 (N_4652,In_1413,In_2088);
nor U4653 (N_4653,In_2421,In_2811);
nor U4654 (N_4654,In_2963,In_1403);
and U4655 (N_4655,In_2391,In_1711);
and U4656 (N_4656,In_989,In_382);
nor U4657 (N_4657,In_318,In_734);
nor U4658 (N_4658,In_2311,In_2599);
or U4659 (N_4659,In_198,In_964);
nor U4660 (N_4660,In_166,In_1667);
nand U4661 (N_4661,In_2995,In_1186);
nor U4662 (N_4662,In_546,In_2562);
nor U4663 (N_4663,In_2310,In_2545);
nand U4664 (N_4664,In_302,In_1448);
xnor U4665 (N_4665,In_2034,In_2089);
or U4666 (N_4666,In_121,In_2032);
nand U4667 (N_4667,In_1104,In_1016);
and U4668 (N_4668,In_2727,In_780);
or U4669 (N_4669,In_2327,In_1099);
nor U4670 (N_4670,In_1677,In_1112);
or U4671 (N_4671,In_457,In_15);
xnor U4672 (N_4672,In_2224,In_2934);
nor U4673 (N_4673,In_1968,In_124);
and U4674 (N_4674,In_1845,In_2735);
and U4675 (N_4675,In_2218,In_1069);
or U4676 (N_4676,In_2089,In_640);
or U4677 (N_4677,In_338,In_1142);
and U4678 (N_4678,In_1238,In_2711);
nor U4679 (N_4679,In_1409,In_1251);
xor U4680 (N_4680,In_233,In_108);
xnor U4681 (N_4681,In_953,In_2570);
nand U4682 (N_4682,In_689,In_1630);
xnor U4683 (N_4683,In_2366,In_903);
or U4684 (N_4684,In_2280,In_2967);
or U4685 (N_4685,In_319,In_2731);
nand U4686 (N_4686,In_1700,In_743);
nor U4687 (N_4687,In_1857,In_2377);
nand U4688 (N_4688,In_527,In_95);
and U4689 (N_4689,In_2900,In_2519);
nor U4690 (N_4690,In_1144,In_298);
or U4691 (N_4691,In_1428,In_2204);
nand U4692 (N_4692,In_1794,In_1881);
nand U4693 (N_4693,In_1047,In_2707);
nand U4694 (N_4694,In_2927,In_478);
and U4695 (N_4695,In_891,In_286);
nand U4696 (N_4696,In_1261,In_918);
and U4697 (N_4697,In_2108,In_1368);
and U4698 (N_4698,In_1240,In_1387);
and U4699 (N_4699,In_1510,In_265);
nand U4700 (N_4700,In_678,In_1265);
xnor U4701 (N_4701,In_1717,In_624);
nand U4702 (N_4702,In_249,In_612);
nor U4703 (N_4703,In_28,In_1485);
nor U4704 (N_4704,In_482,In_2246);
nand U4705 (N_4705,In_1594,In_1098);
xnor U4706 (N_4706,In_2121,In_1909);
and U4707 (N_4707,In_2980,In_2428);
or U4708 (N_4708,In_1632,In_2386);
or U4709 (N_4709,In_2495,In_981);
nor U4710 (N_4710,In_2407,In_1292);
nand U4711 (N_4711,In_2092,In_1909);
or U4712 (N_4712,In_1709,In_1585);
nor U4713 (N_4713,In_2899,In_1404);
xor U4714 (N_4714,In_1798,In_1700);
or U4715 (N_4715,In_2031,In_2105);
nand U4716 (N_4716,In_400,In_453);
and U4717 (N_4717,In_2470,In_2304);
nand U4718 (N_4718,In_757,In_812);
or U4719 (N_4719,In_119,In_2410);
nor U4720 (N_4720,In_1396,In_553);
nand U4721 (N_4721,In_2593,In_997);
xnor U4722 (N_4722,In_1578,In_1471);
or U4723 (N_4723,In_2148,In_1416);
nand U4724 (N_4724,In_1491,In_54);
nor U4725 (N_4725,In_1502,In_1458);
or U4726 (N_4726,In_597,In_2536);
nor U4727 (N_4727,In_40,In_1433);
nor U4728 (N_4728,In_2422,In_443);
nand U4729 (N_4729,In_732,In_423);
or U4730 (N_4730,In_246,In_2535);
or U4731 (N_4731,In_2326,In_2718);
or U4732 (N_4732,In_1682,In_1445);
nor U4733 (N_4733,In_645,In_597);
nand U4734 (N_4734,In_494,In_2454);
nor U4735 (N_4735,In_2215,In_2127);
nand U4736 (N_4736,In_2191,In_1886);
or U4737 (N_4737,In_1803,In_412);
nand U4738 (N_4738,In_1771,In_2862);
nor U4739 (N_4739,In_1562,In_2464);
and U4740 (N_4740,In_811,In_16);
xor U4741 (N_4741,In_2794,In_558);
nor U4742 (N_4742,In_399,In_576);
nor U4743 (N_4743,In_2696,In_1953);
nor U4744 (N_4744,In_940,In_123);
nor U4745 (N_4745,In_2714,In_1008);
xor U4746 (N_4746,In_1745,In_367);
nand U4747 (N_4747,In_573,In_1420);
or U4748 (N_4748,In_955,In_840);
and U4749 (N_4749,In_1507,In_2135);
xor U4750 (N_4750,In_2405,In_2851);
nor U4751 (N_4751,In_1271,In_2948);
and U4752 (N_4752,In_42,In_1740);
nor U4753 (N_4753,In_2043,In_2298);
nor U4754 (N_4754,In_1881,In_912);
nor U4755 (N_4755,In_2353,In_1490);
and U4756 (N_4756,In_1967,In_643);
or U4757 (N_4757,In_2322,In_2656);
and U4758 (N_4758,In_1062,In_1692);
and U4759 (N_4759,In_2317,In_2040);
or U4760 (N_4760,In_2081,In_58);
or U4761 (N_4761,In_2732,In_367);
or U4762 (N_4762,In_798,In_1662);
nor U4763 (N_4763,In_2008,In_235);
nand U4764 (N_4764,In_945,In_1249);
xor U4765 (N_4765,In_721,In_1844);
and U4766 (N_4766,In_2468,In_1158);
and U4767 (N_4767,In_2467,In_2935);
and U4768 (N_4768,In_747,In_1880);
or U4769 (N_4769,In_2550,In_1083);
and U4770 (N_4770,In_2994,In_852);
or U4771 (N_4771,In_2361,In_2359);
nand U4772 (N_4772,In_1589,In_2891);
xnor U4773 (N_4773,In_0,In_564);
nor U4774 (N_4774,In_290,In_1522);
nor U4775 (N_4775,In_339,In_1083);
nor U4776 (N_4776,In_1105,In_709);
nand U4777 (N_4777,In_2707,In_336);
nor U4778 (N_4778,In_1475,In_2848);
or U4779 (N_4779,In_569,In_179);
nor U4780 (N_4780,In_1401,In_1199);
or U4781 (N_4781,In_1151,In_2840);
nand U4782 (N_4782,In_850,In_1398);
or U4783 (N_4783,In_1077,In_2328);
nand U4784 (N_4784,In_2598,In_788);
and U4785 (N_4785,In_2272,In_2777);
or U4786 (N_4786,In_2940,In_2655);
xor U4787 (N_4787,In_2188,In_1776);
xnor U4788 (N_4788,In_557,In_770);
nor U4789 (N_4789,In_126,In_2327);
or U4790 (N_4790,In_2745,In_1863);
nor U4791 (N_4791,In_2853,In_2913);
nor U4792 (N_4792,In_786,In_1461);
nand U4793 (N_4793,In_2267,In_109);
and U4794 (N_4794,In_2771,In_980);
xnor U4795 (N_4795,In_2888,In_2974);
or U4796 (N_4796,In_2566,In_1948);
xnor U4797 (N_4797,In_1993,In_1199);
and U4798 (N_4798,In_1908,In_2777);
and U4799 (N_4799,In_1009,In_892);
or U4800 (N_4800,In_2917,In_2822);
nor U4801 (N_4801,In_1458,In_1641);
and U4802 (N_4802,In_1461,In_2642);
and U4803 (N_4803,In_2138,In_743);
nand U4804 (N_4804,In_1166,In_1690);
nor U4805 (N_4805,In_2699,In_257);
nand U4806 (N_4806,In_1557,In_1311);
or U4807 (N_4807,In_2319,In_2976);
and U4808 (N_4808,In_880,In_680);
nor U4809 (N_4809,In_2651,In_1722);
nand U4810 (N_4810,In_267,In_2763);
nand U4811 (N_4811,In_1773,In_2337);
and U4812 (N_4812,In_2635,In_1782);
nor U4813 (N_4813,In_206,In_662);
and U4814 (N_4814,In_1640,In_1162);
nand U4815 (N_4815,In_688,In_1629);
or U4816 (N_4816,In_1163,In_2195);
and U4817 (N_4817,In_159,In_1395);
and U4818 (N_4818,In_2186,In_2061);
nor U4819 (N_4819,In_824,In_1053);
nand U4820 (N_4820,In_929,In_2302);
nor U4821 (N_4821,In_2853,In_1453);
or U4822 (N_4822,In_1838,In_1812);
xor U4823 (N_4823,In_868,In_1395);
or U4824 (N_4824,In_2288,In_2417);
and U4825 (N_4825,In_205,In_2430);
nor U4826 (N_4826,In_2453,In_816);
xnor U4827 (N_4827,In_1694,In_786);
and U4828 (N_4828,In_1895,In_2857);
and U4829 (N_4829,In_502,In_2060);
nand U4830 (N_4830,In_2397,In_1263);
or U4831 (N_4831,In_1613,In_477);
nand U4832 (N_4832,In_2172,In_348);
nor U4833 (N_4833,In_1022,In_2359);
nand U4834 (N_4834,In_2671,In_428);
nand U4835 (N_4835,In_1158,In_988);
nand U4836 (N_4836,In_53,In_2965);
xnor U4837 (N_4837,In_1984,In_1717);
nand U4838 (N_4838,In_599,In_318);
nand U4839 (N_4839,In_677,In_1675);
and U4840 (N_4840,In_1339,In_2149);
or U4841 (N_4841,In_1917,In_2180);
nor U4842 (N_4842,In_2467,In_1905);
nand U4843 (N_4843,In_1716,In_1678);
or U4844 (N_4844,In_1837,In_1709);
nand U4845 (N_4845,In_709,In_1606);
nand U4846 (N_4846,In_909,In_2882);
nor U4847 (N_4847,In_2497,In_255);
nor U4848 (N_4848,In_1895,In_2913);
nor U4849 (N_4849,In_1185,In_1793);
xor U4850 (N_4850,In_823,In_1287);
or U4851 (N_4851,In_1758,In_2905);
xor U4852 (N_4852,In_2878,In_1022);
nand U4853 (N_4853,In_1043,In_1837);
nand U4854 (N_4854,In_1571,In_862);
and U4855 (N_4855,In_567,In_2925);
or U4856 (N_4856,In_1882,In_1058);
nand U4857 (N_4857,In_2391,In_1885);
or U4858 (N_4858,In_743,In_2160);
nor U4859 (N_4859,In_1640,In_556);
nor U4860 (N_4860,In_2568,In_1589);
or U4861 (N_4861,In_2236,In_541);
or U4862 (N_4862,In_2312,In_2260);
nor U4863 (N_4863,In_381,In_2612);
nand U4864 (N_4864,In_1962,In_1884);
and U4865 (N_4865,In_1312,In_2074);
xor U4866 (N_4866,In_614,In_810);
xor U4867 (N_4867,In_1973,In_1589);
or U4868 (N_4868,In_2472,In_362);
nor U4869 (N_4869,In_913,In_1581);
xnor U4870 (N_4870,In_2435,In_953);
nor U4871 (N_4871,In_2168,In_2928);
and U4872 (N_4872,In_2032,In_1031);
nand U4873 (N_4873,In_1454,In_259);
xnor U4874 (N_4874,In_669,In_1472);
and U4875 (N_4875,In_1133,In_1835);
and U4876 (N_4876,In_2329,In_817);
nand U4877 (N_4877,In_2737,In_2801);
or U4878 (N_4878,In_1927,In_341);
or U4879 (N_4879,In_1758,In_259);
nand U4880 (N_4880,In_2914,In_65);
and U4881 (N_4881,In_396,In_1596);
and U4882 (N_4882,In_61,In_2997);
nand U4883 (N_4883,In_1469,In_2356);
nand U4884 (N_4884,In_2402,In_2463);
or U4885 (N_4885,In_431,In_2101);
and U4886 (N_4886,In_1416,In_1938);
and U4887 (N_4887,In_2034,In_2540);
or U4888 (N_4888,In_1582,In_2468);
nand U4889 (N_4889,In_196,In_1543);
nor U4890 (N_4890,In_548,In_1346);
and U4891 (N_4891,In_1655,In_1047);
or U4892 (N_4892,In_1006,In_2666);
xnor U4893 (N_4893,In_110,In_1119);
and U4894 (N_4894,In_1421,In_1448);
and U4895 (N_4895,In_748,In_2975);
nand U4896 (N_4896,In_1919,In_692);
or U4897 (N_4897,In_2656,In_2924);
nand U4898 (N_4898,In_2915,In_1672);
nor U4899 (N_4899,In_1989,In_1631);
and U4900 (N_4900,In_2352,In_288);
nor U4901 (N_4901,In_1264,In_1420);
nor U4902 (N_4902,In_2553,In_2770);
nor U4903 (N_4903,In_2029,In_335);
nand U4904 (N_4904,In_1280,In_868);
nand U4905 (N_4905,In_2862,In_1953);
nor U4906 (N_4906,In_811,In_1020);
and U4907 (N_4907,In_1906,In_607);
nand U4908 (N_4908,In_2950,In_1999);
nor U4909 (N_4909,In_2557,In_388);
nand U4910 (N_4910,In_2185,In_2368);
nor U4911 (N_4911,In_1864,In_572);
nor U4912 (N_4912,In_2317,In_1554);
nor U4913 (N_4913,In_878,In_1957);
and U4914 (N_4914,In_2406,In_1889);
nor U4915 (N_4915,In_1156,In_1724);
and U4916 (N_4916,In_2318,In_720);
nand U4917 (N_4917,In_1115,In_1224);
and U4918 (N_4918,In_338,In_2617);
nand U4919 (N_4919,In_751,In_1534);
nand U4920 (N_4920,In_2010,In_849);
nand U4921 (N_4921,In_2757,In_1301);
nand U4922 (N_4922,In_1721,In_2617);
and U4923 (N_4923,In_904,In_230);
nor U4924 (N_4924,In_1543,In_1298);
nor U4925 (N_4925,In_795,In_1937);
nand U4926 (N_4926,In_1882,In_2532);
and U4927 (N_4927,In_1864,In_174);
nor U4928 (N_4928,In_2463,In_1563);
or U4929 (N_4929,In_500,In_1698);
and U4930 (N_4930,In_1199,In_840);
or U4931 (N_4931,In_1097,In_2758);
or U4932 (N_4932,In_2467,In_2963);
or U4933 (N_4933,In_939,In_1749);
and U4934 (N_4934,In_295,In_1367);
nand U4935 (N_4935,In_2239,In_745);
xnor U4936 (N_4936,In_2836,In_1989);
nand U4937 (N_4937,In_1666,In_950);
xor U4938 (N_4938,In_1527,In_1737);
or U4939 (N_4939,In_968,In_2016);
or U4940 (N_4940,In_2629,In_1905);
xnor U4941 (N_4941,In_1303,In_1741);
and U4942 (N_4942,In_1599,In_1062);
or U4943 (N_4943,In_2501,In_164);
or U4944 (N_4944,In_186,In_153);
or U4945 (N_4945,In_326,In_456);
nand U4946 (N_4946,In_1888,In_1681);
nor U4947 (N_4947,In_847,In_1296);
nor U4948 (N_4948,In_2171,In_175);
nand U4949 (N_4949,In_1364,In_2449);
nor U4950 (N_4950,In_956,In_72);
or U4951 (N_4951,In_2525,In_1480);
and U4952 (N_4952,In_2948,In_523);
nand U4953 (N_4953,In_2250,In_2840);
nand U4954 (N_4954,In_487,In_992);
nand U4955 (N_4955,In_55,In_1043);
and U4956 (N_4956,In_384,In_614);
or U4957 (N_4957,In_2420,In_2103);
xnor U4958 (N_4958,In_1189,In_2967);
nand U4959 (N_4959,In_2112,In_423);
or U4960 (N_4960,In_1194,In_1523);
or U4961 (N_4961,In_869,In_729);
nor U4962 (N_4962,In_1145,In_2974);
nor U4963 (N_4963,In_539,In_418);
xnor U4964 (N_4964,In_2962,In_2851);
or U4965 (N_4965,In_1678,In_1004);
nor U4966 (N_4966,In_2274,In_2727);
or U4967 (N_4967,In_2402,In_578);
nand U4968 (N_4968,In_666,In_638);
nor U4969 (N_4969,In_1088,In_361);
and U4970 (N_4970,In_2446,In_773);
or U4971 (N_4971,In_1961,In_2758);
nor U4972 (N_4972,In_2973,In_413);
nand U4973 (N_4973,In_1443,In_2770);
and U4974 (N_4974,In_661,In_2561);
xnor U4975 (N_4975,In_2375,In_394);
and U4976 (N_4976,In_1509,In_1921);
nand U4977 (N_4977,In_1523,In_34);
or U4978 (N_4978,In_59,In_391);
nor U4979 (N_4979,In_1720,In_358);
nand U4980 (N_4980,In_858,In_824);
xor U4981 (N_4981,In_219,In_1622);
or U4982 (N_4982,In_2628,In_1383);
xor U4983 (N_4983,In_2714,In_2997);
nor U4984 (N_4984,In_1939,In_1771);
and U4985 (N_4985,In_58,In_760);
or U4986 (N_4986,In_2910,In_2438);
nand U4987 (N_4987,In_2314,In_529);
or U4988 (N_4988,In_452,In_900);
and U4989 (N_4989,In_2636,In_1198);
xnor U4990 (N_4990,In_1123,In_994);
xor U4991 (N_4991,In_1526,In_1186);
and U4992 (N_4992,In_1306,In_2678);
nor U4993 (N_4993,In_2239,In_2915);
nand U4994 (N_4994,In_1720,In_441);
and U4995 (N_4995,In_515,In_1167);
nand U4996 (N_4996,In_476,In_2703);
nand U4997 (N_4997,In_1583,In_2538);
or U4998 (N_4998,In_573,In_2896);
nor U4999 (N_4999,In_1776,In_2611);
nand U5000 (N_5000,In_787,In_1436);
xor U5001 (N_5001,In_1127,In_822);
or U5002 (N_5002,In_200,In_1261);
nand U5003 (N_5003,In_2076,In_1090);
or U5004 (N_5004,In_998,In_2883);
nor U5005 (N_5005,In_804,In_2423);
nor U5006 (N_5006,In_1908,In_134);
nand U5007 (N_5007,In_615,In_1088);
or U5008 (N_5008,In_1526,In_2473);
and U5009 (N_5009,In_1265,In_1673);
nor U5010 (N_5010,In_671,In_1200);
or U5011 (N_5011,In_2212,In_190);
or U5012 (N_5012,In_1714,In_701);
or U5013 (N_5013,In_1899,In_1768);
or U5014 (N_5014,In_130,In_2417);
xor U5015 (N_5015,In_2851,In_1627);
xnor U5016 (N_5016,In_1808,In_845);
or U5017 (N_5017,In_1998,In_1193);
nor U5018 (N_5018,In_654,In_2058);
and U5019 (N_5019,In_2774,In_322);
nor U5020 (N_5020,In_1622,In_1833);
nor U5021 (N_5021,In_1401,In_2186);
or U5022 (N_5022,In_1267,In_795);
or U5023 (N_5023,In_1526,In_568);
xor U5024 (N_5024,In_407,In_258);
nand U5025 (N_5025,In_1414,In_403);
xnor U5026 (N_5026,In_2196,In_152);
xnor U5027 (N_5027,In_344,In_730);
or U5028 (N_5028,In_1408,In_370);
nand U5029 (N_5029,In_636,In_277);
or U5030 (N_5030,In_1032,In_1747);
or U5031 (N_5031,In_1315,In_2228);
nand U5032 (N_5032,In_2639,In_1444);
nand U5033 (N_5033,In_1354,In_2064);
or U5034 (N_5034,In_81,In_1790);
nand U5035 (N_5035,In_2132,In_1766);
nand U5036 (N_5036,In_1517,In_1748);
nor U5037 (N_5037,In_1556,In_1848);
and U5038 (N_5038,In_110,In_1160);
nand U5039 (N_5039,In_1317,In_2732);
and U5040 (N_5040,In_1339,In_582);
nand U5041 (N_5041,In_2172,In_2168);
nand U5042 (N_5042,In_1137,In_0);
nor U5043 (N_5043,In_1412,In_2540);
nor U5044 (N_5044,In_1684,In_183);
xor U5045 (N_5045,In_2174,In_935);
nor U5046 (N_5046,In_962,In_2248);
nor U5047 (N_5047,In_145,In_2080);
and U5048 (N_5048,In_1063,In_919);
nor U5049 (N_5049,In_2724,In_609);
nand U5050 (N_5050,In_1298,In_109);
xnor U5051 (N_5051,In_1226,In_2684);
and U5052 (N_5052,In_2331,In_2277);
nand U5053 (N_5053,In_330,In_338);
nand U5054 (N_5054,In_2642,In_1748);
nand U5055 (N_5055,In_2089,In_2816);
and U5056 (N_5056,In_1442,In_2347);
xor U5057 (N_5057,In_2446,In_2732);
or U5058 (N_5058,In_1167,In_2302);
nor U5059 (N_5059,In_2274,In_603);
xnor U5060 (N_5060,In_461,In_1303);
or U5061 (N_5061,In_576,In_109);
xor U5062 (N_5062,In_1720,In_1011);
nor U5063 (N_5063,In_1299,In_622);
and U5064 (N_5064,In_2524,In_1242);
xor U5065 (N_5065,In_1499,In_1855);
and U5066 (N_5066,In_1309,In_1524);
and U5067 (N_5067,In_1726,In_94);
and U5068 (N_5068,In_1899,In_77);
and U5069 (N_5069,In_1592,In_2156);
nor U5070 (N_5070,In_2802,In_1424);
xnor U5071 (N_5071,In_98,In_267);
or U5072 (N_5072,In_2245,In_1355);
or U5073 (N_5073,In_1406,In_2950);
nor U5074 (N_5074,In_980,In_623);
xnor U5075 (N_5075,In_2579,In_756);
xnor U5076 (N_5076,In_450,In_742);
or U5077 (N_5077,In_370,In_556);
or U5078 (N_5078,In_875,In_734);
or U5079 (N_5079,In_1779,In_2497);
nand U5080 (N_5080,In_1604,In_2654);
or U5081 (N_5081,In_320,In_587);
or U5082 (N_5082,In_1001,In_2723);
nor U5083 (N_5083,In_1741,In_1739);
nand U5084 (N_5084,In_815,In_2621);
or U5085 (N_5085,In_1618,In_637);
or U5086 (N_5086,In_1645,In_2979);
or U5087 (N_5087,In_2289,In_1162);
and U5088 (N_5088,In_2027,In_796);
or U5089 (N_5089,In_2796,In_1664);
or U5090 (N_5090,In_1775,In_269);
nand U5091 (N_5091,In_2514,In_1474);
or U5092 (N_5092,In_1412,In_1868);
nor U5093 (N_5093,In_2716,In_408);
or U5094 (N_5094,In_903,In_201);
or U5095 (N_5095,In_851,In_1822);
or U5096 (N_5096,In_590,In_1451);
and U5097 (N_5097,In_242,In_568);
nand U5098 (N_5098,In_550,In_1570);
and U5099 (N_5099,In_1592,In_2033);
nor U5100 (N_5100,In_2624,In_2269);
or U5101 (N_5101,In_894,In_1060);
nor U5102 (N_5102,In_890,In_2974);
nand U5103 (N_5103,In_542,In_1501);
nor U5104 (N_5104,In_711,In_1888);
and U5105 (N_5105,In_2597,In_1692);
nor U5106 (N_5106,In_2260,In_295);
nand U5107 (N_5107,In_1184,In_1941);
nor U5108 (N_5108,In_1229,In_697);
or U5109 (N_5109,In_698,In_2564);
or U5110 (N_5110,In_1763,In_44);
or U5111 (N_5111,In_899,In_252);
or U5112 (N_5112,In_2575,In_1064);
nor U5113 (N_5113,In_2071,In_1879);
or U5114 (N_5114,In_1528,In_1189);
nand U5115 (N_5115,In_1346,In_2570);
nand U5116 (N_5116,In_594,In_2218);
or U5117 (N_5117,In_2098,In_471);
or U5118 (N_5118,In_2025,In_589);
and U5119 (N_5119,In_1067,In_2816);
xor U5120 (N_5120,In_1626,In_1953);
or U5121 (N_5121,In_232,In_1876);
or U5122 (N_5122,In_1499,In_2182);
nor U5123 (N_5123,In_769,In_1387);
and U5124 (N_5124,In_2180,In_683);
nand U5125 (N_5125,In_1593,In_2985);
and U5126 (N_5126,In_1567,In_1399);
nor U5127 (N_5127,In_2001,In_1032);
nor U5128 (N_5128,In_1791,In_312);
and U5129 (N_5129,In_2245,In_2167);
nor U5130 (N_5130,In_2786,In_1018);
nor U5131 (N_5131,In_2666,In_1810);
xnor U5132 (N_5132,In_39,In_1645);
and U5133 (N_5133,In_2828,In_1167);
xnor U5134 (N_5134,In_1457,In_585);
and U5135 (N_5135,In_2560,In_1697);
nor U5136 (N_5136,In_2599,In_1744);
or U5137 (N_5137,In_2787,In_1711);
and U5138 (N_5138,In_2576,In_2173);
and U5139 (N_5139,In_55,In_1784);
and U5140 (N_5140,In_224,In_1480);
nand U5141 (N_5141,In_498,In_2515);
and U5142 (N_5142,In_450,In_2760);
and U5143 (N_5143,In_1115,In_2665);
xnor U5144 (N_5144,In_808,In_865);
or U5145 (N_5145,In_2814,In_2983);
nand U5146 (N_5146,In_2064,In_542);
nor U5147 (N_5147,In_238,In_1187);
nand U5148 (N_5148,In_410,In_37);
nor U5149 (N_5149,In_527,In_763);
or U5150 (N_5150,In_1434,In_1734);
nor U5151 (N_5151,In_35,In_1928);
nor U5152 (N_5152,In_62,In_57);
and U5153 (N_5153,In_292,In_1302);
or U5154 (N_5154,In_2759,In_604);
xor U5155 (N_5155,In_1655,In_2670);
xnor U5156 (N_5156,In_232,In_2692);
and U5157 (N_5157,In_296,In_2156);
and U5158 (N_5158,In_1735,In_1971);
xor U5159 (N_5159,In_688,In_963);
and U5160 (N_5160,In_816,In_730);
and U5161 (N_5161,In_1179,In_2736);
nand U5162 (N_5162,In_716,In_2714);
or U5163 (N_5163,In_418,In_2940);
nand U5164 (N_5164,In_1012,In_1896);
xor U5165 (N_5165,In_1087,In_2713);
nor U5166 (N_5166,In_2643,In_551);
nand U5167 (N_5167,In_1989,In_1525);
nor U5168 (N_5168,In_1287,In_2374);
and U5169 (N_5169,In_839,In_535);
nor U5170 (N_5170,In_1702,In_589);
and U5171 (N_5171,In_2741,In_1123);
nor U5172 (N_5172,In_2858,In_2197);
nor U5173 (N_5173,In_1575,In_2753);
or U5174 (N_5174,In_1778,In_2972);
and U5175 (N_5175,In_2991,In_443);
nand U5176 (N_5176,In_2738,In_1946);
nand U5177 (N_5177,In_2047,In_225);
and U5178 (N_5178,In_1481,In_2402);
nor U5179 (N_5179,In_1531,In_1497);
xnor U5180 (N_5180,In_1224,In_1648);
or U5181 (N_5181,In_463,In_1114);
or U5182 (N_5182,In_2415,In_929);
and U5183 (N_5183,In_2950,In_246);
nand U5184 (N_5184,In_1613,In_2409);
or U5185 (N_5185,In_1076,In_2316);
or U5186 (N_5186,In_859,In_832);
nor U5187 (N_5187,In_2983,In_1328);
nor U5188 (N_5188,In_339,In_2072);
or U5189 (N_5189,In_1145,In_1637);
nor U5190 (N_5190,In_1566,In_428);
nor U5191 (N_5191,In_1509,In_2875);
or U5192 (N_5192,In_499,In_1407);
or U5193 (N_5193,In_1959,In_509);
nand U5194 (N_5194,In_1470,In_1997);
xor U5195 (N_5195,In_4,In_1620);
nor U5196 (N_5196,In_2511,In_916);
and U5197 (N_5197,In_2187,In_2026);
nor U5198 (N_5198,In_2993,In_2055);
xor U5199 (N_5199,In_1470,In_1958);
and U5200 (N_5200,In_1897,In_1554);
nor U5201 (N_5201,In_2792,In_1693);
and U5202 (N_5202,In_2501,In_2175);
or U5203 (N_5203,In_1529,In_1730);
and U5204 (N_5204,In_276,In_2226);
nor U5205 (N_5205,In_1256,In_154);
nor U5206 (N_5206,In_2643,In_1504);
nand U5207 (N_5207,In_2132,In_632);
nand U5208 (N_5208,In_1936,In_926);
and U5209 (N_5209,In_124,In_1191);
nand U5210 (N_5210,In_1831,In_2997);
or U5211 (N_5211,In_847,In_1739);
nor U5212 (N_5212,In_764,In_988);
nand U5213 (N_5213,In_240,In_1242);
xnor U5214 (N_5214,In_2868,In_2915);
nor U5215 (N_5215,In_1466,In_1870);
nand U5216 (N_5216,In_1487,In_122);
nand U5217 (N_5217,In_2468,In_2197);
nor U5218 (N_5218,In_2907,In_2641);
and U5219 (N_5219,In_1169,In_2098);
nand U5220 (N_5220,In_337,In_1398);
nor U5221 (N_5221,In_2481,In_1183);
nand U5222 (N_5222,In_1807,In_399);
and U5223 (N_5223,In_2248,In_1781);
or U5224 (N_5224,In_873,In_1174);
or U5225 (N_5225,In_2228,In_1029);
or U5226 (N_5226,In_1010,In_1969);
xnor U5227 (N_5227,In_375,In_1835);
nand U5228 (N_5228,In_2603,In_733);
xnor U5229 (N_5229,In_2906,In_1257);
or U5230 (N_5230,In_2175,In_263);
nor U5231 (N_5231,In_2264,In_2430);
or U5232 (N_5232,In_240,In_1311);
or U5233 (N_5233,In_661,In_2315);
and U5234 (N_5234,In_556,In_548);
or U5235 (N_5235,In_1662,In_1993);
xnor U5236 (N_5236,In_2143,In_2109);
nand U5237 (N_5237,In_1698,In_2065);
nor U5238 (N_5238,In_1776,In_365);
or U5239 (N_5239,In_705,In_1365);
or U5240 (N_5240,In_435,In_518);
nand U5241 (N_5241,In_828,In_2617);
nand U5242 (N_5242,In_2033,In_986);
and U5243 (N_5243,In_595,In_495);
and U5244 (N_5244,In_329,In_550);
nand U5245 (N_5245,In_2857,In_46);
nor U5246 (N_5246,In_2781,In_2585);
nor U5247 (N_5247,In_144,In_2895);
xor U5248 (N_5248,In_1374,In_558);
nor U5249 (N_5249,In_1440,In_1516);
or U5250 (N_5250,In_2584,In_833);
and U5251 (N_5251,In_1406,In_794);
nand U5252 (N_5252,In_2969,In_654);
nor U5253 (N_5253,In_1642,In_2130);
and U5254 (N_5254,In_1388,In_2553);
and U5255 (N_5255,In_2239,In_2570);
or U5256 (N_5256,In_887,In_2991);
xnor U5257 (N_5257,In_1980,In_1441);
and U5258 (N_5258,In_1682,In_2479);
or U5259 (N_5259,In_2858,In_1620);
and U5260 (N_5260,In_1857,In_1467);
xnor U5261 (N_5261,In_1706,In_1929);
nand U5262 (N_5262,In_1756,In_668);
or U5263 (N_5263,In_626,In_2390);
nor U5264 (N_5264,In_141,In_1206);
or U5265 (N_5265,In_183,In_2971);
nand U5266 (N_5266,In_2353,In_1598);
nand U5267 (N_5267,In_2731,In_543);
nand U5268 (N_5268,In_2386,In_2395);
or U5269 (N_5269,In_2029,In_1020);
or U5270 (N_5270,In_1247,In_2986);
and U5271 (N_5271,In_297,In_1290);
nand U5272 (N_5272,In_1362,In_2715);
or U5273 (N_5273,In_1248,In_1950);
or U5274 (N_5274,In_1955,In_1927);
or U5275 (N_5275,In_1078,In_537);
and U5276 (N_5276,In_230,In_2184);
and U5277 (N_5277,In_2792,In_1726);
nand U5278 (N_5278,In_2044,In_750);
and U5279 (N_5279,In_389,In_435);
nor U5280 (N_5280,In_1583,In_1157);
xnor U5281 (N_5281,In_451,In_2484);
or U5282 (N_5282,In_1268,In_1056);
xor U5283 (N_5283,In_311,In_1413);
nand U5284 (N_5284,In_1148,In_2122);
and U5285 (N_5285,In_56,In_897);
nor U5286 (N_5286,In_2455,In_4);
nor U5287 (N_5287,In_1578,In_1665);
nand U5288 (N_5288,In_2443,In_682);
or U5289 (N_5289,In_884,In_2791);
nand U5290 (N_5290,In_398,In_429);
xnor U5291 (N_5291,In_2883,In_581);
nand U5292 (N_5292,In_49,In_17);
or U5293 (N_5293,In_1355,In_1944);
and U5294 (N_5294,In_2490,In_2673);
or U5295 (N_5295,In_317,In_938);
xnor U5296 (N_5296,In_2873,In_410);
or U5297 (N_5297,In_2744,In_2208);
nor U5298 (N_5298,In_382,In_1982);
or U5299 (N_5299,In_1281,In_2239);
or U5300 (N_5300,In_1085,In_1034);
nand U5301 (N_5301,In_2751,In_2297);
nand U5302 (N_5302,In_254,In_668);
and U5303 (N_5303,In_2397,In_1426);
and U5304 (N_5304,In_820,In_1356);
or U5305 (N_5305,In_1745,In_274);
and U5306 (N_5306,In_980,In_1412);
and U5307 (N_5307,In_1424,In_341);
nor U5308 (N_5308,In_754,In_2272);
nor U5309 (N_5309,In_2924,In_2761);
or U5310 (N_5310,In_2265,In_1772);
nor U5311 (N_5311,In_2415,In_1510);
xnor U5312 (N_5312,In_85,In_1044);
or U5313 (N_5313,In_2543,In_62);
nand U5314 (N_5314,In_959,In_2891);
nand U5315 (N_5315,In_1836,In_592);
nand U5316 (N_5316,In_7,In_2470);
and U5317 (N_5317,In_272,In_1613);
or U5318 (N_5318,In_1394,In_940);
nor U5319 (N_5319,In_1228,In_645);
or U5320 (N_5320,In_1978,In_602);
nand U5321 (N_5321,In_1220,In_1347);
and U5322 (N_5322,In_1846,In_725);
nor U5323 (N_5323,In_1393,In_234);
nor U5324 (N_5324,In_1160,In_2758);
xnor U5325 (N_5325,In_2558,In_2335);
nor U5326 (N_5326,In_2562,In_2472);
and U5327 (N_5327,In_2606,In_2293);
nand U5328 (N_5328,In_2803,In_2640);
xnor U5329 (N_5329,In_185,In_2703);
nand U5330 (N_5330,In_1927,In_455);
or U5331 (N_5331,In_838,In_313);
xor U5332 (N_5332,In_2583,In_352);
xor U5333 (N_5333,In_1463,In_1444);
nand U5334 (N_5334,In_2166,In_1160);
nor U5335 (N_5335,In_2097,In_1620);
xor U5336 (N_5336,In_941,In_7);
or U5337 (N_5337,In_1759,In_999);
or U5338 (N_5338,In_1328,In_257);
and U5339 (N_5339,In_596,In_2794);
nand U5340 (N_5340,In_2378,In_247);
nor U5341 (N_5341,In_2531,In_2308);
or U5342 (N_5342,In_2497,In_1319);
nand U5343 (N_5343,In_1981,In_888);
or U5344 (N_5344,In_2292,In_1701);
or U5345 (N_5345,In_2440,In_919);
nand U5346 (N_5346,In_2172,In_2229);
nor U5347 (N_5347,In_2556,In_2424);
nor U5348 (N_5348,In_1136,In_2264);
or U5349 (N_5349,In_1377,In_2013);
or U5350 (N_5350,In_330,In_1757);
and U5351 (N_5351,In_2140,In_2275);
nor U5352 (N_5352,In_1334,In_2268);
nor U5353 (N_5353,In_2098,In_927);
xor U5354 (N_5354,In_1604,In_2419);
nand U5355 (N_5355,In_2243,In_834);
and U5356 (N_5356,In_1985,In_352);
or U5357 (N_5357,In_2496,In_1773);
and U5358 (N_5358,In_297,In_2384);
and U5359 (N_5359,In_1044,In_2007);
and U5360 (N_5360,In_821,In_2714);
nand U5361 (N_5361,In_1386,In_1992);
or U5362 (N_5362,In_2408,In_2258);
nor U5363 (N_5363,In_146,In_1981);
nor U5364 (N_5364,In_2954,In_1640);
nor U5365 (N_5365,In_2654,In_2176);
and U5366 (N_5366,In_1344,In_1051);
nand U5367 (N_5367,In_46,In_2313);
or U5368 (N_5368,In_1872,In_1112);
or U5369 (N_5369,In_1235,In_216);
nor U5370 (N_5370,In_2261,In_1315);
nor U5371 (N_5371,In_2760,In_1220);
or U5372 (N_5372,In_2046,In_1312);
nand U5373 (N_5373,In_292,In_1927);
or U5374 (N_5374,In_564,In_2673);
and U5375 (N_5375,In_1601,In_1804);
nand U5376 (N_5376,In_2037,In_1579);
and U5377 (N_5377,In_2179,In_1692);
nand U5378 (N_5378,In_721,In_2350);
nand U5379 (N_5379,In_1940,In_562);
xnor U5380 (N_5380,In_1079,In_2773);
or U5381 (N_5381,In_2990,In_2273);
or U5382 (N_5382,In_385,In_2200);
nor U5383 (N_5383,In_918,In_1154);
and U5384 (N_5384,In_2783,In_2958);
and U5385 (N_5385,In_321,In_2288);
xor U5386 (N_5386,In_2161,In_1318);
or U5387 (N_5387,In_1265,In_1489);
or U5388 (N_5388,In_202,In_1809);
nand U5389 (N_5389,In_134,In_779);
or U5390 (N_5390,In_1765,In_1127);
xnor U5391 (N_5391,In_895,In_1490);
nor U5392 (N_5392,In_2532,In_271);
nor U5393 (N_5393,In_2501,In_1124);
nand U5394 (N_5394,In_627,In_1496);
nand U5395 (N_5395,In_254,In_299);
or U5396 (N_5396,In_2690,In_1829);
and U5397 (N_5397,In_2134,In_1401);
nand U5398 (N_5398,In_1054,In_1926);
and U5399 (N_5399,In_725,In_1833);
nor U5400 (N_5400,In_633,In_417);
xor U5401 (N_5401,In_1010,In_2485);
nand U5402 (N_5402,In_2393,In_1570);
or U5403 (N_5403,In_1523,In_687);
and U5404 (N_5404,In_2541,In_1473);
or U5405 (N_5405,In_1460,In_1704);
xor U5406 (N_5406,In_1428,In_1682);
nand U5407 (N_5407,In_816,In_2925);
nand U5408 (N_5408,In_2641,In_512);
and U5409 (N_5409,In_1297,In_1076);
or U5410 (N_5410,In_39,In_2049);
and U5411 (N_5411,In_1069,In_2983);
nand U5412 (N_5412,In_2061,In_122);
and U5413 (N_5413,In_2177,In_1294);
or U5414 (N_5414,In_2552,In_2896);
nand U5415 (N_5415,In_828,In_893);
nand U5416 (N_5416,In_1120,In_2876);
or U5417 (N_5417,In_204,In_1901);
nor U5418 (N_5418,In_109,In_2325);
or U5419 (N_5419,In_1905,In_214);
or U5420 (N_5420,In_1961,In_1169);
nor U5421 (N_5421,In_1779,In_773);
xor U5422 (N_5422,In_731,In_2651);
or U5423 (N_5423,In_2057,In_2278);
nand U5424 (N_5424,In_1088,In_1962);
or U5425 (N_5425,In_823,In_0);
nand U5426 (N_5426,In_1562,In_2756);
nor U5427 (N_5427,In_2578,In_2383);
xor U5428 (N_5428,In_711,In_161);
nand U5429 (N_5429,In_2932,In_1466);
or U5430 (N_5430,In_2832,In_2605);
and U5431 (N_5431,In_2607,In_2128);
and U5432 (N_5432,In_605,In_2120);
and U5433 (N_5433,In_2329,In_356);
or U5434 (N_5434,In_1698,In_458);
and U5435 (N_5435,In_1059,In_1610);
or U5436 (N_5436,In_2316,In_2497);
nor U5437 (N_5437,In_2200,In_1225);
nand U5438 (N_5438,In_1036,In_591);
or U5439 (N_5439,In_2761,In_8);
xnor U5440 (N_5440,In_396,In_1237);
nor U5441 (N_5441,In_445,In_1136);
nand U5442 (N_5442,In_2903,In_1097);
nor U5443 (N_5443,In_1806,In_1267);
and U5444 (N_5444,In_380,In_2048);
nand U5445 (N_5445,In_548,In_1617);
xor U5446 (N_5446,In_2697,In_539);
nor U5447 (N_5447,In_2139,In_786);
nor U5448 (N_5448,In_968,In_1254);
and U5449 (N_5449,In_2122,In_1179);
or U5450 (N_5450,In_146,In_1315);
or U5451 (N_5451,In_2860,In_645);
nand U5452 (N_5452,In_277,In_2061);
and U5453 (N_5453,In_1795,In_2544);
nand U5454 (N_5454,In_331,In_576);
nor U5455 (N_5455,In_1191,In_1117);
and U5456 (N_5456,In_2661,In_1411);
nand U5457 (N_5457,In_581,In_380);
xor U5458 (N_5458,In_396,In_2317);
and U5459 (N_5459,In_426,In_2127);
xnor U5460 (N_5460,In_2647,In_2349);
or U5461 (N_5461,In_1079,In_2843);
nand U5462 (N_5462,In_2776,In_825);
nand U5463 (N_5463,In_1480,In_2292);
xor U5464 (N_5464,In_1637,In_2287);
and U5465 (N_5465,In_2844,In_1924);
nand U5466 (N_5466,In_254,In_217);
nor U5467 (N_5467,In_294,In_1043);
nor U5468 (N_5468,In_273,In_486);
or U5469 (N_5469,In_2160,In_481);
nand U5470 (N_5470,In_1145,In_1923);
and U5471 (N_5471,In_473,In_132);
and U5472 (N_5472,In_44,In_334);
or U5473 (N_5473,In_852,In_2193);
and U5474 (N_5474,In_2464,In_2524);
nand U5475 (N_5475,In_1083,In_642);
xor U5476 (N_5476,In_81,In_412);
nand U5477 (N_5477,In_2672,In_1988);
nand U5478 (N_5478,In_1494,In_684);
or U5479 (N_5479,In_2564,In_2242);
nor U5480 (N_5480,In_464,In_1498);
xor U5481 (N_5481,In_2087,In_2887);
nand U5482 (N_5482,In_2636,In_1521);
nand U5483 (N_5483,In_2477,In_47);
nor U5484 (N_5484,In_333,In_2984);
nor U5485 (N_5485,In_1706,In_2613);
nor U5486 (N_5486,In_2404,In_2019);
nor U5487 (N_5487,In_973,In_2949);
nand U5488 (N_5488,In_1290,In_707);
or U5489 (N_5489,In_1061,In_2863);
and U5490 (N_5490,In_399,In_1772);
nor U5491 (N_5491,In_2875,In_487);
and U5492 (N_5492,In_1364,In_808);
or U5493 (N_5493,In_683,In_2172);
nand U5494 (N_5494,In_87,In_1362);
or U5495 (N_5495,In_2872,In_282);
nor U5496 (N_5496,In_131,In_1910);
xor U5497 (N_5497,In_2130,In_1133);
nor U5498 (N_5498,In_1073,In_958);
nand U5499 (N_5499,In_525,In_2049);
and U5500 (N_5500,In_1260,In_1407);
nor U5501 (N_5501,In_2422,In_518);
nor U5502 (N_5502,In_2233,In_598);
and U5503 (N_5503,In_634,In_203);
xnor U5504 (N_5504,In_499,In_1654);
or U5505 (N_5505,In_174,In_2913);
nand U5506 (N_5506,In_1341,In_2736);
and U5507 (N_5507,In_2748,In_1799);
or U5508 (N_5508,In_1888,In_1142);
xor U5509 (N_5509,In_2740,In_1519);
or U5510 (N_5510,In_1709,In_1682);
nand U5511 (N_5511,In_1802,In_2352);
nor U5512 (N_5512,In_1395,In_2641);
and U5513 (N_5513,In_2923,In_596);
and U5514 (N_5514,In_422,In_383);
nor U5515 (N_5515,In_623,In_1407);
and U5516 (N_5516,In_1293,In_1498);
nand U5517 (N_5517,In_638,In_2510);
nor U5518 (N_5518,In_1132,In_1850);
or U5519 (N_5519,In_2425,In_435);
and U5520 (N_5520,In_731,In_2711);
or U5521 (N_5521,In_2241,In_2506);
xnor U5522 (N_5522,In_2176,In_196);
nor U5523 (N_5523,In_1108,In_2069);
or U5524 (N_5524,In_1102,In_1908);
and U5525 (N_5525,In_1096,In_36);
and U5526 (N_5526,In_2444,In_2049);
and U5527 (N_5527,In_2711,In_1279);
or U5528 (N_5528,In_567,In_168);
nor U5529 (N_5529,In_1979,In_787);
nor U5530 (N_5530,In_1670,In_141);
or U5531 (N_5531,In_2816,In_895);
nand U5532 (N_5532,In_933,In_2219);
xnor U5533 (N_5533,In_2268,In_2078);
or U5534 (N_5534,In_2842,In_206);
nor U5535 (N_5535,In_1526,In_1510);
nand U5536 (N_5536,In_1805,In_944);
xnor U5537 (N_5537,In_659,In_690);
nand U5538 (N_5538,In_199,In_2544);
or U5539 (N_5539,In_450,In_426);
or U5540 (N_5540,In_313,In_2349);
nand U5541 (N_5541,In_1562,In_2923);
or U5542 (N_5542,In_2247,In_377);
and U5543 (N_5543,In_1462,In_2772);
or U5544 (N_5544,In_2969,In_2867);
nand U5545 (N_5545,In_321,In_2789);
or U5546 (N_5546,In_198,In_2335);
nor U5547 (N_5547,In_264,In_1867);
nor U5548 (N_5548,In_1397,In_1120);
nor U5549 (N_5549,In_1149,In_1413);
nand U5550 (N_5550,In_2920,In_454);
nor U5551 (N_5551,In_346,In_623);
nor U5552 (N_5552,In_1435,In_2704);
nor U5553 (N_5553,In_726,In_1189);
xor U5554 (N_5554,In_1287,In_973);
and U5555 (N_5555,In_2225,In_517);
or U5556 (N_5556,In_2186,In_2291);
nand U5557 (N_5557,In_263,In_1543);
and U5558 (N_5558,In_2714,In_2550);
nor U5559 (N_5559,In_2199,In_1338);
and U5560 (N_5560,In_307,In_702);
nor U5561 (N_5561,In_2068,In_352);
nand U5562 (N_5562,In_1059,In_2963);
xnor U5563 (N_5563,In_2207,In_1625);
or U5564 (N_5564,In_1079,In_2767);
or U5565 (N_5565,In_1383,In_1001);
nor U5566 (N_5566,In_857,In_2291);
nand U5567 (N_5567,In_1752,In_2758);
nor U5568 (N_5568,In_1786,In_894);
nand U5569 (N_5569,In_101,In_2335);
nor U5570 (N_5570,In_1495,In_1305);
nand U5571 (N_5571,In_1995,In_1723);
or U5572 (N_5572,In_1755,In_12);
and U5573 (N_5573,In_2963,In_2232);
nor U5574 (N_5574,In_690,In_1772);
nor U5575 (N_5575,In_2506,In_109);
and U5576 (N_5576,In_1683,In_1302);
nand U5577 (N_5577,In_2232,In_797);
and U5578 (N_5578,In_2598,In_1374);
xnor U5579 (N_5579,In_1884,In_424);
nand U5580 (N_5580,In_2735,In_201);
and U5581 (N_5581,In_1986,In_280);
or U5582 (N_5582,In_2320,In_1032);
or U5583 (N_5583,In_102,In_1126);
xor U5584 (N_5584,In_558,In_830);
and U5585 (N_5585,In_1637,In_1506);
xnor U5586 (N_5586,In_609,In_2263);
nor U5587 (N_5587,In_1257,In_1053);
or U5588 (N_5588,In_2138,In_901);
xnor U5589 (N_5589,In_1131,In_214);
nand U5590 (N_5590,In_2457,In_2218);
and U5591 (N_5591,In_1124,In_1299);
xor U5592 (N_5592,In_2065,In_799);
or U5593 (N_5593,In_132,In_167);
nor U5594 (N_5594,In_2301,In_2634);
and U5595 (N_5595,In_2657,In_2500);
nand U5596 (N_5596,In_2721,In_715);
nor U5597 (N_5597,In_2848,In_1705);
and U5598 (N_5598,In_455,In_2647);
or U5599 (N_5599,In_1130,In_1719);
and U5600 (N_5600,In_1983,In_1383);
or U5601 (N_5601,In_1789,In_885);
nor U5602 (N_5602,In_351,In_1055);
xor U5603 (N_5603,In_2710,In_566);
and U5604 (N_5604,In_1380,In_2780);
nor U5605 (N_5605,In_2401,In_261);
and U5606 (N_5606,In_2902,In_2680);
xnor U5607 (N_5607,In_2204,In_1532);
nor U5608 (N_5608,In_276,In_1352);
nor U5609 (N_5609,In_1357,In_1957);
and U5610 (N_5610,In_1929,In_2217);
nor U5611 (N_5611,In_2654,In_1714);
or U5612 (N_5612,In_839,In_1051);
or U5613 (N_5613,In_899,In_430);
or U5614 (N_5614,In_2461,In_1008);
nand U5615 (N_5615,In_436,In_2223);
nor U5616 (N_5616,In_2409,In_1007);
nand U5617 (N_5617,In_1901,In_933);
or U5618 (N_5618,In_642,In_433);
and U5619 (N_5619,In_2658,In_1027);
nor U5620 (N_5620,In_198,In_233);
and U5621 (N_5621,In_2490,In_1463);
nand U5622 (N_5622,In_2476,In_190);
or U5623 (N_5623,In_2821,In_2874);
nor U5624 (N_5624,In_2213,In_995);
nor U5625 (N_5625,In_1590,In_1676);
or U5626 (N_5626,In_112,In_42);
or U5627 (N_5627,In_2843,In_27);
or U5628 (N_5628,In_659,In_1795);
and U5629 (N_5629,In_8,In_1397);
nand U5630 (N_5630,In_1733,In_655);
or U5631 (N_5631,In_2402,In_332);
nor U5632 (N_5632,In_2761,In_1266);
or U5633 (N_5633,In_1559,In_277);
and U5634 (N_5634,In_988,In_2852);
nor U5635 (N_5635,In_2171,In_13);
nand U5636 (N_5636,In_423,In_1642);
and U5637 (N_5637,In_2335,In_2700);
nor U5638 (N_5638,In_113,In_1317);
or U5639 (N_5639,In_99,In_495);
and U5640 (N_5640,In_1461,In_1884);
or U5641 (N_5641,In_2687,In_2662);
and U5642 (N_5642,In_1799,In_2294);
xnor U5643 (N_5643,In_2546,In_935);
and U5644 (N_5644,In_2062,In_1442);
nand U5645 (N_5645,In_1089,In_2280);
nor U5646 (N_5646,In_2803,In_2098);
xor U5647 (N_5647,In_2467,In_2082);
nor U5648 (N_5648,In_2077,In_976);
nor U5649 (N_5649,In_2880,In_1732);
or U5650 (N_5650,In_2277,In_960);
xor U5651 (N_5651,In_1769,In_887);
or U5652 (N_5652,In_507,In_1895);
nand U5653 (N_5653,In_1276,In_102);
and U5654 (N_5654,In_348,In_1174);
or U5655 (N_5655,In_849,In_955);
and U5656 (N_5656,In_1206,In_750);
or U5657 (N_5657,In_2807,In_378);
nor U5658 (N_5658,In_450,In_2370);
nor U5659 (N_5659,In_2305,In_2124);
xor U5660 (N_5660,In_1484,In_2396);
nand U5661 (N_5661,In_2312,In_2686);
xor U5662 (N_5662,In_814,In_751);
or U5663 (N_5663,In_669,In_1313);
and U5664 (N_5664,In_1755,In_2840);
nand U5665 (N_5665,In_2924,In_2945);
and U5666 (N_5666,In_1336,In_135);
nand U5667 (N_5667,In_2644,In_2065);
nand U5668 (N_5668,In_331,In_1635);
nand U5669 (N_5669,In_399,In_2178);
and U5670 (N_5670,In_860,In_360);
and U5671 (N_5671,In_893,In_2809);
and U5672 (N_5672,In_199,In_2424);
or U5673 (N_5673,In_1988,In_1424);
xor U5674 (N_5674,In_2452,In_336);
xnor U5675 (N_5675,In_1274,In_1910);
nor U5676 (N_5676,In_655,In_2307);
and U5677 (N_5677,In_2427,In_1391);
nand U5678 (N_5678,In_1093,In_574);
and U5679 (N_5679,In_2242,In_2073);
and U5680 (N_5680,In_2873,In_513);
or U5681 (N_5681,In_463,In_1697);
nor U5682 (N_5682,In_185,In_1416);
and U5683 (N_5683,In_1307,In_317);
or U5684 (N_5684,In_2303,In_58);
or U5685 (N_5685,In_2830,In_1641);
or U5686 (N_5686,In_2823,In_2855);
and U5687 (N_5687,In_1160,In_2852);
nand U5688 (N_5688,In_2367,In_2527);
nand U5689 (N_5689,In_1044,In_1002);
nor U5690 (N_5690,In_559,In_666);
nor U5691 (N_5691,In_600,In_2435);
and U5692 (N_5692,In_674,In_700);
nor U5693 (N_5693,In_453,In_2936);
xnor U5694 (N_5694,In_2823,In_1715);
and U5695 (N_5695,In_2360,In_1890);
nor U5696 (N_5696,In_1623,In_2579);
nor U5697 (N_5697,In_2973,In_10);
xnor U5698 (N_5698,In_1763,In_870);
and U5699 (N_5699,In_1778,In_926);
or U5700 (N_5700,In_1334,In_176);
or U5701 (N_5701,In_2402,In_311);
or U5702 (N_5702,In_2372,In_2282);
nor U5703 (N_5703,In_2615,In_105);
nor U5704 (N_5704,In_1255,In_2846);
nor U5705 (N_5705,In_1935,In_1977);
nand U5706 (N_5706,In_1266,In_1237);
nand U5707 (N_5707,In_1082,In_2179);
nand U5708 (N_5708,In_653,In_160);
xor U5709 (N_5709,In_1140,In_177);
and U5710 (N_5710,In_1288,In_2106);
xor U5711 (N_5711,In_561,In_2896);
and U5712 (N_5712,In_1010,In_42);
xor U5713 (N_5713,In_1767,In_2683);
xor U5714 (N_5714,In_2679,In_2357);
and U5715 (N_5715,In_2508,In_2469);
nor U5716 (N_5716,In_1384,In_542);
or U5717 (N_5717,In_1097,In_302);
or U5718 (N_5718,In_2277,In_1960);
nor U5719 (N_5719,In_1950,In_1629);
nor U5720 (N_5720,In_116,In_2304);
nand U5721 (N_5721,In_1233,In_499);
or U5722 (N_5722,In_2985,In_1745);
or U5723 (N_5723,In_1236,In_27);
nor U5724 (N_5724,In_1448,In_1860);
and U5725 (N_5725,In_617,In_1721);
nand U5726 (N_5726,In_881,In_2631);
nor U5727 (N_5727,In_1698,In_1445);
nor U5728 (N_5728,In_2391,In_2759);
nor U5729 (N_5729,In_2417,In_1389);
and U5730 (N_5730,In_2301,In_2658);
nor U5731 (N_5731,In_785,In_2759);
nor U5732 (N_5732,In_1934,In_2842);
or U5733 (N_5733,In_2634,In_2079);
nor U5734 (N_5734,In_1736,In_2933);
or U5735 (N_5735,In_2800,In_1234);
nor U5736 (N_5736,In_1965,In_724);
and U5737 (N_5737,In_2357,In_1069);
nor U5738 (N_5738,In_1284,In_1327);
nand U5739 (N_5739,In_1265,In_22);
or U5740 (N_5740,In_2830,In_995);
nor U5741 (N_5741,In_543,In_9);
or U5742 (N_5742,In_928,In_1098);
or U5743 (N_5743,In_1499,In_480);
or U5744 (N_5744,In_1860,In_2147);
nand U5745 (N_5745,In_2185,In_924);
nand U5746 (N_5746,In_1011,In_1405);
and U5747 (N_5747,In_1819,In_1743);
xor U5748 (N_5748,In_1100,In_1268);
nand U5749 (N_5749,In_2926,In_639);
and U5750 (N_5750,In_360,In_2784);
nand U5751 (N_5751,In_1080,In_1397);
nand U5752 (N_5752,In_788,In_781);
or U5753 (N_5753,In_186,In_983);
or U5754 (N_5754,In_701,In_2063);
nor U5755 (N_5755,In_204,In_2094);
and U5756 (N_5756,In_990,In_866);
xnor U5757 (N_5757,In_211,In_1239);
nor U5758 (N_5758,In_1595,In_2523);
nor U5759 (N_5759,In_1999,In_1165);
or U5760 (N_5760,In_136,In_451);
nor U5761 (N_5761,In_490,In_760);
nor U5762 (N_5762,In_1614,In_2601);
nor U5763 (N_5763,In_2824,In_2635);
and U5764 (N_5764,In_1068,In_2067);
nor U5765 (N_5765,In_2625,In_638);
or U5766 (N_5766,In_2050,In_110);
nand U5767 (N_5767,In_2627,In_2389);
and U5768 (N_5768,In_450,In_1076);
or U5769 (N_5769,In_2737,In_1287);
nor U5770 (N_5770,In_1466,In_1034);
nand U5771 (N_5771,In_1597,In_1599);
nor U5772 (N_5772,In_1294,In_1822);
nor U5773 (N_5773,In_1019,In_1917);
nor U5774 (N_5774,In_2484,In_610);
nand U5775 (N_5775,In_1804,In_855);
xor U5776 (N_5776,In_141,In_229);
and U5777 (N_5777,In_1216,In_2842);
nor U5778 (N_5778,In_2298,In_507);
nand U5779 (N_5779,In_2126,In_1297);
and U5780 (N_5780,In_237,In_2770);
or U5781 (N_5781,In_76,In_2592);
and U5782 (N_5782,In_147,In_2282);
xnor U5783 (N_5783,In_1288,In_295);
or U5784 (N_5784,In_2137,In_181);
nor U5785 (N_5785,In_2653,In_2443);
nand U5786 (N_5786,In_1091,In_560);
and U5787 (N_5787,In_2606,In_855);
or U5788 (N_5788,In_2381,In_2890);
nand U5789 (N_5789,In_2714,In_1244);
nor U5790 (N_5790,In_594,In_1315);
nand U5791 (N_5791,In_821,In_254);
nand U5792 (N_5792,In_732,In_1867);
and U5793 (N_5793,In_791,In_1585);
nor U5794 (N_5794,In_197,In_620);
nor U5795 (N_5795,In_408,In_2535);
and U5796 (N_5796,In_2934,In_2330);
nand U5797 (N_5797,In_2195,In_815);
or U5798 (N_5798,In_1430,In_1714);
xor U5799 (N_5799,In_604,In_1704);
nand U5800 (N_5800,In_1839,In_1459);
nor U5801 (N_5801,In_1590,In_2830);
or U5802 (N_5802,In_890,In_2845);
nand U5803 (N_5803,In_2662,In_2278);
xor U5804 (N_5804,In_1972,In_927);
xor U5805 (N_5805,In_228,In_2947);
and U5806 (N_5806,In_790,In_2955);
xor U5807 (N_5807,In_2541,In_2842);
xnor U5808 (N_5808,In_244,In_999);
nand U5809 (N_5809,In_2172,In_1615);
or U5810 (N_5810,In_97,In_673);
and U5811 (N_5811,In_1518,In_545);
nand U5812 (N_5812,In_2192,In_1753);
nand U5813 (N_5813,In_2817,In_1520);
or U5814 (N_5814,In_1791,In_1977);
or U5815 (N_5815,In_2167,In_2927);
and U5816 (N_5816,In_1586,In_2923);
xnor U5817 (N_5817,In_299,In_1478);
or U5818 (N_5818,In_176,In_254);
xor U5819 (N_5819,In_2923,In_719);
or U5820 (N_5820,In_2153,In_551);
nor U5821 (N_5821,In_2071,In_2259);
nor U5822 (N_5822,In_1568,In_2259);
nor U5823 (N_5823,In_510,In_848);
nand U5824 (N_5824,In_1652,In_1522);
and U5825 (N_5825,In_2845,In_2381);
and U5826 (N_5826,In_75,In_2823);
or U5827 (N_5827,In_1320,In_2506);
or U5828 (N_5828,In_238,In_2555);
nand U5829 (N_5829,In_339,In_23);
or U5830 (N_5830,In_2696,In_2418);
or U5831 (N_5831,In_1048,In_651);
xnor U5832 (N_5832,In_2963,In_2337);
nand U5833 (N_5833,In_1844,In_1462);
nand U5834 (N_5834,In_1532,In_2048);
nor U5835 (N_5835,In_152,In_820);
and U5836 (N_5836,In_2983,In_1518);
and U5837 (N_5837,In_1148,In_294);
and U5838 (N_5838,In_1479,In_2665);
or U5839 (N_5839,In_872,In_308);
nand U5840 (N_5840,In_2886,In_1547);
nor U5841 (N_5841,In_2424,In_441);
or U5842 (N_5842,In_2563,In_2549);
nor U5843 (N_5843,In_1618,In_1564);
or U5844 (N_5844,In_2689,In_35);
or U5845 (N_5845,In_874,In_488);
or U5846 (N_5846,In_2411,In_1280);
nor U5847 (N_5847,In_407,In_1692);
nand U5848 (N_5848,In_1768,In_1367);
or U5849 (N_5849,In_2912,In_2588);
or U5850 (N_5850,In_1035,In_1288);
nor U5851 (N_5851,In_2217,In_367);
nand U5852 (N_5852,In_134,In_1259);
and U5853 (N_5853,In_2504,In_2674);
nand U5854 (N_5854,In_879,In_2340);
nor U5855 (N_5855,In_2799,In_2865);
or U5856 (N_5856,In_1168,In_126);
nor U5857 (N_5857,In_2296,In_1727);
or U5858 (N_5858,In_2807,In_2742);
nand U5859 (N_5859,In_1442,In_108);
xnor U5860 (N_5860,In_459,In_319);
nand U5861 (N_5861,In_1828,In_2812);
and U5862 (N_5862,In_2616,In_2064);
or U5863 (N_5863,In_419,In_187);
and U5864 (N_5864,In_1621,In_142);
or U5865 (N_5865,In_833,In_2194);
nor U5866 (N_5866,In_1906,In_1526);
nor U5867 (N_5867,In_263,In_717);
nand U5868 (N_5868,In_839,In_1009);
nand U5869 (N_5869,In_1153,In_1456);
xnor U5870 (N_5870,In_621,In_490);
nor U5871 (N_5871,In_2957,In_1427);
or U5872 (N_5872,In_455,In_43);
nand U5873 (N_5873,In_1237,In_2763);
nor U5874 (N_5874,In_1035,In_802);
or U5875 (N_5875,In_2179,In_1811);
nor U5876 (N_5876,In_2111,In_1389);
nand U5877 (N_5877,In_501,In_755);
nor U5878 (N_5878,In_1001,In_2772);
nor U5879 (N_5879,In_1156,In_2695);
nand U5880 (N_5880,In_207,In_1183);
or U5881 (N_5881,In_1978,In_616);
nand U5882 (N_5882,In_0,In_2656);
and U5883 (N_5883,In_2350,In_1768);
nand U5884 (N_5884,In_368,In_1132);
and U5885 (N_5885,In_1615,In_1803);
nand U5886 (N_5886,In_2748,In_2792);
nor U5887 (N_5887,In_2493,In_2824);
or U5888 (N_5888,In_545,In_1675);
nand U5889 (N_5889,In_473,In_1340);
nor U5890 (N_5890,In_112,In_2226);
or U5891 (N_5891,In_2954,In_67);
or U5892 (N_5892,In_10,In_1469);
nand U5893 (N_5893,In_884,In_707);
nor U5894 (N_5894,In_2771,In_1952);
nor U5895 (N_5895,In_1567,In_2720);
nand U5896 (N_5896,In_1326,In_593);
or U5897 (N_5897,In_875,In_2500);
nand U5898 (N_5898,In_735,In_2302);
and U5899 (N_5899,In_1555,In_961);
nand U5900 (N_5900,In_1075,In_601);
nand U5901 (N_5901,In_1706,In_2259);
and U5902 (N_5902,In_2777,In_136);
nand U5903 (N_5903,In_2531,In_2465);
and U5904 (N_5904,In_650,In_1838);
or U5905 (N_5905,In_1724,In_2145);
nor U5906 (N_5906,In_2696,In_825);
xnor U5907 (N_5907,In_342,In_1352);
and U5908 (N_5908,In_243,In_1482);
and U5909 (N_5909,In_2030,In_2006);
or U5910 (N_5910,In_1778,In_294);
or U5911 (N_5911,In_1260,In_494);
xnor U5912 (N_5912,In_1164,In_2255);
nand U5913 (N_5913,In_2545,In_348);
and U5914 (N_5914,In_129,In_2080);
xnor U5915 (N_5915,In_459,In_2170);
xnor U5916 (N_5916,In_1191,In_2883);
nor U5917 (N_5917,In_574,In_2997);
or U5918 (N_5918,In_2335,In_1430);
and U5919 (N_5919,In_51,In_1746);
nand U5920 (N_5920,In_1269,In_2584);
nor U5921 (N_5921,In_1044,In_167);
xor U5922 (N_5922,In_1343,In_2558);
or U5923 (N_5923,In_2805,In_2971);
and U5924 (N_5924,In_1418,In_2315);
xor U5925 (N_5925,In_2122,In_2423);
nand U5926 (N_5926,In_496,In_1841);
nand U5927 (N_5927,In_678,In_2287);
or U5928 (N_5928,In_461,In_1813);
nand U5929 (N_5929,In_2505,In_1603);
nor U5930 (N_5930,In_1484,In_1372);
nand U5931 (N_5931,In_1968,In_2910);
nor U5932 (N_5932,In_706,In_89);
and U5933 (N_5933,In_2566,In_2931);
nand U5934 (N_5934,In_2811,In_812);
or U5935 (N_5935,In_127,In_359);
nor U5936 (N_5936,In_1550,In_1897);
nor U5937 (N_5937,In_52,In_935);
or U5938 (N_5938,In_734,In_816);
xnor U5939 (N_5939,In_875,In_215);
nor U5940 (N_5940,In_435,In_340);
and U5941 (N_5941,In_25,In_2546);
nor U5942 (N_5942,In_315,In_543);
nor U5943 (N_5943,In_2494,In_672);
nor U5944 (N_5944,In_2024,In_1517);
nor U5945 (N_5945,In_2445,In_728);
or U5946 (N_5946,In_1369,In_2330);
nor U5947 (N_5947,In_2074,In_1132);
xor U5948 (N_5948,In_1588,In_50);
and U5949 (N_5949,In_1033,In_2638);
and U5950 (N_5950,In_605,In_2460);
nor U5951 (N_5951,In_766,In_2811);
or U5952 (N_5952,In_2629,In_2014);
nand U5953 (N_5953,In_22,In_2779);
or U5954 (N_5954,In_565,In_280);
and U5955 (N_5955,In_2098,In_2759);
nor U5956 (N_5956,In_2326,In_404);
nor U5957 (N_5957,In_1451,In_2762);
nor U5958 (N_5958,In_1307,In_1116);
or U5959 (N_5959,In_2879,In_2442);
or U5960 (N_5960,In_476,In_379);
xor U5961 (N_5961,In_2927,In_535);
and U5962 (N_5962,In_2869,In_1910);
and U5963 (N_5963,In_1580,In_408);
and U5964 (N_5964,In_585,In_1832);
nand U5965 (N_5965,In_354,In_2752);
nor U5966 (N_5966,In_43,In_1196);
nand U5967 (N_5967,In_1704,In_61);
nand U5968 (N_5968,In_2039,In_633);
or U5969 (N_5969,In_1542,In_2579);
nand U5970 (N_5970,In_90,In_170);
nand U5971 (N_5971,In_28,In_776);
and U5972 (N_5972,In_1933,In_16);
or U5973 (N_5973,In_1337,In_733);
nor U5974 (N_5974,In_2415,In_392);
nor U5975 (N_5975,In_935,In_912);
and U5976 (N_5976,In_1849,In_505);
and U5977 (N_5977,In_1223,In_2397);
nand U5978 (N_5978,In_1738,In_2010);
or U5979 (N_5979,In_1672,In_2469);
nor U5980 (N_5980,In_177,In_304);
or U5981 (N_5981,In_1555,In_2936);
or U5982 (N_5982,In_246,In_803);
xnor U5983 (N_5983,In_1275,In_2553);
nor U5984 (N_5984,In_1949,In_538);
nor U5985 (N_5985,In_2580,In_2315);
or U5986 (N_5986,In_1454,In_2803);
nor U5987 (N_5987,In_2052,In_1207);
nor U5988 (N_5988,In_2682,In_1602);
nor U5989 (N_5989,In_1416,In_2285);
and U5990 (N_5990,In_2759,In_2306);
or U5991 (N_5991,In_194,In_2023);
or U5992 (N_5992,In_2152,In_2559);
and U5993 (N_5993,In_940,In_189);
or U5994 (N_5994,In_2860,In_1957);
and U5995 (N_5995,In_1994,In_2865);
nand U5996 (N_5996,In_2429,In_2959);
nand U5997 (N_5997,In_900,In_2403);
or U5998 (N_5998,In_542,In_2885);
nor U5999 (N_5999,In_1523,In_516);
nand U6000 (N_6000,In_1380,In_2321);
nand U6001 (N_6001,In_207,In_2565);
nand U6002 (N_6002,In_880,In_817);
xnor U6003 (N_6003,In_2464,In_1145);
or U6004 (N_6004,In_484,In_2949);
nand U6005 (N_6005,In_2890,In_256);
xnor U6006 (N_6006,In_784,In_16);
nor U6007 (N_6007,In_1164,In_2834);
or U6008 (N_6008,In_235,In_247);
nor U6009 (N_6009,In_711,In_2091);
nor U6010 (N_6010,In_301,In_396);
nand U6011 (N_6011,In_1014,In_2733);
xnor U6012 (N_6012,In_1607,In_453);
and U6013 (N_6013,In_2831,In_1704);
nor U6014 (N_6014,In_1457,In_2986);
or U6015 (N_6015,In_2040,In_1839);
and U6016 (N_6016,In_1019,In_2687);
nor U6017 (N_6017,In_2659,In_1294);
and U6018 (N_6018,In_636,In_1736);
nor U6019 (N_6019,In_1679,In_792);
and U6020 (N_6020,In_836,In_2125);
nor U6021 (N_6021,In_1300,In_1347);
or U6022 (N_6022,In_2046,In_534);
and U6023 (N_6023,In_1626,In_518);
nand U6024 (N_6024,In_265,In_701);
nand U6025 (N_6025,In_1720,In_1595);
and U6026 (N_6026,In_1888,In_1330);
nand U6027 (N_6027,In_277,In_1720);
or U6028 (N_6028,In_406,In_964);
or U6029 (N_6029,In_2525,In_2642);
nand U6030 (N_6030,In_2440,In_2188);
or U6031 (N_6031,In_719,In_2611);
or U6032 (N_6032,In_2750,In_2875);
or U6033 (N_6033,In_729,In_2776);
nand U6034 (N_6034,In_586,In_140);
nand U6035 (N_6035,In_27,In_997);
or U6036 (N_6036,In_2221,In_2589);
and U6037 (N_6037,In_1223,In_1190);
nand U6038 (N_6038,In_784,In_1682);
nor U6039 (N_6039,In_155,In_1798);
and U6040 (N_6040,In_1036,In_2674);
and U6041 (N_6041,In_1355,In_285);
or U6042 (N_6042,In_2162,In_2348);
xnor U6043 (N_6043,In_2586,In_2474);
nand U6044 (N_6044,In_1372,In_1370);
nand U6045 (N_6045,In_682,In_1010);
nor U6046 (N_6046,In_327,In_2476);
xnor U6047 (N_6047,In_765,In_1406);
nand U6048 (N_6048,In_2775,In_31);
nor U6049 (N_6049,In_2225,In_1384);
xnor U6050 (N_6050,In_352,In_292);
and U6051 (N_6051,In_201,In_2789);
and U6052 (N_6052,In_508,In_874);
and U6053 (N_6053,In_2641,In_2825);
nand U6054 (N_6054,In_2323,In_310);
nor U6055 (N_6055,In_32,In_110);
or U6056 (N_6056,In_1725,In_1230);
nand U6057 (N_6057,In_1502,In_2485);
or U6058 (N_6058,In_860,In_1173);
nor U6059 (N_6059,In_176,In_2896);
xor U6060 (N_6060,In_1748,In_1179);
or U6061 (N_6061,In_685,In_2563);
nand U6062 (N_6062,In_2530,In_2788);
and U6063 (N_6063,In_1052,In_873);
xnor U6064 (N_6064,In_120,In_1286);
nor U6065 (N_6065,In_54,In_471);
and U6066 (N_6066,In_140,In_1278);
nand U6067 (N_6067,In_889,In_2595);
or U6068 (N_6068,In_2703,In_2268);
or U6069 (N_6069,In_344,In_925);
and U6070 (N_6070,In_386,In_1264);
or U6071 (N_6071,In_1054,In_442);
nand U6072 (N_6072,In_1117,In_334);
or U6073 (N_6073,In_1373,In_871);
nor U6074 (N_6074,In_815,In_626);
or U6075 (N_6075,In_820,In_1244);
nand U6076 (N_6076,In_816,In_2438);
nor U6077 (N_6077,In_1226,In_485);
nand U6078 (N_6078,In_2854,In_1592);
nor U6079 (N_6079,In_514,In_746);
and U6080 (N_6080,In_1240,In_2380);
and U6081 (N_6081,In_2335,In_2323);
or U6082 (N_6082,In_1853,In_160);
or U6083 (N_6083,In_963,In_1010);
or U6084 (N_6084,In_2301,In_1898);
and U6085 (N_6085,In_1593,In_2452);
nand U6086 (N_6086,In_1158,In_2904);
nand U6087 (N_6087,In_2785,In_1954);
xnor U6088 (N_6088,In_2928,In_2685);
nor U6089 (N_6089,In_1118,In_2202);
nor U6090 (N_6090,In_1107,In_2209);
nand U6091 (N_6091,In_2534,In_2688);
nand U6092 (N_6092,In_694,In_1046);
and U6093 (N_6093,In_1119,In_462);
or U6094 (N_6094,In_2122,In_120);
and U6095 (N_6095,In_2178,In_776);
nor U6096 (N_6096,In_2982,In_2902);
nor U6097 (N_6097,In_1285,In_1216);
xor U6098 (N_6098,In_2931,In_1537);
and U6099 (N_6099,In_2446,In_1165);
nand U6100 (N_6100,In_2966,In_2922);
and U6101 (N_6101,In_1558,In_2963);
and U6102 (N_6102,In_1304,In_1607);
or U6103 (N_6103,In_2285,In_1215);
nand U6104 (N_6104,In_378,In_440);
and U6105 (N_6105,In_476,In_1835);
or U6106 (N_6106,In_2431,In_697);
nor U6107 (N_6107,In_772,In_2115);
xor U6108 (N_6108,In_775,In_1787);
nand U6109 (N_6109,In_380,In_1641);
nor U6110 (N_6110,In_2421,In_287);
nand U6111 (N_6111,In_1552,In_2101);
xor U6112 (N_6112,In_2056,In_2127);
and U6113 (N_6113,In_2202,In_1060);
or U6114 (N_6114,In_1156,In_2739);
or U6115 (N_6115,In_592,In_1482);
and U6116 (N_6116,In_1585,In_1234);
and U6117 (N_6117,In_2738,In_1978);
nand U6118 (N_6118,In_2816,In_2429);
and U6119 (N_6119,In_952,In_2380);
or U6120 (N_6120,In_1840,In_2457);
nand U6121 (N_6121,In_1110,In_1751);
or U6122 (N_6122,In_2764,In_2633);
nand U6123 (N_6123,In_1169,In_1068);
or U6124 (N_6124,In_888,In_139);
and U6125 (N_6125,In_979,In_2704);
or U6126 (N_6126,In_569,In_1510);
nand U6127 (N_6127,In_2442,In_1864);
nor U6128 (N_6128,In_1289,In_616);
or U6129 (N_6129,In_189,In_1283);
nor U6130 (N_6130,In_1005,In_1152);
nor U6131 (N_6131,In_1513,In_142);
or U6132 (N_6132,In_1599,In_1239);
and U6133 (N_6133,In_163,In_1130);
nor U6134 (N_6134,In_139,In_2431);
nand U6135 (N_6135,In_2338,In_1259);
xor U6136 (N_6136,In_1902,In_46);
nor U6137 (N_6137,In_400,In_2325);
or U6138 (N_6138,In_1836,In_1676);
or U6139 (N_6139,In_376,In_2992);
or U6140 (N_6140,In_779,In_2258);
nand U6141 (N_6141,In_453,In_2519);
and U6142 (N_6142,In_1539,In_1434);
nand U6143 (N_6143,In_2075,In_1097);
nand U6144 (N_6144,In_1487,In_912);
or U6145 (N_6145,In_2792,In_1684);
and U6146 (N_6146,In_2780,In_401);
and U6147 (N_6147,In_678,In_684);
nand U6148 (N_6148,In_2242,In_1752);
xor U6149 (N_6149,In_283,In_2470);
and U6150 (N_6150,In_2664,In_945);
nor U6151 (N_6151,In_2054,In_1806);
nor U6152 (N_6152,In_1141,In_1091);
or U6153 (N_6153,In_198,In_2538);
or U6154 (N_6154,In_2035,In_2008);
nand U6155 (N_6155,In_912,In_1661);
nor U6156 (N_6156,In_90,In_2660);
nand U6157 (N_6157,In_2190,In_2655);
nor U6158 (N_6158,In_2867,In_2150);
nor U6159 (N_6159,In_1082,In_2569);
nor U6160 (N_6160,In_2906,In_64);
or U6161 (N_6161,In_1451,In_2360);
nor U6162 (N_6162,In_1159,In_687);
and U6163 (N_6163,In_1124,In_1459);
or U6164 (N_6164,In_981,In_998);
or U6165 (N_6165,In_468,In_650);
nor U6166 (N_6166,In_737,In_2709);
nor U6167 (N_6167,In_2100,In_1301);
or U6168 (N_6168,In_2677,In_2899);
nor U6169 (N_6169,In_1292,In_2994);
nand U6170 (N_6170,In_1981,In_1873);
xor U6171 (N_6171,In_2893,In_745);
and U6172 (N_6172,In_2014,In_424);
nor U6173 (N_6173,In_2319,In_2886);
xnor U6174 (N_6174,In_1442,In_874);
nor U6175 (N_6175,In_783,In_2239);
and U6176 (N_6176,In_2582,In_2824);
nor U6177 (N_6177,In_1342,In_2578);
and U6178 (N_6178,In_230,In_1605);
or U6179 (N_6179,In_284,In_2141);
nor U6180 (N_6180,In_908,In_1156);
nand U6181 (N_6181,In_767,In_26);
nand U6182 (N_6182,In_873,In_55);
or U6183 (N_6183,In_683,In_1727);
xor U6184 (N_6184,In_240,In_2236);
xnor U6185 (N_6185,In_620,In_1726);
nand U6186 (N_6186,In_1225,In_1224);
xnor U6187 (N_6187,In_419,In_132);
nor U6188 (N_6188,In_2944,In_1229);
or U6189 (N_6189,In_1303,In_1246);
nor U6190 (N_6190,In_2812,In_2384);
or U6191 (N_6191,In_649,In_2654);
and U6192 (N_6192,In_1976,In_2912);
or U6193 (N_6193,In_1107,In_203);
nand U6194 (N_6194,In_250,In_115);
xnor U6195 (N_6195,In_1622,In_2018);
xor U6196 (N_6196,In_1855,In_1427);
or U6197 (N_6197,In_1877,In_172);
or U6198 (N_6198,In_1251,In_2224);
nor U6199 (N_6199,In_1830,In_2524);
or U6200 (N_6200,In_1412,In_142);
nor U6201 (N_6201,In_2902,In_2537);
or U6202 (N_6202,In_2771,In_1788);
nor U6203 (N_6203,In_905,In_1587);
and U6204 (N_6204,In_2749,In_2518);
and U6205 (N_6205,In_2445,In_965);
xnor U6206 (N_6206,In_2962,In_1398);
or U6207 (N_6207,In_784,In_2253);
and U6208 (N_6208,In_862,In_198);
and U6209 (N_6209,In_2714,In_2797);
xor U6210 (N_6210,In_1364,In_2638);
nand U6211 (N_6211,In_2078,In_2336);
xnor U6212 (N_6212,In_601,In_133);
nand U6213 (N_6213,In_2378,In_794);
xor U6214 (N_6214,In_1829,In_1002);
nand U6215 (N_6215,In_778,In_2064);
or U6216 (N_6216,In_2796,In_2020);
nand U6217 (N_6217,In_2334,In_2306);
nand U6218 (N_6218,In_1763,In_1098);
nand U6219 (N_6219,In_650,In_715);
or U6220 (N_6220,In_2102,In_35);
or U6221 (N_6221,In_2423,In_2032);
xor U6222 (N_6222,In_2616,In_2318);
and U6223 (N_6223,In_2461,In_169);
nand U6224 (N_6224,In_834,In_1919);
xor U6225 (N_6225,In_572,In_523);
xnor U6226 (N_6226,In_2525,In_1152);
nand U6227 (N_6227,In_960,In_1465);
nand U6228 (N_6228,In_1651,In_2098);
nor U6229 (N_6229,In_1931,In_855);
nor U6230 (N_6230,In_755,In_2703);
nand U6231 (N_6231,In_1200,In_1703);
nand U6232 (N_6232,In_1578,In_2825);
nand U6233 (N_6233,In_825,In_1388);
or U6234 (N_6234,In_1075,In_2164);
nor U6235 (N_6235,In_2379,In_574);
nor U6236 (N_6236,In_2068,In_1185);
and U6237 (N_6237,In_110,In_2035);
or U6238 (N_6238,In_2344,In_1035);
and U6239 (N_6239,In_2195,In_2317);
and U6240 (N_6240,In_578,In_205);
and U6241 (N_6241,In_1481,In_251);
nor U6242 (N_6242,In_2541,In_2564);
and U6243 (N_6243,In_1685,In_1618);
or U6244 (N_6244,In_2614,In_2423);
nor U6245 (N_6245,In_1892,In_1563);
nand U6246 (N_6246,In_83,In_90);
and U6247 (N_6247,In_345,In_1255);
xnor U6248 (N_6248,In_1517,In_717);
nor U6249 (N_6249,In_1107,In_2545);
or U6250 (N_6250,In_2798,In_2126);
nand U6251 (N_6251,In_1380,In_2227);
or U6252 (N_6252,In_1955,In_1735);
xor U6253 (N_6253,In_1770,In_2573);
nand U6254 (N_6254,In_683,In_1447);
nor U6255 (N_6255,In_432,In_2002);
nor U6256 (N_6256,In_246,In_1932);
or U6257 (N_6257,In_695,In_288);
nand U6258 (N_6258,In_2355,In_2814);
nor U6259 (N_6259,In_2957,In_809);
xor U6260 (N_6260,In_2106,In_898);
nor U6261 (N_6261,In_2611,In_2413);
or U6262 (N_6262,In_427,In_2475);
and U6263 (N_6263,In_235,In_2862);
nand U6264 (N_6264,In_1887,In_2357);
or U6265 (N_6265,In_370,In_298);
nand U6266 (N_6266,In_1548,In_1091);
nand U6267 (N_6267,In_484,In_891);
nand U6268 (N_6268,In_1628,In_1929);
nand U6269 (N_6269,In_1051,In_2802);
or U6270 (N_6270,In_96,In_1872);
and U6271 (N_6271,In_2687,In_2096);
nand U6272 (N_6272,In_1686,In_1173);
nand U6273 (N_6273,In_2322,In_1847);
and U6274 (N_6274,In_635,In_1360);
nor U6275 (N_6275,In_37,In_1416);
or U6276 (N_6276,In_913,In_2172);
nand U6277 (N_6277,In_1351,In_364);
and U6278 (N_6278,In_2563,In_2778);
nor U6279 (N_6279,In_951,In_2427);
nand U6280 (N_6280,In_396,In_1658);
or U6281 (N_6281,In_735,In_1968);
xnor U6282 (N_6282,In_604,In_169);
nand U6283 (N_6283,In_1747,In_2785);
nand U6284 (N_6284,In_1241,In_1825);
or U6285 (N_6285,In_897,In_2982);
and U6286 (N_6286,In_2160,In_638);
nand U6287 (N_6287,In_11,In_790);
and U6288 (N_6288,In_74,In_214);
nor U6289 (N_6289,In_2428,In_15);
nor U6290 (N_6290,In_317,In_173);
or U6291 (N_6291,In_2484,In_483);
nand U6292 (N_6292,In_835,In_219);
xnor U6293 (N_6293,In_2916,In_173);
and U6294 (N_6294,In_131,In_16);
or U6295 (N_6295,In_1981,In_1563);
nor U6296 (N_6296,In_1951,In_384);
or U6297 (N_6297,In_625,In_2396);
xnor U6298 (N_6298,In_229,In_151);
or U6299 (N_6299,In_1104,In_1267);
nor U6300 (N_6300,In_332,In_233);
nor U6301 (N_6301,In_1172,In_1073);
and U6302 (N_6302,In_2725,In_1655);
and U6303 (N_6303,In_1954,In_2031);
and U6304 (N_6304,In_2240,In_1317);
or U6305 (N_6305,In_2182,In_41);
nand U6306 (N_6306,In_2263,In_2529);
and U6307 (N_6307,In_7,In_301);
nand U6308 (N_6308,In_2824,In_1116);
or U6309 (N_6309,In_2478,In_774);
or U6310 (N_6310,In_1301,In_2843);
nor U6311 (N_6311,In_2774,In_1565);
nor U6312 (N_6312,In_1569,In_1583);
or U6313 (N_6313,In_790,In_2343);
xnor U6314 (N_6314,In_935,In_2417);
nand U6315 (N_6315,In_330,In_2546);
nor U6316 (N_6316,In_1182,In_2339);
nor U6317 (N_6317,In_2913,In_763);
and U6318 (N_6318,In_1625,In_302);
and U6319 (N_6319,In_1684,In_455);
nand U6320 (N_6320,In_635,In_2543);
nor U6321 (N_6321,In_2060,In_1193);
or U6322 (N_6322,In_2794,In_914);
nor U6323 (N_6323,In_763,In_1327);
xor U6324 (N_6324,In_2546,In_1582);
nand U6325 (N_6325,In_1994,In_2088);
or U6326 (N_6326,In_1231,In_686);
nand U6327 (N_6327,In_1729,In_1449);
or U6328 (N_6328,In_116,In_948);
and U6329 (N_6329,In_1103,In_1318);
xor U6330 (N_6330,In_254,In_2797);
nor U6331 (N_6331,In_2061,In_2207);
and U6332 (N_6332,In_1928,In_1891);
or U6333 (N_6333,In_1211,In_2601);
nand U6334 (N_6334,In_2408,In_2830);
and U6335 (N_6335,In_1712,In_1923);
and U6336 (N_6336,In_2749,In_2276);
or U6337 (N_6337,In_834,In_1992);
nand U6338 (N_6338,In_2251,In_1858);
and U6339 (N_6339,In_359,In_898);
or U6340 (N_6340,In_75,In_783);
nand U6341 (N_6341,In_1673,In_2455);
or U6342 (N_6342,In_695,In_2541);
or U6343 (N_6343,In_2458,In_94);
xnor U6344 (N_6344,In_1766,In_2470);
or U6345 (N_6345,In_2548,In_2635);
xor U6346 (N_6346,In_915,In_417);
nor U6347 (N_6347,In_2451,In_717);
xor U6348 (N_6348,In_721,In_2755);
nand U6349 (N_6349,In_2949,In_1752);
nand U6350 (N_6350,In_680,In_1886);
xnor U6351 (N_6351,In_97,In_2683);
nand U6352 (N_6352,In_1385,In_258);
or U6353 (N_6353,In_2532,In_1116);
or U6354 (N_6354,In_2941,In_1923);
nand U6355 (N_6355,In_2857,In_2346);
nand U6356 (N_6356,In_2784,In_692);
or U6357 (N_6357,In_16,In_1410);
and U6358 (N_6358,In_2257,In_1080);
or U6359 (N_6359,In_1280,In_865);
nor U6360 (N_6360,In_735,In_2491);
nand U6361 (N_6361,In_2697,In_825);
or U6362 (N_6362,In_2519,In_11);
xnor U6363 (N_6363,In_2402,In_2382);
nor U6364 (N_6364,In_1672,In_701);
or U6365 (N_6365,In_2740,In_1816);
and U6366 (N_6366,In_2017,In_498);
nand U6367 (N_6367,In_289,In_1853);
nor U6368 (N_6368,In_867,In_2827);
xnor U6369 (N_6369,In_533,In_1860);
nor U6370 (N_6370,In_22,In_2554);
nor U6371 (N_6371,In_570,In_541);
or U6372 (N_6372,In_1370,In_662);
and U6373 (N_6373,In_1646,In_2375);
xor U6374 (N_6374,In_110,In_473);
or U6375 (N_6375,In_1049,In_718);
and U6376 (N_6376,In_1501,In_1966);
and U6377 (N_6377,In_4,In_2017);
nor U6378 (N_6378,In_302,In_1746);
and U6379 (N_6379,In_1093,In_795);
nor U6380 (N_6380,In_2685,In_2274);
or U6381 (N_6381,In_869,In_1653);
nand U6382 (N_6382,In_2925,In_606);
or U6383 (N_6383,In_15,In_1150);
or U6384 (N_6384,In_1426,In_2949);
xor U6385 (N_6385,In_125,In_701);
xnor U6386 (N_6386,In_2058,In_556);
nor U6387 (N_6387,In_1559,In_1635);
nor U6388 (N_6388,In_836,In_1187);
xnor U6389 (N_6389,In_1549,In_1343);
nand U6390 (N_6390,In_2550,In_2634);
nor U6391 (N_6391,In_2968,In_2896);
nor U6392 (N_6392,In_1897,In_2767);
or U6393 (N_6393,In_1311,In_1078);
nor U6394 (N_6394,In_1469,In_601);
xor U6395 (N_6395,In_334,In_1698);
nand U6396 (N_6396,In_128,In_1626);
nand U6397 (N_6397,In_2311,In_743);
nor U6398 (N_6398,In_2737,In_1067);
or U6399 (N_6399,In_2058,In_2351);
or U6400 (N_6400,In_286,In_97);
nand U6401 (N_6401,In_2727,In_2215);
and U6402 (N_6402,In_144,In_1003);
or U6403 (N_6403,In_1243,In_1917);
and U6404 (N_6404,In_575,In_1670);
and U6405 (N_6405,In_1975,In_291);
nor U6406 (N_6406,In_1595,In_2465);
nand U6407 (N_6407,In_330,In_329);
nor U6408 (N_6408,In_922,In_1673);
or U6409 (N_6409,In_2207,In_2368);
nor U6410 (N_6410,In_2312,In_2522);
nand U6411 (N_6411,In_1244,In_2311);
nor U6412 (N_6412,In_2640,In_1877);
nand U6413 (N_6413,In_1827,In_1466);
and U6414 (N_6414,In_2101,In_2472);
nand U6415 (N_6415,In_2695,In_168);
nor U6416 (N_6416,In_1130,In_1999);
nor U6417 (N_6417,In_1880,In_2028);
nor U6418 (N_6418,In_2720,In_1922);
or U6419 (N_6419,In_1304,In_2382);
and U6420 (N_6420,In_2233,In_1081);
or U6421 (N_6421,In_927,In_2808);
or U6422 (N_6422,In_965,In_466);
xnor U6423 (N_6423,In_230,In_1880);
and U6424 (N_6424,In_1255,In_1116);
and U6425 (N_6425,In_391,In_2563);
nand U6426 (N_6426,In_531,In_1796);
or U6427 (N_6427,In_2859,In_1026);
nand U6428 (N_6428,In_2629,In_1775);
nor U6429 (N_6429,In_1188,In_1236);
nor U6430 (N_6430,In_2894,In_1841);
nor U6431 (N_6431,In_723,In_497);
and U6432 (N_6432,In_103,In_1305);
and U6433 (N_6433,In_2313,In_1938);
or U6434 (N_6434,In_2688,In_1068);
nor U6435 (N_6435,In_1789,In_2337);
and U6436 (N_6436,In_1051,In_1220);
or U6437 (N_6437,In_1380,In_622);
nand U6438 (N_6438,In_2942,In_861);
and U6439 (N_6439,In_2915,In_582);
nor U6440 (N_6440,In_873,In_1442);
or U6441 (N_6441,In_1506,In_1676);
or U6442 (N_6442,In_2689,In_976);
or U6443 (N_6443,In_2559,In_2374);
nor U6444 (N_6444,In_1232,In_2884);
and U6445 (N_6445,In_445,In_1353);
or U6446 (N_6446,In_1089,In_2016);
and U6447 (N_6447,In_658,In_1532);
nand U6448 (N_6448,In_2623,In_328);
nor U6449 (N_6449,In_2150,In_1004);
nor U6450 (N_6450,In_2334,In_2173);
nor U6451 (N_6451,In_156,In_2493);
nand U6452 (N_6452,In_1667,In_1989);
or U6453 (N_6453,In_1015,In_2405);
nor U6454 (N_6454,In_885,In_2233);
and U6455 (N_6455,In_1359,In_2795);
nand U6456 (N_6456,In_1842,In_1849);
nand U6457 (N_6457,In_1366,In_1260);
and U6458 (N_6458,In_2090,In_592);
nor U6459 (N_6459,In_2724,In_408);
and U6460 (N_6460,In_329,In_52);
xor U6461 (N_6461,In_1304,In_338);
or U6462 (N_6462,In_1756,In_2643);
and U6463 (N_6463,In_498,In_643);
or U6464 (N_6464,In_958,In_1804);
xor U6465 (N_6465,In_797,In_2342);
and U6466 (N_6466,In_183,In_2160);
or U6467 (N_6467,In_1677,In_1488);
or U6468 (N_6468,In_2482,In_2688);
and U6469 (N_6469,In_485,In_1094);
nand U6470 (N_6470,In_1941,In_1259);
nor U6471 (N_6471,In_2024,In_2332);
nor U6472 (N_6472,In_1154,In_244);
nand U6473 (N_6473,In_1891,In_1464);
nand U6474 (N_6474,In_105,In_2954);
and U6475 (N_6475,In_2769,In_2467);
and U6476 (N_6476,In_2287,In_2735);
nor U6477 (N_6477,In_1185,In_2964);
or U6478 (N_6478,In_1765,In_305);
or U6479 (N_6479,In_2025,In_290);
xnor U6480 (N_6480,In_2937,In_1951);
nor U6481 (N_6481,In_447,In_518);
and U6482 (N_6482,In_327,In_585);
and U6483 (N_6483,In_1588,In_1355);
nor U6484 (N_6484,In_2172,In_2103);
or U6485 (N_6485,In_1707,In_740);
xor U6486 (N_6486,In_1189,In_1775);
nor U6487 (N_6487,In_170,In_1198);
nand U6488 (N_6488,In_723,In_1832);
nand U6489 (N_6489,In_2386,In_2700);
and U6490 (N_6490,In_1186,In_906);
nand U6491 (N_6491,In_1225,In_511);
nand U6492 (N_6492,In_576,In_2963);
nor U6493 (N_6493,In_1464,In_585);
nand U6494 (N_6494,In_2613,In_2361);
nand U6495 (N_6495,In_2395,In_2347);
nand U6496 (N_6496,In_2358,In_2645);
or U6497 (N_6497,In_1049,In_1085);
or U6498 (N_6498,In_1947,In_2206);
or U6499 (N_6499,In_371,In_714);
or U6500 (N_6500,In_2559,In_1028);
and U6501 (N_6501,In_42,In_41);
and U6502 (N_6502,In_847,In_2403);
nand U6503 (N_6503,In_1430,In_818);
and U6504 (N_6504,In_1826,In_99);
or U6505 (N_6505,In_1214,In_1014);
and U6506 (N_6506,In_2938,In_1078);
nor U6507 (N_6507,In_1493,In_2688);
xor U6508 (N_6508,In_839,In_1503);
and U6509 (N_6509,In_1693,In_2927);
and U6510 (N_6510,In_538,In_1406);
nand U6511 (N_6511,In_2540,In_468);
or U6512 (N_6512,In_1018,In_2111);
or U6513 (N_6513,In_1872,In_2926);
nand U6514 (N_6514,In_1533,In_1918);
nand U6515 (N_6515,In_275,In_2118);
or U6516 (N_6516,In_2022,In_754);
or U6517 (N_6517,In_775,In_809);
nand U6518 (N_6518,In_2206,In_585);
nand U6519 (N_6519,In_1571,In_1618);
nor U6520 (N_6520,In_1758,In_2720);
and U6521 (N_6521,In_2580,In_279);
and U6522 (N_6522,In_517,In_2355);
nor U6523 (N_6523,In_2828,In_2244);
and U6524 (N_6524,In_1002,In_1637);
xnor U6525 (N_6525,In_388,In_2427);
or U6526 (N_6526,In_584,In_2625);
nor U6527 (N_6527,In_639,In_164);
nor U6528 (N_6528,In_983,In_156);
xnor U6529 (N_6529,In_1688,In_2557);
or U6530 (N_6530,In_771,In_2628);
and U6531 (N_6531,In_2495,In_1030);
nor U6532 (N_6532,In_1382,In_460);
nor U6533 (N_6533,In_2650,In_1182);
nor U6534 (N_6534,In_2111,In_2507);
xor U6535 (N_6535,In_475,In_1514);
and U6536 (N_6536,In_2337,In_994);
or U6537 (N_6537,In_1443,In_1203);
or U6538 (N_6538,In_1440,In_527);
or U6539 (N_6539,In_1841,In_1967);
nand U6540 (N_6540,In_273,In_1474);
nand U6541 (N_6541,In_1760,In_607);
or U6542 (N_6542,In_1170,In_2828);
and U6543 (N_6543,In_1169,In_463);
xnor U6544 (N_6544,In_444,In_2064);
nor U6545 (N_6545,In_2664,In_512);
nor U6546 (N_6546,In_2795,In_2939);
and U6547 (N_6547,In_1812,In_938);
nor U6548 (N_6548,In_686,In_1251);
or U6549 (N_6549,In_1473,In_2822);
nand U6550 (N_6550,In_1070,In_2513);
xnor U6551 (N_6551,In_337,In_1562);
nand U6552 (N_6552,In_1403,In_2661);
nor U6553 (N_6553,In_2306,In_1258);
nor U6554 (N_6554,In_487,In_2531);
nand U6555 (N_6555,In_1488,In_2047);
or U6556 (N_6556,In_1398,In_1106);
xor U6557 (N_6557,In_672,In_2730);
nand U6558 (N_6558,In_141,In_854);
nand U6559 (N_6559,In_2105,In_1481);
and U6560 (N_6560,In_44,In_428);
or U6561 (N_6561,In_744,In_1348);
nor U6562 (N_6562,In_2474,In_129);
nand U6563 (N_6563,In_331,In_127);
nand U6564 (N_6564,In_603,In_1551);
nand U6565 (N_6565,In_2142,In_806);
nand U6566 (N_6566,In_2480,In_1986);
nand U6567 (N_6567,In_996,In_2708);
nor U6568 (N_6568,In_2265,In_775);
nor U6569 (N_6569,In_1154,In_496);
nor U6570 (N_6570,In_2449,In_320);
nor U6571 (N_6571,In_1397,In_679);
and U6572 (N_6572,In_2186,In_327);
xor U6573 (N_6573,In_2018,In_2933);
and U6574 (N_6574,In_2612,In_653);
or U6575 (N_6575,In_1145,In_56);
or U6576 (N_6576,In_1201,In_2271);
nand U6577 (N_6577,In_196,In_778);
nand U6578 (N_6578,In_2310,In_508);
or U6579 (N_6579,In_2457,In_1483);
or U6580 (N_6580,In_511,In_2227);
nand U6581 (N_6581,In_965,In_932);
and U6582 (N_6582,In_1243,In_1315);
nand U6583 (N_6583,In_1266,In_527);
nand U6584 (N_6584,In_216,In_2446);
or U6585 (N_6585,In_818,In_2954);
and U6586 (N_6586,In_1882,In_216);
xnor U6587 (N_6587,In_242,In_2624);
and U6588 (N_6588,In_2625,In_2057);
nand U6589 (N_6589,In_2408,In_2502);
nor U6590 (N_6590,In_103,In_278);
nand U6591 (N_6591,In_789,In_2187);
or U6592 (N_6592,In_2324,In_1691);
or U6593 (N_6593,In_2779,In_1574);
nand U6594 (N_6594,In_2645,In_1338);
or U6595 (N_6595,In_889,In_25);
nor U6596 (N_6596,In_554,In_2186);
nand U6597 (N_6597,In_1740,In_2828);
xor U6598 (N_6598,In_209,In_1896);
nor U6599 (N_6599,In_282,In_1246);
and U6600 (N_6600,In_202,In_2841);
nand U6601 (N_6601,In_1529,In_933);
or U6602 (N_6602,In_163,In_1307);
and U6603 (N_6603,In_1074,In_2325);
or U6604 (N_6604,In_807,In_1942);
nor U6605 (N_6605,In_618,In_2019);
and U6606 (N_6606,In_2212,In_426);
and U6607 (N_6607,In_2406,In_1864);
nand U6608 (N_6608,In_1677,In_1619);
nand U6609 (N_6609,In_1976,In_496);
nand U6610 (N_6610,In_1760,In_1201);
xor U6611 (N_6611,In_270,In_1278);
or U6612 (N_6612,In_876,In_1290);
and U6613 (N_6613,In_274,In_1078);
and U6614 (N_6614,In_2927,In_1704);
and U6615 (N_6615,In_1748,In_1719);
nand U6616 (N_6616,In_1087,In_250);
nor U6617 (N_6617,In_1010,In_1692);
or U6618 (N_6618,In_1166,In_896);
or U6619 (N_6619,In_2885,In_2029);
or U6620 (N_6620,In_2782,In_364);
xor U6621 (N_6621,In_2941,In_2878);
nand U6622 (N_6622,In_419,In_2465);
nor U6623 (N_6623,In_38,In_2988);
xor U6624 (N_6624,In_359,In_1999);
nor U6625 (N_6625,In_2470,In_2350);
nor U6626 (N_6626,In_1093,In_349);
nor U6627 (N_6627,In_1185,In_2567);
and U6628 (N_6628,In_1728,In_2183);
nor U6629 (N_6629,In_125,In_755);
or U6630 (N_6630,In_2041,In_951);
nand U6631 (N_6631,In_1825,In_355);
nand U6632 (N_6632,In_1103,In_2332);
nor U6633 (N_6633,In_2603,In_375);
nor U6634 (N_6634,In_230,In_54);
xor U6635 (N_6635,In_900,In_2959);
nand U6636 (N_6636,In_2415,In_2459);
nor U6637 (N_6637,In_2648,In_1847);
nand U6638 (N_6638,In_2219,In_1980);
and U6639 (N_6639,In_575,In_667);
and U6640 (N_6640,In_2600,In_876);
nand U6641 (N_6641,In_1394,In_1665);
nor U6642 (N_6642,In_2632,In_1198);
nor U6643 (N_6643,In_2646,In_210);
and U6644 (N_6644,In_1348,In_149);
and U6645 (N_6645,In_2467,In_2581);
nand U6646 (N_6646,In_2377,In_2082);
nor U6647 (N_6647,In_1677,In_2666);
nand U6648 (N_6648,In_1192,In_2846);
nor U6649 (N_6649,In_1443,In_2764);
and U6650 (N_6650,In_2727,In_2835);
nand U6651 (N_6651,In_2137,In_1790);
nor U6652 (N_6652,In_1824,In_1498);
xor U6653 (N_6653,In_236,In_2671);
and U6654 (N_6654,In_821,In_2379);
nor U6655 (N_6655,In_1364,In_396);
and U6656 (N_6656,In_2635,In_2775);
nand U6657 (N_6657,In_220,In_1983);
and U6658 (N_6658,In_1136,In_1944);
and U6659 (N_6659,In_218,In_2845);
nand U6660 (N_6660,In_1494,In_2022);
nand U6661 (N_6661,In_747,In_305);
nor U6662 (N_6662,In_994,In_1913);
or U6663 (N_6663,In_2134,In_2700);
or U6664 (N_6664,In_530,In_1877);
xnor U6665 (N_6665,In_1952,In_2818);
xor U6666 (N_6666,In_454,In_1484);
xor U6667 (N_6667,In_1159,In_2192);
or U6668 (N_6668,In_2145,In_2268);
nand U6669 (N_6669,In_2804,In_2853);
xnor U6670 (N_6670,In_2213,In_1385);
or U6671 (N_6671,In_364,In_1734);
nand U6672 (N_6672,In_2148,In_853);
and U6673 (N_6673,In_2901,In_2571);
nor U6674 (N_6674,In_911,In_2950);
and U6675 (N_6675,In_1504,In_499);
and U6676 (N_6676,In_177,In_1571);
or U6677 (N_6677,In_2337,In_1524);
nand U6678 (N_6678,In_663,In_1688);
nand U6679 (N_6679,In_1518,In_212);
nand U6680 (N_6680,In_2204,In_2492);
nand U6681 (N_6681,In_526,In_438);
and U6682 (N_6682,In_1016,In_2847);
and U6683 (N_6683,In_2374,In_1006);
or U6684 (N_6684,In_180,In_1622);
nor U6685 (N_6685,In_579,In_2672);
xnor U6686 (N_6686,In_79,In_896);
or U6687 (N_6687,In_1659,In_1798);
and U6688 (N_6688,In_1149,In_1728);
nand U6689 (N_6689,In_1188,In_979);
and U6690 (N_6690,In_2317,In_601);
nor U6691 (N_6691,In_1835,In_1071);
nor U6692 (N_6692,In_440,In_603);
and U6693 (N_6693,In_1652,In_2937);
or U6694 (N_6694,In_2174,In_1374);
xor U6695 (N_6695,In_2260,In_1862);
and U6696 (N_6696,In_315,In_2669);
and U6697 (N_6697,In_2797,In_1403);
and U6698 (N_6698,In_393,In_546);
nand U6699 (N_6699,In_1620,In_1855);
and U6700 (N_6700,In_2225,In_2759);
nor U6701 (N_6701,In_1613,In_2368);
or U6702 (N_6702,In_2027,In_856);
and U6703 (N_6703,In_1007,In_1353);
nand U6704 (N_6704,In_1349,In_155);
and U6705 (N_6705,In_1180,In_812);
xor U6706 (N_6706,In_346,In_2744);
nand U6707 (N_6707,In_291,In_2534);
nand U6708 (N_6708,In_1516,In_1275);
and U6709 (N_6709,In_279,In_843);
and U6710 (N_6710,In_45,In_2872);
or U6711 (N_6711,In_2720,In_354);
nor U6712 (N_6712,In_2265,In_104);
xor U6713 (N_6713,In_408,In_2649);
and U6714 (N_6714,In_1800,In_2450);
nand U6715 (N_6715,In_975,In_1187);
or U6716 (N_6716,In_1437,In_2626);
and U6717 (N_6717,In_1455,In_2805);
or U6718 (N_6718,In_1728,In_2553);
nor U6719 (N_6719,In_800,In_1062);
and U6720 (N_6720,In_1961,In_1671);
xor U6721 (N_6721,In_2203,In_2024);
nor U6722 (N_6722,In_1977,In_660);
and U6723 (N_6723,In_866,In_1246);
or U6724 (N_6724,In_2247,In_2099);
and U6725 (N_6725,In_1267,In_549);
nor U6726 (N_6726,In_1326,In_608);
or U6727 (N_6727,In_826,In_1481);
nor U6728 (N_6728,In_823,In_1669);
and U6729 (N_6729,In_1254,In_1308);
nand U6730 (N_6730,In_2921,In_1406);
and U6731 (N_6731,In_2133,In_469);
nand U6732 (N_6732,In_646,In_1206);
nand U6733 (N_6733,In_207,In_2725);
and U6734 (N_6734,In_177,In_1260);
xnor U6735 (N_6735,In_1660,In_511);
or U6736 (N_6736,In_1432,In_510);
nor U6737 (N_6737,In_1561,In_2755);
or U6738 (N_6738,In_1098,In_1620);
or U6739 (N_6739,In_272,In_1695);
xnor U6740 (N_6740,In_2756,In_2575);
nor U6741 (N_6741,In_2869,In_2635);
nor U6742 (N_6742,In_1039,In_2307);
and U6743 (N_6743,In_990,In_11);
and U6744 (N_6744,In_2178,In_1933);
and U6745 (N_6745,In_1987,In_503);
or U6746 (N_6746,In_2822,In_355);
nand U6747 (N_6747,In_1466,In_2267);
and U6748 (N_6748,In_1582,In_541);
nor U6749 (N_6749,In_1775,In_266);
and U6750 (N_6750,In_2564,In_112);
nand U6751 (N_6751,In_566,In_1096);
and U6752 (N_6752,In_2802,In_1626);
or U6753 (N_6753,In_2753,In_1897);
nor U6754 (N_6754,In_322,In_1307);
and U6755 (N_6755,In_21,In_1314);
and U6756 (N_6756,In_1809,In_1818);
nand U6757 (N_6757,In_797,In_1762);
nor U6758 (N_6758,In_1514,In_191);
and U6759 (N_6759,In_2795,In_727);
and U6760 (N_6760,In_1784,In_776);
xor U6761 (N_6761,In_1501,In_775);
nand U6762 (N_6762,In_1035,In_833);
and U6763 (N_6763,In_972,In_2627);
nand U6764 (N_6764,In_2162,In_1047);
nor U6765 (N_6765,In_245,In_1600);
nor U6766 (N_6766,In_521,In_2095);
nor U6767 (N_6767,In_124,In_2166);
and U6768 (N_6768,In_2095,In_636);
or U6769 (N_6769,In_935,In_247);
nand U6770 (N_6770,In_2507,In_1274);
nor U6771 (N_6771,In_370,In_1075);
or U6772 (N_6772,In_1271,In_2914);
or U6773 (N_6773,In_2477,In_2779);
xor U6774 (N_6774,In_2207,In_1069);
and U6775 (N_6775,In_2635,In_1969);
nor U6776 (N_6776,In_2865,In_1413);
nand U6777 (N_6777,In_2764,In_2844);
nor U6778 (N_6778,In_1226,In_2665);
and U6779 (N_6779,In_1960,In_1742);
nor U6780 (N_6780,In_329,In_624);
and U6781 (N_6781,In_2524,In_554);
nor U6782 (N_6782,In_2864,In_17);
nor U6783 (N_6783,In_2869,In_2908);
and U6784 (N_6784,In_1872,In_2918);
nor U6785 (N_6785,In_2528,In_2852);
nand U6786 (N_6786,In_818,In_1054);
nand U6787 (N_6787,In_2690,In_2641);
and U6788 (N_6788,In_1925,In_2819);
and U6789 (N_6789,In_2807,In_2308);
nand U6790 (N_6790,In_67,In_1157);
nand U6791 (N_6791,In_20,In_1483);
and U6792 (N_6792,In_1673,In_1973);
or U6793 (N_6793,In_2962,In_693);
and U6794 (N_6794,In_612,In_2558);
or U6795 (N_6795,In_636,In_838);
and U6796 (N_6796,In_428,In_473);
xnor U6797 (N_6797,In_1986,In_1663);
and U6798 (N_6798,In_2803,In_2913);
and U6799 (N_6799,In_2260,In_261);
or U6800 (N_6800,In_1384,In_2109);
or U6801 (N_6801,In_2759,In_1303);
or U6802 (N_6802,In_2379,In_2365);
and U6803 (N_6803,In_2260,In_709);
nor U6804 (N_6804,In_360,In_8);
nand U6805 (N_6805,In_887,In_1037);
and U6806 (N_6806,In_1689,In_917);
and U6807 (N_6807,In_1065,In_1355);
nand U6808 (N_6808,In_409,In_827);
nand U6809 (N_6809,In_2313,In_2855);
and U6810 (N_6810,In_510,In_1224);
nand U6811 (N_6811,In_498,In_683);
nor U6812 (N_6812,In_1435,In_945);
nor U6813 (N_6813,In_1771,In_2876);
nand U6814 (N_6814,In_652,In_123);
or U6815 (N_6815,In_1594,In_1947);
nand U6816 (N_6816,In_839,In_172);
and U6817 (N_6817,In_552,In_1214);
nor U6818 (N_6818,In_787,In_1987);
nand U6819 (N_6819,In_2285,In_1901);
xnor U6820 (N_6820,In_824,In_1190);
or U6821 (N_6821,In_36,In_975);
nand U6822 (N_6822,In_2940,In_1359);
and U6823 (N_6823,In_623,In_2481);
and U6824 (N_6824,In_178,In_1366);
nor U6825 (N_6825,In_101,In_1068);
nor U6826 (N_6826,In_1138,In_939);
or U6827 (N_6827,In_96,In_2954);
xor U6828 (N_6828,In_639,In_2502);
nand U6829 (N_6829,In_2648,In_723);
or U6830 (N_6830,In_619,In_872);
and U6831 (N_6831,In_503,In_2114);
or U6832 (N_6832,In_1421,In_391);
and U6833 (N_6833,In_37,In_274);
nor U6834 (N_6834,In_1204,In_582);
nand U6835 (N_6835,In_56,In_2916);
or U6836 (N_6836,In_16,In_2907);
and U6837 (N_6837,In_1758,In_2427);
xnor U6838 (N_6838,In_2018,In_1292);
nand U6839 (N_6839,In_1341,In_2317);
or U6840 (N_6840,In_46,In_979);
xor U6841 (N_6841,In_2720,In_198);
nor U6842 (N_6842,In_2290,In_2733);
nor U6843 (N_6843,In_2672,In_2300);
and U6844 (N_6844,In_264,In_2772);
nand U6845 (N_6845,In_111,In_2058);
nor U6846 (N_6846,In_2720,In_1364);
nand U6847 (N_6847,In_465,In_2356);
and U6848 (N_6848,In_998,In_1715);
nor U6849 (N_6849,In_331,In_539);
nor U6850 (N_6850,In_1746,In_1529);
and U6851 (N_6851,In_1256,In_2002);
or U6852 (N_6852,In_1083,In_1998);
xnor U6853 (N_6853,In_1238,In_2083);
nor U6854 (N_6854,In_1583,In_662);
xor U6855 (N_6855,In_902,In_1581);
nor U6856 (N_6856,In_2074,In_826);
and U6857 (N_6857,In_863,In_868);
xor U6858 (N_6858,In_2094,In_2789);
and U6859 (N_6859,In_2747,In_2366);
or U6860 (N_6860,In_962,In_410);
or U6861 (N_6861,In_524,In_94);
xor U6862 (N_6862,In_883,In_2852);
or U6863 (N_6863,In_441,In_2499);
or U6864 (N_6864,In_2270,In_2110);
xnor U6865 (N_6865,In_1222,In_1987);
nand U6866 (N_6866,In_1332,In_2716);
nor U6867 (N_6867,In_1971,In_2473);
nand U6868 (N_6868,In_1546,In_1773);
nor U6869 (N_6869,In_2439,In_2776);
nand U6870 (N_6870,In_76,In_1861);
nor U6871 (N_6871,In_63,In_2058);
nor U6872 (N_6872,In_1190,In_94);
and U6873 (N_6873,In_2856,In_1313);
xor U6874 (N_6874,In_1981,In_544);
xnor U6875 (N_6875,In_952,In_1629);
and U6876 (N_6876,In_2283,In_268);
and U6877 (N_6877,In_2362,In_2692);
nor U6878 (N_6878,In_1091,In_1568);
nor U6879 (N_6879,In_38,In_2697);
or U6880 (N_6880,In_586,In_274);
and U6881 (N_6881,In_735,In_547);
or U6882 (N_6882,In_2087,In_2965);
nor U6883 (N_6883,In_28,In_1111);
nor U6884 (N_6884,In_2767,In_2362);
nand U6885 (N_6885,In_2978,In_2301);
nor U6886 (N_6886,In_1818,In_1210);
and U6887 (N_6887,In_1874,In_934);
or U6888 (N_6888,In_2607,In_2774);
or U6889 (N_6889,In_1122,In_2268);
nand U6890 (N_6890,In_1235,In_1802);
nand U6891 (N_6891,In_431,In_458);
or U6892 (N_6892,In_2170,In_825);
nor U6893 (N_6893,In_247,In_2121);
nand U6894 (N_6894,In_2755,In_251);
nor U6895 (N_6895,In_1013,In_2406);
nand U6896 (N_6896,In_2369,In_243);
nor U6897 (N_6897,In_2772,In_1581);
nand U6898 (N_6898,In_1618,In_1551);
or U6899 (N_6899,In_1533,In_284);
xnor U6900 (N_6900,In_1807,In_1936);
nand U6901 (N_6901,In_670,In_2423);
xor U6902 (N_6902,In_847,In_2122);
nor U6903 (N_6903,In_17,In_1601);
or U6904 (N_6904,In_2925,In_181);
xor U6905 (N_6905,In_2122,In_1584);
and U6906 (N_6906,In_1153,In_756);
xor U6907 (N_6907,In_15,In_218);
nand U6908 (N_6908,In_1528,In_1311);
nand U6909 (N_6909,In_1705,In_1236);
or U6910 (N_6910,In_59,In_601);
xor U6911 (N_6911,In_2489,In_2843);
xor U6912 (N_6912,In_948,In_1858);
nor U6913 (N_6913,In_2716,In_55);
nor U6914 (N_6914,In_1138,In_1299);
and U6915 (N_6915,In_1262,In_880);
and U6916 (N_6916,In_2259,In_1516);
nor U6917 (N_6917,In_2825,In_430);
nor U6918 (N_6918,In_1090,In_422);
nor U6919 (N_6919,In_2077,In_1208);
or U6920 (N_6920,In_996,In_1322);
xor U6921 (N_6921,In_2474,In_1284);
and U6922 (N_6922,In_630,In_513);
and U6923 (N_6923,In_175,In_493);
nand U6924 (N_6924,In_605,In_1900);
and U6925 (N_6925,In_1110,In_2255);
nand U6926 (N_6926,In_2675,In_818);
nand U6927 (N_6927,In_2023,In_1181);
or U6928 (N_6928,In_2533,In_1249);
or U6929 (N_6929,In_1133,In_2433);
nor U6930 (N_6930,In_1827,In_1579);
nand U6931 (N_6931,In_1005,In_1167);
and U6932 (N_6932,In_1177,In_2403);
nand U6933 (N_6933,In_290,In_2935);
nand U6934 (N_6934,In_1957,In_1805);
or U6935 (N_6935,In_1966,In_2207);
or U6936 (N_6936,In_63,In_803);
nor U6937 (N_6937,In_497,In_1346);
and U6938 (N_6938,In_1314,In_1593);
nand U6939 (N_6939,In_1138,In_384);
nor U6940 (N_6940,In_1942,In_2231);
nor U6941 (N_6941,In_1445,In_2440);
or U6942 (N_6942,In_802,In_1694);
or U6943 (N_6943,In_1748,In_316);
nor U6944 (N_6944,In_354,In_1461);
nand U6945 (N_6945,In_2247,In_1428);
and U6946 (N_6946,In_2719,In_2669);
nor U6947 (N_6947,In_667,In_1962);
or U6948 (N_6948,In_2800,In_1077);
and U6949 (N_6949,In_2244,In_1045);
nor U6950 (N_6950,In_658,In_1809);
nand U6951 (N_6951,In_2434,In_1872);
nor U6952 (N_6952,In_2150,In_168);
nor U6953 (N_6953,In_2403,In_2262);
and U6954 (N_6954,In_1718,In_489);
nand U6955 (N_6955,In_167,In_606);
xor U6956 (N_6956,In_2445,In_1832);
nand U6957 (N_6957,In_1102,In_602);
nor U6958 (N_6958,In_2929,In_1891);
or U6959 (N_6959,In_1526,In_1173);
nand U6960 (N_6960,In_1927,In_1468);
or U6961 (N_6961,In_126,In_61);
nand U6962 (N_6962,In_1252,In_2481);
nand U6963 (N_6963,In_168,In_2630);
nand U6964 (N_6964,In_1123,In_2177);
nor U6965 (N_6965,In_2306,In_1724);
xnor U6966 (N_6966,In_335,In_2522);
nand U6967 (N_6967,In_748,In_1639);
nand U6968 (N_6968,In_1588,In_1818);
or U6969 (N_6969,In_2561,In_2598);
xnor U6970 (N_6970,In_1482,In_1322);
or U6971 (N_6971,In_1699,In_456);
and U6972 (N_6972,In_431,In_2593);
or U6973 (N_6973,In_1552,In_1628);
nor U6974 (N_6974,In_717,In_2804);
or U6975 (N_6975,In_854,In_1691);
and U6976 (N_6976,In_477,In_2166);
xor U6977 (N_6977,In_1057,In_1493);
nor U6978 (N_6978,In_385,In_2440);
and U6979 (N_6979,In_2627,In_2898);
xnor U6980 (N_6980,In_2055,In_2670);
nor U6981 (N_6981,In_1487,In_1270);
nor U6982 (N_6982,In_342,In_28);
nand U6983 (N_6983,In_2999,In_1642);
or U6984 (N_6984,In_1003,In_1531);
or U6985 (N_6985,In_2324,In_2633);
nand U6986 (N_6986,In_2522,In_115);
nor U6987 (N_6987,In_1370,In_1808);
nand U6988 (N_6988,In_719,In_537);
nor U6989 (N_6989,In_2729,In_2085);
nor U6990 (N_6990,In_1243,In_2342);
nand U6991 (N_6991,In_571,In_2199);
nor U6992 (N_6992,In_1359,In_715);
or U6993 (N_6993,In_1712,In_2717);
or U6994 (N_6994,In_2779,In_442);
nor U6995 (N_6995,In_185,In_2907);
and U6996 (N_6996,In_1266,In_2973);
or U6997 (N_6997,In_1579,In_580);
nand U6998 (N_6998,In_1722,In_2199);
and U6999 (N_6999,In_2192,In_1487);
and U7000 (N_7000,In_1475,In_2857);
or U7001 (N_7001,In_2291,In_2147);
nor U7002 (N_7002,In_638,In_2514);
nor U7003 (N_7003,In_901,In_2039);
and U7004 (N_7004,In_2259,In_816);
and U7005 (N_7005,In_1674,In_114);
and U7006 (N_7006,In_50,In_1581);
nand U7007 (N_7007,In_1963,In_1149);
or U7008 (N_7008,In_851,In_2449);
and U7009 (N_7009,In_1553,In_123);
xnor U7010 (N_7010,In_412,In_2090);
nand U7011 (N_7011,In_1696,In_733);
nand U7012 (N_7012,In_179,In_1031);
nand U7013 (N_7013,In_647,In_324);
nand U7014 (N_7014,In_1486,In_1270);
and U7015 (N_7015,In_1752,In_2072);
or U7016 (N_7016,In_726,In_1840);
nor U7017 (N_7017,In_2312,In_2547);
and U7018 (N_7018,In_1597,In_2634);
nor U7019 (N_7019,In_1099,In_2410);
or U7020 (N_7020,In_1066,In_1860);
and U7021 (N_7021,In_331,In_1422);
and U7022 (N_7022,In_1993,In_2382);
xnor U7023 (N_7023,In_2298,In_2028);
nor U7024 (N_7024,In_1142,In_765);
and U7025 (N_7025,In_1286,In_291);
or U7026 (N_7026,In_1908,In_2290);
or U7027 (N_7027,In_1750,In_696);
nor U7028 (N_7028,In_1083,In_740);
and U7029 (N_7029,In_1226,In_1355);
nor U7030 (N_7030,In_2475,In_274);
or U7031 (N_7031,In_728,In_1534);
and U7032 (N_7032,In_1187,In_1165);
nand U7033 (N_7033,In_668,In_1838);
nor U7034 (N_7034,In_1413,In_1617);
nor U7035 (N_7035,In_149,In_2754);
and U7036 (N_7036,In_765,In_2113);
nand U7037 (N_7037,In_1149,In_2677);
nand U7038 (N_7038,In_2732,In_2132);
and U7039 (N_7039,In_2744,In_1724);
nand U7040 (N_7040,In_547,In_2458);
and U7041 (N_7041,In_693,In_1672);
or U7042 (N_7042,In_2156,In_2887);
or U7043 (N_7043,In_2763,In_1382);
nor U7044 (N_7044,In_2906,In_1167);
or U7045 (N_7045,In_981,In_1786);
xor U7046 (N_7046,In_2656,In_2174);
and U7047 (N_7047,In_1445,In_564);
xor U7048 (N_7048,In_125,In_1159);
nand U7049 (N_7049,In_2095,In_2582);
nor U7050 (N_7050,In_1798,In_1368);
nand U7051 (N_7051,In_1158,In_2553);
nor U7052 (N_7052,In_656,In_1819);
and U7053 (N_7053,In_1673,In_2443);
nand U7054 (N_7054,In_2650,In_2952);
nand U7055 (N_7055,In_1263,In_2319);
nand U7056 (N_7056,In_689,In_2493);
nor U7057 (N_7057,In_749,In_2806);
or U7058 (N_7058,In_632,In_1304);
xnor U7059 (N_7059,In_2382,In_641);
nor U7060 (N_7060,In_1105,In_1047);
or U7061 (N_7061,In_517,In_1637);
nand U7062 (N_7062,In_1722,In_1029);
nor U7063 (N_7063,In_2570,In_2103);
xor U7064 (N_7064,In_2787,In_2874);
nor U7065 (N_7065,In_2694,In_510);
nor U7066 (N_7066,In_2728,In_2509);
xor U7067 (N_7067,In_2754,In_1785);
xnor U7068 (N_7068,In_220,In_1927);
xor U7069 (N_7069,In_502,In_2907);
nor U7070 (N_7070,In_1070,In_2497);
and U7071 (N_7071,In_2993,In_1129);
nand U7072 (N_7072,In_2403,In_1791);
nor U7073 (N_7073,In_564,In_995);
nand U7074 (N_7074,In_228,In_2010);
nand U7075 (N_7075,In_2961,In_2850);
or U7076 (N_7076,In_9,In_452);
nor U7077 (N_7077,In_793,In_1484);
nor U7078 (N_7078,In_815,In_655);
nand U7079 (N_7079,In_395,In_361);
and U7080 (N_7080,In_531,In_1286);
nand U7081 (N_7081,In_1899,In_1916);
xor U7082 (N_7082,In_2117,In_2542);
and U7083 (N_7083,In_2489,In_2896);
nor U7084 (N_7084,In_1629,In_2574);
xnor U7085 (N_7085,In_818,In_1456);
and U7086 (N_7086,In_2956,In_613);
nor U7087 (N_7087,In_1084,In_7);
nand U7088 (N_7088,In_2875,In_2619);
nor U7089 (N_7089,In_2594,In_80);
nand U7090 (N_7090,In_1003,In_723);
nand U7091 (N_7091,In_136,In_1086);
and U7092 (N_7092,In_1078,In_2431);
or U7093 (N_7093,In_1559,In_1493);
or U7094 (N_7094,In_1988,In_286);
xnor U7095 (N_7095,In_2040,In_426);
and U7096 (N_7096,In_101,In_1199);
nor U7097 (N_7097,In_670,In_734);
or U7098 (N_7098,In_1600,In_615);
xor U7099 (N_7099,In_1902,In_2857);
and U7100 (N_7100,In_867,In_2657);
nor U7101 (N_7101,In_1119,In_2709);
nand U7102 (N_7102,In_2504,In_1495);
and U7103 (N_7103,In_2765,In_1629);
or U7104 (N_7104,In_1652,In_2076);
nor U7105 (N_7105,In_2016,In_2403);
nor U7106 (N_7106,In_2339,In_2117);
and U7107 (N_7107,In_2980,In_925);
and U7108 (N_7108,In_1882,In_2087);
and U7109 (N_7109,In_2500,In_2069);
nand U7110 (N_7110,In_1005,In_2081);
or U7111 (N_7111,In_622,In_6);
and U7112 (N_7112,In_759,In_1979);
or U7113 (N_7113,In_1462,In_692);
nand U7114 (N_7114,In_1652,In_1426);
or U7115 (N_7115,In_942,In_207);
or U7116 (N_7116,In_1540,In_1608);
xor U7117 (N_7117,In_1845,In_2491);
or U7118 (N_7118,In_2203,In_2646);
or U7119 (N_7119,In_2624,In_1889);
and U7120 (N_7120,In_1117,In_2365);
and U7121 (N_7121,In_727,In_2505);
xnor U7122 (N_7122,In_1441,In_158);
nand U7123 (N_7123,In_326,In_2180);
xor U7124 (N_7124,In_1329,In_2601);
or U7125 (N_7125,In_1368,In_385);
and U7126 (N_7126,In_1549,In_1411);
nor U7127 (N_7127,In_2752,In_1907);
nand U7128 (N_7128,In_2615,In_1053);
nor U7129 (N_7129,In_1995,In_2786);
xnor U7130 (N_7130,In_2455,In_1494);
nor U7131 (N_7131,In_193,In_2798);
nor U7132 (N_7132,In_93,In_2130);
and U7133 (N_7133,In_2282,In_2410);
or U7134 (N_7134,In_2340,In_2893);
or U7135 (N_7135,In_994,In_2459);
xor U7136 (N_7136,In_625,In_2331);
nor U7137 (N_7137,In_1403,In_2387);
xnor U7138 (N_7138,In_2940,In_1545);
nor U7139 (N_7139,In_1962,In_2801);
and U7140 (N_7140,In_226,In_2147);
or U7141 (N_7141,In_667,In_2243);
nand U7142 (N_7142,In_771,In_2905);
xnor U7143 (N_7143,In_1971,In_1555);
nand U7144 (N_7144,In_1984,In_1618);
nor U7145 (N_7145,In_1414,In_1475);
nand U7146 (N_7146,In_890,In_2920);
nand U7147 (N_7147,In_2233,In_2137);
and U7148 (N_7148,In_2315,In_1621);
or U7149 (N_7149,In_1880,In_1849);
nor U7150 (N_7150,In_1004,In_2273);
nor U7151 (N_7151,In_47,In_2201);
and U7152 (N_7152,In_611,In_1406);
nand U7153 (N_7153,In_2155,In_1343);
nand U7154 (N_7154,In_509,In_2494);
nor U7155 (N_7155,In_2428,In_276);
nor U7156 (N_7156,In_2997,In_2083);
xor U7157 (N_7157,In_2940,In_2879);
and U7158 (N_7158,In_325,In_2467);
nand U7159 (N_7159,In_674,In_2585);
nand U7160 (N_7160,In_1222,In_2326);
and U7161 (N_7161,In_1454,In_811);
or U7162 (N_7162,In_2314,In_2194);
and U7163 (N_7163,In_2371,In_926);
and U7164 (N_7164,In_179,In_309);
xor U7165 (N_7165,In_1678,In_2769);
nand U7166 (N_7166,In_860,In_2833);
nor U7167 (N_7167,In_1411,In_2679);
or U7168 (N_7168,In_1553,In_2420);
or U7169 (N_7169,In_546,In_2642);
nor U7170 (N_7170,In_145,In_2625);
and U7171 (N_7171,In_700,In_1161);
nor U7172 (N_7172,In_1401,In_1330);
nor U7173 (N_7173,In_298,In_755);
or U7174 (N_7174,In_1332,In_1548);
xnor U7175 (N_7175,In_1684,In_1265);
and U7176 (N_7176,In_1229,In_656);
xnor U7177 (N_7177,In_1102,In_2286);
and U7178 (N_7178,In_741,In_1117);
nand U7179 (N_7179,In_2014,In_268);
nor U7180 (N_7180,In_2396,In_1122);
nor U7181 (N_7181,In_995,In_2318);
xnor U7182 (N_7182,In_624,In_1146);
nand U7183 (N_7183,In_1864,In_360);
xor U7184 (N_7184,In_2438,In_1332);
or U7185 (N_7185,In_461,In_2934);
nor U7186 (N_7186,In_1316,In_1687);
xnor U7187 (N_7187,In_1676,In_2742);
nand U7188 (N_7188,In_87,In_2322);
and U7189 (N_7189,In_2956,In_1621);
or U7190 (N_7190,In_1066,In_2934);
nor U7191 (N_7191,In_443,In_2070);
nand U7192 (N_7192,In_2529,In_2800);
and U7193 (N_7193,In_671,In_583);
or U7194 (N_7194,In_2352,In_2946);
nand U7195 (N_7195,In_1705,In_2113);
or U7196 (N_7196,In_2399,In_1570);
nand U7197 (N_7197,In_2346,In_412);
and U7198 (N_7198,In_1726,In_1255);
xnor U7199 (N_7199,In_738,In_25);
nor U7200 (N_7200,In_2820,In_2307);
or U7201 (N_7201,In_2884,In_2470);
xnor U7202 (N_7202,In_2481,In_445);
nand U7203 (N_7203,In_2627,In_765);
nor U7204 (N_7204,In_2568,In_1308);
and U7205 (N_7205,In_1178,In_1887);
xor U7206 (N_7206,In_7,In_1733);
or U7207 (N_7207,In_2374,In_2300);
xnor U7208 (N_7208,In_266,In_984);
or U7209 (N_7209,In_115,In_2012);
and U7210 (N_7210,In_519,In_594);
nor U7211 (N_7211,In_2012,In_2622);
or U7212 (N_7212,In_285,In_1219);
xnor U7213 (N_7213,In_697,In_777);
xor U7214 (N_7214,In_2924,In_2916);
xor U7215 (N_7215,In_2728,In_1166);
or U7216 (N_7216,In_989,In_2593);
nand U7217 (N_7217,In_837,In_2887);
or U7218 (N_7218,In_685,In_641);
nor U7219 (N_7219,In_127,In_2958);
nor U7220 (N_7220,In_1268,In_331);
xor U7221 (N_7221,In_1286,In_1394);
nor U7222 (N_7222,In_1607,In_106);
and U7223 (N_7223,In_1438,In_2484);
or U7224 (N_7224,In_2018,In_2559);
or U7225 (N_7225,In_931,In_778);
nand U7226 (N_7226,In_625,In_47);
and U7227 (N_7227,In_1902,In_144);
nand U7228 (N_7228,In_1486,In_236);
xnor U7229 (N_7229,In_272,In_2814);
nand U7230 (N_7230,In_1160,In_105);
and U7231 (N_7231,In_1921,In_1024);
or U7232 (N_7232,In_2520,In_2907);
and U7233 (N_7233,In_1523,In_2984);
or U7234 (N_7234,In_1411,In_869);
and U7235 (N_7235,In_1869,In_2009);
or U7236 (N_7236,In_43,In_1085);
xor U7237 (N_7237,In_2010,In_1631);
or U7238 (N_7238,In_2743,In_1569);
xnor U7239 (N_7239,In_2015,In_902);
nand U7240 (N_7240,In_1961,In_2722);
nor U7241 (N_7241,In_2961,In_1380);
and U7242 (N_7242,In_808,In_2398);
or U7243 (N_7243,In_2174,In_1895);
or U7244 (N_7244,In_2914,In_2955);
nor U7245 (N_7245,In_2373,In_2406);
or U7246 (N_7246,In_402,In_2597);
nor U7247 (N_7247,In_1893,In_1390);
and U7248 (N_7248,In_1295,In_579);
and U7249 (N_7249,In_2578,In_1593);
nand U7250 (N_7250,In_1703,In_2886);
xnor U7251 (N_7251,In_2819,In_1726);
and U7252 (N_7252,In_312,In_113);
or U7253 (N_7253,In_314,In_77);
xor U7254 (N_7254,In_1464,In_1634);
nor U7255 (N_7255,In_621,In_2799);
or U7256 (N_7256,In_1087,In_2835);
nor U7257 (N_7257,In_746,In_572);
or U7258 (N_7258,In_1737,In_2173);
and U7259 (N_7259,In_133,In_2925);
and U7260 (N_7260,In_1742,In_437);
or U7261 (N_7261,In_2295,In_1465);
xnor U7262 (N_7262,In_1088,In_2794);
nor U7263 (N_7263,In_1478,In_388);
or U7264 (N_7264,In_2586,In_2742);
or U7265 (N_7265,In_1335,In_1142);
nor U7266 (N_7266,In_2883,In_746);
or U7267 (N_7267,In_539,In_2276);
xnor U7268 (N_7268,In_147,In_894);
nand U7269 (N_7269,In_499,In_899);
nor U7270 (N_7270,In_939,In_1619);
nor U7271 (N_7271,In_1628,In_989);
and U7272 (N_7272,In_809,In_692);
or U7273 (N_7273,In_1566,In_2646);
or U7274 (N_7274,In_772,In_1377);
nor U7275 (N_7275,In_97,In_1680);
nor U7276 (N_7276,In_2846,In_2602);
or U7277 (N_7277,In_1611,In_1571);
or U7278 (N_7278,In_293,In_2);
or U7279 (N_7279,In_2010,In_2266);
nand U7280 (N_7280,In_1518,In_153);
xor U7281 (N_7281,In_2000,In_1356);
xor U7282 (N_7282,In_2329,In_738);
or U7283 (N_7283,In_1118,In_596);
and U7284 (N_7284,In_383,In_498);
and U7285 (N_7285,In_2835,In_2249);
and U7286 (N_7286,In_796,In_1717);
nand U7287 (N_7287,In_2833,In_522);
nor U7288 (N_7288,In_2623,In_2071);
nand U7289 (N_7289,In_711,In_779);
nand U7290 (N_7290,In_2311,In_1023);
nand U7291 (N_7291,In_421,In_577);
or U7292 (N_7292,In_2891,In_2974);
and U7293 (N_7293,In_2732,In_1600);
nand U7294 (N_7294,In_1041,In_1099);
nor U7295 (N_7295,In_681,In_2944);
nand U7296 (N_7296,In_2380,In_389);
or U7297 (N_7297,In_2668,In_1162);
nor U7298 (N_7298,In_1802,In_1515);
or U7299 (N_7299,In_572,In_224);
and U7300 (N_7300,In_386,In_2826);
nor U7301 (N_7301,In_2830,In_2285);
nor U7302 (N_7302,In_2665,In_79);
xnor U7303 (N_7303,In_2171,In_866);
or U7304 (N_7304,In_922,In_2225);
or U7305 (N_7305,In_2536,In_878);
nand U7306 (N_7306,In_2411,In_633);
or U7307 (N_7307,In_1412,In_1596);
xor U7308 (N_7308,In_2755,In_2711);
nor U7309 (N_7309,In_780,In_643);
and U7310 (N_7310,In_1437,In_105);
xnor U7311 (N_7311,In_2958,In_2397);
nand U7312 (N_7312,In_70,In_2860);
nand U7313 (N_7313,In_2104,In_1182);
nand U7314 (N_7314,In_123,In_2816);
nand U7315 (N_7315,In_645,In_2990);
nand U7316 (N_7316,In_573,In_2917);
nand U7317 (N_7317,In_1302,In_1717);
and U7318 (N_7318,In_886,In_2565);
xnor U7319 (N_7319,In_1566,In_749);
xor U7320 (N_7320,In_2663,In_2390);
xnor U7321 (N_7321,In_1871,In_2599);
or U7322 (N_7322,In_649,In_1007);
or U7323 (N_7323,In_175,In_240);
and U7324 (N_7324,In_2514,In_2377);
nor U7325 (N_7325,In_1679,In_1324);
nor U7326 (N_7326,In_1083,In_1322);
and U7327 (N_7327,In_898,In_548);
nand U7328 (N_7328,In_1771,In_1884);
nand U7329 (N_7329,In_1327,In_521);
nand U7330 (N_7330,In_10,In_1764);
nor U7331 (N_7331,In_1797,In_930);
nand U7332 (N_7332,In_658,In_1366);
nand U7333 (N_7333,In_20,In_2352);
or U7334 (N_7334,In_2425,In_2565);
nand U7335 (N_7335,In_2335,In_2610);
nor U7336 (N_7336,In_2138,In_1925);
nor U7337 (N_7337,In_2976,In_1573);
nor U7338 (N_7338,In_1816,In_795);
xor U7339 (N_7339,In_2443,In_778);
nand U7340 (N_7340,In_2426,In_1513);
nor U7341 (N_7341,In_194,In_221);
nor U7342 (N_7342,In_2620,In_1485);
nand U7343 (N_7343,In_816,In_1488);
nand U7344 (N_7344,In_2282,In_493);
and U7345 (N_7345,In_2327,In_2197);
xnor U7346 (N_7346,In_1538,In_2646);
nor U7347 (N_7347,In_2840,In_474);
nor U7348 (N_7348,In_1388,In_1513);
and U7349 (N_7349,In_2626,In_1402);
and U7350 (N_7350,In_2293,In_402);
and U7351 (N_7351,In_327,In_2091);
nand U7352 (N_7352,In_973,In_1944);
and U7353 (N_7353,In_1948,In_1467);
nor U7354 (N_7354,In_306,In_1468);
xor U7355 (N_7355,In_2902,In_1298);
or U7356 (N_7356,In_853,In_745);
and U7357 (N_7357,In_874,In_865);
or U7358 (N_7358,In_2611,In_674);
nand U7359 (N_7359,In_100,In_1372);
and U7360 (N_7360,In_2317,In_944);
nand U7361 (N_7361,In_2802,In_112);
or U7362 (N_7362,In_2610,In_2249);
nor U7363 (N_7363,In_2604,In_2646);
or U7364 (N_7364,In_1430,In_2715);
nor U7365 (N_7365,In_2863,In_213);
nor U7366 (N_7366,In_2987,In_2599);
and U7367 (N_7367,In_1496,In_102);
nand U7368 (N_7368,In_543,In_763);
nand U7369 (N_7369,In_2706,In_878);
and U7370 (N_7370,In_2243,In_2641);
nand U7371 (N_7371,In_2354,In_2060);
and U7372 (N_7372,In_2116,In_1273);
nor U7373 (N_7373,In_761,In_1244);
nand U7374 (N_7374,In_804,In_363);
nand U7375 (N_7375,In_2539,In_531);
and U7376 (N_7376,In_979,In_1697);
nand U7377 (N_7377,In_884,In_2529);
nand U7378 (N_7378,In_1593,In_159);
and U7379 (N_7379,In_1004,In_2223);
or U7380 (N_7380,In_135,In_2565);
or U7381 (N_7381,In_712,In_1109);
nor U7382 (N_7382,In_758,In_735);
nand U7383 (N_7383,In_1769,In_433);
nand U7384 (N_7384,In_519,In_776);
nor U7385 (N_7385,In_26,In_2191);
nor U7386 (N_7386,In_1468,In_131);
and U7387 (N_7387,In_1866,In_315);
or U7388 (N_7388,In_1438,In_1159);
nor U7389 (N_7389,In_839,In_2903);
xnor U7390 (N_7390,In_1428,In_1050);
nand U7391 (N_7391,In_298,In_1281);
or U7392 (N_7392,In_1158,In_1346);
and U7393 (N_7393,In_115,In_2938);
and U7394 (N_7394,In_483,In_2072);
nor U7395 (N_7395,In_2736,In_2921);
or U7396 (N_7396,In_1505,In_1457);
nor U7397 (N_7397,In_618,In_2427);
nand U7398 (N_7398,In_2429,In_2632);
and U7399 (N_7399,In_943,In_926);
or U7400 (N_7400,In_320,In_1893);
nor U7401 (N_7401,In_2318,In_876);
and U7402 (N_7402,In_1276,In_1162);
or U7403 (N_7403,In_1208,In_867);
nor U7404 (N_7404,In_1791,In_264);
nor U7405 (N_7405,In_555,In_2532);
nand U7406 (N_7406,In_2462,In_761);
nand U7407 (N_7407,In_1281,In_1657);
or U7408 (N_7408,In_478,In_2947);
nor U7409 (N_7409,In_1990,In_2926);
or U7410 (N_7410,In_2319,In_2576);
or U7411 (N_7411,In_2217,In_875);
nand U7412 (N_7412,In_51,In_1983);
xor U7413 (N_7413,In_57,In_1220);
nor U7414 (N_7414,In_899,In_2081);
nor U7415 (N_7415,In_126,In_134);
nand U7416 (N_7416,In_2227,In_2368);
or U7417 (N_7417,In_1408,In_1794);
and U7418 (N_7418,In_418,In_1988);
or U7419 (N_7419,In_2252,In_1452);
and U7420 (N_7420,In_2747,In_1660);
nor U7421 (N_7421,In_945,In_1245);
nor U7422 (N_7422,In_202,In_1993);
and U7423 (N_7423,In_2960,In_187);
or U7424 (N_7424,In_1128,In_2796);
and U7425 (N_7425,In_1082,In_2715);
nor U7426 (N_7426,In_1327,In_2565);
or U7427 (N_7427,In_2867,In_606);
nor U7428 (N_7428,In_1946,In_787);
and U7429 (N_7429,In_1770,In_1427);
nand U7430 (N_7430,In_2826,In_2312);
xor U7431 (N_7431,In_2378,In_2186);
xor U7432 (N_7432,In_2069,In_1373);
or U7433 (N_7433,In_715,In_163);
and U7434 (N_7434,In_2702,In_1421);
nand U7435 (N_7435,In_2623,In_136);
xnor U7436 (N_7436,In_2091,In_1009);
or U7437 (N_7437,In_2352,In_298);
nand U7438 (N_7438,In_2305,In_1010);
or U7439 (N_7439,In_2886,In_1177);
nand U7440 (N_7440,In_2131,In_1342);
or U7441 (N_7441,In_2741,In_1719);
and U7442 (N_7442,In_876,In_1628);
nand U7443 (N_7443,In_2516,In_961);
and U7444 (N_7444,In_459,In_1028);
xor U7445 (N_7445,In_469,In_2619);
xnor U7446 (N_7446,In_1503,In_616);
or U7447 (N_7447,In_180,In_453);
or U7448 (N_7448,In_1962,In_1484);
or U7449 (N_7449,In_102,In_2000);
nand U7450 (N_7450,In_59,In_2467);
nor U7451 (N_7451,In_1843,In_1417);
xnor U7452 (N_7452,In_90,In_2879);
xnor U7453 (N_7453,In_1856,In_2720);
or U7454 (N_7454,In_580,In_1736);
and U7455 (N_7455,In_2265,In_1618);
nor U7456 (N_7456,In_2984,In_2691);
nor U7457 (N_7457,In_1087,In_2604);
xnor U7458 (N_7458,In_2641,In_798);
or U7459 (N_7459,In_2899,In_784);
or U7460 (N_7460,In_1819,In_2568);
and U7461 (N_7461,In_1398,In_2943);
nand U7462 (N_7462,In_1154,In_1530);
nand U7463 (N_7463,In_1455,In_681);
or U7464 (N_7464,In_35,In_113);
nor U7465 (N_7465,In_249,In_1354);
nand U7466 (N_7466,In_486,In_1044);
and U7467 (N_7467,In_2045,In_2936);
nor U7468 (N_7468,In_2960,In_1015);
or U7469 (N_7469,In_2102,In_1031);
and U7470 (N_7470,In_266,In_2408);
or U7471 (N_7471,In_2189,In_2935);
xor U7472 (N_7472,In_1763,In_856);
nor U7473 (N_7473,In_188,In_1523);
or U7474 (N_7474,In_2212,In_757);
nand U7475 (N_7475,In_285,In_2457);
nand U7476 (N_7476,In_2540,In_662);
and U7477 (N_7477,In_999,In_1071);
or U7478 (N_7478,In_560,In_1326);
xor U7479 (N_7479,In_1113,In_2487);
xor U7480 (N_7480,In_338,In_2122);
or U7481 (N_7481,In_1117,In_2567);
xor U7482 (N_7482,In_1187,In_682);
or U7483 (N_7483,In_1925,In_1907);
and U7484 (N_7484,In_1875,In_762);
nor U7485 (N_7485,In_1415,In_1968);
nand U7486 (N_7486,In_782,In_860);
or U7487 (N_7487,In_2583,In_2762);
and U7488 (N_7488,In_795,In_2892);
and U7489 (N_7489,In_199,In_2295);
or U7490 (N_7490,In_2943,In_2255);
or U7491 (N_7491,In_2495,In_2519);
or U7492 (N_7492,In_2825,In_406);
nor U7493 (N_7493,In_267,In_2366);
or U7494 (N_7494,In_517,In_1872);
nor U7495 (N_7495,In_779,In_369);
nor U7496 (N_7496,In_921,In_1017);
nor U7497 (N_7497,In_1751,In_462);
or U7498 (N_7498,In_2614,In_2557);
nor U7499 (N_7499,In_1963,In_2936);
and U7500 (N_7500,In_2847,In_1532);
nand U7501 (N_7501,In_431,In_2294);
nand U7502 (N_7502,In_1784,In_2974);
or U7503 (N_7503,In_171,In_346);
or U7504 (N_7504,In_2565,In_91);
nor U7505 (N_7505,In_607,In_1981);
nor U7506 (N_7506,In_655,In_2662);
nor U7507 (N_7507,In_2918,In_826);
nand U7508 (N_7508,In_2046,In_2798);
and U7509 (N_7509,In_1278,In_638);
and U7510 (N_7510,In_1174,In_757);
and U7511 (N_7511,In_213,In_564);
nand U7512 (N_7512,In_1161,In_2108);
xor U7513 (N_7513,In_2601,In_2586);
xnor U7514 (N_7514,In_1016,In_2059);
or U7515 (N_7515,In_2784,In_2363);
nor U7516 (N_7516,In_2331,In_1539);
nand U7517 (N_7517,In_165,In_322);
and U7518 (N_7518,In_556,In_1167);
or U7519 (N_7519,In_1576,In_2117);
or U7520 (N_7520,In_1490,In_2861);
nand U7521 (N_7521,In_553,In_1686);
and U7522 (N_7522,In_1032,In_2671);
nor U7523 (N_7523,In_275,In_2855);
nor U7524 (N_7524,In_363,In_2510);
and U7525 (N_7525,In_2015,In_1033);
nand U7526 (N_7526,In_811,In_621);
or U7527 (N_7527,In_2411,In_2160);
or U7528 (N_7528,In_1850,In_928);
and U7529 (N_7529,In_1983,In_2922);
and U7530 (N_7530,In_1819,In_1538);
or U7531 (N_7531,In_1939,In_1596);
nand U7532 (N_7532,In_963,In_505);
and U7533 (N_7533,In_130,In_2054);
or U7534 (N_7534,In_924,In_1758);
nand U7535 (N_7535,In_492,In_2517);
nand U7536 (N_7536,In_590,In_1020);
nand U7537 (N_7537,In_2750,In_2392);
and U7538 (N_7538,In_70,In_1031);
nor U7539 (N_7539,In_691,In_1342);
and U7540 (N_7540,In_1227,In_2956);
nand U7541 (N_7541,In_1796,In_1815);
xnor U7542 (N_7542,In_1551,In_951);
and U7543 (N_7543,In_1326,In_576);
nor U7544 (N_7544,In_2438,In_1732);
nor U7545 (N_7545,In_637,In_2120);
nand U7546 (N_7546,In_1317,In_2613);
nand U7547 (N_7547,In_693,In_1121);
nand U7548 (N_7548,In_1870,In_1212);
or U7549 (N_7549,In_2305,In_1378);
or U7550 (N_7550,In_1310,In_387);
or U7551 (N_7551,In_675,In_599);
nand U7552 (N_7552,In_2633,In_816);
or U7553 (N_7553,In_2854,In_516);
nand U7554 (N_7554,In_1727,In_837);
and U7555 (N_7555,In_2154,In_2730);
and U7556 (N_7556,In_388,In_209);
and U7557 (N_7557,In_2108,In_2413);
nor U7558 (N_7558,In_242,In_1062);
nor U7559 (N_7559,In_824,In_1643);
nor U7560 (N_7560,In_218,In_2588);
nor U7561 (N_7561,In_1679,In_96);
nor U7562 (N_7562,In_1132,In_1225);
nand U7563 (N_7563,In_488,In_219);
nand U7564 (N_7564,In_2748,In_188);
nor U7565 (N_7565,In_2674,In_1269);
nand U7566 (N_7566,In_2000,In_993);
or U7567 (N_7567,In_822,In_1744);
nand U7568 (N_7568,In_1579,In_2872);
nand U7569 (N_7569,In_823,In_1182);
or U7570 (N_7570,In_2413,In_1863);
nor U7571 (N_7571,In_1261,In_1206);
nor U7572 (N_7572,In_1024,In_2500);
nor U7573 (N_7573,In_1692,In_2290);
xnor U7574 (N_7574,In_2353,In_932);
nand U7575 (N_7575,In_820,In_1418);
nand U7576 (N_7576,In_799,In_2129);
nor U7577 (N_7577,In_1161,In_2820);
or U7578 (N_7578,In_2579,In_2125);
nor U7579 (N_7579,In_1316,In_1291);
and U7580 (N_7580,In_257,In_679);
or U7581 (N_7581,In_729,In_1748);
nor U7582 (N_7582,In_268,In_563);
xor U7583 (N_7583,In_1327,In_1142);
nor U7584 (N_7584,In_392,In_1168);
or U7585 (N_7585,In_2387,In_771);
nor U7586 (N_7586,In_2539,In_1646);
and U7587 (N_7587,In_1192,In_240);
and U7588 (N_7588,In_1860,In_1484);
and U7589 (N_7589,In_2413,In_2741);
or U7590 (N_7590,In_2099,In_1739);
and U7591 (N_7591,In_2023,In_1745);
nand U7592 (N_7592,In_2425,In_2139);
and U7593 (N_7593,In_1555,In_2462);
and U7594 (N_7594,In_1969,In_1872);
nand U7595 (N_7595,In_2177,In_2831);
or U7596 (N_7596,In_2702,In_1817);
or U7597 (N_7597,In_2121,In_1662);
and U7598 (N_7598,In_2337,In_765);
or U7599 (N_7599,In_2690,In_1161);
nand U7600 (N_7600,In_1164,In_2066);
or U7601 (N_7601,In_157,In_224);
or U7602 (N_7602,In_227,In_1232);
nand U7603 (N_7603,In_2079,In_141);
nor U7604 (N_7604,In_148,In_1908);
nor U7605 (N_7605,In_515,In_302);
nor U7606 (N_7606,In_1261,In_528);
nor U7607 (N_7607,In_1130,In_269);
xnor U7608 (N_7608,In_437,In_1529);
or U7609 (N_7609,In_472,In_2588);
nor U7610 (N_7610,In_2606,In_2307);
and U7611 (N_7611,In_1643,In_555);
or U7612 (N_7612,In_1090,In_2793);
or U7613 (N_7613,In_2913,In_391);
nand U7614 (N_7614,In_225,In_1789);
and U7615 (N_7615,In_2810,In_1317);
and U7616 (N_7616,In_1619,In_918);
and U7617 (N_7617,In_342,In_2393);
nand U7618 (N_7618,In_289,In_6);
or U7619 (N_7619,In_2971,In_1915);
nor U7620 (N_7620,In_1799,In_1286);
nand U7621 (N_7621,In_1698,In_1935);
xnor U7622 (N_7622,In_2681,In_1212);
and U7623 (N_7623,In_2798,In_997);
nand U7624 (N_7624,In_2242,In_2537);
or U7625 (N_7625,In_1624,In_1378);
nor U7626 (N_7626,In_2457,In_2069);
and U7627 (N_7627,In_2487,In_202);
nor U7628 (N_7628,In_2699,In_1825);
or U7629 (N_7629,In_1422,In_2152);
or U7630 (N_7630,In_253,In_474);
or U7631 (N_7631,In_670,In_1966);
or U7632 (N_7632,In_433,In_324);
nor U7633 (N_7633,In_1408,In_1470);
and U7634 (N_7634,In_1792,In_2696);
nor U7635 (N_7635,In_2246,In_374);
xor U7636 (N_7636,In_1987,In_2289);
xnor U7637 (N_7637,In_2725,In_2450);
and U7638 (N_7638,In_70,In_1233);
nor U7639 (N_7639,In_370,In_1856);
nor U7640 (N_7640,In_1871,In_2023);
and U7641 (N_7641,In_2580,In_146);
nand U7642 (N_7642,In_479,In_580);
nor U7643 (N_7643,In_2340,In_2944);
nor U7644 (N_7644,In_1819,In_1599);
or U7645 (N_7645,In_870,In_702);
xor U7646 (N_7646,In_1028,In_410);
nand U7647 (N_7647,In_2698,In_31);
nor U7648 (N_7648,In_965,In_1531);
and U7649 (N_7649,In_2183,In_2742);
or U7650 (N_7650,In_1019,In_1250);
and U7651 (N_7651,In_2175,In_2664);
nand U7652 (N_7652,In_498,In_1087);
nand U7653 (N_7653,In_535,In_2690);
and U7654 (N_7654,In_1760,In_2074);
nand U7655 (N_7655,In_1928,In_1748);
nor U7656 (N_7656,In_1897,In_742);
and U7657 (N_7657,In_2204,In_1897);
nor U7658 (N_7658,In_1223,In_783);
or U7659 (N_7659,In_2411,In_905);
nand U7660 (N_7660,In_2720,In_2115);
nand U7661 (N_7661,In_414,In_899);
nand U7662 (N_7662,In_1015,In_6);
nand U7663 (N_7663,In_780,In_2875);
xor U7664 (N_7664,In_2883,In_2705);
or U7665 (N_7665,In_1517,In_102);
nor U7666 (N_7666,In_2164,In_2989);
or U7667 (N_7667,In_867,In_1292);
or U7668 (N_7668,In_1471,In_2738);
and U7669 (N_7669,In_2108,In_1653);
nand U7670 (N_7670,In_2682,In_2806);
xor U7671 (N_7671,In_1169,In_2786);
and U7672 (N_7672,In_1371,In_303);
nand U7673 (N_7673,In_1333,In_2912);
or U7674 (N_7674,In_2613,In_28);
nand U7675 (N_7675,In_564,In_1786);
and U7676 (N_7676,In_2079,In_1734);
xor U7677 (N_7677,In_290,In_1696);
and U7678 (N_7678,In_446,In_2856);
nand U7679 (N_7679,In_993,In_2069);
and U7680 (N_7680,In_2718,In_1984);
nand U7681 (N_7681,In_2348,In_1615);
nor U7682 (N_7682,In_2137,In_940);
or U7683 (N_7683,In_1116,In_1560);
xor U7684 (N_7684,In_1265,In_2190);
nand U7685 (N_7685,In_142,In_2693);
or U7686 (N_7686,In_930,In_339);
xnor U7687 (N_7687,In_343,In_2628);
nand U7688 (N_7688,In_687,In_660);
nor U7689 (N_7689,In_1443,In_2187);
nand U7690 (N_7690,In_166,In_2602);
nand U7691 (N_7691,In_1180,In_1099);
nand U7692 (N_7692,In_2834,In_1606);
and U7693 (N_7693,In_1662,In_124);
or U7694 (N_7694,In_1606,In_687);
nand U7695 (N_7695,In_259,In_1501);
nor U7696 (N_7696,In_2536,In_1819);
nand U7697 (N_7697,In_1719,In_1475);
nand U7698 (N_7698,In_752,In_1329);
or U7699 (N_7699,In_1460,In_1836);
nor U7700 (N_7700,In_355,In_2294);
and U7701 (N_7701,In_655,In_1307);
or U7702 (N_7702,In_840,In_418);
or U7703 (N_7703,In_2795,In_2892);
nor U7704 (N_7704,In_1428,In_2577);
xnor U7705 (N_7705,In_1006,In_732);
nand U7706 (N_7706,In_2528,In_66);
or U7707 (N_7707,In_2695,In_197);
or U7708 (N_7708,In_562,In_2057);
nor U7709 (N_7709,In_731,In_1690);
nor U7710 (N_7710,In_2394,In_919);
and U7711 (N_7711,In_2295,In_2899);
or U7712 (N_7712,In_461,In_1089);
and U7713 (N_7713,In_279,In_2194);
nand U7714 (N_7714,In_1625,In_1670);
xnor U7715 (N_7715,In_901,In_2405);
xnor U7716 (N_7716,In_1565,In_1895);
or U7717 (N_7717,In_1377,In_263);
nand U7718 (N_7718,In_645,In_632);
nand U7719 (N_7719,In_1511,In_1911);
nand U7720 (N_7720,In_2849,In_2414);
or U7721 (N_7721,In_2695,In_596);
and U7722 (N_7722,In_1541,In_1282);
or U7723 (N_7723,In_1566,In_452);
xnor U7724 (N_7724,In_2438,In_1648);
and U7725 (N_7725,In_1445,In_114);
xnor U7726 (N_7726,In_899,In_1205);
nor U7727 (N_7727,In_2592,In_339);
nor U7728 (N_7728,In_1568,In_1872);
nand U7729 (N_7729,In_323,In_527);
nand U7730 (N_7730,In_2656,In_655);
nand U7731 (N_7731,In_423,In_257);
nand U7732 (N_7732,In_2509,In_1749);
nor U7733 (N_7733,In_83,In_291);
and U7734 (N_7734,In_1375,In_1974);
nor U7735 (N_7735,In_1908,In_608);
or U7736 (N_7736,In_2278,In_837);
or U7737 (N_7737,In_2685,In_1964);
or U7738 (N_7738,In_731,In_2791);
or U7739 (N_7739,In_289,In_2096);
nor U7740 (N_7740,In_19,In_2012);
nor U7741 (N_7741,In_174,In_285);
and U7742 (N_7742,In_1030,In_669);
and U7743 (N_7743,In_2221,In_2491);
nand U7744 (N_7744,In_1949,In_2731);
nor U7745 (N_7745,In_1652,In_1821);
nor U7746 (N_7746,In_1516,In_47);
and U7747 (N_7747,In_309,In_2226);
nand U7748 (N_7748,In_2594,In_1822);
or U7749 (N_7749,In_1343,In_1851);
nor U7750 (N_7750,In_1145,In_2488);
and U7751 (N_7751,In_592,In_281);
or U7752 (N_7752,In_864,In_2378);
or U7753 (N_7753,In_1671,In_1443);
xor U7754 (N_7754,In_1286,In_2077);
xor U7755 (N_7755,In_353,In_2415);
xor U7756 (N_7756,In_211,In_2368);
and U7757 (N_7757,In_1558,In_2925);
xor U7758 (N_7758,In_223,In_1072);
or U7759 (N_7759,In_182,In_751);
and U7760 (N_7760,In_1376,In_1676);
xnor U7761 (N_7761,In_310,In_2207);
nor U7762 (N_7762,In_1863,In_1666);
and U7763 (N_7763,In_2569,In_1035);
and U7764 (N_7764,In_767,In_2645);
nor U7765 (N_7765,In_963,In_2545);
and U7766 (N_7766,In_381,In_2390);
and U7767 (N_7767,In_364,In_1302);
and U7768 (N_7768,In_1390,In_3);
nand U7769 (N_7769,In_2379,In_258);
or U7770 (N_7770,In_780,In_1056);
nand U7771 (N_7771,In_711,In_2490);
and U7772 (N_7772,In_2910,In_2413);
and U7773 (N_7773,In_832,In_693);
and U7774 (N_7774,In_1104,In_1753);
or U7775 (N_7775,In_526,In_2824);
nand U7776 (N_7776,In_2803,In_1895);
or U7777 (N_7777,In_2006,In_762);
and U7778 (N_7778,In_1046,In_2456);
nor U7779 (N_7779,In_2376,In_778);
nor U7780 (N_7780,In_2036,In_589);
xor U7781 (N_7781,In_759,In_1111);
nor U7782 (N_7782,In_800,In_386);
and U7783 (N_7783,In_1248,In_743);
nand U7784 (N_7784,In_2512,In_2144);
xor U7785 (N_7785,In_1410,In_1187);
and U7786 (N_7786,In_43,In_1019);
or U7787 (N_7787,In_957,In_1336);
nand U7788 (N_7788,In_500,In_111);
nor U7789 (N_7789,In_2763,In_2774);
nor U7790 (N_7790,In_2138,In_1470);
nand U7791 (N_7791,In_1852,In_1703);
nor U7792 (N_7792,In_1438,In_798);
nand U7793 (N_7793,In_2040,In_1256);
nand U7794 (N_7794,In_1349,In_1704);
xnor U7795 (N_7795,In_2957,In_2197);
nand U7796 (N_7796,In_2363,In_1380);
nor U7797 (N_7797,In_2565,In_611);
and U7798 (N_7798,In_343,In_164);
nor U7799 (N_7799,In_951,In_1575);
nor U7800 (N_7800,In_1517,In_1065);
nor U7801 (N_7801,In_469,In_1465);
and U7802 (N_7802,In_1695,In_1530);
or U7803 (N_7803,In_2587,In_2828);
xnor U7804 (N_7804,In_226,In_1381);
nor U7805 (N_7805,In_38,In_1719);
xnor U7806 (N_7806,In_1240,In_2650);
and U7807 (N_7807,In_2546,In_2215);
nor U7808 (N_7808,In_2130,In_327);
or U7809 (N_7809,In_1393,In_1654);
or U7810 (N_7810,In_2058,In_221);
and U7811 (N_7811,In_380,In_2504);
or U7812 (N_7812,In_374,In_2439);
nand U7813 (N_7813,In_1484,In_1233);
or U7814 (N_7814,In_2605,In_1230);
nand U7815 (N_7815,In_501,In_1237);
nor U7816 (N_7816,In_2015,In_19);
and U7817 (N_7817,In_1360,In_683);
and U7818 (N_7818,In_1204,In_2559);
nand U7819 (N_7819,In_2271,In_1949);
or U7820 (N_7820,In_186,In_31);
nor U7821 (N_7821,In_757,In_1402);
nor U7822 (N_7822,In_2124,In_1167);
or U7823 (N_7823,In_2571,In_376);
and U7824 (N_7824,In_611,In_761);
nor U7825 (N_7825,In_1934,In_1475);
nor U7826 (N_7826,In_2218,In_73);
nand U7827 (N_7827,In_1527,In_735);
nor U7828 (N_7828,In_1648,In_2269);
and U7829 (N_7829,In_1270,In_2656);
nand U7830 (N_7830,In_17,In_596);
nor U7831 (N_7831,In_2659,In_503);
nand U7832 (N_7832,In_2717,In_726);
nor U7833 (N_7833,In_2769,In_1307);
nand U7834 (N_7834,In_267,In_1394);
or U7835 (N_7835,In_1855,In_2739);
or U7836 (N_7836,In_1172,In_1440);
or U7837 (N_7837,In_369,In_587);
or U7838 (N_7838,In_1150,In_341);
and U7839 (N_7839,In_2378,In_2992);
nor U7840 (N_7840,In_1698,In_1773);
or U7841 (N_7841,In_2618,In_1323);
and U7842 (N_7842,In_1560,In_38);
and U7843 (N_7843,In_222,In_2417);
and U7844 (N_7844,In_2580,In_1907);
or U7845 (N_7845,In_1458,In_973);
or U7846 (N_7846,In_1173,In_471);
nand U7847 (N_7847,In_1030,In_2825);
nand U7848 (N_7848,In_1539,In_115);
nand U7849 (N_7849,In_457,In_1172);
nand U7850 (N_7850,In_1265,In_1139);
xor U7851 (N_7851,In_668,In_751);
and U7852 (N_7852,In_1304,In_383);
and U7853 (N_7853,In_2123,In_1513);
or U7854 (N_7854,In_2003,In_2780);
nor U7855 (N_7855,In_1049,In_2419);
or U7856 (N_7856,In_2640,In_407);
and U7857 (N_7857,In_370,In_1080);
and U7858 (N_7858,In_1015,In_2275);
and U7859 (N_7859,In_515,In_2068);
and U7860 (N_7860,In_2205,In_2315);
nand U7861 (N_7861,In_558,In_288);
and U7862 (N_7862,In_2750,In_2301);
and U7863 (N_7863,In_1162,In_131);
xnor U7864 (N_7864,In_2210,In_2885);
and U7865 (N_7865,In_2573,In_933);
and U7866 (N_7866,In_97,In_2688);
nand U7867 (N_7867,In_2482,In_491);
and U7868 (N_7868,In_171,In_2927);
and U7869 (N_7869,In_656,In_1745);
nor U7870 (N_7870,In_745,In_2895);
nand U7871 (N_7871,In_1011,In_2388);
nor U7872 (N_7872,In_803,In_1706);
xnor U7873 (N_7873,In_2998,In_2893);
or U7874 (N_7874,In_2435,In_696);
nand U7875 (N_7875,In_2363,In_1097);
nor U7876 (N_7876,In_2974,In_2651);
nor U7877 (N_7877,In_160,In_2249);
or U7878 (N_7878,In_1041,In_2177);
and U7879 (N_7879,In_264,In_1186);
nand U7880 (N_7880,In_298,In_1870);
and U7881 (N_7881,In_1797,In_316);
nor U7882 (N_7882,In_2287,In_2123);
or U7883 (N_7883,In_1892,In_242);
nor U7884 (N_7884,In_812,In_1686);
nand U7885 (N_7885,In_1513,In_1506);
or U7886 (N_7886,In_1360,In_518);
nand U7887 (N_7887,In_2150,In_727);
and U7888 (N_7888,In_67,In_1315);
and U7889 (N_7889,In_668,In_1552);
and U7890 (N_7890,In_2076,In_645);
nand U7891 (N_7891,In_2478,In_1419);
nor U7892 (N_7892,In_85,In_2721);
and U7893 (N_7893,In_886,In_2466);
or U7894 (N_7894,In_496,In_129);
or U7895 (N_7895,In_156,In_1355);
or U7896 (N_7896,In_397,In_1391);
and U7897 (N_7897,In_145,In_1730);
nor U7898 (N_7898,In_1129,In_176);
or U7899 (N_7899,In_2391,In_2995);
or U7900 (N_7900,In_207,In_1787);
and U7901 (N_7901,In_1601,In_453);
or U7902 (N_7902,In_1276,In_725);
or U7903 (N_7903,In_1708,In_204);
and U7904 (N_7904,In_2532,In_566);
nor U7905 (N_7905,In_1403,In_1028);
nor U7906 (N_7906,In_2487,In_1160);
and U7907 (N_7907,In_597,In_613);
xor U7908 (N_7908,In_2740,In_1043);
or U7909 (N_7909,In_178,In_2582);
nand U7910 (N_7910,In_1114,In_2311);
and U7911 (N_7911,In_732,In_900);
nor U7912 (N_7912,In_2927,In_437);
and U7913 (N_7913,In_1898,In_1315);
nor U7914 (N_7914,In_1364,In_2588);
or U7915 (N_7915,In_771,In_2038);
or U7916 (N_7916,In_1289,In_2629);
nand U7917 (N_7917,In_2581,In_775);
nand U7918 (N_7918,In_1456,In_1085);
nand U7919 (N_7919,In_715,In_412);
or U7920 (N_7920,In_73,In_1561);
or U7921 (N_7921,In_1842,In_686);
nand U7922 (N_7922,In_2087,In_977);
nand U7923 (N_7923,In_1539,In_2124);
nand U7924 (N_7924,In_2720,In_1012);
or U7925 (N_7925,In_2444,In_205);
xnor U7926 (N_7926,In_1480,In_1737);
nor U7927 (N_7927,In_1578,In_1017);
nand U7928 (N_7928,In_1848,In_950);
or U7929 (N_7929,In_2650,In_72);
nand U7930 (N_7930,In_983,In_106);
and U7931 (N_7931,In_7,In_2006);
and U7932 (N_7932,In_1387,In_2799);
or U7933 (N_7933,In_2304,In_989);
nand U7934 (N_7934,In_415,In_1016);
or U7935 (N_7935,In_240,In_88);
nor U7936 (N_7936,In_2547,In_249);
or U7937 (N_7937,In_2765,In_523);
and U7938 (N_7938,In_766,In_866);
nand U7939 (N_7939,In_1689,In_1005);
nor U7940 (N_7940,In_2899,In_2676);
nor U7941 (N_7941,In_1893,In_2482);
and U7942 (N_7942,In_2166,In_2187);
or U7943 (N_7943,In_2321,In_555);
or U7944 (N_7944,In_1762,In_738);
xor U7945 (N_7945,In_475,In_221);
or U7946 (N_7946,In_1071,In_133);
or U7947 (N_7947,In_1875,In_2937);
and U7948 (N_7948,In_2876,In_1412);
nor U7949 (N_7949,In_214,In_2211);
xor U7950 (N_7950,In_1519,In_540);
nand U7951 (N_7951,In_2452,In_2829);
nand U7952 (N_7952,In_1884,In_1486);
nand U7953 (N_7953,In_2620,In_2889);
nand U7954 (N_7954,In_725,In_167);
and U7955 (N_7955,In_2003,In_2042);
or U7956 (N_7956,In_2382,In_2270);
or U7957 (N_7957,In_151,In_2929);
nand U7958 (N_7958,In_1570,In_2897);
nand U7959 (N_7959,In_2385,In_187);
nor U7960 (N_7960,In_2256,In_1451);
xnor U7961 (N_7961,In_2563,In_1665);
or U7962 (N_7962,In_1768,In_2745);
or U7963 (N_7963,In_2114,In_2360);
nor U7964 (N_7964,In_6,In_1350);
and U7965 (N_7965,In_1530,In_691);
nand U7966 (N_7966,In_2168,In_1116);
nor U7967 (N_7967,In_2160,In_2308);
xnor U7968 (N_7968,In_828,In_2695);
nand U7969 (N_7969,In_2430,In_2181);
nor U7970 (N_7970,In_823,In_2961);
or U7971 (N_7971,In_2305,In_2669);
nand U7972 (N_7972,In_566,In_2615);
and U7973 (N_7973,In_72,In_2926);
nand U7974 (N_7974,In_2961,In_1092);
xor U7975 (N_7975,In_601,In_1741);
nand U7976 (N_7976,In_1174,In_2307);
or U7977 (N_7977,In_444,In_2519);
and U7978 (N_7978,In_2828,In_2530);
nor U7979 (N_7979,In_853,In_885);
nand U7980 (N_7980,In_95,In_1656);
xnor U7981 (N_7981,In_2704,In_1024);
and U7982 (N_7982,In_2142,In_733);
and U7983 (N_7983,In_938,In_1385);
nand U7984 (N_7984,In_416,In_678);
and U7985 (N_7985,In_874,In_1981);
nand U7986 (N_7986,In_1328,In_1460);
nor U7987 (N_7987,In_1775,In_2899);
or U7988 (N_7988,In_1464,In_2357);
and U7989 (N_7989,In_2085,In_1710);
xnor U7990 (N_7990,In_1727,In_1882);
nand U7991 (N_7991,In_1079,In_533);
nor U7992 (N_7992,In_1885,In_54);
and U7993 (N_7993,In_2066,In_2872);
nand U7994 (N_7994,In_811,In_2354);
nor U7995 (N_7995,In_711,In_1673);
nand U7996 (N_7996,In_427,In_2202);
nand U7997 (N_7997,In_873,In_1575);
and U7998 (N_7998,In_827,In_763);
or U7999 (N_7999,In_1673,In_2802);
nor U8000 (N_8000,In_552,In_113);
nor U8001 (N_8001,In_854,In_1283);
xor U8002 (N_8002,In_2207,In_1875);
nand U8003 (N_8003,In_689,In_1897);
nand U8004 (N_8004,In_2280,In_2506);
nand U8005 (N_8005,In_489,In_1710);
and U8006 (N_8006,In_776,In_183);
and U8007 (N_8007,In_1617,In_2962);
nor U8008 (N_8008,In_2829,In_1331);
nand U8009 (N_8009,In_2604,In_2746);
or U8010 (N_8010,In_1597,In_337);
nor U8011 (N_8011,In_2605,In_2516);
nand U8012 (N_8012,In_2609,In_992);
and U8013 (N_8013,In_1805,In_1341);
nor U8014 (N_8014,In_1890,In_749);
nand U8015 (N_8015,In_1926,In_2626);
or U8016 (N_8016,In_2534,In_1813);
xnor U8017 (N_8017,In_1659,In_808);
nor U8018 (N_8018,In_128,In_2439);
nor U8019 (N_8019,In_574,In_2410);
nand U8020 (N_8020,In_2787,In_778);
and U8021 (N_8021,In_2293,In_414);
nand U8022 (N_8022,In_2231,In_1348);
nand U8023 (N_8023,In_492,In_672);
nor U8024 (N_8024,In_1508,In_2235);
or U8025 (N_8025,In_2300,In_1504);
or U8026 (N_8026,In_2521,In_645);
xnor U8027 (N_8027,In_2634,In_2590);
nor U8028 (N_8028,In_1564,In_708);
or U8029 (N_8029,In_2083,In_1524);
nand U8030 (N_8030,In_1478,In_776);
and U8031 (N_8031,In_1586,In_2875);
nor U8032 (N_8032,In_2022,In_2471);
nand U8033 (N_8033,In_39,In_828);
or U8034 (N_8034,In_2465,In_2947);
nor U8035 (N_8035,In_2612,In_697);
or U8036 (N_8036,In_2130,In_1616);
nor U8037 (N_8037,In_577,In_1772);
or U8038 (N_8038,In_128,In_651);
nand U8039 (N_8039,In_2010,In_2639);
nand U8040 (N_8040,In_2955,In_2205);
or U8041 (N_8041,In_803,In_37);
xnor U8042 (N_8042,In_1535,In_1930);
nor U8043 (N_8043,In_2539,In_1714);
nor U8044 (N_8044,In_1529,In_2104);
and U8045 (N_8045,In_2335,In_1450);
xnor U8046 (N_8046,In_801,In_2457);
nand U8047 (N_8047,In_1311,In_1106);
and U8048 (N_8048,In_107,In_108);
or U8049 (N_8049,In_2556,In_1418);
and U8050 (N_8050,In_761,In_2416);
and U8051 (N_8051,In_2361,In_1852);
and U8052 (N_8052,In_2576,In_1425);
and U8053 (N_8053,In_475,In_650);
or U8054 (N_8054,In_2286,In_1025);
nor U8055 (N_8055,In_1653,In_1984);
nor U8056 (N_8056,In_860,In_1056);
nand U8057 (N_8057,In_232,In_869);
and U8058 (N_8058,In_581,In_2831);
and U8059 (N_8059,In_1622,In_1940);
and U8060 (N_8060,In_530,In_2828);
nand U8061 (N_8061,In_2061,In_2779);
and U8062 (N_8062,In_2789,In_770);
nor U8063 (N_8063,In_771,In_198);
or U8064 (N_8064,In_2098,In_1771);
nor U8065 (N_8065,In_152,In_1294);
xor U8066 (N_8066,In_2200,In_2597);
or U8067 (N_8067,In_2770,In_1384);
or U8068 (N_8068,In_2092,In_2091);
nor U8069 (N_8069,In_1253,In_2849);
and U8070 (N_8070,In_576,In_2150);
xnor U8071 (N_8071,In_1675,In_1617);
nor U8072 (N_8072,In_2,In_616);
nor U8073 (N_8073,In_1138,In_1350);
or U8074 (N_8074,In_1044,In_1039);
nand U8075 (N_8075,In_1925,In_728);
nor U8076 (N_8076,In_2657,In_438);
and U8077 (N_8077,In_1740,In_2160);
nor U8078 (N_8078,In_1177,In_1883);
or U8079 (N_8079,In_946,In_2936);
or U8080 (N_8080,In_364,In_2977);
or U8081 (N_8081,In_49,In_2720);
or U8082 (N_8082,In_940,In_2839);
nand U8083 (N_8083,In_2998,In_1366);
nand U8084 (N_8084,In_1902,In_2717);
and U8085 (N_8085,In_540,In_515);
nor U8086 (N_8086,In_2022,In_1624);
nand U8087 (N_8087,In_2611,In_2117);
nor U8088 (N_8088,In_2198,In_32);
nand U8089 (N_8089,In_2992,In_818);
or U8090 (N_8090,In_134,In_2095);
nand U8091 (N_8091,In_521,In_1233);
or U8092 (N_8092,In_292,In_2322);
nor U8093 (N_8093,In_2376,In_1629);
or U8094 (N_8094,In_958,In_830);
or U8095 (N_8095,In_1076,In_573);
or U8096 (N_8096,In_904,In_2486);
xnor U8097 (N_8097,In_1557,In_555);
or U8098 (N_8098,In_2028,In_1576);
nand U8099 (N_8099,In_18,In_989);
nand U8100 (N_8100,In_2359,In_2864);
nor U8101 (N_8101,In_2320,In_834);
xnor U8102 (N_8102,In_2726,In_653);
nor U8103 (N_8103,In_2915,In_2630);
nand U8104 (N_8104,In_2761,In_2588);
or U8105 (N_8105,In_454,In_255);
and U8106 (N_8106,In_1894,In_2496);
nor U8107 (N_8107,In_1085,In_1964);
nor U8108 (N_8108,In_738,In_1037);
nand U8109 (N_8109,In_156,In_2199);
xor U8110 (N_8110,In_9,In_2540);
and U8111 (N_8111,In_2784,In_381);
or U8112 (N_8112,In_1542,In_1833);
or U8113 (N_8113,In_2722,In_253);
nor U8114 (N_8114,In_824,In_464);
xnor U8115 (N_8115,In_2658,In_2078);
and U8116 (N_8116,In_606,In_1913);
or U8117 (N_8117,In_1052,In_96);
and U8118 (N_8118,In_1007,In_32);
nand U8119 (N_8119,In_2930,In_2676);
or U8120 (N_8120,In_1013,In_54);
nor U8121 (N_8121,In_31,In_1396);
or U8122 (N_8122,In_1414,In_1426);
and U8123 (N_8123,In_265,In_1141);
xnor U8124 (N_8124,In_319,In_191);
nor U8125 (N_8125,In_36,In_2960);
nand U8126 (N_8126,In_2367,In_173);
nand U8127 (N_8127,In_2681,In_2361);
nand U8128 (N_8128,In_542,In_2904);
or U8129 (N_8129,In_183,In_2432);
nand U8130 (N_8130,In_1646,In_1785);
nand U8131 (N_8131,In_2438,In_1833);
xnor U8132 (N_8132,In_2536,In_540);
nand U8133 (N_8133,In_2651,In_2330);
nor U8134 (N_8134,In_2702,In_2776);
nand U8135 (N_8135,In_1149,In_2987);
nor U8136 (N_8136,In_1296,In_1799);
or U8137 (N_8137,In_412,In_1182);
and U8138 (N_8138,In_2481,In_2121);
nor U8139 (N_8139,In_520,In_2620);
nand U8140 (N_8140,In_2965,In_2073);
and U8141 (N_8141,In_2654,In_202);
nand U8142 (N_8142,In_2272,In_2046);
nor U8143 (N_8143,In_1012,In_680);
nand U8144 (N_8144,In_791,In_2473);
and U8145 (N_8145,In_565,In_2165);
or U8146 (N_8146,In_1984,In_1609);
xnor U8147 (N_8147,In_588,In_1616);
xnor U8148 (N_8148,In_1387,In_2526);
nand U8149 (N_8149,In_2751,In_20);
xor U8150 (N_8150,In_2107,In_2935);
xnor U8151 (N_8151,In_381,In_239);
nor U8152 (N_8152,In_292,In_2241);
or U8153 (N_8153,In_442,In_1738);
and U8154 (N_8154,In_694,In_102);
or U8155 (N_8155,In_597,In_799);
and U8156 (N_8156,In_530,In_1608);
and U8157 (N_8157,In_2229,In_2571);
or U8158 (N_8158,In_1454,In_1643);
nand U8159 (N_8159,In_772,In_2708);
and U8160 (N_8160,In_323,In_110);
or U8161 (N_8161,In_2665,In_2945);
nor U8162 (N_8162,In_672,In_684);
nand U8163 (N_8163,In_2079,In_980);
and U8164 (N_8164,In_1109,In_1597);
or U8165 (N_8165,In_32,In_1455);
and U8166 (N_8166,In_708,In_963);
and U8167 (N_8167,In_2513,In_1885);
nand U8168 (N_8168,In_2388,In_1652);
or U8169 (N_8169,In_2141,In_2429);
or U8170 (N_8170,In_2407,In_2950);
nand U8171 (N_8171,In_81,In_1638);
and U8172 (N_8172,In_1626,In_1205);
and U8173 (N_8173,In_1803,In_298);
nand U8174 (N_8174,In_2207,In_87);
and U8175 (N_8175,In_1250,In_1464);
nand U8176 (N_8176,In_2023,In_2490);
and U8177 (N_8177,In_2804,In_2790);
or U8178 (N_8178,In_2013,In_1641);
nor U8179 (N_8179,In_2436,In_735);
xnor U8180 (N_8180,In_229,In_1797);
or U8181 (N_8181,In_627,In_1165);
nand U8182 (N_8182,In_410,In_2492);
nand U8183 (N_8183,In_168,In_2581);
nand U8184 (N_8184,In_1665,In_2379);
nor U8185 (N_8185,In_2716,In_2113);
and U8186 (N_8186,In_508,In_2950);
and U8187 (N_8187,In_2212,In_2557);
nand U8188 (N_8188,In_1646,In_276);
nor U8189 (N_8189,In_403,In_2108);
nor U8190 (N_8190,In_1654,In_386);
and U8191 (N_8191,In_2166,In_2427);
or U8192 (N_8192,In_72,In_2065);
nor U8193 (N_8193,In_1990,In_1625);
nor U8194 (N_8194,In_712,In_2653);
nor U8195 (N_8195,In_2608,In_1130);
nor U8196 (N_8196,In_1909,In_1516);
and U8197 (N_8197,In_852,In_105);
xnor U8198 (N_8198,In_2087,In_1379);
nor U8199 (N_8199,In_1978,In_36);
nand U8200 (N_8200,In_106,In_2371);
or U8201 (N_8201,In_828,In_701);
nor U8202 (N_8202,In_646,In_1078);
or U8203 (N_8203,In_2883,In_1612);
nor U8204 (N_8204,In_1380,In_1080);
nand U8205 (N_8205,In_1831,In_1060);
and U8206 (N_8206,In_1001,In_2737);
and U8207 (N_8207,In_2312,In_1912);
and U8208 (N_8208,In_1650,In_1255);
xnor U8209 (N_8209,In_910,In_2830);
nand U8210 (N_8210,In_1579,In_234);
nand U8211 (N_8211,In_952,In_2341);
nand U8212 (N_8212,In_1028,In_672);
and U8213 (N_8213,In_1765,In_66);
nor U8214 (N_8214,In_2178,In_1091);
or U8215 (N_8215,In_1996,In_122);
nor U8216 (N_8216,In_1768,In_1690);
or U8217 (N_8217,In_240,In_2187);
nand U8218 (N_8218,In_264,In_886);
nor U8219 (N_8219,In_2275,In_76);
and U8220 (N_8220,In_384,In_2144);
nand U8221 (N_8221,In_1018,In_1226);
nor U8222 (N_8222,In_2593,In_168);
or U8223 (N_8223,In_1435,In_1471);
nand U8224 (N_8224,In_2917,In_2482);
nor U8225 (N_8225,In_896,In_1175);
nand U8226 (N_8226,In_2979,In_1903);
and U8227 (N_8227,In_2080,In_2174);
or U8228 (N_8228,In_303,In_2009);
or U8229 (N_8229,In_2632,In_1145);
nand U8230 (N_8230,In_841,In_798);
or U8231 (N_8231,In_1758,In_1656);
nand U8232 (N_8232,In_318,In_2935);
or U8233 (N_8233,In_674,In_2);
nor U8234 (N_8234,In_2052,In_1112);
and U8235 (N_8235,In_2435,In_2781);
xor U8236 (N_8236,In_373,In_1238);
and U8237 (N_8237,In_588,In_1149);
nor U8238 (N_8238,In_1340,In_685);
nor U8239 (N_8239,In_1567,In_787);
nor U8240 (N_8240,In_308,In_1154);
or U8241 (N_8241,In_1727,In_1143);
nand U8242 (N_8242,In_555,In_299);
nand U8243 (N_8243,In_2772,In_2316);
or U8244 (N_8244,In_2145,In_164);
and U8245 (N_8245,In_152,In_2191);
or U8246 (N_8246,In_2749,In_919);
and U8247 (N_8247,In_2228,In_323);
nor U8248 (N_8248,In_1280,In_1556);
nand U8249 (N_8249,In_2804,In_666);
nand U8250 (N_8250,In_1520,In_1566);
nor U8251 (N_8251,In_2259,In_678);
xor U8252 (N_8252,In_2933,In_643);
xnor U8253 (N_8253,In_254,In_1525);
nor U8254 (N_8254,In_2715,In_959);
xor U8255 (N_8255,In_2465,In_2754);
xnor U8256 (N_8256,In_2929,In_1938);
or U8257 (N_8257,In_2310,In_2198);
or U8258 (N_8258,In_1439,In_2220);
nand U8259 (N_8259,In_461,In_1044);
and U8260 (N_8260,In_728,In_2440);
nor U8261 (N_8261,In_2150,In_960);
nor U8262 (N_8262,In_769,In_1788);
nand U8263 (N_8263,In_1712,In_1371);
nor U8264 (N_8264,In_2691,In_2336);
or U8265 (N_8265,In_2040,In_2961);
nor U8266 (N_8266,In_2411,In_150);
and U8267 (N_8267,In_2512,In_752);
and U8268 (N_8268,In_2928,In_1879);
and U8269 (N_8269,In_2626,In_404);
or U8270 (N_8270,In_1787,In_148);
nor U8271 (N_8271,In_842,In_1521);
nand U8272 (N_8272,In_1225,In_58);
nor U8273 (N_8273,In_1822,In_105);
nor U8274 (N_8274,In_2810,In_1017);
or U8275 (N_8275,In_770,In_2982);
and U8276 (N_8276,In_238,In_297);
and U8277 (N_8277,In_2681,In_916);
xor U8278 (N_8278,In_13,In_1630);
nand U8279 (N_8279,In_2264,In_1805);
nor U8280 (N_8280,In_1844,In_1924);
nor U8281 (N_8281,In_2962,In_1219);
nor U8282 (N_8282,In_2395,In_1137);
or U8283 (N_8283,In_2066,In_2268);
nand U8284 (N_8284,In_2310,In_1802);
nor U8285 (N_8285,In_2193,In_2509);
and U8286 (N_8286,In_1359,In_1879);
nor U8287 (N_8287,In_552,In_1058);
or U8288 (N_8288,In_1702,In_2155);
nor U8289 (N_8289,In_281,In_1166);
nand U8290 (N_8290,In_1972,In_774);
nor U8291 (N_8291,In_1754,In_1486);
nor U8292 (N_8292,In_1607,In_1945);
nand U8293 (N_8293,In_2075,In_1158);
or U8294 (N_8294,In_2727,In_1837);
nand U8295 (N_8295,In_1409,In_1560);
or U8296 (N_8296,In_623,In_1703);
or U8297 (N_8297,In_11,In_924);
nand U8298 (N_8298,In_564,In_2473);
nand U8299 (N_8299,In_1970,In_2548);
nor U8300 (N_8300,In_615,In_1428);
or U8301 (N_8301,In_777,In_1285);
xor U8302 (N_8302,In_2536,In_440);
xor U8303 (N_8303,In_1708,In_2957);
and U8304 (N_8304,In_371,In_2995);
or U8305 (N_8305,In_1195,In_864);
nor U8306 (N_8306,In_451,In_842);
nor U8307 (N_8307,In_1543,In_2180);
nor U8308 (N_8308,In_692,In_1687);
nand U8309 (N_8309,In_2790,In_1598);
and U8310 (N_8310,In_397,In_2896);
xnor U8311 (N_8311,In_1027,In_708);
nand U8312 (N_8312,In_1086,In_1989);
and U8313 (N_8313,In_1624,In_1319);
nand U8314 (N_8314,In_97,In_920);
nor U8315 (N_8315,In_2147,In_1192);
nand U8316 (N_8316,In_2965,In_1688);
or U8317 (N_8317,In_2379,In_1940);
nor U8318 (N_8318,In_924,In_1004);
nand U8319 (N_8319,In_438,In_550);
and U8320 (N_8320,In_284,In_1187);
xor U8321 (N_8321,In_647,In_2640);
nand U8322 (N_8322,In_826,In_465);
nor U8323 (N_8323,In_1816,In_1008);
nand U8324 (N_8324,In_1630,In_1334);
nor U8325 (N_8325,In_2461,In_2620);
or U8326 (N_8326,In_2660,In_790);
and U8327 (N_8327,In_1770,In_2515);
or U8328 (N_8328,In_1547,In_2218);
nor U8329 (N_8329,In_63,In_1078);
or U8330 (N_8330,In_327,In_1800);
or U8331 (N_8331,In_2526,In_1522);
and U8332 (N_8332,In_159,In_2361);
or U8333 (N_8333,In_1953,In_1776);
or U8334 (N_8334,In_129,In_2733);
xor U8335 (N_8335,In_2269,In_2008);
and U8336 (N_8336,In_2816,In_160);
xor U8337 (N_8337,In_104,In_728);
and U8338 (N_8338,In_241,In_2656);
xor U8339 (N_8339,In_130,In_1607);
nor U8340 (N_8340,In_1279,In_2928);
and U8341 (N_8341,In_433,In_1571);
xor U8342 (N_8342,In_2640,In_2154);
and U8343 (N_8343,In_2976,In_2988);
or U8344 (N_8344,In_675,In_2469);
nand U8345 (N_8345,In_466,In_1699);
or U8346 (N_8346,In_1505,In_1363);
xor U8347 (N_8347,In_2243,In_1476);
nor U8348 (N_8348,In_990,In_962);
and U8349 (N_8349,In_465,In_1503);
xnor U8350 (N_8350,In_432,In_2585);
or U8351 (N_8351,In_609,In_676);
nand U8352 (N_8352,In_1585,In_1319);
and U8353 (N_8353,In_1677,In_1874);
nor U8354 (N_8354,In_862,In_440);
nor U8355 (N_8355,In_714,In_72);
nor U8356 (N_8356,In_2939,In_363);
or U8357 (N_8357,In_2052,In_871);
nor U8358 (N_8358,In_1162,In_1265);
or U8359 (N_8359,In_1459,In_2112);
nor U8360 (N_8360,In_1862,In_987);
nand U8361 (N_8361,In_598,In_2180);
and U8362 (N_8362,In_268,In_488);
and U8363 (N_8363,In_1828,In_1299);
and U8364 (N_8364,In_2068,In_2097);
nor U8365 (N_8365,In_217,In_2945);
or U8366 (N_8366,In_1409,In_1339);
nor U8367 (N_8367,In_2923,In_2974);
nor U8368 (N_8368,In_2888,In_2473);
nand U8369 (N_8369,In_1258,In_2406);
and U8370 (N_8370,In_2856,In_2247);
nand U8371 (N_8371,In_1070,In_1496);
xor U8372 (N_8372,In_1228,In_1231);
and U8373 (N_8373,In_1017,In_2835);
nand U8374 (N_8374,In_2220,In_685);
or U8375 (N_8375,In_1940,In_2629);
nor U8376 (N_8376,In_1075,In_1615);
or U8377 (N_8377,In_795,In_2351);
nor U8378 (N_8378,In_1584,In_198);
or U8379 (N_8379,In_2086,In_1036);
or U8380 (N_8380,In_2399,In_2195);
nor U8381 (N_8381,In_1075,In_2277);
and U8382 (N_8382,In_1511,In_1886);
xnor U8383 (N_8383,In_44,In_498);
nor U8384 (N_8384,In_1574,In_1825);
and U8385 (N_8385,In_1468,In_520);
or U8386 (N_8386,In_2245,In_2686);
nor U8387 (N_8387,In_201,In_2054);
or U8388 (N_8388,In_743,In_1078);
and U8389 (N_8389,In_1147,In_2667);
xor U8390 (N_8390,In_2127,In_998);
and U8391 (N_8391,In_2762,In_2531);
nand U8392 (N_8392,In_988,In_972);
nand U8393 (N_8393,In_1115,In_1240);
xor U8394 (N_8394,In_147,In_712);
nor U8395 (N_8395,In_2352,In_1739);
or U8396 (N_8396,In_1788,In_813);
or U8397 (N_8397,In_954,In_1382);
or U8398 (N_8398,In_824,In_1316);
and U8399 (N_8399,In_584,In_2817);
xnor U8400 (N_8400,In_2631,In_2061);
nand U8401 (N_8401,In_1666,In_1780);
or U8402 (N_8402,In_2973,In_623);
or U8403 (N_8403,In_1384,In_2606);
xnor U8404 (N_8404,In_297,In_1641);
or U8405 (N_8405,In_39,In_2776);
nand U8406 (N_8406,In_1590,In_505);
and U8407 (N_8407,In_1979,In_457);
nand U8408 (N_8408,In_2276,In_865);
and U8409 (N_8409,In_59,In_190);
nand U8410 (N_8410,In_1678,In_617);
and U8411 (N_8411,In_153,In_1012);
and U8412 (N_8412,In_1561,In_2235);
nor U8413 (N_8413,In_2345,In_1234);
and U8414 (N_8414,In_617,In_987);
nor U8415 (N_8415,In_2467,In_1033);
nor U8416 (N_8416,In_450,In_120);
nor U8417 (N_8417,In_2135,In_2247);
and U8418 (N_8418,In_1401,In_877);
and U8419 (N_8419,In_1008,In_1711);
nor U8420 (N_8420,In_1301,In_2393);
nor U8421 (N_8421,In_2262,In_932);
or U8422 (N_8422,In_1120,In_1737);
nand U8423 (N_8423,In_1088,In_371);
and U8424 (N_8424,In_671,In_2618);
nor U8425 (N_8425,In_1867,In_132);
and U8426 (N_8426,In_1687,In_2651);
xor U8427 (N_8427,In_1354,In_697);
xnor U8428 (N_8428,In_2770,In_2799);
nor U8429 (N_8429,In_517,In_172);
nand U8430 (N_8430,In_1466,In_1057);
nor U8431 (N_8431,In_873,In_1418);
nor U8432 (N_8432,In_1038,In_232);
and U8433 (N_8433,In_1313,In_2302);
nor U8434 (N_8434,In_971,In_1169);
nor U8435 (N_8435,In_2054,In_2270);
nor U8436 (N_8436,In_1090,In_482);
xor U8437 (N_8437,In_532,In_1088);
nand U8438 (N_8438,In_1786,In_1331);
nand U8439 (N_8439,In_1525,In_1742);
nor U8440 (N_8440,In_1278,In_2652);
nand U8441 (N_8441,In_2430,In_1048);
nand U8442 (N_8442,In_664,In_521);
or U8443 (N_8443,In_1910,In_917);
and U8444 (N_8444,In_1919,In_2160);
xnor U8445 (N_8445,In_2891,In_2357);
and U8446 (N_8446,In_1443,In_931);
and U8447 (N_8447,In_46,In_664);
or U8448 (N_8448,In_2722,In_1750);
nand U8449 (N_8449,In_2740,In_1852);
nand U8450 (N_8450,In_2518,In_200);
xnor U8451 (N_8451,In_309,In_1758);
nand U8452 (N_8452,In_1672,In_2720);
and U8453 (N_8453,In_2589,In_1652);
or U8454 (N_8454,In_1232,In_1038);
and U8455 (N_8455,In_1218,In_2169);
nor U8456 (N_8456,In_2667,In_2548);
nand U8457 (N_8457,In_1940,In_844);
or U8458 (N_8458,In_917,In_1854);
nor U8459 (N_8459,In_2880,In_1758);
or U8460 (N_8460,In_1695,In_132);
nor U8461 (N_8461,In_387,In_2487);
nand U8462 (N_8462,In_89,In_1786);
nand U8463 (N_8463,In_1736,In_1565);
xor U8464 (N_8464,In_1941,In_2156);
and U8465 (N_8465,In_786,In_2552);
and U8466 (N_8466,In_2649,In_2058);
or U8467 (N_8467,In_741,In_2865);
or U8468 (N_8468,In_396,In_2171);
nor U8469 (N_8469,In_1671,In_2580);
and U8470 (N_8470,In_2050,In_666);
or U8471 (N_8471,In_2081,In_1483);
or U8472 (N_8472,In_645,In_2136);
xnor U8473 (N_8473,In_247,In_1651);
nand U8474 (N_8474,In_199,In_2012);
xor U8475 (N_8475,In_2384,In_593);
xor U8476 (N_8476,In_1849,In_2605);
or U8477 (N_8477,In_357,In_1258);
and U8478 (N_8478,In_1686,In_2300);
and U8479 (N_8479,In_2914,In_2598);
or U8480 (N_8480,In_1350,In_434);
nand U8481 (N_8481,In_2271,In_313);
and U8482 (N_8482,In_2987,In_2043);
nor U8483 (N_8483,In_2443,In_886);
or U8484 (N_8484,In_833,In_2014);
and U8485 (N_8485,In_168,In_2292);
nor U8486 (N_8486,In_912,In_395);
and U8487 (N_8487,In_421,In_2510);
nor U8488 (N_8488,In_1563,In_2708);
or U8489 (N_8489,In_476,In_890);
or U8490 (N_8490,In_941,In_2077);
nor U8491 (N_8491,In_530,In_171);
or U8492 (N_8492,In_938,In_1527);
or U8493 (N_8493,In_820,In_2672);
and U8494 (N_8494,In_1958,In_2193);
or U8495 (N_8495,In_748,In_1282);
or U8496 (N_8496,In_1041,In_519);
or U8497 (N_8497,In_321,In_137);
or U8498 (N_8498,In_1991,In_62);
and U8499 (N_8499,In_537,In_1456);
or U8500 (N_8500,In_2999,In_1707);
nand U8501 (N_8501,In_739,In_1573);
or U8502 (N_8502,In_1200,In_2335);
and U8503 (N_8503,In_2951,In_2691);
and U8504 (N_8504,In_1605,In_719);
or U8505 (N_8505,In_813,In_553);
or U8506 (N_8506,In_1799,In_1552);
or U8507 (N_8507,In_868,In_390);
nor U8508 (N_8508,In_356,In_549);
nand U8509 (N_8509,In_772,In_2660);
nand U8510 (N_8510,In_942,In_2065);
and U8511 (N_8511,In_18,In_283);
nor U8512 (N_8512,In_1864,In_2324);
or U8513 (N_8513,In_1583,In_1481);
xor U8514 (N_8514,In_2488,In_2447);
nor U8515 (N_8515,In_487,In_1459);
nor U8516 (N_8516,In_1408,In_1699);
and U8517 (N_8517,In_135,In_913);
and U8518 (N_8518,In_1580,In_50);
nand U8519 (N_8519,In_1255,In_1506);
nand U8520 (N_8520,In_2204,In_2711);
nand U8521 (N_8521,In_1909,In_842);
or U8522 (N_8522,In_1096,In_1252);
nand U8523 (N_8523,In_48,In_1798);
nand U8524 (N_8524,In_2664,In_2136);
or U8525 (N_8525,In_1663,In_1461);
nor U8526 (N_8526,In_869,In_486);
nor U8527 (N_8527,In_581,In_42);
nor U8528 (N_8528,In_112,In_1519);
nand U8529 (N_8529,In_2642,In_1943);
nor U8530 (N_8530,In_818,In_949);
or U8531 (N_8531,In_1496,In_2172);
and U8532 (N_8532,In_784,In_786);
and U8533 (N_8533,In_2828,In_2067);
and U8534 (N_8534,In_2947,In_506);
or U8535 (N_8535,In_146,In_2479);
and U8536 (N_8536,In_1516,In_1142);
and U8537 (N_8537,In_951,In_1298);
and U8538 (N_8538,In_2571,In_2787);
nand U8539 (N_8539,In_2003,In_1723);
and U8540 (N_8540,In_1892,In_137);
and U8541 (N_8541,In_418,In_14);
and U8542 (N_8542,In_1872,In_1812);
nor U8543 (N_8543,In_1464,In_2345);
or U8544 (N_8544,In_1623,In_2606);
and U8545 (N_8545,In_1161,In_1404);
nand U8546 (N_8546,In_1838,In_762);
nor U8547 (N_8547,In_1855,In_2838);
xnor U8548 (N_8548,In_100,In_717);
and U8549 (N_8549,In_2252,In_1891);
and U8550 (N_8550,In_2265,In_908);
xor U8551 (N_8551,In_2369,In_2877);
nor U8552 (N_8552,In_2726,In_2361);
nor U8553 (N_8553,In_84,In_2272);
nand U8554 (N_8554,In_2281,In_2406);
or U8555 (N_8555,In_2195,In_1123);
and U8556 (N_8556,In_2630,In_2804);
or U8557 (N_8557,In_1112,In_873);
nor U8558 (N_8558,In_1290,In_931);
and U8559 (N_8559,In_2861,In_1686);
nor U8560 (N_8560,In_440,In_1444);
nand U8561 (N_8561,In_134,In_1329);
nand U8562 (N_8562,In_326,In_2209);
nand U8563 (N_8563,In_1858,In_1988);
or U8564 (N_8564,In_1407,In_1342);
nor U8565 (N_8565,In_2428,In_440);
or U8566 (N_8566,In_1879,In_1688);
and U8567 (N_8567,In_1882,In_2591);
nand U8568 (N_8568,In_1936,In_1410);
nand U8569 (N_8569,In_1655,In_2831);
and U8570 (N_8570,In_354,In_1739);
nor U8571 (N_8571,In_327,In_1180);
and U8572 (N_8572,In_2738,In_1442);
or U8573 (N_8573,In_132,In_2342);
xnor U8574 (N_8574,In_397,In_1381);
nor U8575 (N_8575,In_334,In_2435);
nand U8576 (N_8576,In_2873,In_1349);
nand U8577 (N_8577,In_537,In_2250);
nand U8578 (N_8578,In_1588,In_1917);
nand U8579 (N_8579,In_947,In_1327);
nor U8580 (N_8580,In_2032,In_1803);
nand U8581 (N_8581,In_16,In_2005);
nand U8582 (N_8582,In_603,In_281);
or U8583 (N_8583,In_2568,In_2129);
nand U8584 (N_8584,In_2555,In_2526);
nand U8585 (N_8585,In_2558,In_1622);
and U8586 (N_8586,In_2702,In_2993);
or U8587 (N_8587,In_1039,In_860);
and U8588 (N_8588,In_1661,In_2894);
or U8589 (N_8589,In_553,In_1694);
nand U8590 (N_8590,In_2099,In_528);
or U8591 (N_8591,In_1760,In_1282);
or U8592 (N_8592,In_2008,In_681);
or U8593 (N_8593,In_2392,In_1370);
or U8594 (N_8594,In_1672,In_1559);
nor U8595 (N_8595,In_465,In_292);
and U8596 (N_8596,In_2474,In_2977);
nand U8597 (N_8597,In_1160,In_76);
and U8598 (N_8598,In_2066,In_1592);
nand U8599 (N_8599,In_1265,In_2177);
xor U8600 (N_8600,In_433,In_2601);
xnor U8601 (N_8601,In_25,In_1155);
or U8602 (N_8602,In_2841,In_2250);
and U8603 (N_8603,In_1465,In_1390);
nand U8604 (N_8604,In_1548,In_994);
nor U8605 (N_8605,In_2809,In_1425);
nor U8606 (N_8606,In_2942,In_2154);
nor U8607 (N_8607,In_438,In_2711);
nand U8608 (N_8608,In_1587,In_1568);
nor U8609 (N_8609,In_1193,In_2350);
and U8610 (N_8610,In_1789,In_1448);
and U8611 (N_8611,In_2815,In_762);
nand U8612 (N_8612,In_160,In_2594);
and U8613 (N_8613,In_310,In_1976);
and U8614 (N_8614,In_1793,In_2900);
nand U8615 (N_8615,In_972,In_1080);
or U8616 (N_8616,In_2712,In_1640);
and U8617 (N_8617,In_143,In_2419);
nor U8618 (N_8618,In_1986,In_2288);
or U8619 (N_8619,In_93,In_2035);
xor U8620 (N_8620,In_2202,In_1901);
or U8621 (N_8621,In_2471,In_1654);
nor U8622 (N_8622,In_709,In_1233);
or U8623 (N_8623,In_2092,In_1769);
nor U8624 (N_8624,In_1389,In_1678);
and U8625 (N_8625,In_2461,In_1293);
nand U8626 (N_8626,In_2970,In_1323);
and U8627 (N_8627,In_541,In_1706);
and U8628 (N_8628,In_1415,In_2954);
nor U8629 (N_8629,In_1301,In_1809);
nand U8630 (N_8630,In_2807,In_1735);
nor U8631 (N_8631,In_1580,In_1084);
nor U8632 (N_8632,In_850,In_2588);
nor U8633 (N_8633,In_1757,In_101);
xnor U8634 (N_8634,In_1493,In_2761);
and U8635 (N_8635,In_178,In_1947);
nor U8636 (N_8636,In_2374,In_476);
nand U8637 (N_8637,In_1663,In_123);
or U8638 (N_8638,In_1403,In_2270);
nor U8639 (N_8639,In_2082,In_978);
nand U8640 (N_8640,In_1525,In_2204);
nor U8641 (N_8641,In_439,In_2984);
or U8642 (N_8642,In_2202,In_651);
xor U8643 (N_8643,In_72,In_2978);
xor U8644 (N_8644,In_1848,In_1915);
xnor U8645 (N_8645,In_1285,In_1549);
nor U8646 (N_8646,In_1397,In_2818);
and U8647 (N_8647,In_2826,In_1167);
nand U8648 (N_8648,In_1402,In_2869);
nand U8649 (N_8649,In_2174,In_150);
and U8650 (N_8650,In_82,In_138);
and U8651 (N_8651,In_372,In_2295);
and U8652 (N_8652,In_231,In_2305);
nor U8653 (N_8653,In_1996,In_1765);
nor U8654 (N_8654,In_1736,In_1106);
nand U8655 (N_8655,In_1238,In_2571);
nand U8656 (N_8656,In_21,In_843);
or U8657 (N_8657,In_2460,In_456);
xor U8658 (N_8658,In_2107,In_2133);
nand U8659 (N_8659,In_2763,In_450);
nand U8660 (N_8660,In_613,In_1639);
nand U8661 (N_8661,In_2899,In_487);
nand U8662 (N_8662,In_2665,In_1433);
and U8663 (N_8663,In_2832,In_770);
and U8664 (N_8664,In_130,In_2523);
or U8665 (N_8665,In_2616,In_449);
nor U8666 (N_8666,In_1771,In_2026);
nand U8667 (N_8667,In_209,In_1190);
or U8668 (N_8668,In_1165,In_1330);
xnor U8669 (N_8669,In_2684,In_182);
nand U8670 (N_8670,In_2845,In_151);
and U8671 (N_8671,In_2362,In_2765);
xnor U8672 (N_8672,In_125,In_999);
or U8673 (N_8673,In_2448,In_962);
or U8674 (N_8674,In_1543,In_2052);
nand U8675 (N_8675,In_1910,In_2561);
or U8676 (N_8676,In_1245,In_273);
nor U8677 (N_8677,In_1503,In_1284);
nand U8678 (N_8678,In_2091,In_1611);
xor U8679 (N_8679,In_49,In_262);
nor U8680 (N_8680,In_252,In_1631);
or U8681 (N_8681,In_2224,In_2433);
nor U8682 (N_8682,In_1113,In_2077);
and U8683 (N_8683,In_2804,In_973);
or U8684 (N_8684,In_1067,In_222);
nor U8685 (N_8685,In_2455,In_1950);
and U8686 (N_8686,In_387,In_2228);
nor U8687 (N_8687,In_543,In_2743);
nor U8688 (N_8688,In_1515,In_2070);
nand U8689 (N_8689,In_2293,In_726);
and U8690 (N_8690,In_166,In_1354);
nand U8691 (N_8691,In_388,In_2975);
or U8692 (N_8692,In_657,In_2837);
or U8693 (N_8693,In_2772,In_1975);
nand U8694 (N_8694,In_1116,In_603);
nand U8695 (N_8695,In_2724,In_534);
and U8696 (N_8696,In_2816,In_2294);
xor U8697 (N_8697,In_1224,In_737);
nor U8698 (N_8698,In_1621,In_1704);
and U8699 (N_8699,In_1505,In_1561);
nor U8700 (N_8700,In_2904,In_1372);
nor U8701 (N_8701,In_1577,In_2708);
nor U8702 (N_8702,In_20,In_142);
nor U8703 (N_8703,In_2620,In_371);
and U8704 (N_8704,In_1337,In_1818);
nor U8705 (N_8705,In_480,In_443);
nand U8706 (N_8706,In_915,In_844);
nand U8707 (N_8707,In_1483,In_711);
or U8708 (N_8708,In_1088,In_2649);
nor U8709 (N_8709,In_2084,In_664);
and U8710 (N_8710,In_462,In_556);
nand U8711 (N_8711,In_2766,In_2702);
or U8712 (N_8712,In_108,In_314);
xnor U8713 (N_8713,In_315,In_2397);
nor U8714 (N_8714,In_2996,In_444);
nand U8715 (N_8715,In_1873,In_108);
nand U8716 (N_8716,In_1445,In_553);
and U8717 (N_8717,In_2470,In_892);
or U8718 (N_8718,In_988,In_537);
or U8719 (N_8719,In_148,In_1495);
and U8720 (N_8720,In_1459,In_2376);
nand U8721 (N_8721,In_1830,In_175);
nor U8722 (N_8722,In_514,In_2012);
nand U8723 (N_8723,In_2594,In_2140);
or U8724 (N_8724,In_2694,In_1224);
nor U8725 (N_8725,In_2209,In_1180);
and U8726 (N_8726,In_812,In_2349);
nor U8727 (N_8727,In_2347,In_2896);
and U8728 (N_8728,In_223,In_2594);
nand U8729 (N_8729,In_1750,In_2305);
nor U8730 (N_8730,In_1819,In_2429);
nand U8731 (N_8731,In_660,In_2319);
nor U8732 (N_8732,In_1984,In_1766);
nand U8733 (N_8733,In_420,In_430);
nand U8734 (N_8734,In_233,In_1163);
nor U8735 (N_8735,In_301,In_632);
nand U8736 (N_8736,In_318,In_557);
and U8737 (N_8737,In_901,In_1065);
xor U8738 (N_8738,In_676,In_778);
nand U8739 (N_8739,In_2633,In_1964);
nand U8740 (N_8740,In_358,In_553);
nor U8741 (N_8741,In_260,In_1545);
or U8742 (N_8742,In_549,In_2563);
or U8743 (N_8743,In_453,In_2431);
or U8744 (N_8744,In_799,In_960);
or U8745 (N_8745,In_1357,In_834);
or U8746 (N_8746,In_2368,In_536);
nand U8747 (N_8747,In_1699,In_1948);
xnor U8748 (N_8748,In_566,In_496);
xnor U8749 (N_8749,In_646,In_2216);
or U8750 (N_8750,In_1190,In_96);
nand U8751 (N_8751,In_128,In_2824);
xnor U8752 (N_8752,In_2119,In_11);
or U8753 (N_8753,In_777,In_316);
nand U8754 (N_8754,In_826,In_2295);
nand U8755 (N_8755,In_416,In_772);
or U8756 (N_8756,In_350,In_2905);
or U8757 (N_8757,In_2367,In_2102);
and U8758 (N_8758,In_2298,In_1254);
xnor U8759 (N_8759,In_1074,In_2395);
nor U8760 (N_8760,In_2596,In_93);
or U8761 (N_8761,In_2257,In_1349);
or U8762 (N_8762,In_2349,In_831);
and U8763 (N_8763,In_2196,In_2563);
nor U8764 (N_8764,In_2189,In_1717);
nor U8765 (N_8765,In_2881,In_1584);
nand U8766 (N_8766,In_918,In_2144);
xnor U8767 (N_8767,In_2974,In_1691);
nand U8768 (N_8768,In_562,In_2067);
or U8769 (N_8769,In_2017,In_476);
nor U8770 (N_8770,In_2035,In_74);
nor U8771 (N_8771,In_1428,In_917);
or U8772 (N_8772,In_1819,In_2845);
nand U8773 (N_8773,In_908,In_73);
or U8774 (N_8774,In_727,In_2180);
and U8775 (N_8775,In_2310,In_45);
and U8776 (N_8776,In_259,In_451);
or U8777 (N_8777,In_606,In_2892);
and U8778 (N_8778,In_126,In_2319);
nand U8779 (N_8779,In_771,In_2441);
or U8780 (N_8780,In_2707,In_2455);
and U8781 (N_8781,In_355,In_340);
or U8782 (N_8782,In_1564,In_639);
nand U8783 (N_8783,In_445,In_1808);
nand U8784 (N_8784,In_883,In_2628);
nor U8785 (N_8785,In_1919,In_2644);
and U8786 (N_8786,In_1655,In_2107);
nor U8787 (N_8787,In_1973,In_429);
nor U8788 (N_8788,In_1409,In_724);
and U8789 (N_8789,In_2687,In_2112);
nor U8790 (N_8790,In_1677,In_2589);
nand U8791 (N_8791,In_2214,In_2363);
nand U8792 (N_8792,In_2677,In_2822);
and U8793 (N_8793,In_1490,In_266);
nand U8794 (N_8794,In_420,In_1147);
nand U8795 (N_8795,In_1795,In_554);
nor U8796 (N_8796,In_2319,In_1947);
nor U8797 (N_8797,In_1128,In_1768);
or U8798 (N_8798,In_2517,In_193);
or U8799 (N_8799,In_1824,In_1364);
nor U8800 (N_8800,In_1214,In_509);
nor U8801 (N_8801,In_2334,In_1594);
and U8802 (N_8802,In_1015,In_2584);
and U8803 (N_8803,In_1472,In_581);
or U8804 (N_8804,In_608,In_2566);
nor U8805 (N_8805,In_1826,In_2746);
nand U8806 (N_8806,In_1083,In_1249);
and U8807 (N_8807,In_834,In_734);
xor U8808 (N_8808,In_2833,In_631);
nor U8809 (N_8809,In_1114,In_515);
nand U8810 (N_8810,In_1212,In_459);
nor U8811 (N_8811,In_428,In_1549);
nor U8812 (N_8812,In_2904,In_409);
nand U8813 (N_8813,In_210,In_2386);
nand U8814 (N_8814,In_912,In_2248);
nor U8815 (N_8815,In_1753,In_2442);
and U8816 (N_8816,In_512,In_1794);
or U8817 (N_8817,In_1902,In_1973);
nor U8818 (N_8818,In_1728,In_2695);
and U8819 (N_8819,In_1999,In_2428);
or U8820 (N_8820,In_2081,In_2224);
or U8821 (N_8821,In_151,In_2434);
or U8822 (N_8822,In_481,In_2152);
and U8823 (N_8823,In_861,In_2745);
and U8824 (N_8824,In_2550,In_1674);
nor U8825 (N_8825,In_2474,In_565);
or U8826 (N_8826,In_386,In_41);
or U8827 (N_8827,In_389,In_2289);
nand U8828 (N_8828,In_1948,In_2046);
nor U8829 (N_8829,In_1139,In_223);
xor U8830 (N_8830,In_1043,In_228);
or U8831 (N_8831,In_2954,In_1885);
and U8832 (N_8832,In_2295,In_1641);
or U8833 (N_8833,In_1042,In_1048);
xnor U8834 (N_8834,In_2865,In_377);
nand U8835 (N_8835,In_2577,In_992);
nor U8836 (N_8836,In_889,In_2117);
and U8837 (N_8837,In_609,In_2400);
nor U8838 (N_8838,In_2744,In_2473);
and U8839 (N_8839,In_384,In_773);
nor U8840 (N_8840,In_2958,In_133);
and U8841 (N_8841,In_1491,In_2454);
nor U8842 (N_8842,In_169,In_2501);
or U8843 (N_8843,In_640,In_2534);
or U8844 (N_8844,In_2535,In_720);
nor U8845 (N_8845,In_2464,In_1328);
and U8846 (N_8846,In_96,In_666);
or U8847 (N_8847,In_797,In_1453);
nor U8848 (N_8848,In_507,In_1984);
or U8849 (N_8849,In_516,In_986);
or U8850 (N_8850,In_425,In_1111);
and U8851 (N_8851,In_354,In_1249);
and U8852 (N_8852,In_759,In_2116);
and U8853 (N_8853,In_2346,In_2672);
nand U8854 (N_8854,In_2657,In_1087);
nor U8855 (N_8855,In_698,In_2008);
or U8856 (N_8856,In_1955,In_2369);
and U8857 (N_8857,In_2808,In_342);
nor U8858 (N_8858,In_1451,In_688);
nand U8859 (N_8859,In_308,In_1604);
nor U8860 (N_8860,In_2079,In_626);
or U8861 (N_8861,In_1692,In_2938);
xnor U8862 (N_8862,In_1294,In_1411);
or U8863 (N_8863,In_2544,In_220);
and U8864 (N_8864,In_1621,In_99);
or U8865 (N_8865,In_892,In_1980);
nor U8866 (N_8866,In_2078,In_2496);
nor U8867 (N_8867,In_1579,In_2148);
nor U8868 (N_8868,In_456,In_2722);
nor U8869 (N_8869,In_1658,In_1213);
or U8870 (N_8870,In_611,In_990);
nor U8871 (N_8871,In_1054,In_2339);
nand U8872 (N_8872,In_2157,In_1453);
nand U8873 (N_8873,In_106,In_1739);
and U8874 (N_8874,In_1903,In_2261);
xnor U8875 (N_8875,In_2169,In_2205);
xor U8876 (N_8876,In_1113,In_2485);
nand U8877 (N_8877,In_876,In_1278);
or U8878 (N_8878,In_136,In_1201);
nor U8879 (N_8879,In_2859,In_310);
nor U8880 (N_8880,In_220,In_131);
nor U8881 (N_8881,In_1765,In_2102);
or U8882 (N_8882,In_1637,In_600);
nand U8883 (N_8883,In_133,In_2168);
nand U8884 (N_8884,In_1636,In_2575);
and U8885 (N_8885,In_806,In_2421);
nand U8886 (N_8886,In_2761,In_2765);
and U8887 (N_8887,In_2484,In_1961);
nor U8888 (N_8888,In_2875,In_107);
nor U8889 (N_8889,In_2277,In_2529);
xor U8890 (N_8890,In_2688,In_2563);
and U8891 (N_8891,In_2723,In_1031);
nor U8892 (N_8892,In_2697,In_743);
or U8893 (N_8893,In_2517,In_1584);
or U8894 (N_8894,In_1597,In_762);
nand U8895 (N_8895,In_1752,In_1513);
nand U8896 (N_8896,In_188,In_1509);
and U8897 (N_8897,In_216,In_2014);
or U8898 (N_8898,In_2593,In_1011);
and U8899 (N_8899,In_1212,In_2539);
nor U8900 (N_8900,In_2220,In_2481);
and U8901 (N_8901,In_2749,In_2772);
xnor U8902 (N_8902,In_724,In_1423);
nor U8903 (N_8903,In_1086,In_2511);
xor U8904 (N_8904,In_1168,In_1253);
nor U8905 (N_8905,In_704,In_484);
nor U8906 (N_8906,In_153,In_1997);
nor U8907 (N_8907,In_2059,In_1638);
nand U8908 (N_8908,In_695,In_1463);
xor U8909 (N_8909,In_2760,In_1992);
nand U8910 (N_8910,In_544,In_1437);
nand U8911 (N_8911,In_617,In_1161);
and U8912 (N_8912,In_1391,In_2322);
nor U8913 (N_8913,In_1027,In_1939);
or U8914 (N_8914,In_1048,In_1061);
xor U8915 (N_8915,In_2349,In_1606);
nand U8916 (N_8916,In_2371,In_2871);
nand U8917 (N_8917,In_1186,In_1245);
nand U8918 (N_8918,In_1546,In_2408);
nand U8919 (N_8919,In_1428,In_1384);
or U8920 (N_8920,In_2472,In_2590);
xor U8921 (N_8921,In_343,In_1543);
or U8922 (N_8922,In_2098,In_1352);
or U8923 (N_8923,In_2386,In_1362);
and U8924 (N_8924,In_795,In_2955);
nor U8925 (N_8925,In_282,In_2006);
nor U8926 (N_8926,In_341,In_567);
nor U8927 (N_8927,In_2301,In_464);
nor U8928 (N_8928,In_288,In_2636);
or U8929 (N_8929,In_623,In_1958);
xor U8930 (N_8930,In_1723,In_2653);
and U8931 (N_8931,In_2747,In_2009);
nor U8932 (N_8932,In_1969,In_2149);
nor U8933 (N_8933,In_229,In_1034);
nand U8934 (N_8934,In_2681,In_1209);
and U8935 (N_8935,In_1790,In_1483);
nand U8936 (N_8936,In_2874,In_2516);
xnor U8937 (N_8937,In_916,In_1425);
nor U8938 (N_8938,In_2417,In_2006);
nand U8939 (N_8939,In_486,In_922);
or U8940 (N_8940,In_2723,In_282);
and U8941 (N_8941,In_283,In_2802);
nand U8942 (N_8942,In_977,In_2919);
nand U8943 (N_8943,In_2195,In_18);
nor U8944 (N_8944,In_2227,In_1786);
xnor U8945 (N_8945,In_692,In_2941);
nand U8946 (N_8946,In_2159,In_342);
nand U8947 (N_8947,In_2672,In_2656);
or U8948 (N_8948,In_2774,In_2312);
or U8949 (N_8949,In_2045,In_898);
nand U8950 (N_8950,In_2371,In_2883);
nor U8951 (N_8951,In_1434,In_908);
nand U8952 (N_8952,In_1873,In_2221);
or U8953 (N_8953,In_2152,In_1975);
xnor U8954 (N_8954,In_1231,In_1299);
nand U8955 (N_8955,In_1149,In_524);
and U8956 (N_8956,In_1405,In_1815);
nand U8957 (N_8957,In_2960,In_1826);
nand U8958 (N_8958,In_2632,In_272);
nor U8959 (N_8959,In_1522,In_1689);
and U8960 (N_8960,In_2741,In_2978);
and U8961 (N_8961,In_1163,In_1151);
nand U8962 (N_8962,In_2722,In_2668);
or U8963 (N_8963,In_298,In_2292);
nor U8964 (N_8964,In_944,In_2982);
nor U8965 (N_8965,In_1637,In_1280);
nand U8966 (N_8966,In_2857,In_283);
and U8967 (N_8967,In_2955,In_547);
nand U8968 (N_8968,In_1582,In_499);
and U8969 (N_8969,In_2577,In_2505);
or U8970 (N_8970,In_2701,In_148);
or U8971 (N_8971,In_1307,In_2433);
nand U8972 (N_8972,In_614,In_466);
nand U8973 (N_8973,In_925,In_350);
nor U8974 (N_8974,In_1243,In_10);
or U8975 (N_8975,In_2705,In_1734);
and U8976 (N_8976,In_1213,In_2171);
xor U8977 (N_8977,In_2258,In_1685);
nand U8978 (N_8978,In_2012,In_2627);
xor U8979 (N_8979,In_1941,In_1212);
nand U8980 (N_8980,In_2698,In_2146);
or U8981 (N_8981,In_2043,In_1689);
and U8982 (N_8982,In_1842,In_2887);
nor U8983 (N_8983,In_1012,In_500);
nand U8984 (N_8984,In_151,In_4);
nand U8985 (N_8985,In_1034,In_1457);
or U8986 (N_8986,In_1885,In_20);
nor U8987 (N_8987,In_1984,In_8);
or U8988 (N_8988,In_2815,In_945);
nand U8989 (N_8989,In_1637,In_2685);
nor U8990 (N_8990,In_1453,In_2838);
and U8991 (N_8991,In_1556,In_2917);
and U8992 (N_8992,In_8,In_409);
nor U8993 (N_8993,In_2377,In_2919);
or U8994 (N_8994,In_721,In_1695);
nand U8995 (N_8995,In_2534,In_970);
nand U8996 (N_8996,In_2457,In_340);
or U8997 (N_8997,In_1726,In_2382);
nor U8998 (N_8998,In_1268,In_883);
or U8999 (N_8999,In_133,In_2053);
or U9000 (N_9000,In_2288,In_1908);
and U9001 (N_9001,In_2135,In_890);
nand U9002 (N_9002,In_980,In_2379);
nor U9003 (N_9003,In_272,In_2157);
xor U9004 (N_9004,In_2751,In_81);
nand U9005 (N_9005,In_1247,In_1384);
or U9006 (N_9006,In_1862,In_1374);
and U9007 (N_9007,In_196,In_1378);
and U9008 (N_9008,In_503,In_1189);
nor U9009 (N_9009,In_1866,In_2096);
nor U9010 (N_9010,In_106,In_2117);
or U9011 (N_9011,In_1502,In_377);
or U9012 (N_9012,In_1765,In_1149);
or U9013 (N_9013,In_1327,In_2316);
or U9014 (N_9014,In_2497,In_2806);
nand U9015 (N_9015,In_2135,In_2439);
nand U9016 (N_9016,In_1954,In_792);
or U9017 (N_9017,In_2868,In_2224);
nor U9018 (N_9018,In_2515,In_1559);
nor U9019 (N_9019,In_2850,In_2895);
nand U9020 (N_9020,In_224,In_624);
and U9021 (N_9021,In_1495,In_903);
nand U9022 (N_9022,In_1076,In_1237);
or U9023 (N_9023,In_1309,In_1282);
or U9024 (N_9024,In_2808,In_484);
and U9025 (N_9025,In_384,In_1234);
nand U9026 (N_9026,In_1352,In_623);
nor U9027 (N_9027,In_1378,In_2910);
or U9028 (N_9028,In_419,In_2793);
nor U9029 (N_9029,In_1518,In_2464);
nand U9030 (N_9030,In_2486,In_1508);
and U9031 (N_9031,In_1646,In_1823);
nor U9032 (N_9032,In_2459,In_2444);
nor U9033 (N_9033,In_724,In_2809);
or U9034 (N_9034,In_913,In_2450);
nand U9035 (N_9035,In_1005,In_903);
xor U9036 (N_9036,In_2813,In_2022);
nor U9037 (N_9037,In_2125,In_720);
nand U9038 (N_9038,In_440,In_23);
and U9039 (N_9039,In_1749,In_1702);
nand U9040 (N_9040,In_222,In_117);
nor U9041 (N_9041,In_2743,In_1548);
and U9042 (N_9042,In_2258,In_1705);
nand U9043 (N_9043,In_2014,In_84);
nand U9044 (N_9044,In_293,In_902);
or U9045 (N_9045,In_1785,In_1877);
nor U9046 (N_9046,In_170,In_606);
or U9047 (N_9047,In_2000,In_1745);
xnor U9048 (N_9048,In_2468,In_1229);
or U9049 (N_9049,In_2367,In_31);
and U9050 (N_9050,In_2623,In_654);
or U9051 (N_9051,In_1928,In_924);
nor U9052 (N_9052,In_712,In_1489);
or U9053 (N_9053,In_2320,In_185);
nor U9054 (N_9054,In_477,In_2968);
or U9055 (N_9055,In_1719,In_881);
or U9056 (N_9056,In_2762,In_1463);
nand U9057 (N_9057,In_354,In_1852);
nor U9058 (N_9058,In_2300,In_1821);
nor U9059 (N_9059,In_2547,In_250);
nand U9060 (N_9060,In_1028,In_1019);
nor U9061 (N_9061,In_2685,In_742);
and U9062 (N_9062,In_1900,In_692);
and U9063 (N_9063,In_1620,In_2076);
or U9064 (N_9064,In_2506,In_2358);
and U9065 (N_9065,In_1726,In_261);
xor U9066 (N_9066,In_1533,In_2416);
and U9067 (N_9067,In_9,In_403);
xor U9068 (N_9068,In_602,In_1398);
or U9069 (N_9069,In_2159,In_2205);
or U9070 (N_9070,In_771,In_2065);
xor U9071 (N_9071,In_1437,In_446);
nor U9072 (N_9072,In_2002,In_1279);
xnor U9073 (N_9073,In_1399,In_114);
nand U9074 (N_9074,In_1423,In_2885);
xnor U9075 (N_9075,In_1927,In_53);
nand U9076 (N_9076,In_630,In_456);
nand U9077 (N_9077,In_2006,In_1702);
and U9078 (N_9078,In_2157,In_2328);
and U9079 (N_9079,In_2824,In_2309);
nand U9080 (N_9080,In_2308,In_1648);
nor U9081 (N_9081,In_604,In_2610);
or U9082 (N_9082,In_2841,In_1648);
nor U9083 (N_9083,In_656,In_2336);
nand U9084 (N_9084,In_2189,In_1055);
nor U9085 (N_9085,In_2481,In_2782);
or U9086 (N_9086,In_1315,In_770);
nand U9087 (N_9087,In_2000,In_1316);
or U9088 (N_9088,In_108,In_1174);
and U9089 (N_9089,In_841,In_1279);
xor U9090 (N_9090,In_2506,In_1340);
nand U9091 (N_9091,In_404,In_2189);
nor U9092 (N_9092,In_2409,In_1480);
nand U9093 (N_9093,In_2605,In_2020);
nor U9094 (N_9094,In_2603,In_0);
nor U9095 (N_9095,In_23,In_1649);
nor U9096 (N_9096,In_199,In_1715);
nor U9097 (N_9097,In_2240,In_2222);
nor U9098 (N_9098,In_1479,In_2874);
nor U9099 (N_9099,In_167,In_2479);
nand U9100 (N_9100,In_128,In_60);
and U9101 (N_9101,In_465,In_200);
nand U9102 (N_9102,In_2459,In_2665);
nor U9103 (N_9103,In_826,In_1365);
nand U9104 (N_9104,In_2110,In_2414);
nor U9105 (N_9105,In_29,In_1606);
and U9106 (N_9106,In_886,In_80);
and U9107 (N_9107,In_2662,In_1330);
or U9108 (N_9108,In_2006,In_513);
and U9109 (N_9109,In_1927,In_916);
nor U9110 (N_9110,In_2142,In_2290);
and U9111 (N_9111,In_24,In_1849);
nor U9112 (N_9112,In_2366,In_654);
nand U9113 (N_9113,In_1151,In_1422);
nor U9114 (N_9114,In_542,In_904);
nand U9115 (N_9115,In_2612,In_1935);
nor U9116 (N_9116,In_1475,In_2940);
nor U9117 (N_9117,In_1804,In_1733);
or U9118 (N_9118,In_1713,In_2325);
nand U9119 (N_9119,In_790,In_950);
or U9120 (N_9120,In_1956,In_287);
xor U9121 (N_9121,In_2456,In_1221);
and U9122 (N_9122,In_462,In_1019);
nor U9123 (N_9123,In_1691,In_1611);
or U9124 (N_9124,In_631,In_887);
nand U9125 (N_9125,In_2956,In_432);
and U9126 (N_9126,In_2871,In_1315);
nand U9127 (N_9127,In_2776,In_2068);
and U9128 (N_9128,In_330,In_1074);
or U9129 (N_9129,In_2636,In_2042);
or U9130 (N_9130,In_740,In_2653);
or U9131 (N_9131,In_340,In_1613);
nor U9132 (N_9132,In_30,In_2301);
nand U9133 (N_9133,In_919,In_1384);
nor U9134 (N_9134,In_1488,In_710);
and U9135 (N_9135,In_405,In_916);
or U9136 (N_9136,In_26,In_1603);
or U9137 (N_9137,In_1184,In_1065);
or U9138 (N_9138,In_1108,In_2920);
or U9139 (N_9139,In_1097,In_1043);
nor U9140 (N_9140,In_365,In_1374);
and U9141 (N_9141,In_2275,In_988);
or U9142 (N_9142,In_1133,In_2481);
nor U9143 (N_9143,In_2581,In_1514);
or U9144 (N_9144,In_2600,In_2893);
nand U9145 (N_9145,In_1376,In_1713);
or U9146 (N_9146,In_842,In_1578);
and U9147 (N_9147,In_317,In_2400);
and U9148 (N_9148,In_1790,In_2715);
nor U9149 (N_9149,In_1013,In_1277);
and U9150 (N_9150,In_581,In_2375);
and U9151 (N_9151,In_285,In_1095);
nor U9152 (N_9152,In_2284,In_1380);
nand U9153 (N_9153,In_2337,In_191);
xnor U9154 (N_9154,In_1357,In_2892);
or U9155 (N_9155,In_1051,In_2206);
or U9156 (N_9156,In_37,In_50);
nand U9157 (N_9157,In_419,In_1168);
nand U9158 (N_9158,In_565,In_1695);
and U9159 (N_9159,In_1604,In_695);
nor U9160 (N_9160,In_1066,In_2131);
xor U9161 (N_9161,In_1665,In_397);
nor U9162 (N_9162,In_2844,In_968);
xnor U9163 (N_9163,In_1781,In_341);
nand U9164 (N_9164,In_1628,In_476);
and U9165 (N_9165,In_1958,In_2640);
xnor U9166 (N_9166,In_1508,In_1880);
nor U9167 (N_9167,In_2501,In_1284);
nand U9168 (N_9168,In_303,In_2467);
nand U9169 (N_9169,In_1730,In_2134);
nand U9170 (N_9170,In_1115,In_1095);
and U9171 (N_9171,In_2757,In_1633);
nand U9172 (N_9172,In_1238,In_2194);
nor U9173 (N_9173,In_1600,In_617);
nand U9174 (N_9174,In_1467,In_2683);
xor U9175 (N_9175,In_2129,In_1710);
nand U9176 (N_9176,In_74,In_1386);
nor U9177 (N_9177,In_1164,In_566);
or U9178 (N_9178,In_825,In_2949);
nor U9179 (N_9179,In_1579,In_2175);
and U9180 (N_9180,In_1753,In_2338);
nand U9181 (N_9181,In_1314,In_213);
or U9182 (N_9182,In_2668,In_2482);
or U9183 (N_9183,In_2601,In_2129);
nand U9184 (N_9184,In_1985,In_2679);
and U9185 (N_9185,In_528,In_140);
and U9186 (N_9186,In_1607,In_2310);
nand U9187 (N_9187,In_642,In_1351);
or U9188 (N_9188,In_830,In_317);
and U9189 (N_9189,In_1187,In_530);
or U9190 (N_9190,In_1936,In_454);
nand U9191 (N_9191,In_854,In_2801);
xnor U9192 (N_9192,In_2530,In_2284);
xnor U9193 (N_9193,In_2156,In_2511);
nand U9194 (N_9194,In_2539,In_1249);
and U9195 (N_9195,In_693,In_1830);
nor U9196 (N_9196,In_2895,In_1953);
or U9197 (N_9197,In_2458,In_2292);
xor U9198 (N_9198,In_1810,In_63);
and U9199 (N_9199,In_1708,In_2619);
and U9200 (N_9200,In_2623,In_2776);
and U9201 (N_9201,In_2176,In_1442);
xnor U9202 (N_9202,In_1091,In_2522);
and U9203 (N_9203,In_1003,In_863);
nand U9204 (N_9204,In_350,In_886);
nand U9205 (N_9205,In_2625,In_946);
xnor U9206 (N_9206,In_1526,In_278);
nor U9207 (N_9207,In_1997,In_2168);
nand U9208 (N_9208,In_69,In_1383);
nand U9209 (N_9209,In_1031,In_1231);
nand U9210 (N_9210,In_2954,In_835);
nor U9211 (N_9211,In_2592,In_1668);
or U9212 (N_9212,In_509,In_2432);
nand U9213 (N_9213,In_361,In_169);
and U9214 (N_9214,In_2548,In_839);
nor U9215 (N_9215,In_2888,In_1982);
or U9216 (N_9216,In_716,In_224);
or U9217 (N_9217,In_1424,In_2569);
nor U9218 (N_9218,In_2242,In_1757);
nand U9219 (N_9219,In_2560,In_1154);
or U9220 (N_9220,In_139,In_1360);
and U9221 (N_9221,In_2019,In_995);
and U9222 (N_9222,In_1253,In_501);
or U9223 (N_9223,In_2973,In_2708);
and U9224 (N_9224,In_1316,In_2990);
or U9225 (N_9225,In_2423,In_105);
nand U9226 (N_9226,In_2856,In_140);
or U9227 (N_9227,In_2890,In_2653);
and U9228 (N_9228,In_2983,In_434);
or U9229 (N_9229,In_2524,In_385);
or U9230 (N_9230,In_628,In_2054);
or U9231 (N_9231,In_832,In_1366);
nand U9232 (N_9232,In_1343,In_81);
and U9233 (N_9233,In_1512,In_1034);
xor U9234 (N_9234,In_2645,In_168);
nand U9235 (N_9235,In_2125,In_2703);
and U9236 (N_9236,In_1122,In_2509);
nand U9237 (N_9237,In_323,In_2378);
nand U9238 (N_9238,In_960,In_1515);
or U9239 (N_9239,In_2094,In_2615);
or U9240 (N_9240,In_2791,In_382);
nor U9241 (N_9241,In_2121,In_1623);
or U9242 (N_9242,In_223,In_51);
and U9243 (N_9243,In_62,In_1508);
nor U9244 (N_9244,In_2483,In_983);
nand U9245 (N_9245,In_2491,In_762);
or U9246 (N_9246,In_1774,In_2628);
nand U9247 (N_9247,In_423,In_295);
xor U9248 (N_9248,In_2491,In_2843);
and U9249 (N_9249,In_364,In_601);
nor U9250 (N_9250,In_2685,In_483);
nor U9251 (N_9251,In_2052,In_2764);
and U9252 (N_9252,In_1879,In_1053);
or U9253 (N_9253,In_2600,In_2320);
nand U9254 (N_9254,In_591,In_2338);
nand U9255 (N_9255,In_640,In_1035);
nand U9256 (N_9256,In_2622,In_2103);
and U9257 (N_9257,In_1052,In_550);
nand U9258 (N_9258,In_2967,In_1981);
and U9259 (N_9259,In_1544,In_2134);
nor U9260 (N_9260,In_1782,In_2834);
and U9261 (N_9261,In_813,In_741);
nand U9262 (N_9262,In_1176,In_2446);
nor U9263 (N_9263,In_108,In_1785);
or U9264 (N_9264,In_680,In_2177);
nand U9265 (N_9265,In_1200,In_2311);
nand U9266 (N_9266,In_353,In_1080);
nor U9267 (N_9267,In_10,In_707);
or U9268 (N_9268,In_2208,In_395);
and U9269 (N_9269,In_51,In_624);
nand U9270 (N_9270,In_1807,In_1591);
or U9271 (N_9271,In_812,In_2865);
nor U9272 (N_9272,In_1806,In_769);
nand U9273 (N_9273,In_1606,In_1208);
nand U9274 (N_9274,In_1076,In_2212);
and U9275 (N_9275,In_2840,In_586);
and U9276 (N_9276,In_1340,In_1555);
nor U9277 (N_9277,In_2900,In_1528);
xor U9278 (N_9278,In_948,In_1170);
or U9279 (N_9279,In_1163,In_1218);
nor U9280 (N_9280,In_2368,In_175);
nand U9281 (N_9281,In_2027,In_2452);
or U9282 (N_9282,In_2651,In_1880);
nor U9283 (N_9283,In_2373,In_2107);
nand U9284 (N_9284,In_743,In_1385);
and U9285 (N_9285,In_1481,In_1762);
xor U9286 (N_9286,In_49,In_2903);
and U9287 (N_9287,In_2646,In_2818);
and U9288 (N_9288,In_838,In_677);
nand U9289 (N_9289,In_2398,In_515);
nor U9290 (N_9290,In_321,In_2026);
nand U9291 (N_9291,In_2366,In_2711);
nand U9292 (N_9292,In_2619,In_1926);
nand U9293 (N_9293,In_985,In_2124);
or U9294 (N_9294,In_1579,In_2767);
or U9295 (N_9295,In_329,In_2576);
or U9296 (N_9296,In_2102,In_764);
or U9297 (N_9297,In_637,In_1168);
and U9298 (N_9298,In_1027,In_750);
and U9299 (N_9299,In_2844,In_2425);
or U9300 (N_9300,In_2249,In_1706);
nand U9301 (N_9301,In_1893,In_1998);
or U9302 (N_9302,In_1736,In_794);
nor U9303 (N_9303,In_228,In_684);
xor U9304 (N_9304,In_2645,In_814);
nand U9305 (N_9305,In_2386,In_668);
or U9306 (N_9306,In_435,In_1466);
nand U9307 (N_9307,In_1319,In_301);
or U9308 (N_9308,In_2669,In_2973);
nand U9309 (N_9309,In_290,In_2883);
and U9310 (N_9310,In_2410,In_2032);
nor U9311 (N_9311,In_357,In_2829);
or U9312 (N_9312,In_2618,In_2435);
and U9313 (N_9313,In_2756,In_189);
nor U9314 (N_9314,In_317,In_1512);
nor U9315 (N_9315,In_659,In_792);
nand U9316 (N_9316,In_2246,In_2218);
or U9317 (N_9317,In_2763,In_1456);
and U9318 (N_9318,In_621,In_1535);
nand U9319 (N_9319,In_967,In_1317);
or U9320 (N_9320,In_1020,In_601);
or U9321 (N_9321,In_614,In_1161);
xnor U9322 (N_9322,In_2224,In_197);
nor U9323 (N_9323,In_2406,In_2830);
nand U9324 (N_9324,In_62,In_1417);
and U9325 (N_9325,In_2671,In_539);
nand U9326 (N_9326,In_728,In_2286);
and U9327 (N_9327,In_2366,In_834);
nor U9328 (N_9328,In_1281,In_2853);
or U9329 (N_9329,In_1415,In_2453);
and U9330 (N_9330,In_1279,In_1497);
xnor U9331 (N_9331,In_2385,In_1998);
nor U9332 (N_9332,In_1476,In_1944);
xor U9333 (N_9333,In_505,In_525);
nand U9334 (N_9334,In_2598,In_1348);
nor U9335 (N_9335,In_2335,In_610);
xnor U9336 (N_9336,In_1975,In_285);
xor U9337 (N_9337,In_602,In_28);
xnor U9338 (N_9338,In_2588,In_983);
or U9339 (N_9339,In_117,In_1422);
nor U9340 (N_9340,In_331,In_513);
nor U9341 (N_9341,In_1826,In_950);
xor U9342 (N_9342,In_1354,In_2513);
xor U9343 (N_9343,In_1135,In_2025);
and U9344 (N_9344,In_343,In_1196);
and U9345 (N_9345,In_1307,In_2876);
or U9346 (N_9346,In_1073,In_2989);
and U9347 (N_9347,In_2466,In_1130);
and U9348 (N_9348,In_1565,In_2056);
and U9349 (N_9349,In_440,In_1669);
and U9350 (N_9350,In_1757,In_2890);
nor U9351 (N_9351,In_338,In_2101);
nor U9352 (N_9352,In_760,In_445);
nand U9353 (N_9353,In_83,In_2419);
and U9354 (N_9354,In_64,In_802);
and U9355 (N_9355,In_1036,In_1552);
or U9356 (N_9356,In_2820,In_2202);
nand U9357 (N_9357,In_2487,In_21);
and U9358 (N_9358,In_1613,In_795);
xor U9359 (N_9359,In_2231,In_2274);
nand U9360 (N_9360,In_175,In_2461);
and U9361 (N_9361,In_2601,In_1802);
or U9362 (N_9362,In_1990,In_374);
and U9363 (N_9363,In_243,In_1566);
and U9364 (N_9364,In_515,In_1131);
nor U9365 (N_9365,In_2735,In_159);
and U9366 (N_9366,In_2009,In_720);
nand U9367 (N_9367,In_380,In_2234);
xor U9368 (N_9368,In_2179,In_2139);
xor U9369 (N_9369,In_2609,In_340);
nor U9370 (N_9370,In_178,In_1117);
or U9371 (N_9371,In_70,In_2490);
or U9372 (N_9372,In_2831,In_425);
and U9373 (N_9373,In_1140,In_130);
or U9374 (N_9374,In_1821,In_2703);
xor U9375 (N_9375,In_1535,In_1794);
xnor U9376 (N_9376,In_608,In_1038);
nor U9377 (N_9377,In_2938,In_1801);
nand U9378 (N_9378,In_2296,In_1522);
nor U9379 (N_9379,In_809,In_307);
nor U9380 (N_9380,In_1971,In_2619);
and U9381 (N_9381,In_951,In_1382);
and U9382 (N_9382,In_1353,In_2873);
and U9383 (N_9383,In_1367,In_666);
and U9384 (N_9384,In_337,In_1247);
nor U9385 (N_9385,In_922,In_2453);
and U9386 (N_9386,In_2421,In_314);
or U9387 (N_9387,In_1018,In_1017);
nand U9388 (N_9388,In_2416,In_789);
or U9389 (N_9389,In_732,In_2075);
nor U9390 (N_9390,In_1893,In_90);
and U9391 (N_9391,In_2793,In_2503);
or U9392 (N_9392,In_1659,In_396);
nor U9393 (N_9393,In_1955,In_154);
or U9394 (N_9394,In_377,In_2743);
or U9395 (N_9395,In_2767,In_1978);
and U9396 (N_9396,In_2527,In_1110);
nor U9397 (N_9397,In_1189,In_2401);
or U9398 (N_9398,In_2565,In_2885);
and U9399 (N_9399,In_1854,In_2269);
xnor U9400 (N_9400,In_1637,In_2862);
xor U9401 (N_9401,In_722,In_989);
nand U9402 (N_9402,In_906,In_1038);
or U9403 (N_9403,In_2845,In_2541);
nand U9404 (N_9404,In_1757,In_2038);
and U9405 (N_9405,In_2867,In_191);
or U9406 (N_9406,In_2152,In_1048);
xnor U9407 (N_9407,In_784,In_2036);
nand U9408 (N_9408,In_1599,In_1953);
nand U9409 (N_9409,In_2897,In_1863);
nand U9410 (N_9410,In_1605,In_2356);
nor U9411 (N_9411,In_1094,In_1867);
nand U9412 (N_9412,In_549,In_662);
or U9413 (N_9413,In_2842,In_119);
nand U9414 (N_9414,In_758,In_847);
or U9415 (N_9415,In_2264,In_271);
or U9416 (N_9416,In_2669,In_599);
nor U9417 (N_9417,In_2404,In_2390);
nor U9418 (N_9418,In_2461,In_2350);
and U9419 (N_9419,In_375,In_668);
nand U9420 (N_9420,In_1529,In_1416);
or U9421 (N_9421,In_887,In_794);
or U9422 (N_9422,In_2249,In_2742);
and U9423 (N_9423,In_535,In_1687);
and U9424 (N_9424,In_505,In_1269);
nand U9425 (N_9425,In_1148,In_1206);
and U9426 (N_9426,In_177,In_2058);
or U9427 (N_9427,In_1695,In_394);
xor U9428 (N_9428,In_2405,In_115);
and U9429 (N_9429,In_1555,In_1025);
nand U9430 (N_9430,In_1289,In_1574);
nand U9431 (N_9431,In_213,In_308);
and U9432 (N_9432,In_2963,In_915);
or U9433 (N_9433,In_1872,In_545);
and U9434 (N_9434,In_2835,In_836);
nand U9435 (N_9435,In_254,In_283);
and U9436 (N_9436,In_325,In_955);
xor U9437 (N_9437,In_1661,In_212);
and U9438 (N_9438,In_1274,In_2608);
xnor U9439 (N_9439,In_1608,In_2770);
xor U9440 (N_9440,In_2928,In_973);
xnor U9441 (N_9441,In_808,In_1033);
nand U9442 (N_9442,In_980,In_149);
or U9443 (N_9443,In_785,In_429);
nor U9444 (N_9444,In_2286,In_2315);
nand U9445 (N_9445,In_503,In_2146);
nor U9446 (N_9446,In_1589,In_1840);
or U9447 (N_9447,In_1209,In_2564);
xnor U9448 (N_9448,In_430,In_1973);
nor U9449 (N_9449,In_1500,In_882);
nand U9450 (N_9450,In_1928,In_2002);
nand U9451 (N_9451,In_2927,In_1160);
nor U9452 (N_9452,In_2913,In_2329);
and U9453 (N_9453,In_1115,In_1082);
nand U9454 (N_9454,In_1160,In_1263);
or U9455 (N_9455,In_1815,In_2668);
and U9456 (N_9456,In_2325,In_654);
nor U9457 (N_9457,In_68,In_1471);
or U9458 (N_9458,In_1985,In_2161);
nand U9459 (N_9459,In_286,In_136);
nand U9460 (N_9460,In_2876,In_1338);
nor U9461 (N_9461,In_338,In_640);
nor U9462 (N_9462,In_1998,In_2889);
and U9463 (N_9463,In_1372,In_1333);
and U9464 (N_9464,In_472,In_514);
nand U9465 (N_9465,In_2324,In_964);
nand U9466 (N_9466,In_2636,In_2217);
nand U9467 (N_9467,In_2934,In_1537);
xnor U9468 (N_9468,In_2017,In_2954);
or U9469 (N_9469,In_1700,In_284);
nand U9470 (N_9470,In_2242,In_2416);
nand U9471 (N_9471,In_738,In_2255);
xnor U9472 (N_9472,In_2655,In_2906);
or U9473 (N_9473,In_2095,In_1179);
and U9474 (N_9474,In_2026,In_1430);
or U9475 (N_9475,In_1835,In_2564);
nor U9476 (N_9476,In_2081,In_314);
nor U9477 (N_9477,In_1072,In_684);
or U9478 (N_9478,In_2000,In_556);
nor U9479 (N_9479,In_2090,In_1743);
nor U9480 (N_9480,In_189,In_1541);
nor U9481 (N_9481,In_261,In_2952);
and U9482 (N_9482,In_2597,In_1676);
nand U9483 (N_9483,In_2981,In_159);
nand U9484 (N_9484,In_2466,In_1591);
and U9485 (N_9485,In_1784,In_2954);
nand U9486 (N_9486,In_1351,In_950);
and U9487 (N_9487,In_2699,In_1980);
nor U9488 (N_9488,In_605,In_2229);
nand U9489 (N_9489,In_1064,In_2290);
or U9490 (N_9490,In_1656,In_1307);
xor U9491 (N_9491,In_1362,In_1094);
xnor U9492 (N_9492,In_2110,In_2741);
or U9493 (N_9493,In_2533,In_1781);
nor U9494 (N_9494,In_104,In_2692);
nand U9495 (N_9495,In_2203,In_640);
nand U9496 (N_9496,In_1470,In_1448);
nor U9497 (N_9497,In_814,In_2367);
nand U9498 (N_9498,In_112,In_2417);
nand U9499 (N_9499,In_1654,In_534);
nor U9500 (N_9500,In_470,In_2084);
or U9501 (N_9501,In_1082,In_884);
and U9502 (N_9502,In_2363,In_2369);
nand U9503 (N_9503,In_2263,In_2292);
nand U9504 (N_9504,In_830,In_1646);
and U9505 (N_9505,In_1392,In_1068);
nor U9506 (N_9506,In_344,In_1080);
or U9507 (N_9507,In_328,In_1140);
nand U9508 (N_9508,In_1050,In_1870);
and U9509 (N_9509,In_362,In_2052);
xnor U9510 (N_9510,In_1214,In_2707);
and U9511 (N_9511,In_1141,In_277);
nor U9512 (N_9512,In_455,In_2574);
and U9513 (N_9513,In_1392,In_734);
and U9514 (N_9514,In_906,In_2843);
and U9515 (N_9515,In_2231,In_1814);
nand U9516 (N_9516,In_945,In_1348);
xor U9517 (N_9517,In_617,In_138);
xor U9518 (N_9518,In_1915,In_2150);
nand U9519 (N_9519,In_2708,In_1906);
and U9520 (N_9520,In_2953,In_2869);
and U9521 (N_9521,In_2271,In_1220);
nor U9522 (N_9522,In_1679,In_2174);
and U9523 (N_9523,In_1387,In_2615);
nor U9524 (N_9524,In_2683,In_1454);
or U9525 (N_9525,In_85,In_862);
nor U9526 (N_9526,In_2480,In_836);
or U9527 (N_9527,In_2427,In_681);
nand U9528 (N_9528,In_918,In_288);
nor U9529 (N_9529,In_617,In_1221);
and U9530 (N_9530,In_282,In_800);
nor U9531 (N_9531,In_1069,In_2608);
and U9532 (N_9532,In_2534,In_344);
and U9533 (N_9533,In_488,In_577);
or U9534 (N_9534,In_209,In_155);
nor U9535 (N_9535,In_1026,In_41);
or U9536 (N_9536,In_270,In_295);
nand U9537 (N_9537,In_2807,In_877);
nor U9538 (N_9538,In_1038,In_2763);
nor U9539 (N_9539,In_574,In_232);
or U9540 (N_9540,In_2139,In_1512);
and U9541 (N_9541,In_2111,In_2560);
nor U9542 (N_9542,In_609,In_2551);
and U9543 (N_9543,In_1591,In_2819);
xnor U9544 (N_9544,In_961,In_476);
nor U9545 (N_9545,In_633,In_2472);
and U9546 (N_9546,In_40,In_251);
nor U9547 (N_9547,In_895,In_2290);
xor U9548 (N_9548,In_2143,In_1573);
and U9549 (N_9549,In_1455,In_1424);
nand U9550 (N_9550,In_1729,In_612);
or U9551 (N_9551,In_1176,In_2221);
and U9552 (N_9552,In_2305,In_2032);
nor U9553 (N_9553,In_156,In_719);
nand U9554 (N_9554,In_1838,In_268);
nor U9555 (N_9555,In_2969,In_2941);
nand U9556 (N_9556,In_1369,In_1237);
nand U9557 (N_9557,In_2744,In_1234);
nand U9558 (N_9558,In_401,In_2041);
nor U9559 (N_9559,In_492,In_861);
and U9560 (N_9560,In_958,In_2253);
xor U9561 (N_9561,In_1087,In_1310);
nand U9562 (N_9562,In_111,In_2041);
xnor U9563 (N_9563,In_2591,In_117);
or U9564 (N_9564,In_1220,In_1890);
xor U9565 (N_9565,In_2578,In_50);
nor U9566 (N_9566,In_1859,In_41);
nand U9567 (N_9567,In_945,In_154);
nor U9568 (N_9568,In_353,In_2676);
nand U9569 (N_9569,In_1374,In_2291);
and U9570 (N_9570,In_1755,In_1829);
nor U9571 (N_9571,In_1279,In_214);
nor U9572 (N_9572,In_1530,In_1634);
and U9573 (N_9573,In_2697,In_1863);
nor U9574 (N_9574,In_1883,In_2941);
or U9575 (N_9575,In_2491,In_1910);
or U9576 (N_9576,In_2997,In_2182);
nor U9577 (N_9577,In_1976,In_313);
nor U9578 (N_9578,In_1044,In_705);
or U9579 (N_9579,In_1629,In_777);
nor U9580 (N_9580,In_427,In_2236);
nand U9581 (N_9581,In_493,In_174);
nand U9582 (N_9582,In_1637,In_1620);
nor U9583 (N_9583,In_1870,In_680);
and U9584 (N_9584,In_42,In_142);
and U9585 (N_9585,In_2698,In_453);
nand U9586 (N_9586,In_1035,In_2328);
nor U9587 (N_9587,In_730,In_1964);
and U9588 (N_9588,In_2826,In_1970);
xnor U9589 (N_9589,In_6,In_2663);
or U9590 (N_9590,In_1153,In_1732);
nand U9591 (N_9591,In_2548,In_2198);
or U9592 (N_9592,In_2792,In_1219);
or U9593 (N_9593,In_603,In_1215);
nand U9594 (N_9594,In_2094,In_2326);
xnor U9595 (N_9595,In_2138,In_1655);
or U9596 (N_9596,In_2277,In_1799);
nand U9597 (N_9597,In_1591,In_553);
nand U9598 (N_9598,In_978,In_1253);
nand U9599 (N_9599,In_2080,In_548);
nand U9600 (N_9600,In_242,In_850);
nor U9601 (N_9601,In_1441,In_1532);
nand U9602 (N_9602,In_1833,In_2953);
nand U9603 (N_9603,In_804,In_738);
nand U9604 (N_9604,In_2997,In_1429);
and U9605 (N_9605,In_2113,In_1225);
nand U9606 (N_9606,In_188,In_1480);
nand U9607 (N_9607,In_2986,In_2071);
or U9608 (N_9608,In_1626,In_1731);
or U9609 (N_9609,In_1975,In_2555);
and U9610 (N_9610,In_954,In_1046);
nor U9611 (N_9611,In_2645,In_183);
or U9612 (N_9612,In_1493,In_2863);
nand U9613 (N_9613,In_2538,In_2609);
xor U9614 (N_9614,In_157,In_507);
or U9615 (N_9615,In_162,In_1751);
nor U9616 (N_9616,In_2190,In_1322);
or U9617 (N_9617,In_1211,In_1729);
and U9618 (N_9618,In_601,In_681);
or U9619 (N_9619,In_46,In_1898);
nand U9620 (N_9620,In_1506,In_2180);
or U9621 (N_9621,In_2497,In_2783);
and U9622 (N_9622,In_431,In_285);
nand U9623 (N_9623,In_2023,In_522);
nand U9624 (N_9624,In_2034,In_2130);
nor U9625 (N_9625,In_1636,In_2005);
nor U9626 (N_9626,In_2860,In_2285);
xnor U9627 (N_9627,In_1920,In_2703);
or U9628 (N_9628,In_2384,In_1681);
or U9629 (N_9629,In_1266,In_2510);
nor U9630 (N_9630,In_202,In_2771);
nor U9631 (N_9631,In_1900,In_1459);
nand U9632 (N_9632,In_870,In_2912);
and U9633 (N_9633,In_2037,In_2959);
and U9634 (N_9634,In_1713,In_2159);
nand U9635 (N_9635,In_375,In_839);
or U9636 (N_9636,In_2772,In_403);
or U9637 (N_9637,In_1040,In_555);
nor U9638 (N_9638,In_934,In_2450);
nand U9639 (N_9639,In_602,In_2871);
nand U9640 (N_9640,In_794,In_1136);
or U9641 (N_9641,In_588,In_1641);
or U9642 (N_9642,In_707,In_2569);
or U9643 (N_9643,In_963,In_722);
or U9644 (N_9644,In_1761,In_694);
and U9645 (N_9645,In_33,In_256);
nand U9646 (N_9646,In_2465,In_616);
xor U9647 (N_9647,In_1096,In_70);
and U9648 (N_9648,In_2401,In_158);
nor U9649 (N_9649,In_264,In_1596);
xor U9650 (N_9650,In_1946,In_1482);
nor U9651 (N_9651,In_191,In_2721);
or U9652 (N_9652,In_929,In_308);
or U9653 (N_9653,In_210,In_2288);
xor U9654 (N_9654,In_2597,In_2477);
or U9655 (N_9655,In_2513,In_29);
or U9656 (N_9656,In_1977,In_1329);
and U9657 (N_9657,In_110,In_1470);
nand U9658 (N_9658,In_2297,In_1294);
xnor U9659 (N_9659,In_2112,In_2757);
nor U9660 (N_9660,In_455,In_2535);
nand U9661 (N_9661,In_2042,In_369);
nor U9662 (N_9662,In_491,In_2642);
or U9663 (N_9663,In_2235,In_267);
and U9664 (N_9664,In_964,In_2304);
or U9665 (N_9665,In_1910,In_2972);
and U9666 (N_9666,In_1029,In_890);
and U9667 (N_9667,In_2343,In_1833);
or U9668 (N_9668,In_1132,In_668);
or U9669 (N_9669,In_205,In_641);
xor U9670 (N_9670,In_1769,In_316);
nor U9671 (N_9671,In_879,In_1980);
nor U9672 (N_9672,In_1214,In_30);
and U9673 (N_9673,In_2457,In_120);
or U9674 (N_9674,In_849,In_2209);
and U9675 (N_9675,In_181,In_2428);
nor U9676 (N_9676,In_2088,In_346);
and U9677 (N_9677,In_1445,In_1180);
and U9678 (N_9678,In_397,In_483);
xnor U9679 (N_9679,In_2547,In_354);
or U9680 (N_9680,In_2828,In_1686);
nor U9681 (N_9681,In_147,In_2528);
xnor U9682 (N_9682,In_576,In_755);
and U9683 (N_9683,In_2426,In_2023);
xor U9684 (N_9684,In_1103,In_1714);
nand U9685 (N_9685,In_620,In_1781);
nor U9686 (N_9686,In_2858,In_2827);
or U9687 (N_9687,In_2139,In_1694);
and U9688 (N_9688,In_871,In_151);
and U9689 (N_9689,In_1796,In_1186);
or U9690 (N_9690,In_371,In_2403);
nand U9691 (N_9691,In_2375,In_1976);
nand U9692 (N_9692,In_2330,In_2392);
nand U9693 (N_9693,In_799,In_1925);
and U9694 (N_9694,In_2425,In_988);
xnor U9695 (N_9695,In_2551,In_1563);
nand U9696 (N_9696,In_2167,In_637);
or U9697 (N_9697,In_1783,In_2179);
or U9698 (N_9698,In_1648,In_1080);
and U9699 (N_9699,In_661,In_54);
nand U9700 (N_9700,In_1334,In_1975);
nand U9701 (N_9701,In_2912,In_1453);
nand U9702 (N_9702,In_2040,In_99);
nor U9703 (N_9703,In_1438,In_655);
or U9704 (N_9704,In_1550,In_2060);
nand U9705 (N_9705,In_2959,In_1822);
and U9706 (N_9706,In_720,In_748);
or U9707 (N_9707,In_2217,In_2334);
and U9708 (N_9708,In_1252,In_1820);
nand U9709 (N_9709,In_1798,In_518);
nor U9710 (N_9710,In_2398,In_1437);
nor U9711 (N_9711,In_991,In_2265);
and U9712 (N_9712,In_1243,In_2194);
nand U9713 (N_9713,In_925,In_2578);
and U9714 (N_9714,In_222,In_1394);
nor U9715 (N_9715,In_2437,In_2102);
nor U9716 (N_9716,In_2776,In_596);
nor U9717 (N_9717,In_2279,In_2402);
nand U9718 (N_9718,In_1956,In_1442);
nor U9719 (N_9719,In_1082,In_974);
and U9720 (N_9720,In_1262,In_591);
nand U9721 (N_9721,In_2764,In_1824);
or U9722 (N_9722,In_1933,In_978);
nand U9723 (N_9723,In_2284,In_829);
nor U9724 (N_9724,In_88,In_1718);
xor U9725 (N_9725,In_1307,In_2390);
nor U9726 (N_9726,In_1144,In_154);
nand U9727 (N_9727,In_2955,In_2999);
nor U9728 (N_9728,In_1659,In_2486);
nand U9729 (N_9729,In_1657,In_1309);
and U9730 (N_9730,In_2562,In_2304);
nand U9731 (N_9731,In_102,In_603);
nor U9732 (N_9732,In_1258,In_1822);
nor U9733 (N_9733,In_778,In_121);
nand U9734 (N_9734,In_538,In_2051);
or U9735 (N_9735,In_370,In_1040);
and U9736 (N_9736,In_2711,In_583);
nor U9737 (N_9737,In_1900,In_2919);
nand U9738 (N_9738,In_2681,In_579);
and U9739 (N_9739,In_1943,In_1642);
nor U9740 (N_9740,In_1349,In_2069);
nand U9741 (N_9741,In_224,In_2554);
nor U9742 (N_9742,In_342,In_2800);
or U9743 (N_9743,In_2219,In_770);
or U9744 (N_9744,In_2723,In_1570);
or U9745 (N_9745,In_1612,In_1080);
and U9746 (N_9746,In_2226,In_1064);
nand U9747 (N_9747,In_2575,In_1042);
and U9748 (N_9748,In_8,In_1285);
nor U9749 (N_9749,In_55,In_768);
nand U9750 (N_9750,In_988,In_2276);
or U9751 (N_9751,In_2359,In_2101);
or U9752 (N_9752,In_1204,In_212);
and U9753 (N_9753,In_1758,In_537);
and U9754 (N_9754,In_95,In_676);
and U9755 (N_9755,In_640,In_2159);
and U9756 (N_9756,In_590,In_2434);
nor U9757 (N_9757,In_1500,In_2231);
nor U9758 (N_9758,In_2026,In_1704);
or U9759 (N_9759,In_1362,In_1343);
or U9760 (N_9760,In_89,In_2307);
or U9761 (N_9761,In_1750,In_2070);
nand U9762 (N_9762,In_1589,In_1329);
nor U9763 (N_9763,In_1560,In_210);
nand U9764 (N_9764,In_194,In_742);
nor U9765 (N_9765,In_2962,In_551);
or U9766 (N_9766,In_1662,In_437);
nand U9767 (N_9767,In_1944,In_58);
nand U9768 (N_9768,In_2542,In_2859);
or U9769 (N_9769,In_1071,In_2255);
nand U9770 (N_9770,In_2854,In_1559);
nor U9771 (N_9771,In_886,In_527);
xnor U9772 (N_9772,In_525,In_2735);
and U9773 (N_9773,In_288,In_1893);
and U9774 (N_9774,In_21,In_2879);
and U9775 (N_9775,In_1835,In_2958);
nand U9776 (N_9776,In_2805,In_175);
and U9777 (N_9777,In_2672,In_902);
nor U9778 (N_9778,In_1207,In_457);
nand U9779 (N_9779,In_2128,In_1502);
nor U9780 (N_9780,In_1051,In_2415);
nand U9781 (N_9781,In_2741,In_565);
and U9782 (N_9782,In_1543,In_814);
and U9783 (N_9783,In_1566,In_2005);
nand U9784 (N_9784,In_2444,In_271);
nor U9785 (N_9785,In_2773,In_921);
or U9786 (N_9786,In_850,In_2543);
nand U9787 (N_9787,In_2103,In_92);
nand U9788 (N_9788,In_2496,In_1069);
nand U9789 (N_9789,In_1444,In_2568);
or U9790 (N_9790,In_904,In_1884);
and U9791 (N_9791,In_2116,In_2525);
nor U9792 (N_9792,In_2236,In_2174);
nand U9793 (N_9793,In_1331,In_696);
xor U9794 (N_9794,In_866,In_890);
nor U9795 (N_9795,In_588,In_2502);
or U9796 (N_9796,In_2843,In_1782);
nor U9797 (N_9797,In_1319,In_1876);
or U9798 (N_9798,In_206,In_1830);
or U9799 (N_9799,In_1541,In_1557);
nor U9800 (N_9800,In_2353,In_2798);
and U9801 (N_9801,In_1585,In_1104);
nor U9802 (N_9802,In_402,In_1561);
or U9803 (N_9803,In_2858,In_2544);
nor U9804 (N_9804,In_966,In_1947);
or U9805 (N_9805,In_2290,In_1785);
or U9806 (N_9806,In_627,In_1128);
nor U9807 (N_9807,In_18,In_1198);
and U9808 (N_9808,In_554,In_454);
nor U9809 (N_9809,In_11,In_1736);
nor U9810 (N_9810,In_1639,In_1448);
and U9811 (N_9811,In_2636,In_625);
nand U9812 (N_9812,In_2535,In_288);
and U9813 (N_9813,In_1318,In_21);
nand U9814 (N_9814,In_1702,In_441);
or U9815 (N_9815,In_326,In_382);
nor U9816 (N_9816,In_2098,In_473);
or U9817 (N_9817,In_1052,In_2185);
or U9818 (N_9818,In_85,In_803);
and U9819 (N_9819,In_93,In_1744);
nand U9820 (N_9820,In_2710,In_1990);
xor U9821 (N_9821,In_1060,In_2490);
or U9822 (N_9822,In_92,In_804);
nand U9823 (N_9823,In_2078,In_528);
and U9824 (N_9824,In_215,In_1100);
or U9825 (N_9825,In_601,In_919);
nor U9826 (N_9826,In_164,In_2627);
or U9827 (N_9827,In_652,In_94);
nand U9828 (N_9828,In_982,In_2148);
xnor U9829 (N_9829,In_2460,In_1566);
and U9830 (N_9830,In_1877,In_2885);
nor U9831 (N_9831,In_2316,In_2507);
nand U9832 (N_9832,In_2749,In_324);
or U9833 (N_9833,In_1149,In_2816);
nor U9834 (N_9834,In_2370,In_2359);
nand U9835 (N_9835,In_227,In_797);
nand U9836 (N_9836,In_2973,In_2013);
and U9837 (N_9837,In_2133,In_34);
or U9838 (N_9838,In_304,In_54);
nor U9839 (N_9839,In_2090,In_2943);
nor U9840 (N_9840,In_2734,In_134);
nor U9841 (N_9841,In_66,In_432);
or U9842 (N_9842,In_1771,In_163);
and U9843 (N_9843,In_2484,In_718);
or U9844 (N_9844,In_584,In_29);
or U9845 (N_9845,In_2247,In_1677);
nor U9846 (N_9846,In_2307,In_1044);
and U9847 (N_9847,In_792,In_2365);
or U9848 (N_9848,In_489,In_2060);
xor U9849 (N_9849,In_770,In_1340);
or U9850 (N_9850,In_1368,In_1401);
nor U9851 (N_9851,In_2295,In_2460);
and U9852 (N_9852,In_1856,In_870);
and U9853 (N_9853,In_2843,In_1994);
nand U9854 (N_9854,In_1685,In_265);
nor U9855 (N_9855,In_1160,In_2090);
and U9856 (N_9856,In_998,In_2484);
or U9857 (N_9857,In_1317,In_1549);
and U9858 (N_9858,In_695,In_1843);
or U9859 (N_9859,In_1575,In_2916);
nand U9860 (N_9860,In_845,In_1286);
and U9861 (N_9861,In_704,In_428);
nand U9862 (N_9862,In_2860,In_260);
xor U9863 (N_9863,In_1018,In_1641);
and U9864 (N_9864,In_29,In_1577);
xor U9865 (N_9865,In_2398,In_318);
nand U9866 (N_9866,In_858,In_18);
and U9867 (N_9867,In_1845,In_742);
nor U9868 (N_9868,In_1784,In_1176);
and U9869 (N_9869,In_2419,In_967);
xnor U9870 (N_9870,In_2117,In_914);
nand U9871 (N_9871,In_1930,In_1447);
or U9872 (N_9872,In_251,In_976);
nor U9873 (N_9873,In_491,In_1001);
and U9874 (N_9874,In_1190,In_2108);
nor U9875 (N_9875,In_2814,In_1028);
xnor U9876 (N_9876,In_581,In_2350);
or U9877 (N_9877,In_1688,In_556);
and U9878 (N_9878,In_1601,In_2270);
nand U9879 (N_9879,In_2554,In_1061);
or U9880 (N_9880,In_899,In_2041);
nor U9881 (N_9881,In_875,In_1452);
and U9882 (N_9882,In_1075,In_1048);
and U9883 (N_9883,In_168,In_2032);
nor U9884 (N_9884,In_495,In_2090);
or U9885 (N_9885,In_2454,In_2353);
nor U9886 (N_9886,In_909,In_2524);
or U9887 (N_9887,In_1992,In_2955);
nor U9888 (N_9888,In_767,In_2088);
or U9889 (N_9889,In_2165,In_2191);
nand U9890 (N_9890,In_173,In_603);
xnor U9891 (N_9891,In_1474,In_2788);
nor U9892 (N_9892,In_1301,In_1095);
nor U9893 (N_9893,In_1741,In_2595);
or U9894 (N_9894,In_1515,In_2245);
or U9895 (N_9895,In_2101,In_1475);
and U9896 (N_9896,In_2416,In_2348);
nand U9897 (N_9897,In_2025,In_1681);
nand U9898 (N_9898,In_2013,In_1399);
or U9899 (N_9899,In_1028,In_2097);
and U9900 (N_9900,In_138,In_2246);
or U9901 (N_9901,In_351,In_1287);
or U9902 (N_9902,In_888,In_106);
nor U9903 (N_9903,In_784,In_2025);
nor U9904 (N_9904,In_2842,In_295);
nor U9905 (N_9905,In_282,In_1548);
nand U9906 (N_9906,In_1729,In_533);
or U9907 (N_9907,In_2674,In_1741);
xnor U9908 (N_9908,In_2001,In_2895);
and U9909 (N_9909,In_1803,In_2502);
and U9910 (N_9910,In_934,In_2700);
nor U9911 (N_9911,In_102,In_2401);
nand U9912 (N_9912,In_29,In_2076);
nand U9913 (N_9913,In_321,In_63);
xor U9914 (N_9914,In_2905,In_1551);
or U9915 (N_9915,In_857,In_55);
nor U9916 (N_9916,In_2592,In_2278);
nand U9917 (N_9917,In_235,In_2485);
or U9918 (N_9918,In_2651,In_2499);
nand U9919 (N_9919,In_866,In_2311);
and U9920 (N_9920,In_67,In_521);
nor U9921 (N_9921,In_747,In_625);
and U9922 (N_9922,In_1693,In_2629);
and U9923 (N_9923,In_2322,In_2693);
xnor U9924 (N_9924,In_2247,In_215);
and U9925 (N_9925,In_1158,In_999);
nand U9926 (N_9926,In_1703,In_2455);
and U9927 (N_9927,In_67,In_1483);
nand U9928 (N_9928,In_1686,In_1261);
or U9929 (N_9929,In_1425,In_1598);
nor U9930 (N_9930,In_2078,In_956);
nor U9931 (N_9931,In_2505,In_953);
xnor U9932 (N_9932,In_1238,In_1607);
nand U9933 (N_9933,In_1906,In_195);
xor U9934 (N_9934,In_2404,In_237);
or U9935 (N_9935,In_2216,In_1964);
or U9936 (N_9936,In_1597,In_183);
and U9937 (N_9937,In_832,In_2355);
nor U9938 (N_9938,In_1961,In_184);
xor U9939 (N_9939,In_330,In_1318);
or U9940 (N_9940,In_1742,In_1830);
nor U9941 (N_9941,In_2426,In_2955);
xor U9942 (N_9942,In_92,In_1974);
nor U9943 (N_9943,In_91,In_455);
and U9944 (N_9944,In_738,In_362);
or U9945 (N_9945,In_671,In_2203);
nor U9946 (N_9946,In_373,In_2300);
nand U9947 (N_9947,In_750,In_598);
nor U9948 (N_9948,In_1550,In_1385);
xor U9949 (N_9949,In_1462,In_77);
and U9950 (N_9950,In_385,In_486);
and U9951 (N_9951,In_554,In_2482);
and U9952 (N_9952,In_2897,In_546);
and U9953 (N_9953,In_2132,In_447);
nor U9954 (N_9954,In_1874,In_1977);
nor U9955 (N_9955,In_2387,In_1335);
and U9956 (N_9956,In_701,In_496);
or U9957 (N_9957,In_30,In_579);
nor U9958 (N_9958,In_1107,In_2013);
or U9959 (N_9959,In_436,In_2235);
nand U9960 (N_9960,In_963,In_1898);
and U9961 (N_9961,In_357,In_1094);
nor U9962 (N_9962,In_774,In_2927);
or U9963 (N_9963,In_350,In_2036);
nor U9964 (N_9964,In_309,In_2895);
xor U9965 (N_9965,In_1684,In_847);
and U9966 (N_9966,In_746,In_2727);
and U9967 (N_9967,In_12,In_2003);
nor U9968 (N_9968,In_4,In_1152);
nand U9969 (N_9969,In_439,In_2061);
nor U9970 (N_9970,In_1412,In_108);
or U9971 (N_9971,In_2295,In_893);
or U9972 (N_9972,In_207,In_2211);
nor U9973 (N_9973,In_8,In_2274);
nand U9974 (N_9974,In_2608,In_2435);
or U9975 (N_9975,In_2812,In_1478);
or U9976 (N_9976,In_639,In_1234);
nand U9977 (N_9977,In_2441,In_2371);
xor U9978 (N_9978,In_1492,In_2733);
nand U9979 (N_9979,In_2973,In_1446);
or U9980 (N_9980,In_472,In_1551);
nand U9981 (N_9981,In_1688,In_2090);
or U9982 (N_9982,In_2991,In_2689);
and U9983 (N_9983,In_16,In_1862);
nor U9984 (N_9984,In_2780,In_91);
xnor U9985 (N_9985,In_2133,In_448);
or U9986 (N_9986,In_1934,In_1332);
or U9987 (N_9987,In_1922,In_1848);
and U9988 (N_9988,In_437,In_2997);
nand U9989 (N_9989,In_1835,In_2849);
or U9990 (N_9990,In_689,In_185);
nor U9991 (N_9991,In_223,In_2050);
and U9992 (N_9992,In_2527,In_1079);
or U9993 (N_9993,In_2323,In_2670);
xor U9994 (N_9994,In_1894,In_1152);
nand U9995 (N_9995,In_2610,In_2072);
nor U9996 (N_9996,In_130,In_1894);
nor U9997 (N_9997,In_443,In_1442);
and U9998 (N_9998,In_2544,In_967);
nand U9999 (N_9999,In_1793,In_1930);
nand U10000 (N_10000,N_8307,N_212);
or U10001 (N_10001,N_9754,N_4063);
nor U10002 (N_10002,N_7707,N_5406);
and U10003 (N_10003,N_7740,N_7331);
nor U10004 (N_10004,N_5660,N_2471);
and U10005 (N_10005,N_7163,N_5918);
xnor U10006 (N_10006,N_787,N_8709);
nor U10007 (N_10007,N_9808,N_1944);
nor U10008 (N_10008,N_240,N_7678);
nand U10009 (N_10009,N_3802,N_7757);
nand U10010 (N_10010,N_439,N_2307);
nand U10011 (N_10011,N_9122,N_5617);
xnor U10012 (N_10012,N_6599,N_969);
xnor U10013 (N_10013,N_2881,N_7866);
nor U10014 (N_10014,N_2227,N_1673);
nor U10015 (N_10015,N_3786,N_9080);
nand U10016 (N_10016,N_6899,N_9397);
nand U10017 (N_10017,N_1819,N_8653);
or U10018 (N_10018,N_6700,N_2714);
nand U10019 (N_10019,N_5117,N_6866);
nand U10020 (N_10020,N_9686,N_21);
nor U10021 (N_10021,N_9757,N_8453);
or U10022 (N_10022,N_5319,N_5059);
or U10023 (N_10023,N_3125,N_2679);
and U10024 (N_10024,N_1799,N_9094);
nor U10025 (N_10025,N_5884,N_8640);
xor U10026 (N_10026,N_5475,N_2545);
and U10027 (N_10027,N_7861,N_1757);
nand U10028 (N_10028,N_4742,N_5831);
or U10029 (N_10029,N_8589,N_9087);
nand U10030 (N_10030,N_1120,N_3626);
nand U10031 (N_10031,N_3092,N_4762);
nor U10032 (N_10032,N_5885,N_5904);
nor U10033 (N_10033,N_9371,N_8702);
and U10034 (N_10034,N_2889,N_7122);
nor U10035 (N_10035,N_4938,N_462);
and U10036 (N_10036,N_31,N_4022);
nor U10037 (N_10037,N_1561,N_126);
nand U10038 (N_10038,N_3957,N_6260);
or U10039 (N_10039,N_7726,N_1386);
nor U10040 (N_10040,N_5632,N_1192);
or U10041 (N_10041,N_5735,N_4327);
nand U10042 (N_10042,N_3034,N_7074);
or U10043 (N_10043,N_215,N_1103);
nand U10044 (N_10044,N_4065,N_943);
or U10045 (N_10045,N_7324,N_2981);
nor U10046 (N_10046,N_2111,N_3378);
and U10047 (N_10047,N_8907,N_2984);
and U10048 (N_10048,N_8260,N_6058);
nor U10049 (N_10049,N_7061,N_2280);
and U10050 (N_10050,N_5925,N_9652);
nand U10051 (N_10051,N_3598,N_8673);
and U10052 (N_10052,N_2461,N_5381);
nor U10053 (N_10053,N_2396,N_291);
nor U10054 (N_10054,N_5242,N_9509);
or U10055 (N_10055,N_568,N_6887);
nand U10056 (N_10056,N_7064,N_7858);
or U10057 (N_10057,N_5569,N_9255);
and U10058 (N_10058,N_5961,N_2053);
and U10059 (N_10059,N_7106,N_8201);
nand U10060 (N_10060,N_4399,N_9515);
nand U10061 (N_10061,N_2433,N_3989);
nand U10062 (N_10062,N_6013,N_1579);
or U10063 (N_10063,N_1572,N_705);
nand U10064 (N_10064,N_1491,N_2359);
nor U10065 (N_10065,N_1224,N_4530);
nand U10066 (N_10066,N_5626,N_4945);
xor U10067 (N_10067,N_8835,N_3245);
nand U10068 (N_10068,N_5757,N_9793);
or U10069 (N_10069,N_5678,N_4823);
and U10070 (N_10070,N_8197,N_1328);
xor U10071 (N_10071,N_1980,N_3352);
nor U10072 (N_10072,N_7268,N_1054);
nor U10073 (N_10073,N_4102,N_2482);
nor U10074 (N_10074,N_6881,N_9385);
and U10075 (N_10075,N_5267,N_9548);
xor U10076 (N_10076,N_2872,N_2963);
or U10077 (N_10077,N_3912,N_3816);
nor U10078 (N_10078,N_1449,N_607);
and U10079 (N_10079,N_2397,N_3451);
or U10080 (N_10080,N_5517,N_9843);
nand U10081 (N_10081,N_528,N_4208);
xor U10082 (N_10082,N_3376,N_3562);
xor U10083 (N_10083,N_4278,N_394);
nor U10084 (N_10084,N_4370,N_4750);
nor U10085 (N_10085,N_3143,N_915);
nor U10086 (N_10086,N_4169,N_1680);
and U10087 (N_10087,N_2052,N_4857);
or U10088 (N_10088,N_2116,N_3917);
nor U10089 (N_10089,N_7865,N_898);
and U10090 (N_10090,N_1719,N_4377);
nand U10091 (N_10091,N_1765,N_629);
xor U10092 (N_10092,N_2692,N_8927);
and U10093 (N_10093,N_8394,N_3906);
nand U10094 (N_10094,N_9677,N_2896);
or U10095 (N_10095,N_498,N_2999);
or U10096 (N_10096,N_1649,N_177);
nand U10097 (N_10097,N_6506,N_7665);
nor U10098 (N_10098,N_7084,N_4747);
nand U10099 (N_10099,N_4196,N_5848);
and U10100 (N_10100,N_8172,N_8754);
and U10101 (N_10101,N_9797,N_414);
and U10102 (N_10102,N_2712,N_2312);
or U10103 (N_10103,N_2731,N_2214);
and U10104 (N_10104,N_3889,N_4570);
or U10105 (N_10105,N_7519,N_1911);
and U10106 (N_10106,N_1418,N_1621);
nand U10107 (N_10107,N_6863,N_2757);
and U10108 (N_10108,N_6499,N_4287);
nor U10109 (N_10109,N_6782,N_9322);
and U10110 (N_10110,N_1310,N_604);
nor U10111 (N_10111,N_2842,N_9767);
nand U10112 (N_10112,N_8795,N_5328);
and U10113 (N_10113,N_504,N_259);
or U10114 (N_10114,N_2969,N_1315);
and U10115 (N_10115,N_8928,N_1422);
or U10116 (N_10116,N_3702,N_9526);
and U10117 (N_10117,N_3777,N_6318);
nor U10118 (N_10118,N_4581,N_7774);
nor U10119 (N_10119,N_4357,N_6624);
and U10120 (N_10120,N_5285,N_2763);
nand U10121 (N_10121,N_9406,N_7225);
and U10122 (N_10122,N_7343,N_315);
and U10123 (N_10123,N_3808,N_7816);
nand U10124 (N_10124,N_9824,N_2220);
nor U10125 (N_10125,N_5808,N_260);
nor U10126 (N_10126,N_2733,N_1075);
nor U10127 (N_10127,N_6463,N_2498);
nand U10128 (N_10128,N_6750,N_1909);
and U10129 (N_10129,N_5384,N_2418);
or U10130 (N_10130,N_3051,N_4703);
nor U10131 (N_10131,N_2125,N_756);
and U10132 (N_10132,N_5086,N_9773);
and U10133 (N_10133,N_9533,N_7638);
or U10134 (N_10134,N_1287,N_8265);
and U10135 (N_10135,N_168,N_5582);
nor U10136 (N_10136,N_7885,N_6213);
and U10137 (N_10137,N_636,N_5671);
nand U10138 (N_10138,N_2103,N_5623);
nor U10139 (N_10139,N_7920,N_3190);
and U10140 (N_10140,N_51,N_4461);
or U10141 (N_10141,N_6534,N_1634);
or U10142 (N_10142,N_5295,N_2010);
nand U10143 (N_10143,N_9204,N_3054);
nand U10144 (N_10144,N_6016,N_4586);
nor U10145 (N_10145,N_8430,N_3028);
or U10146 (N_10146,N_2940,N_3470);
nor U10147 (N_10147,N_9071,N_8501);
nand U10148 (N_10148,N_3605,N_3088);
xor U10149 (N_10149,N_870,N_9193);
and U10150 (N_10150,N_6989,N_984);
nor U10151 (N_10151,N_495,N_6482);
nand U10152 (N_10152,N_2862,N_2172);
and U10153 (N_10153,N_3428,N_4215);
or U10154 (N_10154,N_8091,N_5585);
or U10155 (N_10155,N_7203,N_779);
and U10156 (N_10156,N_3840,N_8002);
xnor U10157 (N_10157,N_9577,N_380);
or U10158 (N_10158,N_7512,N_3586);
nand U10159 (N_10159,N_4211,N_9092);
or U10160 (N_10160,N_3818,N_1732);
and U10161 (N_10161,N_6042,N_7206);
nand U10162 (N_10162,N_5291,N_5046);
or U10163 (N_10163,N_4415,N_3550);
and U10164 (N_10164,N_4179,N_9540);
xnor U10165 (N_10165,N_7506,N_9524);
nand U10166 (N_10166,N_4716,N_931);
or U10167 (N_10167,N_4470,N_8144);
and U10168 (N_10168,N_1949,N_1193);
nand U10169 (N_10169,N_8960,N_6731);
and U10170 (N_10170,N_9194,N_4212);
xor U10171 (N_10171,N_7109,N_7894);
xnor U10172 (N_10172,N_5587,N_1678);
nand U10173 (N_10173,N_7040,N_6931);
xnor U10174 (N_10174,N_5902,N_7712);
or U10175 (N_10175,N_1356,N_601);
or U10176 (N_10176,N_9735,N_2541);
nand U10177 (N_10177,N_7263,N_9414);
nor U10178 (N_10178,N_3518,N_7391);
and U10179 (N_10179,N_4761,N_4243);
or U10180 (N_10180,N_2023,N_3096);
nand U10181 (N_10181,N_5986,N_3899);
and U10182 (N_10182,N_4781,N_9026);
and U10183 (N_10183,N_4092,N_1772);
or U10184 (N_10184,N_4442,N_1783);
and U10185 (N_10185,N_8827,N_4804);
nor U10186 (N_10186,N_2056,N_8275);
and U10187 (N_10187,N_4558,N_4411);
nor U10188 (N_10188,N_2208,N_9552);
or U10189 (N_10189,N_2645,N_1487);
and U10190 (N_10190,N_5891,N_1974);
nor U10191 (N_10191,N_1037,N_9520);
nor U10192 (N_10192,N_1872,N_9403);
nor U10193 (N_10193,N_4512,N_4932);
nand U10194 (N_10194,N_2639,N_791);
or U10195 (N_10195,N_1601,N_6633);
nor U10196 (N_10196,N_7035,N_612);
nor U10197 (N_10197,N_3979,N_2738);
nand U10198 (N_10198,N_36,N_6230);
nor U10199 (N_10199,N_8151,N_2887);
or U10200 (N_10200,N_2577,N_2252);
or U10201 (N_10201,N_8713,N_7776);
and U10202 (N_10202,N_7448,N_4293);
or U10203 (N_10203,N_9007,N_1696);
and U10204 (N_10204,N_2070,N_2538);
and U10205 (N_10205,N_9234,N_3113);
xnor U10206 (N_10206,N_9318,N_2860);
nor U10207 (N_10207,N_4994,N_7250);
or U10208 (N_10208,N_4682,N_5203);
nor U10209 (N_10209,N_3983,N_2664);
nor U10210 (N_10210,N_8121,N_84);
nor U10211 (N_10211,N_2138,N_9489);
nor U10212 (N_10212,N_6855,N_4509);
or U10213 (N_10213,N_2580,N_7713);
nand U10214 (N_10214,N_7627,N_9813);
nor U10215 (N_10215,N_6541,N_5476);
and U10216 (N_10216,N_8328,N_6626);
or U10217 (N_10217,N_7424,N_6142);
nand U10218 (N_10218,N_8398,N_8469);
xnor U10219 (N_10219,N_4005,N_5854);
and U10220 (N_10220,N_1286,N_3938);
and U10221 (N_10221,N_3978,N_1584);
nand U10222 (N_10222,N_3279,N_18);
xor U10223 (N_10223,N_6363,N_9389);
nor U10224 (N_10224,N_1822,N_3888);
nand U10225 (N_10225,N_4156,N_6273);
and U10226 (N_10226,N_2115,N_1672);
or U10227 (N_10227,N_1902,N_9165);
xor U10228 (N_10228,N_9067,N_3966);
and U10229 (N_10229,N_7633,N_9706);
and U10230 (N_10230,N_744,N_7398);
nor U10231 (N_10231,N_5132,N_1425);
or U10232 (N_10232,N_7741,N_6780);
nand U10233 (N_10233,N_3952,N_4027);
or U10234 (N_10234,N_6919,N_9881);
or U10235 (N_10235,N_8286,N_6449);
or U10236 (N_10236,N_9140,N_3872);
or U10237 (N_10237,N_917,N_718);
or U10238 (N_10238,N_2951,N_6345);
nor U10239 (N_10239,N_5140,N_871);
xnor U10240 (N_10240,N_1162,N_5561);
and U10241 (N_10241,N_3811,N_5572);
and U10242 (N_10242,N_5622,N_7044);
or U10243 (N_10243,N_4659,N_3568);
nor U10244 (N_10244,N_1982,N_304);
and U10245 (N_10245,N_581,N_2879);
nand U10246 (N_10246,N_1829,N_8459);
or U10247 (N_10247,N_691,N_8438);
and U10248 (N_10248,N_8508,N_7418);
nor U10249 (N_10249,N_109,N_4867);
nand U10250 (N_10250,N_2950,N_2764);
nor U10251 (N_10251,N_4784,N_7188);
nand U10252 (N_10252,N_2921,N_9294);
nor U10253 (N_10253,N_8740,N_8413);
nand U10254 (N_10254,N_2836,N_417);
nand U10255 (N_10255,N_8068,N_6953);
nand U10256 (N_10256,N_4872,N_8364);
nand U10257 (N_10257,N_169,N_9812);
nor U10258 (N_10258,N_5625,N_4381);
and U10259 (N_10259,N_5021,N_3993);
and U10260 (N_10260,N_9572,N_9909);
or U10261 (N_10261,N_4889,N_5698);
and U10262 (N_10262,N_7195,N_6299);
nand U10263 (N_10263,N_3110,N_4058);
and U10264 (N_10264,N_9674,N_6166);
nor U10265 (N_10265,N_8972,N_9596);
nand U10266 (N_10266,N_7834,N_2630);
xor U10267 (N_10267,N_8171,N_9830);
nand U10268 (N_10268,N_221,N_6758);
or U10269 (N_10269,N_5564,N_4817);
nor U10270 (N_10270,N_4201,N_2583);
nand U10271 (N_10271,N_1107,N_7499);
nor U10272 (N_10272,N_6583,N_5967);
and U10273 (N_10273,N_9369,N_1860);
nand U10274 (N_10274,N_7168,N_337);
and U10275 (N_10275,N_8001,N_8076);
xnor U10276 (N_10276,N_4839,N_8473);
nor U10277 (N_10277,N_3967,N_5189);
nand U10278 (N_10278,N_9921,N_4319);
nand U10279 (N_10279,N_2027,N_5847);
or U10280 (N_10280,N_9278,N_6338);
nand U10281 (N_10281,N_7590,N_9077);
or U10282 (N_10282,N_9607,N_6153);
nor U10283 (N_10283,N_541,N_7682);
xor U10284 (N_10284,N_6477,N_8886);
or U10285 (N_10285,N_8034,N_9438);
nand U10286 (N_10286,N_1014,N_9593);
and U10287 (N_10287,N_5283,N_9857);
nand U10288 (N_10288,N_157,N_3929);
nand U10289 (N_10289,N_1709,N_4246);
nor U10290 (N_10290,N_2104,N_5290);
and U10291 (N_10291,N_5579,N_3314);
nand U10292 (N_10292,N_5802,N_9151);
and U10293 (N_10293,N_1919,N_3910);
nand U10294 (N_10294,N_4308,N_7642);
or U10295 (N_10295,N_3537,N_6031);
and U10296 (N_10296,N_6389,N_865);
and U10297 (N_10297,N_7801,N_3831);
nor U10298 (N_10298,N_6003,N_5809);
nand U10299 (N_10299,N_4059,N_709);
nand U10300 (N_10300,N_1085,N_5525);
and U10301 (N_10301,N_2505,N_5674);
nand U10302 (N_10302,N_9115,N_9619);
nand U10303 (N_10303,N_1726,N_6261);
nor U10304 (N_10304,N_595,N_1762);
or U10305 (N_10305,N_603,N_1987);
or U10306 (N_10306,N_2586,N_2225);
xnor U10307 (N_10307,N_9452,N_4134);
and U10308 (N_10308,N_1801,N_204);
nand U10309 (N_10309,N_2196,N_985);
nand U10310 (N_10310,N_5684,N_6029);
nand U10311 (N_10311,N_5062,N_1185);
and U10312 (N_10312,N_3104,N_1414);
and U10313 (N_10313,N_876,N_79);
nor U10314 (N_10314,N_7651,N_5003);
nand U10315 (N_10315,N_3366,N_1111);
nor U10316 (N_10316,N_3436,N_7259);
and U10317 (N_10317,N_5177,N_2722);
and U10318 (N_10318,N_8466,N_4503);
xnor U10319 (N_10319,N_6489,N_1301);
nor U10320 (N_10320,N_4090,N_6883);
or U10321 (N_10321,N_2633,N_672);
or U10322 (N_10322,N_2991,N_7676);
or U10323 (N_10323,N_2055,N_6958);
nor U10324 (N_10324,N_7221,N_8667);
and U10325 (N_10325,N_8272,N_7775);
nand U10326 (N_10326,N_2568,N_7284);
and U10327 (N_10327,N_8449,N_9110);
nand U10328 (N_10328,N_6717,N_2448);
nor U10329 (N_10329,N_8896,N_8029);
or U10330 (N_10330,N_1530,N_8582);
and U10331 (N_10331,N_9642,N_2624);
and U10332 (N_10332,N_6817,N_2222);
or U10333 (N_10333,N_4299,N_4680);
nor U10334 (N_10334,N_3812,N_4748);
xnor U10335 (N_10335,N_1546,N_9437);
nor U10336 (N_10336,N_1473,N_1392);
or U10337 (N_10337,N_5714,N_9055);
nor U10338 (N_10338,N_2118,N_9034);
or U10339 (N_10339,N_3707,N_8203);
and U10340 (N_10340,N_2365,N_9632);
or U10341 (N_10341,N_3915,N_2786);
and U10342 (N_10342,N_9542,N_6436);
xor U10343 (N_10343,N_8601,N_7932);
nand U10344 (N_10344,N_8780,N_1397);
nor U10345 (N_10345,N_9675,N_8958);
nor U10346 (N_10346,N_4136,N_184);
nor U10347 (N_10347,N_6041,N_3992);
xnor U10348 (N_10348,N_8490,N_197);
nor U10349 (N_10349,N_213,N_9175);
nand U10350 (N_10350,N_6146,N_5708);
nand U10351 (N_10351,N_4637,N_4041);
or U10352 (N_10352,N_2736,N_6425);
or U10353 (N_10353,N_7632,N_7677);
or U10354 (N_10354,N_957,N_4292);
nand U10355 (N_10355,N_3542,N_4921);
nand U10356 (N_10356,N_6571,N_4219);
nand U10357 (N_10357,N_349,N_6942);
nor U10358 (N_10358,N_17,N_1060);
or U10359 (N_10359,N_1666,N_7732);
and U10360 (N_10360,N_1493,N_7728);
nand U10361 (N_10361,N_4683,N_4489);
nand U10362 (N_10362,N_2597,N_5098);
xor U10363 (N_10363,N_3463,N_5194);
nor U10364 (N_10364,N_777,N_1019);
or U10365 (N_10365,N_579,N_4729);
nand U10366 (N_10366,N_6017,N_5134);
xnor U10367 (N_10367,N_8761,N_4266);
and U10368 (N_10368,N_4176,N_4900);
and U10369 (N_10369,N_9011,N_5301);
nor U10370 (N_10370,N_7285,N_5131);
nand U10371 (N_10371,N_6563,N_8805);
nor U10372 (N_10372,N_6136,N_7960);
and U10373 (N_10373,N_9459,N_3071);
nand U10374 (N_10374,N_5498,N_1331);
and U10375 (N_10375,N_5022,N_1250);
and U10376 (N_10376,N_9015,N_963);
and U10377 (N_10377,N_5262,N_1888);
nand U10378 (N_10378,N_4105,N_2144);
or U10379 (N_10379,N_4012,N_307);
nand U10380 (N_10380,N_6391,N_3907);
nor U10381 (N_10381,N_5772,N_4960);
nor U10382 (N_10382,N_9212,N_8753);
or U10383 (N_10383,N_9990,N_698);
nand U10384 (N_10384,N_2746,N_2837);
nor U10385 (N_10385,N_4796,N_820);
or U10386 (N_10386,N_2644,N_8989);
nand U10387 (N_10387,N_6638,N_5634);
and U10388 (N_10388,N_3359,N_2952);
nor U10389 (N_10389,N_7395,N_9924);
nand U10390 (N_10390,N_338,N_2354);
nand U10391 (N_10391,N_8297,N_5326);
or U10392 (N_10392,N_5064,N_4643);
or U10393 (N_10393,N_7486,N_7379);
nand U10394 (N_10394,N_4967,N_8357);
nand U10395 (N_10395,N_1953,N_2296);
and U10396 (N_10396,N_9153,N_4192);
or U10397 (N_10397,N_3047,N_8039);
or U10398 (N_10398,N_6418,N_8696);
nand U10399 (N_10399,N_6205,N_7289);
or U10400 (N_10400,N_7274,N_970);
xnor U10401 (N_10401,N_2966,N_6258);
nor U10402 (N_10402,N_4644,N_7631);
and U10403 (N_10403,N_1995,N_7294);
and U10404 (N_10404,N_1190,N_8193);
nor U10405 (N_10405,N_3180,N_9276);
or U10406 (N_10406,N_5769,N_8196);
or U10407 (N_10407,N_1376,N_5388);
or U10408 (N_10408,N_356,N_2360);
nand U10409 (N_10409,N_2537,N_2900);
or U10410 (N_10410,N_1813,N_5182);
or U10411 (N_10411,N_1237,N_118);
and U10412 (N_10412,N_5996,N_5245);
or U10413 (N_10413,N_586,N_1238);
nand U10414 (N_10414,N_7224,N_3927);
and U10415 (N_10415,N_8157,N_7852);
and U10416 (N_10416,N_1394,N_7027);
and U10417 (N_10417,N_2841,N_8758);
nor U10418 (N_10418,N_9474,N_8098);
or U10419 (N_10419,N_6343,N_9684);
and U10420 (N_10420,N_8145,N_2275);
or U10421 (N_10421,N_296,N_3412);
or U10422 (N_10422,N_3078,N_6649);
and U10423 (N_10423,N_1938,N_7969);
nand U10424 (N_10424,N_443,N_331);
nand U10425 (N_10425,N_7514,N_1086);
nand U10426 (N_10426,N_3822,N_4431);
xor U10427 (N_10427,N_885,N_7468);
nand U10428 (N_10428,N_9666,N_7217);
or U10429 (N_10429,N_6228,N_6966);
and U10430 (N_10430,N_1307,N_4147);
nor U10431 (N_10431,N_489,N_7081);
or U10432 (N_10432,N_7098,N_8917);
and U10433 (N_10433,N_9396,N_628);
nor U10434 (N_10434,N_9394,N_5739);
nand U10435 (N_10435,N_8094,N_6487);
and U10436 (N_10436,N_6116,N_6876);
nor U10437 (N_10437,N_428,N_5559);
or U10438 (N_10438,N_2798,N_8544);
nand U10439 (N_10439,N_590,N_4999);
and U10440 (N_10440,N_7002,N_6242);
and U10441 (N_10441,N_936,N_4153);
nand U10442 (N_10442,N_3491,N_2855);
nand U10443 (N_10443,N_3505,N_1255);
and U10444 (N_10444,N_1635,N_642);
nor U10445 (N_10445,N_235,N_4401);
xor U10446 (N_10446,N_5318,N_9595);
nand U10447 (N_10447,N_1859,N_4014);
nor U10448 (N_10448,N_8392,N_6006);
xnor U10449 (N_10449,N_2655,N_8683);
nand U10450 (N_10450,N_8726,N_3538);
and U10451 (N_10451,N_7891,N_7412);
and U10452 (N_10452,N_7513,N_8055);
or U10453 (N_10453,N_9494,N_2124);
or U10454 (N_10454,N_5689,N_343);
nor U10455 (N_10455,N_6945,N_2421);
xor U10456 (N_10456,N_7029,N_928);
nand U10457 (N_10457,N_5038,N_9847);
xnor U10458 (N_10458,N_3229,N_6304);
nand U10459 (N_10459,N_6212,N_3291);
nor U10460 (N_10460,N_5067,N_8672);
nand U10461 (N_10461,N_2885,N_8909);
nand U10462 (N_10462,N_7786,N_2004);
nor U10463 (N_10463,N_3798,N_4195);
xor U10464 (N_10464,N_3189,N_6083);
nor U10465 (N_10465,N_2120,N_8778);
or U10466 (N_10466,N_7771,N_1912);
nand U10467 (N_10467,N_9488,N_1102);
nand U10468 (N_10468,N_4818,N_2000);
or U10469 (N_10469,N_518,N_4406);
and U10470 (N_10470,N_4977,N_2198);
nor U10471 (N_10471,N_6977,N_1878);
or U10472 (N_10472,N_6473,N_9724);
or U10473 (N_10473,N_7384,N_2665);
nor U10474 (N_10474,N_4478,N_6347);
and U10475 (N_10475,N_4048,N_4930);
nand U10476 (N_10476,N_8823,N_9400);
or U10477 (N_10477,N_9436,N_4556);
and U10478 (N_10478,N_5125,N_3619);
and U10479 (N_10479,N_8895,N_9829);
nor U10480 (N_10480,N_3541,N_3928);
xnor U10481 (N_10481,N_6239,N_5873);
and U10482 (N_10482,N_4886,N_9364);
nand U10483 (N_10483,N_9703,N_2635);
or U10484 (N_10484,N_4206,N_9183);
nor U10485 (N_10485,N_6464,N_3453);
and U10486 (N_10486,N_3030,N_6074);
or U10487 (N_10487,N_5520,N_9424);
or U10488 (N_10488,N_1797,N_8798);
nand U10489 (N_10489,N_8208,N_1825);
or U10490 (N_10490,N_2302,N_6714);
and U10491 (N_10491,N_491,N_4053);
and U10492 (N_10492,N_8111,N_8137);
and U10493 (N_10493,N_6396,N_9744);
and U10494 (N_10494,N_9688,N_2835);
or U10495 (N_10495,N_1985,N_5822);
or U10496 (N_10496,N_6572,N_2525);
xor U10497 (N_10497,N_2877,N_3221);
or U10498 (N_10498,N_5836,N_9851);
nor U10499 (N_10499,N_1724,N_8868);
xor U10500 (N_10500,N_2241,N_7878);
xnor U10501 (N_10501,N_3079,N_9263);
or U10502 (N_10502,N_2364,N_7790);
and U10503 (N_10503,N_6685,N_6829);
nor U10504 (N_10504,N_9314,N_4238);
nand U10505 (N_10505,N_2709,N_2257);
nand U10506 (N_10506,N_3860,N_3994);
and U10507 (N_10507,N_1737,N_9074);
and U10508 (N_10508,N_4151,N_8736);
and U10509 (N_10509,N_7314,N_8477);
nand U10510 (N_10510,N_3617,N_1759);
nand U10511 (N_10511,N_1862,N_302);
nor U10512 (N_10512,N_8417,N_3852);
xnor U10513 (N_10513,N_1913,N_9029);
xor U10514 (N_10514,N_188,N_6628);
nand U10515 (N_10515,N_9907,N_887);
nand U10516 (N_10516,N_9315,N_6913);
xor U10517 (N_10517,N_7416,N_3021);
and U10518 (N_10518,N_9682,N_8335);
nand U10519 (N_10519,N_7592,N_9722);
or U10520 (N_10520,N_9466,N_4848);
and U10521 (N_10521,N_8147,N_9640);
nor U10522 (N_10522,N_771,N_3526);
nand U10523 (N_10523,N_5765,N_3884);
nor U10524 (N_10524,N_4903,N_4820);
xnor U10525 (N_10525,N_5400,N_8507);
or U10526 (N_10526,N_2935,N_7952);
nor U10527 (N_10527,N_6770,N_1364);
and U10528 (N_10528,N_8520,N_6203);
or U10529 (N_10529,N_2084,N_6063);
nand U10530 (N_10530,N_8181,N_5812);
nand U10531 (N_10531,N_3782,N_3918);
or U10532 (N_10532,N_7888,N_8178);
nor U10533 (N_10533,N_1626,N_395);
nand U10534 (N_10534,N_5544,N_9734);
or U10535 (N_10535,N_2730,N_2672);
and U10536 (N_10536,N_5447,N_9521);
nor U10537 (N_10537,N_2799,N_2200);
nor U10538 (N_10538,N_6591,N_6822);
or U10539 (N_10539,N_9645,N_6936);
nand U10540 (N_10540,N_1475,N_7430);
or U10541 (N_10541,N_2033,N_135);
and U10542 (N_10542,N_7198,N_9020);
nor U10543 (N_10543,N_2890,N_2007);
xnor U10544 (N_10544,N_8604,N_9776);
xnor U10545 (N_10545,N_7721,N_2423);
nand U10546 (N_10546,N_8655,N_3581);
nand U10547 (N_10547,N_421,N_4037);
nor U10548 (N_10548,N_1769,N_7619);
nor U10549 (N_10549,N_1627,N_6007);
and U10550 (N_10550,N_7090,N_9357);
and U10551 (N_10551,N_8067,N_65);
nor U10552 (N_10552,N_7146,N_7287);
and U10553 (N_10553,N_1650,N_1536);
nor U10554 (N_10554,N_2399,N_7591);
nand U10555 (N_10555,N_9742,N_167);
nand U10556 (N_10556,N_9362,N_2316);
nand U10557 (N_10557,N_9781,N_1395);
nand U10558 (N_10558,N_1297,N_9119);
or U10559 (N_10559,N_1676,N_5342);
nand U10560 (N_10560,N_6812,N_163);
nor U10561 (N_10561,N_7419,N_6695);
nand U10562 (N_10562,N_3681,N_1201);
nor U10563 (N_10563,N_1999,N_4397);
xor U10564 (N_10564,N_4573,N_1226);
or U10565 (N_10565,N_7515,N_5310);
nand U10566 (N_10566,N_1353,N_9625);
and U10567 (N_10567,N_566,N_6924);
nor U10568 (N_10568,N_8551,N_6381);
and U10569 (N_10569,N_1682,N_276);
nand U10570 (N_10570,N_34,N_7432);
nand U10571 (N_10571,N_5351,N_2983);
nor U10572 (N_10572,N_1450,N_1570);
nand U10573 (N_10573,N_8123,N_4394);
and U10574 (N_10574,N_1889,N_9925);
nor U10575 (N_10575,N_7093,N_3085);
nor U10576 (N_10576,N_4487,N_573);
xnor U10577 (N_10577,N_5361,N_3570);
and U10578 (N_10578,N_2187,N_6590);
or U10579 (N_10579,N_5604,N_7743);
nand U10580 (N_10580,N_9585,N_6704);
and U10581 (N_10581,N_2049,N_5951);
nand U10582 (N_10582,N_6502,N_6963);
nor U10583 (N_10583,N_509,N_4662);
or U10584 (N_10584,N_8112,N_6178);
or U10585 (N_10585,N_5049,N_8996);
or U10586 (N_10586,N_9356,N_4849);
or U10587 (N_10587,N_623,N_4162);
nor U10588 (N_10588,N_195,N_9911);
nor U10589 (N_10589,N_4913,N_6901);
and U10590 (N_10590,N_2516,N_4207);
and U10591 (N_10591,N_933,N_9177);
or U10592 (N_10592,N_7849,N_275);
xnor U10593 (N_10593,N_6814,N_9696);
and U10594 (N_10594,N_9181,N_9929);
or U10595 (N_10595,N_7421,N_2492);
nand U10596 (N_10596,N_6641,N_1308);
xnor U10597 (N_10597,N_4700,N_9731);
nor U10598 (N_10598,N_4517,N_5457);
nor U10599 (N_10599,N_8161,N_5233);
nand U10600 (N_10600,N_8024,N_982);
nor U10601 (N_10601,N_6432,N_1808);
and U10602 (N_10602,N_7055,N_8385);
nand U10603 (N_10603,N_6067,N_1031);
and U10604 (N_10604,N_7930,N_7264);
nor U10605 (N_10605,N_6501,N_2895);
xor U10606 (N_10606,N_6595,N_924);
nand U10607 (N_10607,N_6043,N_735);
nand U10608 (N_10608,N_1661,N_4837);
nand U10609 (N_10609,N_5783,N_633);
or U10610 (N_10610,N_8743,N_8467);
nand U10611 (N_10611,N_5998,N_2077);
and U10612 (N_10612,N_6891,N_4519);
nor U10613 (N_10613,N_5759,N_3951);
nand U10614 (N_10614,N_971,N_7022);
nor U10615 (N_10615,N_316,N_8221);
or U10616 (N_10616,N_1677,N_8062);
nor U10617 (N_10617,N_2022,N_2481);
or U10618 (N_10618,N_7308,N_3830);
and U10619 (N_10619,N_9979,N_9848);
and U10620 (N_10620,N_1600,N_4402);
nor U10621 (N_10621,N_9811,N_1657);
or U10622 (N_10622,N_5425,N_8234);
xor U10623 (N_10623,N_5667,N_7295);
nor U10624 (N_10624,N_6252,N_1865);
xnor U10625 (N_10625,N_2533,N_4840);
nand U10626 (N_10626,N_6483,N_2854);
or U10627 (N_10627,N_6460,N_7010);
xor U10628 (N_10628,N_3897,N_1437);
or U10629 (N_10629,N_4770,N_8256);
or U10630 (N_10630,N_4099,N_6708);
nor U10631 (N_10631,N_2034,N_5421);
nor U10632 (N_10632,N_3044,N_5641);
nand U10633 (N_10633,N_8729,N_3867);
nand U10634 (N_10634,N_1374,N_3266);
nand U10635 (N_10635,N_7269,N_5562);
or U10636 (N_10636,N_3594,N_3925);
and U10637 (N_10637,N_7358,N_7043);
nor U10638 (N_10638,N_9599,N_2372);
nor U10639 (N_10639,N_6323,N_2151);
nand U10640 (N_10640,N_5428,N_5664);
or U10641 (N_10641,N_7401,N_2338);
and U10642 (N_10642,N_7851,N_8813);
nand U10643 (N_10643,N_4190,N_1110);
nand U10644 (N_10644,N_2829,N_4916);
or U10645 (N_10645,N_4917,N_3678);
or U10646 (N_10646,N_867,N_5017);
nor U10647 (N_10647,N_8334,N_490);
and U10648 (N_10648,N_6716,N_849);
nor U10649 (N_10649,N_1388,N_375);
nor U10650 (N_10650,N_7661,N_8591);
xnor U10651 (N_10651,N_1628,N_6879);
or U10652 (N_10652,N_1513,N_6289);
nand U10653 (N_10653,N_330,N_1670);
nor U10654 (N_10654,N_6129,N_4398);
and U10655 (N_10655,N_3126,N_2087);
xnor U10656 (N_10656,N_1613,N_3148);
and U10657 (N_10657,N_6551,N_1932);
xnor U10658 (N_10658,N_6393,N_8635);
nor U10659 (N_10659,N_5792,N_1605);
and U10660 (N_10660,N_6790,N_5528);
or U10661 (N_10661,N_23,N_5914);
or U10662 (N_10662,N_3488,N_5713);
and U10663 (N_10663,N_7141,N_1137);
nand U10664 (N_10664,N_7570,N_411);
or U10665 (N_10665,N_1363,N_2643);
or U10666 (N_10666,N_4002,N_1257);
nand U10667 (N_10667,N_8744,N_3548);
nor U10668 (N_10668,N_3371,N_681);
nor U10669 (N_10669,N_4744,N_6218);
and U10670 (N_10670,N_8444,N_3280);
or U10671 (N_10671,N_9603,N_631);
nand U10672 (N_10672,N_6311,N_7617);
nor U10673 (N_10673,N_9449,N_1061);
nor U10674 (N_10674,N_6734,N_7100);
nand U10675 (N_10675,N_4507,N_3642);
xor U10676 (N_10676,N_9701,N_4484);
nand U10677 (N_10677,N_7273,N_8497);
or U10678 (N_10678,N_7905,N_2479);
nor U10679 (N_10679,N_1890,N_110);
or U10680 (N_10680,N_3954,N_3270);
and U10681 (N_10681,N_1429,N_6785);
or U10682 (N_10682,N_3657,N_5706);
and U10683 (N_10683,N_9537,N_710);
nor U10684 (N_10684,N_8479,N_3406);
or U10685 (N_10685,N_8028,N_8033);
nand U10686 (N_10686,N_9353,N_9286);
xor U10687 (N_10687,N_4922,N_3536);
nand U10688 (N_10688,N_1849,N_3424);
nor U10689 (N_10689,N_7154,N_1906);
nor U10690 (N_10690,N_7152,N_2164);
nand U10691 (N_10691,N_2748,N_7664);
and U10692 (N_10692,N_9901,N_1186);
or U10693 (N_10693,N_2467,N_6360);
or U10694 (N_10694,N_5309,N_1327);
and U10695 (N_10695,N_4342,N_151);
and U10696 (N_10696,N_2849,N_9874);
or U10697 (N_10697,N_7604,N_7306);
and U10698 (N_10698,N_8177,N_6890);
xnor U10699 (N_10699,N_9541,N_5187);
nand U10700 (N_10700,N_3864,N_8666);
nand U10701 (N_10701,N_1321,N_9308);
or U10702 (N_10702,N_1707,N_2487);
and U10703 (N_10703,N_4578,N_1771);
or U10704 (N_10704,N_5500,N_5206);
nand U10705 (N_10705,N_2347,N_4465);
nor U10706 (N_10706,N_7440,N_2542);
nand U10707 (N_10707,N_4253,N_9419);
and U10708 (N_10708,N_5596,N_2976);
xnor U10709 (N_10709,N_1140,N_9347);
nor U10710 (N_10710,N_9935,N_2389);
or U10711 (N_10711,N_9636,N_6361);
nand U10712 (N_10712,N_9501,N_368);
and U10713 (N_10713,N_2958,N_3692);
nand U10714 (N_10714,N_9553,N_9031);
and U10715 (N_10715,N_3481,N_4695);
nor U10716 (N_10716,N_5459,N_7919);
xor U10717 (N_10717,N_9021,N_1464);
nand U10718 (N_10718,N_5896,N_5247);
nor U10719 (N_10719,N_683,N_4685);
nor U10720 (N_10720,N_4490,N_9594);
xor U10721 (N_10721,N_6034,N_3972);
and U10722 (N_10722,N_794,N_5166);
and U10723 (N_10723,N_3610,N_1905);
nor U10724 (N_10724,N_3974,N_369);
or U10725 (N_10725,N_3640,N_6004);
or U10726 (N_10726,N_9482,N_521);
or U10727 (N_10727,N_8363,N_6609);
and U10728 (N_10728,N_1961,N_562);
and U10729 (N_10729,N_9864,N_6181);
nor U10730 (N_10730,N_5719,N_9457);
nor U10731 (N_10731,N_3667,N_3252);
and U10732 (N_10732,N_7436,N_7303);
nor U10733 (N_10733,N_7829,N_946);
or U10734 (N_10734,N_4975,N_5736);
nand U10735 (N_10735,N_9787,N_1994);
nand U10736 (N_10736,N_2923,N_587);
and U10737 (N_10737,N_3742,N_2783);
or U10738 (N_10738,N_1752,N_3963);
and U10739 (N_10739,N_3555,N_7356);
nor U10740 (N_10740,N_664,N_9551);
and U10741 (N_10741,N_1175,N_686);
nor U10742 (N_10742,N_8173,N_5070);
nor U10743 (N_10743,N_4521,N_9772);
nor U10744 (N_10744,N_6813,N_7176);
nor U10745 (N_10745,N_3813,N_3469);
or U10746 (N_10746,N_1496,N_2519);
and U10747 (N_10747,N_9498,N_4710);
nor U10748 (N_10748,N_2961,N_5341);
or U10749 (N_10749,N_7305,N_9836);
and U10750 (N_10750,N_8336,N_3235);
nor U10751 (N_10751,N_2604,N_2340);
and U10752 (N_10752,N_8542,N_9309);
or U10753 (N_10753,N_5815,N_4813);
nor U10754 (N_10754,N_9514,N_2810);
or U10755 (N_10755,N_1393,N_9288);
nor U10756 (N_10756,N_2908,N_4291);
and U10757 (N_10757,N_6545,N_5963);
nand U10758 (N_10758,N_6503,N_7539);
nand U10759 (N_10759,N_4137,N_8636);
nor U10760 (N_10760,N_5453,N_1177);
xor U10761 (N_10761,N_7695,N_2996);
nand U10762 (N_10762,N_2042,N_3857);
nor U10763 (N_10763,N_4705,N_7179);
and U10764 (N_10764,N_6632,N_1055);
nor U10765 (N_10765,N_271,N_137);
nand U10766 (N_10766,N_8419,N_9127);
and U10767 (N_10767,N_7954,N_7341);
and U10768 (N_10768,N_9510,N_4463);
nand U10769 (N_10769,N_9507,N_3485);
nor U10770 (N_10770,N_1280,N_4175);
and U10771 (N_10771,N_6922,N_2486);
nand U10772 (N_10772,N_6607,N_5010);
or U10773 (N_10773,N_1631,N_486);
or U10774 (N_10774,N_4446,N_3762);
nand U10775 (N_10775,N_8911,N_205);
or U10776 (N_10776,N_4275,N_8769);
or U10777 (N_10777,N_9512,N_4878);
nor U10778 (N_10778,N_3207,N_6461);
nand U10779 (N_10779,N_7899,N_2021);
or U10780 (N_10780,N_7625,N_9199);
or U10781 (N_10781,N_3820,N_6808);
or U10782 (N_10782,N_622,N_895);
or U10783 (N_10783,N_1370,N_513);
or U10784 (N_10784,N_7173,N_4720);
or U10785 (N_10785,N_8931,N_8472);
or U10786 (N_10786,N_832,N_1291);
xnor U10787 (N_10787,N_8615,N_8766);
or U10788 (N_10788,N_2267,N_3422);
nor U10789 (N_10789,N_5109,N_6558);
xor U10790 (N_10790,N_2662,N_7149);
xor U10791 (N_10791,N_5325,N_2256);
nor U10792 (N_10792,N_437,N_465);
or U10793 (N_10793,N_5006,N_8058);
or U10794 (N_10794,N_1882,N_652);
or U10795 (N_10795,N_2464,N_5908);
and U10796 (N_10796,N_7639,N_8943);
nor U10797 (N_10797,N_1092,N_3036);
or U10798 (N_10798,N_3045,N_3020);
or U10799 (N_10799,N_55,N_2146);
nand U10800 (N_10800,N_5580,N_7733);
or U10801 (N_10801,N_3108,N_1390);
or U10802 (N_10802,N_4625,N_1832);
and U10803 (N_10803,N_6241,N_8997);
or U10804 (N_10804,N_9952,N_1992);
and U10805 (N_10805,N_8462,N_2357);
nand U10806 (N_10806,N_1147,N_4335);
xnor U10807 (N_10807,N_3004,N_5041);
nor U10808 (N_10808,N_2432,N_746);
xor U10809 (N_10809,N_4550,N_87);
nor U10810 (N_10810,N_6762,N_4907);
and U10811 (N_10811,N_2013,N_5997);
xor U10812 (N_10812,N_5794,N_1811);
nor U10813 (N_10813,N_3216,N_2293);
nand U10814 (N_10814,N_2826,N_2611);
nor U10815 (N_10815,N_1415,N_429);
or U10816 (N_10816,N_7737,N_7595);
or U10817 (N_10817,N_2755,N_8369);
nor U10818 (N_10818,N_2844,N_8155);
nand U10819 (N_10819,N_5892,N_85);
and U10820 (N_10820,N_5373,N_6696);
nor U10821 (N_10821,N_9957,N_7875);
nand U10822 (N_10822,N_3065,N_5950);
and U10823 (N_10823,N_2616,N_7744);
xor U10824 (N_10824,N_8822,N_7659);
xor U10825 (N_10825,N_733,N_57);
nand U10826 (N_10826,N_9368,N_9262);
xnor U10827 (N_10827,N_2845,N_4574);
nand U10828 (N_10828,N_1578,N_3388);
and U10829 (N_10829,N_3213,N_4684);
nand U10830 (N_10830,N_5965,N_7111);
nand U10831 (N_10831,N_2501,N_1270);
or U10832 (N_10832,N_9359,N_2422);
or U10833 (N_10833,N_2093,N_3191);
xnor U10834 (N_10834,N_5537,N_385);
nor U10835 (N_10835,N_2326,N_4746);
or U10836 (N_10836,N_5120,N_880);
nand U10837 (N_10837,N_6699,N_5101);
nor U10838 (N_10838,N_8291,N_1157);
or U10839 (N_10839,N_6961,N_1778);
nor U10840 (N_10840,N_2210,N_6211);
nor U10841 (N_10841,N_6214,N_935);
nor U10842 (N_10842,N_8214,N_2590);
nand U10843 (N_10843,N_9481,N_7482);
nor U10844 (N_10844,N_8947,N_8802);
and U10845 (N_10845,N_9219,N_7406);
nor U10846 (N_10846,N_5380,N_4130);
or U10847 (N_10847,N_3164,N_7957);
xnor U10848 (N_10848,N_1172,N_6661);
or U10849 (N_10849,N_9272,N_5534);
nor U10850 (N_10850,N_336,N_1560);
and U10851 (N_10851,N_8215,N_9882);
nor U10852 (N_10852,N_5843,N_6842);
nor U10853 (N_10853,N_492,N_4594);
and U10854 (N_10854,N_3698,N_389);
nor U10855 (N_10855,N_7753,N_4616);
or U10856 (N_10856,N_677,N_6656);
and U10857 (N_10857,N_5232,N_7756);
nor U10858 (N_10858,N_96,N_3418);
or U10859 (N_10859,N_7014,N_7843);
and U10860 (N_10860,N_1684,N_6438);
nor U10861 (N_10861,N_6157,N_9791);
nand U10862 (N_10862,N_1423,N_2261);
nand U10863 (N_10863,N_7577,N_8568);
and U10864 (N_10864,N_7876,N_7385);
nand U10865 (N_10865,N_949,N_1482);
nor U10866 (N_10866,N_6327,N_6616);
nor U10867 (N_10867,N_529,N_9350);
and U10868 (N_10868,N_3752,N_9729);
xnor U10869 (N_10869,N_4111,N_2570);
or U10870 (N_10870,N_5084,N_7452);
xor U10871 (N_10871,N_6982,N_9500);
nor U10872 (N_10872,N_4325,N_3838);
nor U10873 (N_10873,N_2194,N_7808);
nand U10874 (N_10874,N_2179,N_392);
and U10875 (N_10875,N_6752,N_6328);
xor U10876 (N_10876,N_3448,N_4107);
nor U10877 (N_10877,N_10,N_6933);
nand U10878 (N_10878,N_3663,N_1833);
or U10879 (N_10879,N_108,N_6906);
or U10880 (N_10880,N_5369,N_8889);
xor U10881 (N_10881,N_1435,N_5718);
and U10882 (N_10882,N_2629,N_4160);
nor U10883 (N_10883,N_8274,N_5366);
xor U10884 (N_10884,N_2856,N_1563);
or U10885 (N_10885,N_1343,N_7117);
xnor U10886 (N_10886,N_9173,N_7438);
nor U10887 (N_10887,N_1768,N_5910);
xor U10888 (N_10888,N_702,N_7525);
nor U10889 (N_10889,N_716,N_9855);
xnor U10890 (N_10890,N_5880,N_1633);
xor U10891 (N_10891,N_5516,N_9346);
and U10892 (N_10892,N_7877,N_9663);
and U10893 (N_10893,N_8499,N_1541);
nor U10894 (N_10894,N_8955,N_9499);
nor U10895 (N_10895,N_3240,N_3686);
nand U10896 (N_10896,N_6430,N_9342);
nor U10897 (N_10897,N_4518,N_3363);
nor U10898 (N_10898,N_766,N_7917);
and U10899 (N_10899,N_8498,N_335);
or U10900 (N_10900,N_5103,N_8562);
and U10901 (N_10901,N_5092,N_1115);
nand U10902 (N_10902,N_4966,N_2589);
nand U10903 (N_10903,N_1296,N_4632);
or U10904 (N_10904,N_420,N_3624);
or U10905 (N_10905,N_7126,N_9008);
and U10906 (N_10906,N_8165,N_571);
or U10907 (N_10907,N_9853,N_9623);
and U10908 (N_10908,N_1,N_1034);
and U10909 (N_10909,N_9785,N_7359);
nand U10910 (N_10910,N_7380,N_6198);
and U10911 (N_10911,N_7102,N_7864);
nand U10912 (N_10912,N_6555,N_9422);
and U10913 (N_10913,N_6366,N_4962);
or U10914 (N_10914,N_9679,N_9260);
or U10915 (N_10915,N_862,N_5451);
and U10916 (N_10916,N_7900,N_4283);
and U10917 (N_10917,N_7780,N_1454);
nand U10918 (N_10918,N_8862,N_7994);
xnor U10919 (N_10919,N_231,N_5007);
nor U10920 (N_10920,N_2778,N_9620);
nor U10921 (N_10921,N_7000,N_3655);
and U10922 (N_10922,N_1951,N_404);
nor U10923 (N_10923,N_5814,N_2489);
and U10924 (N_10924,N_1858,N_8382);
and U10925 (N_10925,N_9867,N_5479);
xnor U10926 (N_10926,N_3615,N_8390);
and U10927 (N_10927,N_9846,N_6151);
nand U10928 (N_10928,N_1543,N_7764);
and U10929 (N_10929,N_6466,N_3850);
nor U10930 (N_10930,N_4376,N_1512);
nand U10931 (N_10931,N_4668,N_7666);
nand U10932 (N_10932,N_4629,N_4624);
or U10933 (N_10933,N_6562,N_5779);
nand U10934 (N_10934,N_4665,N_9012);
nor U10935 (N_10935,N_3227,N_2503);
and U10936 (N_10936,N_2440,N_8512);
nand U10937 (N_10937,N_4426,N_6160);
and U10938 (N_10938,N_6072,N_140);
nand U10939 (N_10939,N_3441,N_1335);
or U10940 (N_10940,N_4093,N_9230);
nor U10941 (N_10941,N_7560,N_1052);
and U10942 (N_10942,N_152,N_83);
or U10943 (N_10943,N_4936,N_5050);
nor U10944 (N_10944,N_7998,N_7862);
nand U10945 (N_10945,N_8547,N_3362);
nor U10946 (N_10946,N_9697,N_1163);
nor U10947 (N_10947,N_5523,N_3287);
or U10948 (N_10948,N_7328,N_5359);
or U10949 (N_10949,N_960,N_6237);
or U10950 (N_10950,N_1743,N_2130);
nor U10951 (N_10951,N_952,N_1033);
nand U10952 (N_10952,N_35,N_2030);
or U10953 (N_10953,N_9566,N_9704);
or U10954 (N_10954,N_2411,N_1908);
nor U10955 (N_10955,N_8788,N_5368);
nand U10956 (N_10956,N_3218,N_5820);
nor U10957 (N_10957,N_1733,N_726);
or U10958 (N_10958,N_3124,N_978);
nand U10959 (N_10959,N_9390,N_8424);
or U10960 (N_10960,N_6668,N_6023);
or U10961 (N_10961,N_3837,N_5162);
or U10962 (N_10962,N_4645,N_1013);
nor U10963 (N_10963,N_4429,N_911);
nor U10964 (N_10964,N_3271,N_3935);
nand U10965 (N_10965,N_6739,N_893);
and U10966 (N_10966,N_6411,N_3669);
nand U10967 (N_10967,N_2540,N_8093);
and U10968 (N_10968,N_2276,N_1997);
or U10969 (N_10969,N_4679,N_7530);
and U10970 (N_10970,N_9375,N_5367);
or U10971 (N_10971,N_4870,N_5390);
nor U10972 (N_10972,N_9819,N_7311);
nor U10973 (N_10973,N_8720,N_2699);
and U10974 (N_10974,N_7605,N_2609);
or U10975 (N_10975,N_3704,N_7476);
or U10976 (N_10976,N_2792,N_9713);
or U10977 (N_10977,N_9267,N_6424);
nor U10978 (N_10978,N_1842,N_6233);
nor U10979 (N_10979,N_9550,N_765);
and U10980 (N_10980,N_5921,N_3263);
and U10981 (N_10981,N_4595,N_624);
and U10982 (N_10982,N_9064,N_9852);
nand U10983 (N_10983,N_2694,N_1896);
and U10984 (N_10984,N_727,N_4996);
nor U10985 (N_10985,N_8643,N_7483);
nor U10986 (N_10986,N_7671,N_8027);
and U10987 (N_10987,N_5826,N_9254);
and U10988 (N_10988,N_1253,N_7094);
or U10989 (N_10989,N_7873,N_2818);
or U10990 (N_10990,N_4187,N_4393);
xor U10991 (N_10991,N_5100,N_7811);
nand U10992 (N_10992,N_8326,N_543);
nand U10993 (N_10993,N_5966,N_6446);
xnor U10994 (N_10994,N_803,N_775);
or U10995 (N_10995,N_8942,N_1948);
xor U10996 (N_10996,N_3650,N_8628);
or U10997 (N_10997,N_2726,N_2274);
nor U10998 (N_10998,N_5304,N_7983);
and U10999 (N_10999,N_4905,N_3690);
and U11000 (N_11000,N_995,N_7518);
or U11001 (N_11001,N_5174,N_2691);
and U11002 (N_11002,N_9966,N_7747);
nand U11003 (N_11003,N_2324,N_5455);
and U11004 (N_11004,N_2301,N_4015);
nand U11005 (N_11005,N_3530,N_4709);
xor U11006 (N_11006,N_2898,N_7562);
nor U11007 (N_11007,N_5355,N_9949);
nor U11008 (N_11008,N_4547,N_8321);
and U11009 (N_11009,N_1045,N_5796);
nor U11010 (N_11010,N_2894,N_5218);
and U11011 (N_11011,N_1597,N_4054);
and U11012 (N_11012,N_9777,N_1977);
or U11013 (N_11013,N_1593,N_5266);
and U11014 (N_11014,N_6759,N_1871);
nor U11015 (N_11015,N_6186,N_7101);
nand U11016 (N_11016,N_4576,N_1119);
xnor U11017 (N_11017,N_6159,N_6447);
or U11018 (N_11018,N_3260,N_6015);
and U11019 (N_11019,N_4069,N_3894);
nor U11020 (N_11020,N_9421,N_2801);
xor U11021 (N_11021,N_1169,N_598);
nor U11022 (N_11022,N_3400,N_4775);
xor U11023 (N_11023,N_6715,N_8433);
nor U11024 (N_11024,N_6589,N_3732);
nand U11025 (N_11025,N_4231,N_8509);
xor U11026 (N_11026,N_3933,N_2287);
nor U11027 (N_11027,N_5465,N_4488);
and U11028 (N_11028,N_979,N_4953);
xor U11029 (N_11029,N_8688,N_7978);
and U11030 (N_11030,N_2245,N_5450);
xor U11031 (N_11031,N_7729,N_7646);
and U11032 (N_11032,N_644,N_6227);
nand U11033 (N_11033,N_4112,N_8142);
nor U11034 (N_11034,N_7788,N_8271);
or U11035 (N_11035,N_1306,N_786);
nor U11036 (N_11036,N_1665,N_7769);
nand U11037 (N_11037,N_4864,N_1248);
or U11038 (N_11038,N_5346,N_2970);
or U11039 (N_11039,N_1223,N_9939);
xor U11040 (N_11040,N_2477,N_8432);
nand U11041 (N_11041,N_7365,N_5458);
and U11042 (N_11042,N_6646,N_5350);
and U11043 (N_11043,N_5954,N_1514);
or U11044 (N_11044,N_625,N_8983);
nor U11045 (N_11045,N_3401,N_8423);
and U11046 (N_11046,N_3038,N_9741);
nand U11047 (N_11047,N_1863,N_115);
and U11048 (N_11048,N_5710,N_8421);
nand U11049 (N_11049,N_4792,N_6926);
xor U11050 (N_11050,N_9622,N_1794);
and U11051 (N_11051,N_8590,N_347);
nand U11052 (N_11052,N_7615,N_4620);
and U11053 (N_11053,N_357,N_846);
xnor U11054 (N_11054,N_9462,N_807);
and U11055 (N_11055,N_2438,N_6335);
nand U11056 (N_11056,N_8082,N_3172);
nor U11057 (N_11057,N_899,N_3276);
xnor U11058 (N_11058,N_4835,N_2332);
nand U11059 (N_11059,N_9513,N_3736);
and U11060 (N_11060,N_8757,N_5741);
or U11061 (N_11061,N_1659,N_6301);
nand U11062 (N_11062,N_8042,N_584);
nor U11063 (N_11063,N_968,N_1501);
xnor U11064 (N_11064,N_2016,N_5649);
xnor U11065 (N_11065,N_3597,N_6351);
nand U11066 (N_11066,N_5874,N_8206);
nor U11067 (N_11067,N_2453,N_2957);
nor U11068 (N_11068,N_2192,N_986);
and U11069 (N_11069,N_6594,N_7537);
nand U11070 (N_11070,N_3785,N_4094);
nor U11071 (N_11071,N_976,N_9828);
nand U11072 (N_11072,N_6722,N_6009);
or U11073 (N_11073,N_7545,N_2494);
nor U11074 (N_11074,N_7088,N_3565);
nand U11075 (N_11075,N_9050,N_4158);
nand U11076 (N_11076,N_5347,N_7688);
nand U11077 (N_11077,N_1518,N_8313);
nand U11078 (N_11078,N_4694,N_7887);
nand U11079 (N_11079,N_4961,N_7062);
nand U11080 (N_11080,N_6681,N_2457);
nand U11081 (N_11081,N_4017,N_7817);
nor U11082 (N_11082,N_9017,N_8725);
nor U11083 (N_11083,N_7603,N_107);
nand U11084 (N_11084,N_4242,N_1017);
nor U11085 (N_11085,N_5141,N_1018);
or U11086 (N_11086,N_1897,N_8877);
or U11087 (N_11087,N_4329,N_7946);
nor U11088 (N_11088,N_4453,N_708);
nand U11089 (N_11089,N_1814,N_2658);
or U11090 (N_11090,N_7320,N_8204);
nand U11091 (N_11091,N_7197,N_6912);
nor U11092 (N_11092,N_4428,N_8346);
or U11093 (N_11093,N_7767,N_2980);
nor U11094 (N_11094,N_4998,N_663);
nand U11095 (N_11095,N_6869,N_5543);
nand U11096 (N_11096,N_9150,N_537);
nor U11097 (N_11097,N_3636,N_3544);
and U11098 (N_11098,N_2884,N_6459);
and U11099 (N_11099,N_6274,N_481);
nand U11100 (N_11100,N_1324,N_9442);
xnor U11101 (N_11101,N_560,N_2282);
and U11102 (N_11102,N_1146,N_6312);
nor U11103 (N_11103,N_5211,N_9156);
or U11104 (N_11104,N_3904,N_6799);
nand U11105 (N_11105,N_7734,N_6535);
nor U11106 (N_11106,N_2249,N_5935);
nand U11107 (N_11107,N_7897,N_8079);
nand U11108 (N_11108,N_8607,N_1867);
nor U11109 (N_11109,N_309,N_2839);
or U11110 (N_11110,N_3111,N_621);
nand U11111 (N_11111,N_8162,N_539);
or U11112 (N_11112,N_3368,N_9331);
and U11113 (N_11113,N_3236,N_2406);
or U11114 (N_11114,N_2766,N_8060);
or U11115 (N_11115,N_4635,N_5988);
and U11116 (N_11116,N_3309,N_1225);
nand U11117 (N_11117,N_8777,N_7820);
or U11118 (N_11118,N_53,N_6119);
and U11119 (N_11119,N_2430,N_2223);
or U11120 (N_11120,N_2719,N_9337);
nand U11121 (N_11121,N_9582,N_8704);
nand U11122 (N_11122,N_5990,N_5576);
nor U11123 (N_11123,N_6834,N_5253);
and U11124 (N_11124,N_9664,N_7933);
or U11125 (N_11125,N_7235,N_5821);
nor U11126 (N_11126,N_2617,N_742);
or U11127 (N_11127,N_4188,N_8654);
and U11128 (N_11128,N_6544,N_1222);
and U11129 (N_11129,N_3308,N_1924);
nand U11130 (N_11130,N_9106,N_6576);
xnor U11131 (N_11131,N_5687,N_9086);
nand U11132 (N_11132,N_3665,N_1329);
and U11133 (N_11133,N_5065,N_4413);
or U11134 (N_11134,N_9648,N_7833);
nor U11135 (N_11135,N_7302,N_1483);
xnor U11136 (N_11136,N_2977,N_3756);
xor U11137 (N_11137,N_1469,N_3516);
xnor U11138 (N_11138,N_2912,N_92);
nor U11139 (N_11139,N_9631,N_4634);
nand U11140 (N_11140,N_944,N_3596);
nand U11141 (N_11141,N_8071,N_546);
and U11142 (N_11142,N_2383,N_7496);
nor U11143 (N_11143,N_5829,N_7869);
and U11144 (N_11144,N_7019,N_3173);
nand U11145 (N_11145,N_2075,N_3497);
or U11146 (N_11146,N_6388,N_3572);
nand U11147 (N_11147,N_3415,N_2068);
and U11148 (N_11148,N_3931,N_1520);
nand U11149 (N_11149,N_8340,N_6107);
nand U11150 (N_11150,N_9126,N_478);
nor U11151 (N_11151,N_8858,N_77);
or U11152 (N_11152,N_3552,N_7720);
and U11153 (N_11153,N_5924,N_3341);
or U11154 (N_11154,N_1869,N_1020);
and U11155 (N_11155,N_2689,N_1369);
or U11156 (N_11156,N_2713,N_1910);
nand U11157 (N_11157,N_1149,N_728);
xnor U11158 (N_11158,N_8646,N_7312);
or U11159 (N_11159,N_7386,N_5241);
and U11160 (N_11160,N_9922,N_2169);
and U11161 (N_11161,N_8048,N_5803);
nand U11162 (N_11162,N_1389,N_9059);
and U11163 (N_11163,N_3192,N_7987);
nand U11164 (N_11164,N_1362,N_1686);
nand U11165 (N_11165,N_2646,N_5707);
or U11166 (N_11166,N_1498,N_9559);
nor U11167 (N_11167,N_4630,N_7832);
or U11168 (N_11168,N_570,N_2956);
or U11169 (N_11169,N_5960,N_1132);
nand U11170 (N_11170,N_1332,N_7748);
and U11171 (N_11171,N_3962,N_4923);
nor U11172 (N_11172,N_3675,N_3275);
or U11173 (N_11173,N_1342,N_918);
and U11174 (N_11174,N_287,N_6878);
or U11175 (N_11175,N_3558,N_1962);
or U11176 (N_11176,N_5526,N_7120);
nor U11177 (N_11177,N_5762,N_2562);
or U11178 (N_11178,N_2160,N_9967);
xor U11179 (N_11179,N_4892,N_7770);
nand U11180 (N_11180,N_164,N_2019);
nor U11181 (N_11181,N_9191,N_160);
and U11182 (N_11182,N_9612,N_6346);
nand U11183 (N_11183,N_3389,N_7679);
nor U11184 (N_11184,N_5657,N_4321);
nor U11185 (N_11185,N_9019,N_5694);
or U11186 (N_11186,N_7366,N_706);
or U11187 (N_11187,N_1533,N_2333);
nand U11188 (N_11188,N_6358,N_6600);
or U11189 (N_11189,N_5944,N_4464);
nand U11190 (N_11190,N_4121,N_7704);
and U11191 (N_11191,N_344,N_1026);
or U11192 (N_11192,N_8657,N_5717);
nor U11193 (N_11193,N_7066,N_4165);
xor U11194 (N_11194,N_4713,N_4968);
nand U11195 (N_11195,N_3922,N_3506);
or U11196 (N_11196,N_6944,N_881);
nor U11197 (N_11197,N_5605,N_6614);
nor U11198 (N_11198,N_9384,N_2044);
and U11199 (N_11199,N_1488,N_758);
or U11200 (N_11200,N_3981,N_3824);
nor U11201 (N_11201,N_3289,N_2289);
nand U11202 (N_11202,N_7460,N_6450);
nor U11203 (N_11203,N_7879,N_2313);
nand U11204 (N_11204,N_1524,N_2251);
xor U11205 (N_11205,N_9918,N_3416);
or U11206 (N_11206,N_6150,N_9936);
nand U11207 (N_11207,N_398,N_2510);
xor U11208 (N_11208,N_5506,N_4830);
nand U11209 (N_11209,N_7199,N_1748);
nor U11210 (N_11210,N_7428,N_1215);
and U11211 (N_11211,N_909,N_4025);
xnor U11212 (N_11212,N_3529,N_9339);
or U11213 (N_11213,N_5175,N_2166);
and U11214 (N_11214,N_2888,N_6885);
and U11215 (N_11215,N_8114,N_6893);
and U11216 (N_11216,N_5619,N_3699);
or U11217 (N_11217,N_6278,N_4898);
or U11218 (N_11218,N_5782,N_7971);
nand U11219 (N_11219,N_9885,N_2684);
nand U11220 (N_11220,N_9661,N_2371);
nor U11221 (N_11221,N_5108,N_3440);
or U11222 (N_11222,N_165,N_121);
or U11223 (N_11223,N_7777,N_6801);
and U11224 (N_11224,N_818,N_211);
nand U11225 (N_11225,N_3312,N_1404);
xnor U11226 (N_11226,N_4222,N_2745);
nand U11227 (N_11227,N_1127,N_2002);
or U11228 (N_11228,N_9043,N_6636);
nand U11229 (N_11229,N_5592,N_3579);
or U11230 (N_11230,N_7508,N_3013);
nor U11231 (N_11231,N_9025,N_3634);
nand U11232 (N_11232,N_2349,N_8748);
nand U11233 (N_11233,N_2739,N_8912);
nor U11234 (N_11234,N_6280,N_980);
or U11235 (N_11235,N_6703,N_7528);
xnor U11236 (N_11236,N_9849,N_5229);
nand U11237 (N_11237,N_7768,N_6495);
nand U11238 (N_11238,N_2468,N_5467);
nor U11239 (N_11239,N_5833,N_8259);
nor U11240 (N_11240,N_4873,N_1194);
nor U11241 (N_11241,N_9100,N_5705);
nor U11242 (N_11242,N_3128,N_7142);
xor U11243 (N_11243,N_6336,N_8663);
and U11244 (N_11244,N_8837,N_9539);
or U11245 (N_11245,N_8102,N_4888);
or U11246 (N_11246,N_2780,N_6443);
xor U11247 (N_11247,N_5446,N_2253);
or U11248 (N_11248,N_5612,N_7426);
xnor U11249 (N_11249,N_9676,N_2931);
and U11250 (N_11250,N_7439,N_9154);
or U11251 (N_11251,N_4172,N_5243);
and U11252 (N_11252,N_9471,N_835);
or U11253 (N_11253,N_9899,N_9377);
or U11254 (N_11254,N_9614,N_6823);
xnor U11255 (N_11255,N_2741,N_243);
and U11256 (N_11256,N_8723,N_9892);
and U11257 (N_11257,N_300,N_8536);
and U11258 (N_11258,N_7404,N_8010);
nor U11259 (N_11259,N_6065,N_280);
and U11260 (N_11260,N_4115,N_9993);
or U11261 (N_11261,N_2824,N_7868);
and U11262 (N_11262,N_2735,N_2734);
and U11263 (N_11263,N_459,N_4452);
nand U11264 (N_11264,N_9030,N_4186);
nand U11265 (N_11265,N_2401,N_8238);
nand U11266 (N_11266,N_6666,N_5398);
nor U11267 (N_11267,N_9084,N_2094);
or U11268 (N_11268,N_2229,N_7698);
nand U11269 (N_11269,N_6952,N_4232);
nand U11270 (N_11270,N_9678,N_6914);
and U11271 (N_11271,N_7655,N_7230);
nor U11272 (N_11272,N_8103,N_9736);
and U11273 (N_11273,N_8198,N_5886);
nor U11274 (N_11274,N_4228,N_4726);
nor U11275 (N_11275,N_3290,N_9027);
nand U11276 (N_11276,N_3445,N_4954);
xor U11277 (N_11277,N_1259,N_9923);
nand U11278 (N_11278,N_4899,N_8110);
nand U11279 (N_11279,N_4286,N_180);
xor U11280 (N_11280,N_8941,N_3204);
xor U11281 (N_11281,N_9780,N_894);
nor U11282 (N_11282,N_3528,N_3129);
xnor U11283 (N_11283,N_3833,N_502);
or U11284 (N_11284,N_4262,N_526);
and U11285 (N_11285,N_5472,N_8668);
and U11286 (N_11286,N_3157,N_6130);
nor U11287 (N_11287,N_762,N_6880);
nor U11288 (N_11288,N_6484,N_5248);
xnor U11289 (N_11289,N_737,N_7995);
or U11290 (N_11290,N_693,N_6217);
and U11291 (N_11291,N_1461,N_1097);
xor U11292 (N_11292,N_210,N_503);
nand U11293 (N_11293,N_69,N_9037);
xnor U11294 (N_11294,N_68,N_5607);
and U11295 (N_11295,N_4313,N_6747);
nand U11296 (N_11296,N_5978,N_229);
or U11297 (N_11297,N_5284,N_5644);
and U11298 (N_11298,N_9839,N_1548);
nand U11299 (N_11299,N_6478,N_6971);
or U11300 (N_11300,N_7114,N_295);
nor U11301 (N_11301,N_1441,N_3576);
or U11302 (N_11302,N_8160,N_7478);
or U11303 (N_11303,N_222,N_6909);
or U11304 (N_11304,N_9048,N_5805);
nor U11305 (N_11305,N_4280,N_7039);
xnor U11306 (N_11306,N_2747,N_4569);
nor U11307 (N_11307,N_4969,N_8913);
xnor U11308 (N_11308,N_9296,N_6753);
and U11309 (N_11309,N_3519,N_8268);
and U11310 (N_11310,N_5225,N_2123);
and U11311 (N_11311,N_8990,N_2162);
nand U11312 (N_11312,N_2408,N_383);
nand U11313 (N_11313,N_8096,N_9078);
or U11314 (N_11314,N_7407,N_9529);
nor U11315 (N_11315,N_5330,N_5430);
xnor U11316 (N_11316,N_1426,N_487);
nor U11317 (N_11317,N_6827,N_8288);
nor U11318 (N_11318,N_9345,N_9195);
nand U11319 (N_11319,N_3573,N_6637);
nand U11320 (N_11320,N_3140,N_379);
nand U11321 (N_11321,N_3609,N_7079);
nor U11322 (N_11322,N_4611,N_3687);
nand U11323 (N_11323,N_8930,N_3131);
or U11324 (N_11324,N_1134,N_4995);
nor U11325 (N_11325,N_2078,N_324);
or U11326 (N_11326,N_6485,N_3408);
xor U11327 (N_11327,N_9076,N_8391);
or U11328 (N_11328,N_4367,N_9306);
xnor U11329 (N_11329,N_2091,N_9601);
nor U11330 (N_11330,N_3858,N_5606);
and U11331 (N_11331,N_4171,N_8353);
xnor U11332 (N_11332,N_6172,N_1112);
nand U11333 (N_11333,N_4626,N_2627);
nor U11334 (N_11334,N_2727,N_8567);
xnor U11335 (N_11335,N_7472,N_4731);
nor U11336 (N_11336,N_9089,N_1099);
nor U11337 (N_11337,N_5420,N_6907);
nand U11338 (N_11338,N_3251,N_3975);
and U11339 (N_11339,N_7628,N_3017);
or U11340 (N_11340,N_7965,N_5317);
nand U11341 (N_11341,N_4943,N_5165);
xor U11342 (N_11342,N_4391,N_37);
or U11343 (N_11343,N_9799,N_6617);
nor U11344 (N_11344,N_2939,N_8718);
nand U11345 (N_11345,N_6140,N_6111);
or U11346 (N_11346,N_370,N_3940);
and U11347 (N_11347,N_1152,N_8991);
nor U11348 (N_11348,N_9558,N_5353);
xnor U11349 (N_11349,N_5372,N_2535);
or U11350 (N_11350,N_4500,N_3431);
xnor U11351 (N_11351,N_3799,N_6292);
nor U11352 (N_11352,N_886,N_6713);
and U11353 (N_11353,N_6005,N_6220);
and U11354 (N_11354,N_7982,N_6778);
or U11355 (N_11355,N_6505,N_1656);
or U11356 (N_11356,N_4052,N_5588);
xnor U11357 (N_11357,N_2634,N_5478);
or U11358 (N_11358,N_8097,N_7091);
xnor U11359 (N_11359,N_6567,N_8105);
and U11360 (N_11360,N_7158,N_8349);
nand U11361 (N_11361,N_7571,N_3575);
nor U11362 (N_11362,N_5026,N_7554);
nand U11363 (N_11363,N_7219,N_8381);
nor U11364 (N_11364,N_199,N_6222);
and U11365 (N_11365,N_6531,N_8705);
and U11366 (N_11366,N_220,N_1508);
or U11367 (N_11367,N_4163,N_8159);
nand U11368 (N_11368,N_1767,N_30);
or U11369 (N_11369,N_3313,N_850);
nor U11370 (N_11370,N_2153,N_4730);
nand U11371 (N_11371,N_6075,N_2874);
nand U11372 (N_11372,N_4858,N_1760);
nand U11373 (N_11373,N_6516,N_3623);
xnor U11374 (N_11374,N_208,N_6674);
or U11375 (N_11375,N_6421,N_217);
or U11376 (N_11376,N_5845,N_8892);
nor U11377 (N_11377,N_5665,N_7574);
and U11378 (N_11378,N_4603,N_9470);
nand U11379 (N_11379,N_6984,N_1290);
nand U11380 (N_11380,N_7076,N_7961);
xor U11381 (N_11381,N_5315,N_6342);
nor U11382 (N_11382,N_9042,N_182);
and U11383 (N_11383,N_1722,N_5172);
nor U11384 (N_11384,N_888,N_8826);
nor U11385 (N_11385,N_7610,N_6658);
nand U11386 (N_11386,N_5201,N_9798);
nor U11387 (N_11387,N_1840,N_8018);
xor U11388 (N_11388,N_919,N_7650);
nand U11389 (N_11389,N_1590,N_6768);
nand U11390 (N_11390,N_1334,N_11);
or U11391 (N_11391,N_7362,N_6281);
and U11392 (N_11392,N_7523,N_6298);
nor U11393 (N_11393,N_9716,N_334);
nor U11394 (N_11394,N_614,N_7660);
nand U11395 (N_11395,N_5655,N_650);
nor U11396 (N_11396,N_2504,N_4361);
xor U11397 (N_11397,N_768,N_4177);
or U11398 (N_11398,N_7714,N_6001);
and U11399 (N_11399,N_9516,N_5603);
nand U11400 (N_11400,N_2190,N_7433);
nor U11401 (N_11401,N_3122,N_86);
and U11402 (N_11402,N_4476,N_9950);
nor U11403 (N_11403,N_7614,N_9568);
xnor U11404 (N_11404,N_7021,N_2638);
or U11405 (N_11405,N_1692,N_8523);
xnor U11406 (N_11406,N_5035,N_4141);
nor U11407 (N_11407,N_3411,N_3025);
and U11408 (N_11408,N_7802,N_332);
or U11409 (N_11409,N_5042,N_9984);
nand U11410 (N_11410,N_403,N_855);
xor U11411 (N_11411,N_610,N_4633);
or U11412 (N_11412,N_7883,N_8914);
nand U11413 (N_11413,N_1667,N_1609);
and U11414 (N_11414,N_8641,N_8377);
nor U11415 (N_11415,N_5157,N_3439);
nor U11416 (N_11416,N_4561,N_2328);
and U11417 (N_11417,N_40,N_1581);
or U11418 (N_11418,N_1925,N_8436);
or U11419 (N_11419,N_5111,N_1644);
nor U11420 (N_11420,N_3379,N_9382);
nand U11421 (N_11421,N_9279,N_1571);
or U11422 (N_11422,N_3583,N_7921);
nand U11423 (N_11423,N_1080,N_9253);
and U11424 (N_11424,N_2949,N_5608);
nor U11425 (N_11425,N_8658,N_9841);
nor U11426 (N_11426,N_2804,N_7618);
or U11427 (N_11427,N_7470,N_8677);
nor U11428 (N_11428,N_9605,N_549);
nor U11429 (N_11429,N_8087,N_9915);
nor U11430 (N_11430,N_4439,N_4987);
xnor U11431 (N_11431,N_8999,N_2614);
nand U11432 (N_11432,N_7456,N_3328);
and U11433 (N_11433,N_5941,N_9913);
xor U11434 (N_11434,N_839,N_4032);
or U11435 (N_11435,N_8020,N_4765);
or U11436 (N_11436,N_1689,N_9047);
nor U11437 (N_11437,N_3244,N_9142);
xnor U11438 (N_11438,N_2317,N_7675);
or U11439 (N_11439,N_6192,N_1028);
xor U11440 (N_11440,N_7160,N_5090);
nor U11441 (N_11441,N_3112,N_1515);
or U11442 (N_11442,N_2959,N_1935);
nand U11443 (N_11443,N_953,N_814);
nand U11444 (N_11444,N_3549,N_8708);
or U11445 (N_11445,N_6451,N_690);
and U11446 (N_11446,N_9878,N_6056);
nor U11447 (N_11447,N_7422,N_8348);
xnor U11448 (N_11448,N_218,N_6452);
and U11449 (N_11449,N_7200,N_6117);
or U11450 (N_11450,N_8529,N_1352);
nand U11451 (N_11451,N_7007,N_9535);
and U11452 (N_11452,N_9440,N_4984);
nor U11453 (N_11453,N_2563,N_8331);
nand U11454 (N_11454,N_7150,N_5868);
or U11455 (N_11455,N_2150,N_9668);
and U11456 (N_11456,N_3391,N_2803);
nor U11457 (N_11457,N_1168,N_6087);
nor U11458 (N_11458,N_3825,N_3118);
or U11459 (N_11459,N_3214,N_9247);
nand U11460 (N_11460,N_9598,N_9687);
nand U11461 (N_11461,N_5142,N_3627);
or U11462 (N_11462,N_1809,N_1442);
nor U11463 (N_11463,N_2476,N_9914);
or U11464 (N_11464,N_7831,N_2685);
and U11465 (N_11465,N_1065,N_3807);
and U11466 (N_11466,N_9650,N_29);
xor U11467 (N_11467,N_3996,N_9180);
nor U11468 (N_11468,N_747,N_8387);
nand U11469 (N_11469,N_1114,N_9653);
and U11470 (N_11470,N_889,N_7075);
nor U11471 (N_11471,N_3590,N_7569);
nand U11472 (N_11472,N_8066,N_6179);
nor U11473 (N_11473,N_9128,N_7327);
nand U11474 (N_11474,N_2573,N_2145);
or U11475 (N_11475,N_9814,N_1774);
nor U11476 (N_11476,N_1746,N_2518);
nor U11477 (N_11477,N_9139,N_2009);
xnor U11478 (N_11478,N_13,N_185);
or U11479 (N_11479,N_1595,N_5502);
and U11480 (N_11480,N_1749,N_2591);
nor U11481 (N_11481,N_1632,N_3525);
nand U11482 (N_11482,N_7121,N_5823);
nor U11483 (N_11483,N_8863,N_3304);
and U11484 (N_11484,N_1641,N_872);
or U11485 (N_11485,N_3396,N_9134);
or U11486 (N_11486,N_1282,N_9323);
or U11487 (N_11487,N_6190,N_8388);
and U11488 (N_11488,N_3700,N_1141);
nor U11489 (N_11489,N_6928,N_5240);
or U11490 (N_11490,N_3046,N_1525);
nand U11491 (N_11491,N_8182,N_1036);
or U11492 (N_11492,N_6486,N_6108);
or U11493 (N_11493,N_6552,N_8008);
nor U11494 (N_11494,N_5764,N_5397);
or U11495 (N_11495,N_5431,N_6776);
nand U11496 (N_11496,N_5018,N_1607);
nand U11497 (N_11497,N_3517,N_4976);
nand U11498 (N_11498,N_3344,N_4653);
nor U11499 (N_11499,N_7925,N_4693);
and U11500 (N_11500,N_9958,N_8416);
xor U11501 (N_11501,N_4418,N_1411);
nand U11502 (N_11502,N_630,N_5477);
or U11503 (N_11503,N_1077,N_285);
nor U11504 (N_11504,N_278,N_99);
or U11505 (N_11505,N_4350,N_3133);
xor U11506 (N_11506,N_458,N_4800);
nor U11507 (N_11507,N_4203,N_5969);
or U11508 (N_11508,N_6743,N_7005);
nor U11509 (N_11509,N_46,N_9721);
nor U11510 (N_11510,N_2632,N_1489);
or U11511 (N_11511,N_7175,N_9751);
nand U11512 (N_11512,N_5293,N_9820);
or U11513 (N_11513,N_2306,N_132);
nor U11514 (N_11514,N_5734,N_853);
and U11515 (N_11515,N_5075,N_582);
or U11516 (N_11516,N_9239,N_6536);
xor U11517 (N_11517,N_171,N_2793);
nand U11518 (N_11518,N_6481,N_2265);
and U11519 (N_11519,N_8278,N_534);
or U11520 (N_11520,N_5264,N_187);
nand U11521 (N_11521,N_4066,N_1870);
or U11522 (N_11522,N_5863,N_4062);
nand U11523 (N_11523,N_4125,N_308);
nor U11524 (N_11524,N_9880,N_5044);
nor U11525 (N_11525,N_540,N_5013);
and U11526 (N_11526,N_3003,N_7481);
nor U11527 (N_11527,N_4970,N_6373);
xnor U11528 (N_11528,N_9376,N_6103);
nand U11529 (N_11529,N_362,N_494);
and U11530 (N_11530,N_1660,N_7129);
xnor U11531 (N_11531,N_9399,N_6382);
or U11532 (N_11532,N_162,N_7955);
nor U11533 (N_11533,N_100,N_7836);
nor U11534 (N_11534,N_1056,N_9053);
or U11535 (N_11535,N_3694,N_4097);
and U11536 (N_11536,N_1246,N_5709);
nor U11537 (N_11537,N_6548,N_6020);
or U11538 (N_11538,N_2246,N_8505);
or U11539 (N_11539,N_6811,N_5269);
or U11540 (N_11540,N_4675,N_4660);
nand U11541 (N_11541,N_8707,N_6296);
and U11542 (N_11542,N_6940,N_9249);
xnor U11543 (N_11543,N_7454,N_4264);
nor U11544 (N_11544,N_3127,N_2964);
nand U11545 (N_11545,N_7248,N_7761);
xor U11546 (N_11546,N_4193,N_7333);
or U11547 (N_11547,N_1939,N_2167);
nand U11548 (N_11548,N_1675,N_1373);
and U11549 (N_11549,N_4499,N_3696);
or U11550 (N_11550,N_2121,N_202);
nor U11551 (N_11551,N_6184,N_6102);
xnor U11552 (N_11552,N_4042,N_4471);
nor U11553 (N_11553,N_8825,N_2036);
and U11554 (N_11554,N_3523,N_3397);
or U11555 (N_11555,N_1318,N_131);
or U11556 (N_11556,N_3161,N_6476);
nand U11557 (N_11557,N_3641,N_6399);
or U11558 (N_11558,N_8434,N_2782);
and U11559 (N_11559,N_5677,N_7859);
and U11560 (N_11560,N_134,N_4825);
nor U11561 (N_11561,N_7466,N_4483);
and U11562 (N_11562,N_4288,N_377);
and U11563 (N_11563,N_8973,N_8447);
or U11564 (N_11564,N_3613,N_9113);
or U11565 (N_11565,N_1717,N_6251);
and U11566 (N_11566,N_8158,N_155);
and U11567 (N_11567,N_3602,N_499);
nand U11568 (N_11568,N_7409,N_7953);
nand U11569 (N_11569,N_2915,N_3821);
nand U11570 (N_11570,N_5663,N_2381);
or U11571 (N_11571,N_4245,N_4405);
nand U11572 (N_11572,N_1547,N_2690);
xnor U11573 (N_11573,N_8189,N_2385);
nand U11574 (N_11574,N_5991,N_5703);
or U11575 (N_11575,N_183,N_1753);
and U11576 (N_11576,N_3950,N_7271);
nor U11577 (N_11577,N_7099,N_1828);
or U11578 (N_11578,N_1010,N_7477);
nor U11579 (N_11579,N_2564,N_8807);
and U11580 (N_11580,N_4098,N_8207);
nand U11581 (N_11581,N_4013,N_4400);
nor U11582 (N_11582,N_5071,N_5219);
nor U11583 (N_11583,N_1347,N_9206);
and U11584 (N_11584,N_8122,N_6262);
and U11585 (N_11585,N_9065,N_3500);
nand U11586 (N_11586,N_3299,N_6692);
nor U11587 (N_11587,N_496,N_6066);
nand U11588 (N_11588,N_9638,N_5437);
xnor U11589 (N_11589,N_7368,N_2260);
or U11590 (N_11590,N_9522,N_8674);
xor U11591 (N_11591,N_1420,N_3220);
nand U11592 (N_11592,N_9426,N_4774);
and U11593 (N_11593,N_1494,N_2199);
or U11594 (N_11594,N_3600,N_6679);
xnor U11595 (N_11595,N_1218,N_4323);
and U11596 (N_11596,N_7890,N_8302);
nor U11597 (N_11597,N_5492,N_8299);
nor U11598 (N_11598,N_6309,N_9378);
nor U11599 (N_11599,N_1179,N_1564);
nor U11600 (N_11600,N_2270,N_4880);
nand U11601 (N_11601,N_6560,N_8441);
xnor U11602 (N_11602,N_453,N_2445);
xor U11603 (N_11603,N_7566,N_2035);
nor U11604 (N_11604,N_9766,N_4769);
nor U11605 (N_11605,N_3490,N_7968);
nor U11606 (N_11606,N_9995,N_9784);
xor U11607 (N_11607,N_3222,N_3333);
nand U11608 (N_11608,N_7555,N_1359);
and U11609 (N_11609,N_649,N_580);
xor U11610 (N_11610,N_225,N_5146);
xnor U11611 (N_11611,N_9208,N_7784);
nor U11612 (N_11612,N_2846,N_6270);
or U11613 (N_11613,N_9136,N_3874);
or U11614 (N_11614,N_2237,N_6987);
nor U11615 (N_11615,N_2045,N_7755);
and U11616 (N_11616,N_7167,N_884);
or U11617 (N_11617,N_6904,N_2737);
or U11618 (N_11618,N_9289,N_8452);
nor U11619 (N_11619,N_1658,N_455);
and U11620 (N_11620,N_5343,N_6092);
or U11621 (N_11621,N_8052,N_551);
or U11622 (N_11622,N_655,N_1432);
nor U11623 (N_11623,N_1424,N_4702);
nand U11624 (N_11624,N_1463,N_6861);
nand U11625 (N_11625,N_2663,N_474);
or U11626 (N_11626,N_8154,N_8534);
and U11627 (N_11627,N_6394,N_5601);
nor U11628 (N_11628,N_9410,N_9144);
xor U11629 (N_11629,N_5581,N_8675);
and U11630 (N_11630,N_1934,N_5609);
xor U11631 (N_11631,N_806,N_95);
nor U11632 (N_11632,N_6727,N_0);
and U11633 (N_11633,N_9495,N_3960);
and U11634 (N_11634,N_4852,N_9530);
and U11635 (N_11635,N_1326,N_4379);
nor U11636 (N_11636,N_6915,N_5445);
and U11637 (N_11637,N_2297,N_6886);
nor U11638 (N_11638,N_8386,N_8064);
or U11639 (N_11639,N_339,N_7813);
nor U11640 (N_11640,N_3182,N_3987);
and U11641 (N_11641,N_3399,N_3589);
xor U11642 (N_11642,N_6864,N_1181);
and U11643 (N_11643,N_9409,N_5512);
or U11644 (N_11644,N_9182,N_1073);
nand U11645 (N_11645,N_6611,N_8);
nand U11646 (N_11646,N_128,N_371);
nor U11647 (N_11647,N_1142,N_3701);
nor U11648 (N_11648,N_8782,N_2850);
nor U11649 (N_11649,N_721,N_416);
nand U11650 (N_11650,N_9417,N_6200);
or U11651 (N_11651,N_6935,N_1782);
xor U11652 (N_11652,N_554,N_3306);
and U11653 (N_11653,N_9010,N_5188);
nand U11654 (N_11654,N_2756,N_9961);
nand U11655 (N_11655,N_4185,N_4906);
and U11656 (N_11656,N_8543,N_9049);
nor U11657 (N_11657,N_5780,N_9222);
nor U11658 (N_11658,N_9511,N_1113);
and U11659 (N_11659,N_2460,N_5312);
nand U11660 (N_11660,N_4749,N_9738);
or U11661 (N_11661,N_6575,N_8305);
nor U11662 (N_11662,N_1642,N_759);
nand U11663 (N_11663,N_1540,N_2221);
and U11664 (N_11664,N_9765,N_4524);
or U11665 (N_11665,N_5440,N_4591);
nand U11666 (N_11666,N_2188,N_8450);
nor U11667 (N_11667,N_9006,N_7361);
and U11668 (N_11668,N_983,N_578);
and U11669 (N_11669,N_8047,N_9691);
nor U11670 (N_11670,N_6168,N_3513);
or U11671 (N_11671,N_8843,N_4587);
and U11672 (N_11672,N_6938,N_1339);
and U11673 (N_11673,N_4336,N_9480);
and U11674 (N_11674,N_2452,N_2300);
and U11675 (N_11675,N_266,N_1950);
or U11676 (N_11676,N_9497,N_8595);
nand U11677 (N_11677,N_4006,N_9231);
or U11678 (N_11678,N_2647,N_7457);
xor U11679 (N_11679,N_6784,N_9671);
and U11680 (N_11680,N_5195,N_8482);
and U11681 (N_11681,N_588,N_5515);
nor U11682 (N_11682,N_1592,N_6135);
and U11683 (N_11683,N_9694,N_4460);
nor U11684 (N_11684,N_3049,N_9700);
xor U11685 (N_11685,N_9277,N_4664);
or U11686 (N_11686,N_4440,N_1283);
nand U11687 (N_11687,N_320,N_80);
nor U11688 (N_11688,N_8376,N_2413);
xnor U11689 (N_11689,N_1723,N_7279);
nand U11690 (N_11690,N_868,N_3137);
nand U11691 (N_11691,N_6161,N_2811);
nand U11692 (N_11692,N_6824,N_3511);
nand U11693 (N_11693,N_4123,N_3081);
or U11694 (N_11694,N_2495,N_2226);
or U11695 (N_11695,N_4167,N_7606);
and U11696 (N_11696,N_7237,N_772);
nand U11697 (N_11697,N_788,N_3357);
nor U11698 (N_11698,N_2496,N_6375);
nor U11699 (N_11699,N_7068,N_1921);
nor U11700 (N_11700,N_2596,N_3670);
nor U11701 (N_11701,N_9117,N_3188);
and U11702 (N_11702,N_5375,N_1245);
and U11703 (N_11703,N_5584,N_5340);
nor U11704 (N_11704,N_8303,N_5259);
nor U11705 (N_11705,N_6219,N_1647);
and U11706 (N_11706,N_3307,N_200);
and U11707 (N_11707,N_5473,N_7735);
or U11708 (N_11708,N_8884,N_8090);
and U11709 (N_11709,N_8599,N_8936);
nor U11710 (N_11710,N_3336,N_569);
nor U11711 (N_11711,N_533,N_6441);
or U11712 (N_11712,N_9833,N_4758);
or U11713 (N_11713,N_2018,N_3225);
or U11714 (N_11714,N_422,N_3348);
nand U11715 (N_11715,N_9575,N_667);
or U11716 (N_11716,N_2509,N_9391);
nor U11717 (N_11717,N_440,N_3768);
and U11718 (N_11718,N_3574,N_3338);
nand U11719 (N_11719,N_1391,N_4285);
and U11720 (N_11720,N_977,N_6630);
and U11721 (N_11721,N_6098,N_8961);
nand U11722 (N_11722,N_5480,N_5371);
nor U11723 (N_11723,N_3740,N_2209);
nand U11724 (N_11724,N_3052,N_1128);
nor U11725 (N_11725,N_407,N_9455);
or U11726 (N_11726,N_2700,N_9365);
and U11727 (N_11727,N_9804,N_1577);
or U11728 (N_11728,N_2141,N_5560);
and U11729 (N_11729,N_7585,N_4639);
nor U11730 (N_11730,N_9166,N_684);
or U11731 (N_11731,N_1824,N_6027);
xor U11732 (N_11732,N_4301,N_3385);
or U11733 (N_11733,N_9876,N_2680);
and U11734 (N_11734,N_1289,N_1016);
or U11735 (N_11735,N_7193,N_6413);
nand U11736 (N_11736,N_7923,N_6354);
nor U11737 (N_11737,N_1589,N_916);
or U11738 (N_11738,N_130,N_7531);
nor U11739 (N_11739,N_2776,N_3349);
or U11740 (N_11740,N_3082,N_6310);
xnor U11741 (N_11741,N_1211,N_9118);
nand U11742 (N_11742,N_1143,N_6314);
nand U11743 (N_11743,N_6070,N_4706);
or U11744 (N_11744,N_967,N_3067);
nor U11745 (N_11745,N_736,N_156);
and U11746 (N_11746,N_2934,N_1171);
nor U11747 (N_11747,N_7003,N_1969);
and U11748 (N_11748,N_565,N_8631);
nor U11749 (N_11749,N_7926,N_3682);
nand U11750 (N_11750,N_5859,N_4847);
or U11751 (N_11751,N_9250,N_9806);
nor U11752 (N_11752,N_7213,N_1955);
nor U11753 (N_11753,N_6401,N_5410);
nor U11754 (N_11754,N_2729,N_6474);
nor U11755 (N_11755,N_695,N_8077);
or U11756 (N_11756,N_9838,N_7181);
xnor U11757 (N_11757,N_3345,N_6726);
or U11758 (N_11758,N_778,N_5939);
nor U11759 (N_11759,N_5872,N_5239);
or U11760 (N_11760,N_1275,N_2808);
xnor U11761 (N_11761,N_7414,N_2717);
nor U11762 (N_11762,N_856,N_148);
xnor U11763 (N_11763,N_2515,N_6613);
and U11764 (N_11764,N_4711,N_2038);
nand U11765 (N_11765,N_7637,N_5214);
nand U11766 (N_11766,N_2772,N_5995);
or U11767 (N_11767,N_9883,N_8481);
nand U11768 (N_11768,N_2901,N_8700);
or U11769 (N_11769,N_67,N_8712);
and U11770 (N_11770,N_1357,N_4078);
nor U11771 (N_11771,N_4064,N_4646);
and U11772 (N_11772,N_8403,N_1763);
and U11773 (N_11773,N_774,N_4166);
nor U11774 (N_11774,N_1539,N_4734);
or U11775 (N_11775,N_5009,N_6990);
and U11776 (N_11776,N_1164,N_545);
xnor U11777 (N_11777,N_9483,N_4384);
nand U11778 (N_11778,N_4824,N_8475);
and U11779 (N_11779,N_1361,N_4914);
xor U11780 (N_11780,N_8210,N_9075);
nor U11781 (N_11781,N_372,N_8304);
and U11782 (N_11782,N_5583,N_1041);
or U11783 (N_11783,N_2974,N_8174);
xor U11784 (N_11784,N_4941,N_9473);
nand U11785 (N_11785,N_959,N_1272);
or U11786 (N_11786,N_4885,N_9085);
xor U11787 (N_11787,N_3608,N_7435);
nor U11788 (N_11788,N_5629,N_9448);
nand U11789 (N_11789,N_3733,N_1941);
nor U11790 (N_11790,N_7290,N_9699);
and U11791 (N_11791,N_172,N_4244);
nand U11792 (N_11792,N_9955,N_2916);
nand U11793 (N_11793,N_653,N_5483);
nand U11794 (N_11794,N_1519,N_2184);
nor U11795 (N_11795,N_2648,N_2762);
and U11796 (N_11796,N_258,N_7394);
xnor U11797 (N_11797,N_7689,N_5791);
nor U11798 (N_11798,N_4759,N_7405);
and U11799 (N_11799,N_9805,N_4035);
and U11800 (N_11800,N_7280,N_8231);
or U11801 (N_11801,N_4315,N_7251);
nand U11802 (N_11802,N_4248,N_7020);
or U11803 (N_11803,N_145,N_5840);
nand U11804 (N_11804,N_2314,N_268);
or U11805 (N_11805,N_1587,N_2669);
nand U11806 (N_11806,N_6353,N_8493);
nand U11807 (N_11807,N_5533,N_7038);
nor U11808 (N_11808,N_2784,N_3423);
or U11809 (N_11809,N_2149,N_7174);
xor U11810 (N_11810,N_4387,N_3806);
nor U11811 (N_11811,N_4735,N_785);
nor U11812 (N_11812,N_9137,N_9536);
nor U11813 (N_11813,N_1313,N_2759);
nand U11814 (N_11814,N_8742,N_9649);
or U11815 (N_11815,N_7948,N_5499);
nand U11816 (N_11816,N_7680,N_5391);
xor U11817 (N_11817,N_9273,N_1022);
or U11818 (N_11818,N_8373,N_9561);
nand U11819 (N_11819,N_5020,N_6676);
nand U11820 (N_11820,N_7162,N_3176);
nand U11821 (N_11821,N_1039,N_4474);
nand U11822 (N_11822,N_6494,N_5828);
nand U11823 (N_11823,N_838,N_6740);
nand U11824 (N_11824,N_9461,N_3427);
nand U11825 (N_11825,N_7071,N_4663);
and U11826 (N_11826,N_6517,N_6177);
or U11827 (N_11827,N_9665,N_3616);
nand U11828 (N_11828,N_7956,N_1788);
nand U11829 (N_11829,N_5798,N_2907);
and U11830 (N_11830,N_1798,N_8410);
nand U11831 (N_11831,N_5767,N_5488);
or U11832 (N_11832,N_9360,N_4777);
xor U11833 (N_11833,N_638,N_9660);
or U11834 (N_11834,N_9441,N_6417);
or U11835 (N_11835,N_1229,N_3503);
nor U11836 (N_11836,N_7727,N_1810);
nor U11837 (N_11837,N_5501,N_9131);
or U11838 (N_11838,N_1981,N_4106);
nor U11839 (N_11839,N_4184,N_3557);
or U11840 (N_11840,N_8710,N_4148);
or U11841 (N_11841,N_4110,N_9644);
nand U11842 (N_11842,N_1049,N_8824);
nand U11843 (N_11843,N_8962,N_8796);
or U11844 (N_11844,N_5680,N_433);
or U11845 (N_11845,N_3196,N_5721);
or U11846 (N_11846,N_7227,N_3714);
nor U11847 (N_11847,N_9827,N_8081);
nand U11848 (N_11848,N_9870,N_5530);
and U11849 (N_11849,N_4601,N_1124);
nor U11850 (N_11850,N_444,N_4443);
or U11851 (N_11851,N_9528,N_3895);
and U11852 (N_11852,N_6433,N_9689);
nor U11853 (N_11853,N_4138,N_3298);
nand U11854 (N_11854,N_4420,N_9891);
or U11855 (N_11855,N_7557,N_2929);
nor U11856 (N_11856,N_63,N_6405);
or U11857 (N_11857,N_6775,N_5549);
or U11858 (N_11858,N_3355,N_9472);
nor U11859 (N_11859,N_423,N_8169);
nand U11860 (N_11860,N_3827,N_216);
and U11861 (N_11861,N_6686,N_5);
nor U11862 (N_11862,N_9850,N_9072);
or U11863 (N_11863,N_415,N_2174);
or U11864 (N_11864,N_8956,N_609);
nand U11865 (N_11865,N_1135,N_2102);
nor U11866 (N_11866,N_719,N_1456);
nand U11867 (N_11867,N_5673,N_4223);
and U11868 (N_11868,N_8574,N_9771);
or U11869 (N_11869,N_927,N_801);
or U11870 (N_11870,N_923,N_8850);
nor U11871 (N_11871,N_6341,N_4249);
and U11872 (N_11872,N_6490,N_4600);
nand U11873 (N_11873,N_9908,N_9588);
nor U11874 (N_11874,N_448,N_7123);
nor U11875 (N_11875,N_666,N_159);
nand U11876 (N_11876,N_6047,N_4129);
nand U11877 (N_11877,N_2059,N_3535);
nor U11878 (N_11878,N_3194,N_9920);
and U11879 (N_11879,N_7645,N_5545);
xor U11880 (N_11880,N_3645,N_866);
and U11881 (N_11881,N_1917,N_9657);
nand U11882 (N_11882,N_9783,N_7363);
or U11883 (N_11883,N_3486,N_1854);
nand U11884 (N_11884,N_3622,N_4571);
nor U11885 (N_11885,N_5830,N_6243);
nand U11886 (N_11886,N_7854,N_4562);
nor U11887 (N_11887,N_8608,N_3010);
nand U11888 (N_11888,N_1943,N_1087);
and U11889 (N_11889,N_6719,N_7032);
nor U11890 (N_11890,N_56,N_5699);
and U11891 (N_11891,N_597,N_1942);
or U11892 (N_11892,N_3764,N_2651);
xnor U11893 (N_11893,N_2703,N_6078);
xnor U11894 (N_11894,N_8908,N_8075);
nor U11895 (N_11895,N_2667,N_2882);
nand U11896 (N_11896,N_8401,N_7818);
and U11897 (N_11897,N_2906,N_2851);
nand U11898 (N_11898,N_3437,N_4);
and U11899 (N_11899,N_1213,N_6090);
nand U11900 (N_11900,N_4884,N_9753);
and U11901 (N_11901,N_7931,N_6826);
nand U11902 (N_11902,N_3556,N_5114);
nand U11903 (N_11903,N_5595,N_9301);
nand U11904 (N_11904,N_2769,N_9956);
and U11905 (N_11905,N_7872,N_8285);
nand U11906 (N_11906,N_4505,N_4145);
or U11907 (N_11907,N_5402,N_8492);
and U11908 (N_11908,N_9366,N_1812);
nor U11909 (N_11909,N_5320,N_1184);
and U11910 (N_11910,N_274,N_1209);
xnor U11911 (N_11911,N_7643,N_559);
nand U11912 (N_11912,N_4599,N_1183);
nor U11913 (N_11913,N_1611,N_7082);
or U11914 (N_11914,N_6348,N_1182);
nor U11915 (N_11915,N_9326,N_6331);
and U11916 (N_11916,N_2263,N_1550);
and U11917 (N_11917,N_7509,N_4544);
xor U11918 (N_11918,N_261,N_2382);
nor U11919 (N_11919,N_770,N_1837);
nand U11920 (N_11920,N_5933,N_619);
or U11921 (N_11921,N_3614,N_2230);
nor U11922 (N_11922,N_5666,N_6605);
xor U11923 (N_11923,N_5546,N_2337);
nor U11924 (N_11924,N_9344,N_2707);
or U11925 (N_11925,N_2922,N_1900);
nand U11926 (N_11926,N_4545,N_1947);
or U11927 (N_11927,N_1445,N_3117);
or U11928 (N_11928,N_2673,N_6706);
or U11929 (N_11929,N_3845,N_9487);
nor U11930 (N_11930,N_6247,N_7589);
nor U11931 (N_11931,N_7586,N_3727);
or U11932 (N_11932,N_1302,N_8057);
nand U11933 (N_11933,N_784,N_2903);
and U11934 (N_11934,N_1406,N_9792);
and U11935 (N_11935,N_9018,N_8293);
xor U11936 (N_11936,N_4579,N_6777);
or U11937 (N_11937,N_8372,N_1264);
and U11938 (N_11938,N_5513,N_6860);
nand U11939 (N_11939,N_2377,N_4120);
nor U11940 (N_11940,N_7182,N_510);
or U11941 (N_11941,N_2704,N_5093);
nor U11942 (N_11942,N_1894,N_8613);
and U11943 (N_11943,N_3672,N_214);
xnor U11944 (N_11944,N_9534,N_7616);
or U11945 (N_11945,N_2771,N_9863);
xor U11946 (N_11946,N_9430,N_2303);
and U11947 (N_11947,N_2420,N_5594);
or U11948 (N_11948,N_3932,N_5568);
nand U11949 (N_11949,N_1559,N_9790);
and U11950 (N_11950,N_7556,N_6350);
and U11951 (N_11951,N_2682,N_5773);
nor U11952 (N_11952,N_7841,N_6574);
or U11953 (N_11953,N_2339,N_8448);
nand U11954 (N_11954,N_3793,N_3988);
nor U11955 (N_11955,N_9980,N_4829);
and U11956 (N_11956,N_5180,N_6781);
and U11957 (N_11957,N_7323,N_7943);
and U11958 (N_11958,N_5314,N_9759);
and U11959 (N_11959,N_8295,N_8446);
nor U11960 (N_11960,N_7489,N_3452);
nor U11961 (N_11961,N_9770,N_2193);
nand U11962 (N_11962,N_4213,N_9335);
nor U11963 (N_11963,N_9002,N_6510);
nor U11964 (N_11964,N_310,N_1800);
nand U11965 (N_11965,N_3924,N_9016);
nand U11966 (N_11966,N_9723,N_1244);
nand U11967 (N_11967,N_5974,N_3628);
or U11968 (N_11968,N_5171,N_4372);
or U11969 (N_11969,N_8616,N_5651);
and U11970 (N_11970,N_1576,N_634);
nor U11971 (N_11971,N_2132,N_9099);
nand U11972 (N_11972,N_1792,N_2960);
or U11973 (N_11973,N_4879,N_6053);
nor U11974 (N_11974,N_5321,N_6427);
or U11975 (N_11975,N_3774,N_4127);
and U11976 (N_11976,N_9491,N_996);
or U11977 (N_11977,N_1261,N_9114);
and U11978 (N_11978,N_9184,N_4297);
xor U11979 (N_11979,N_7985,N_9951);
nand U11980 (N_11980,N_1029,N_111);
nor U11981 (N_11981,N_6968,N_1516);
nor U11982 (N_11982,N_4104,N_9865);
and U11983 (N_11983,N_9768,N_1467);
and U11984 (N_11984,N_7441,N_847);
nand U11985 (N_11985,N_4904,N_1081);
nand U11986 (N_11986,N_2350,N_6664);
nor U11987 (N_11987,N_8056,N_5727);
and U11988 (N_11988,N_7739,N_3353);
xnor U11989 (N_11989,N_6672,N_438);
and U11990 (N_11990,N_7253,N_3902);
and U11991 (N_11991,N_98,N_997);
or U11992 (N_11992,N_2628,N_8527);
nor U11993 (N_11993,N_9373,N_9172);
nand U11994 (N_11994,N_7104,N_851);
nand U11995 (N_11995,N_8439,N_8803);
nor U11996 (N_11996,N_311,N_4338);
nor U11997 (N_11997,N_3991,N_3495);
nand U11998 (N_11998,N_8923,N_2017);
or U11999 (N_11999,N_9815,N_1098);
nor U12000 (N_12000,N_5503,N_1351);
nor U12001 (N_12001,N_981,N_2520);
and U12002 (N_12002,N_8070,N_142);
xnor U12003 (N_12003,N_4785,N_6085);
and U12004 (N_12004,N_7451,N_7568);
nor U12005 (N_12005,N_1986,N_5127);
and U12006 (N_12006,N_7485,N_8532);
or U12007 (N_12007,N_2765,N_4239);
or U12008 (N_12008,N_8195,N_524);
and U12009 (N_12009,N_9643,N_6932);
or U12010 (N_12010,N_4468,N_7417);
and U12011 (N_12011,N_3239,N_227);
nand U12012 (N_12012,N_427,N_405);
or U12013 (N_12013,N_5414,N_5883);
nand U12014 (N_12014,N_8888,N_8371);
and U12015 (N_12015,N_3326,N_7387);
nand U12016 (N_12016,N_6507,N_1133);
nor U12017 (N_12017,N_5403,N_5079);
and U12018 (N_12018,N_5254,N_9464);
nand U12019 (N_12019,N_5276,N_6766);
and U12020 (N_12020,N_9998,N_3185);
xnor U12021 (N_12021,N_1377,N_8333);
and U12022 (N_12022,N_3000,N_6833);
or U12023 (N_12023,N_2315,N_2060);
xnor U12024 (N_12024,N_6745,N_4320);
nand U12025 (N_12025,N_6069,N_793);
nor U12026 (N_12026,N_7540,N_685);
and U12027 (N_12027,N_1956,N_1663);
nand U12028 (N_12028,N_678,N_1568);
nor U12029 (N_12029,N_1305,N_2954);
nand U12030 (N_12030,N_2695,N_6377);
nor U12031 (N_12031,N_9502,N_3668);
nor U12032 (N_12032,N_1203,N_3268);
and U12033 (N_12033,N_7453,N_8294);
xor U12034 (N_12034,N_2473,N_9456);
and U12035 (N_12035,N_9917,N_2136);
nor U12036 (N_12036,N_293,N_692);
or U12037 (N_12037,N_671,N_9235);
or U12038 (N_12038,N_6515,N_5379);
and U12039 (N_12039,N_9229,N_3257);
or U12040 (N_12040,N_8224,N_4502);
or U12041 (N_12041,N_1780,N_8915);
nor U12042 (N_12042,N_567,N_751);
nor U12043 (N_12043,N_5557,N_4077);
nor U12044 (N_12044,N_5618,N_5987);
or U12045 (N_12045,N_1412,N_5456);
or U12046 (N_12046,N_9994,N_5048);
nor U12047 (N_12047,N_7716,N_2129);
nor U12048 (N_12048,N_2243,N_2204);
xnor U12049 (N_12049,N_1413,N_6581);
nand U12050 (N_12050,N_4991,N_4331);
and U12051 (N_12051,N_2788,N_7718);
nor U12052 (N_12052,N_7773,N_2472);
and U12053 (N_12053,N_639,N_4043);
nor U12054 (N_12054,N_8987,N_9213);
nand U12055 (N_12055,N_2582,N_1251);
or U12056 (N_12056,N_8059,N_4740);
or U12057 (N_12057,N_2117,N_776);
and U12058 (N_12058,N_1852,N_5574);
nor U12059 (N_12059,N_1816,N_2972);
nand U12060 (N_12060,N_9840,N_7201);
xor U12061 (N_12061,N_3791,N_7838);
nor U12062 (N_12062,N_4979,N_2913);
or U12063 (N_12063,N_408,N_5496);
or U12064 (N_12064,N_6077,N_4833);
nor U12065 (N_12065,N_9712,N_7103);
and U12066 (N_12066,N_7963,N_1926);
nand U12067 (N_12067,N_8474,N_7423);
and U12068 (N_12068,N_6764,N_907);
nor U12069 (N_12069,N_1790,N_4771);
or U12070 (N_12070,N_2933,N_3779);
or U12071 (N_12071,N_6873,N_2168);
nand U12072 (N_12072,N_9299,N_75);
or U12073 (N_12073,N_7543,N_732);
xnor U12074 (N_12074,N_4170,N_8588);
or U12075 (N_12075,N_3731,N_7630);
nor U12076 (N_12076,N_8578,N_6297);
or U12077 (N_12077,N_284,N_7077);
and U12078 (N_12078,N_3320,N_7973);
and U12079 (N_12079,N_2925,N_9203);
nand U12080 (N_12080,N_902,N_2833);
xnor U12081 (N_12081,N_3386,N_8695);
or U12082 (N_12082,N_6409,N_4745);
and U12083 (N_12083,N_262,N_7125);
nor U12084 (N_12084,N_5917,N_7480);
xor U12085 (N_12085,N_2832,N_8977);
and U12086 (N_12086,N_5593,N_2085);
or U12087 (N_12087,N_9884,N_4414);
nand U12088 (N_12088,N_1148,N_3429);
nand U12089 (N_12089,N_8901,N_5407);
nand U12090 (N_12090,N_9241,N_8352);
and U12091 (N_12091,N_4973,N_5610);
or U12092 (N_12092,N_8864,N_1101);
or U12093 (N_12093,N_3618,N_7979);
and U12094 (N_12094,N_2455,N_861);
or U12095 (N_12095,N_7056,N_247);
or U12096 (N_12096,N_9576,N_2488);
or U12097 (N_12097,N_5662,N_4592);
nand U12098 (N_12098,N_1710,N_7880);
and U12099 (N_12099,N_7434,N_6746);
and U12100 (N_12100,N_618,N_2156);
and U12101 (N_12101,N_7794,N_2773);
and U12102 (N_12102,N_4846,N_6175);
xnor U12103 (N_12103,N_9587,N_934);
xnor U12104 (N_12104,N_7709,N_1945);
and U12105 (N_12105,N_3032,N_6606);
or U12106 (N_12106,N_4265,N_2502);
nand U12107 (N_12107,N_3210,N_2011);
or U12108 (N_12108,N_3551,N_4896);
or U12109 (N_12109,N_6038,N_7231);
nand U12110 (N_12110,N_4454,N_277);
and U12111 (N_12111,N_2224,N_1653);
or U12112 (N_12112,N_6838,N_2674);
or U12113 (N_12113,N_841,N_472);
and U12114 (N_12114,N_1585,N_4806);
or U12115 (N_12115,N_9941,N_5136);
nor U12116 (N_12116,N_2605,N_1721);
nor U12117 (N_12117,N_1354,N_2025);
nor U12118 (N_12118,N_4383,N_9887);
or U12119 (N_12119,N_1622,N_5238);
nand U12120 (N_12120,N_4753,N_9316);
and U12121 (N_12121,N_6208,N_1843);
xnor U12122 (N_12122,N_3310,N_8134);
and U12123 (N_12123,N_2566,N_5069);
and U12124 (N_12124,N_4963,N_9869);
xor U12125 (N_12125,N_8361,N_7840);
or U12126 (N_12126,N_5758,N_181);
nor U12127 (N_12127,N_1786,N_9354);
or U12128 (N_12128,N_4087,N_9358);
or U12129 (N_12129,N_7980,N_8185);
or U12130 (N_12130,N_7458,N_2711);
nor U12131 (N_12131,N_2552,N_9968);
nand U12132 (N_12132,N_8869,N_72);
or U12133 (N_12133,N_1791,N_1625);
and U12134 (N_12134,N_8787,N_5161);
xnor U12135 (N_12135,N_998,N_9101);
xnor U12136 (N_12136,N_2320,N_687);
nand U12137 (N_12137,N_8457,N_3315);
nand U12138 (N_12138,N_2048,N_1457);
or U12139 (N_12139,N_2902,N_5522);
or U12140 (N_12140,N_1920,N_6384);
and U12141 (N_12141,N_4318,N_6858);
nand U12142 (N_12142,N_987,N_5135);
nand U12143 (N_12143,N_1025,N_6959);
and U12144 (N_12144,N_5422,N_5911);
xor U12145 (N_12145,N_3892,N_8699);
or U12146 (N_12146,N_2715,N_8138);
and U12147 (N_12147,N_9890,N_9287);
and U12148 (N_12148,N_8676,N_7330);
or U12149 (N_12149,N_2288,N_9976);
nor U12150 (N_12150,N_8809,N_670);
nand U12151 (N_12151,N_4743,N_6269);
xor U12152 (N_12152,N_6224,N_7635);
and U12153 (N_12153,N_515,N_7692);
nor U12154 (N_12154,N_5763,N_1243);
nand U12155 (N_12155,N_3183,N_4159);
and U12156 (N_12156,N_4230,N_5128);
and U12157 (N_12157,N_7374,N_9446);
nor U12158 (N_12158,N_8685,N_8541);
or U12159 (N_12159,N_3296,N_5849);
nand U12160 (N_12160,N_3800,N_2355);
nand U12161 (N_12161,N_2796,N_1344);
and U12162 (N_12162,N_3848,N_4210);
xnor U12163 (N_12163,N_5280,N_6655);
nor U12164 (N_12164,N_9970,N_3162);
xnor U12165 (N_12165,N_9463,N_8925);
nand U12166 (N_12166,N_3097,N_1030);
nand U12167 (N_12167,N_9202,N_7937);
or U12168 (N_12168,N_9164,N_2965);
nor U12169 (N_12169,N_593,N_2171);
and U12170 (N_12170,N_4268,N_6749);
nor U12171 (N_12171,N_7848,N_2446);
nor U12172 (N_12172,N_5357,N_5577);
or U12173 (N_12173,N_8455,N_2254);
nand U12174 (N_12174,N_826,N_5077);
xor U12175 (N_12175,N_4791,N_7309);
xor U12176 (N_12176,N_9261,N_9581);
nor U12177 (N_12177,N_3566,N_6789);
or U12178 (N_12178,N_7166,N_6123);
or U12179 (N_12179,N_8944,N_5019);
nand U12180 (N_12180,N_9035,N_3649);
nand U12181 (N_12181,N_8319,N_2753);
and U12182 (N_12182,N_1174,N_5862);
nand U12183 (N_12183,N_6818,N_1937);
or U12184 (N_12184,N_97,N_256);
and U12185 (N_12185,N_4445,N_3713);
nand U12186 (N_12186,N_7348,N_4142);
or U12187 (N_12187,N_3202,N_738);
nor U12188 (N_12188,N_2812,N_688);
nor U12189 (N_12189,N_8175,N_5541);
or U12190 (N_12190,N_5216,N_8853);
nand U12191 (N_12191,N_2529,N_4779);
nor U12192 (N_12192,N_7674,N_6303);
nand U12193 (N_12193,N_3968,N_2134);
nor U12194 (N_12194,N_7249,N_406);
nor U12195 (N_12195,N_233,N_9570);
or U12196 (N_12196,N_1477,N_6282);
nand U12197 (N_12197,N_3703,N_1070);
or U12198 (N_12198,N_6253,N_4940);
nand U12199 (N_12199,N_382,N_1345);
nand U12200 (N_12200,N_7806,N_7143);
nor U12201 (N_12201,N_8135,N_9709);
and U12202 (N_12202,N_9611,N_7779);
nand U12203 (N_12203,N_780,N_5096);
nor U12204 (N_12204,N_2767,N_4122);
xor U12205 (N_12205,N_5316,N_7161);
nand U12206 (N_12206,N_4358,N_7369);
nor U12207 (N_12207,N_2191,N_5514);
or U12208 (N_12208,N_3199,N_7752);
nor U12209 (N_12209,N_7050,N_5011);
or U12210 (N_12210,N_3828,N_9467);
nor U12211 (N_12211,N_2112,N_9725);
or U12212 (N_12212,N_1807,N_5441);
or U12213 (N_12213,N_1038,N_1382);
nor U12214 (N_12214,N_4200,N_4955);
or U12215 (N_12215,N_2216,N_4209);
nand U12216 (N_12216,N_2625,N_5221);
xnor U12217 (N_12217,N_8998,N_119);
and U12218 (N_12218,N_3387,N_1368);
xor U12219 (N_12219,N_6011,N_6122);
nand U12220 (N_12220,N_7583,N_6765);
or U12221 (N_12221,N_5748,N_8152);
and U12222 (N_12222,N_6850,N_144);
and U12223 (N_12223,N_470,N_1785);
nor U12224 (N_12224,N_6453,N_8127);
nor U12225 (N_12225,N_6825,N_1309);
nor U12226 (N_12226,N_6528,N_1265);
xor U12227 (N_12227,N_620,N_6908);
or U12228 (N_12228,N_1711,N_2202);
nand U12229 (N_12229,N_1643,N_3585);
nand U12230 (N_12230,N_2631,N_2374);
and U12231 (N_12231,N_2065,N_1573);
nand U12232 (N_12232,N_1744,N_4951);
nand U12233 (N_12233,N_8871,N_7793);
nand U12234 (N_12234,N_483,N_9224);
or U12235 (N_12235,N_4007,N_1903);
nor U12236 (N_12236,N_5246,N_7907);
or U12237 (N_12237,N_9251,N_5834);
nor U12238 (N_12238,N_3417,N_6566);
or U12239 (N_12239,N_2683,N_4944);
nor U12240 (N_12240,N_1455,N_1618);
nand U12241 (N_12241,N_3877,N_7471);
xnor U12242 (N_12242,N_3262,N_7215);
or U12243 (N_12243,N_3170,N_9439);
nand U12244 (N_12244,N_6514,N_4149);
or U12245 (N_12245,N_3846,N_4859);
nor U12246 (N_12246,N_9702,N_6621);
xor U12247 (N_12247,N_825,N_2660);
nor U12248 (N_12248,N_5073,N_9786);
nand U12249 (N_12249,N_173,N_585);
and U12250 (N_12250,N_8344,N_722);
nor U12251 (N_12251,N_6229,N_125);
nand U12252 (N_12252,N_3747,N_6120);
and U12253 (N_12253,N_3947,N_9868);
xor U12254 (N_12254,N_1781,N_3392);
nand U12255 (N_12255,N_7553,N_1285);
xnor U12256 (N_12256,N_713,N_4831);
or U12257 (N_12257,N_47,N_508);
and U12258 (N_12258,N_4667,N_7296);
or U12259 (N_12259,N_8360,N_8656);
or U12260 (N_12260,N_827,N_9349);
nor U12261 (N_12261,N_412,N_2905);
nand U12262 (N_12262,N_544,N_1598);
or U12263 (N_12263,N_9104,N_2414);
and U12264 (N_12264,N_5256,N_5470);
and U12265 (N_12265,N_1716,N_9726);
nor U12266 (N_12266,N_4893,N_2840);
and U12267 (N_12267,N_9381,N_5565);
nor U12268 (N_12268,N_2255,N_8485);
xnor U12269 (N_12269,N_1804,N_4496);
and U12270 (N_12270,N_9,N_4617);
and U12271 (N_12271,N_9407,N_9268);
and U12272 (N_12272,N_1695,N_8848);
or U12273 (N_12273,N_3797,N_8443);
and U12274 (N_12274,N_8580,N_3267);
nand U12275 (N_12275,N_8228,N_209);
nand U12276 (N_12276,N_6055,N_8235);
and U12277 (N_12277,N_2114,N_6018);
xor U12278 (N_12278,N_3063,N_101);
and U12279 (N_12279,N_8425,N_9662);
nand U12280 (N_12280,N_2331,N_3760);
and U12281 (N_12281,N_2513,N_5099);
nand U12282 (N_12282,N_9600,N_366);
and U12283 (N_12283,N_9800,N_5220);
or U12284 (N_12284,N_8202,N_4799);
and U12285 (N_12285,N_9420,N_8484);
nor U12286 (N_12286,N_5004,N_4378);
nand U12287 (N_12287,N_4199,N_6126);
nand U12288 (N_12288,N_7187,N_8651);
or U12289 (N_12289,N_410,N_8218);
and U12290 (N_12290,N_4295,N_8496);
and U12291 (N_12291,N_2852,N_8876);
nor U12292 (N_12292,N_4927,N_3849);
and U12293 (N_12293,N_6073,N_8856);
or U12294 (N_12294,N_9300,N_9519);
nor U12295 (N_12295,N_8793,N_6996);
nand U12296 (N_12296,N_8129,N_1617);
nand U12297 (N_12297,N_5597,N_8017);
nand U12298 (N_12298,N_7345,N_2319);
nand U12299 (N_12299,N_4728,N_7572);
or U12300 (N_12300,N_161,N_2968);
or U12301 (N_12301,N_6603,N_3457);
or U12302 (N_12302,N_3784,N_3653);
or U12303 (N_12303,N_4303,N_4543);
xor U12304 (N_12304,N_1230,N_8652);
and U12305 (N_12305,N_9068,N_4908);
and U12306 (N_12306,N_3896,N_5438);
nor U12307 (N_12307,N_5060,N_7372);
and U12308 (N_12308,N_6965,N_9341);
nand U12309 (N_12309,N_7503,N_2871);
or U12310 (N_12310,N_796,N_4214);
nand U12311 (N_12311,N_9412,N_2659);
or U12312 (N_12312,N_1341,N_5237);
nor U12313 (N_12313,N_2238,N_2781);
nor U12314 (N_12314,N_4843,N_7766);
nand U12315 (N_12315,N_8072,N_3024);
and U12316 (N_12316,N_3726,N_4807);
nor U12317 (N_12317,N_5033,N_8686);
xnor U12318 (N_12318,N_1040,N_3419);
or U12319 (N_12319,N_9763,N_8184);
nand U12320 (N_12320,N_2361,N_4410);
or U12321 (N_12321,N_9415,N_9832);
nand U12322 (N_12322,N_1679,N_1288);
nor U12323 (N_12323,N_6974,N_9141);
xor U12324 (N_12324,N_3587,N_1740);
nor U12325 (N_12325,N_8141,N_4026);
nor U12326 (N_12326,N_6889,N_2547);
nor U12327 (N_12327,N_234,N_3920);
nand U12328 (N_12328,N_9453,N_4375);
and U12329 (N_12329,N_9931,N_7559);
nor U12330 (N_12330,N_2656,N_6033);
nand U12331 (N_12331,N_8200,N_9835);
nand U12332 (N_12332,N_9987,N_3120);
nand U12333 (N_12333,N_9290,N_8875);
and U12334 (N_12334,N_7609,N_2868);
and U12335 (N_12335,N_6385,N_8974);
or U12336 (N_12336,N_4348,N_8186);
or U12337 (N_12337,N_5306,N_2675);
nor U12338 (N_12338,N_8164,N_3639);
and U12339 (N_12339,N_1591,N_4306);
or U12340 (N_12340,N_5015,N_3660);
and U12341 (N_12341,N_6052,N_8222);
nand U12342 (N_12342,N_5023,N_592);
or U12343 (N_12343,N_4085,N_5106);
xor U12344 (N_12344,N_1480,N_6201);
nor U12345 (N_12345,N_3683,N_844);
and U12346 (N_12346,N_5554,N_9311);
xnor U12347 (N_12347,N_2927,N_2318);
xor U12348 (N_12348,N_8584,N_2066);
nand U12349 (N_12349,N_8703,N_7867);
xnor U12350 (N_12350,N_2006,N_7803);
or U12351 (N_12351,N_9275,N_7072);
and U12352 (N_12352,N_9989,N_7058);
and U12353 (N_12353,N_3916,N_8981);
nand U12354 (N_12354,N_8687,N_8339);
nand U12355 (N_12355,N_3763,N_3919);
nor U12356 (N_12356,N_1993,N_5190);
or U12357 (N_12357,N_7781,N_7511);
or U12358 (N_12358,N_1952,N_6927);
or U12359 (N_12359,N_9896,N_7778);
nor U12360 (N_12360,N_9609,N_4764);
nand U12361 (N_12361,N_5728,N_6618);
and U12362 (N_12362,N_8269,N_4354);
nor U12363 (N_12363,N_8300,N_3167);
nor U12364 (N_12364,N_6964,N_9673);
nand U12365 (N_12365,N_9690,N_6690);
or U12366 (N_12366,N_1983,N_555);
nand U12367 (N_12367,N_2451,N_8660);
xor U12368 (N_12368,N_8812,N_1431);
nor U12369 (N_12369,N_9056,N_9475);
or U12370 (N_12370,N_2918,N_3862);
nor U12371 (N_12371,N_3937,N_5578);
xor U12372 (N_12372,N_3165,N_9372);
or U12373 (N_12373,N_6691,N_2155);
nor U12374 (N_12374,N_6080,N_958);
and U12375 (N_12375,N_2409,N_8559);
xnor U12376 (N_12376,N_1918,N_9589);
nand U12377 (N_12377,N_869,N_808);
nor U12378 (N_12378,N_4385,N_3303);
or U12379 (N_12379,N_3462,N_8647);
or U12380 (N_12380,N_5345,N_3680);
nand U12381 (N_12381,N_2524,N_4146);
xor U12382 (N_12382,N_2932,N_2914);
nor U12383 (N_12383,N_5877,N_6437);
nor U12384 (N_12384,N_8623,N_9179);
nand U12385 (N_12385,N_8829,N_1990);
nor U12386 (N_12386,N_1427,N_7844);
and U12387 (N_12387,N_1730,N_5832);
and U12388 (N_12388,N_1850,N_668);
and U12389 (N_12389,N_6554,N_203);
xor U12390 (N_12390,N_9045,N_1360);
or U12391 (N_12391,N_6049,N_5570);
nand U12392 (N_12392,N_1505,N_8012);
and U12393 (N_12393,N_3432,N_8587);
xor U12394 (N_12394,N_2173,N_2143);
xnor U12395 (N_12395,N_6082,N_2930);
and U12396 (N_12396,N_4948,N_7962);
nor U12397 (N_12397,N_193,N_3109);
or U12398 (N_12398,N_6132,N_5994);
and U12399 (N_12399,N_2853,N_3905);
nand U12400 (N_12400,N_2284,N_4427);
nor U12401 (N_12401,N_9842,N_1443);
and U12402 (N_12402,N_8750,N_4117);
nor U12403 (N_12403,N_6498,N_435);
nand U12404 (N_12404,N_4448,N_4103);
and U12405 (N_12405,N_8828,N_514);
xor U12406 (N_12406,N_1651,N_7083);
xnor U12407 (N_12407,N_575,N_3767);
nand U12408 (N_12408,N_4563,N_5553);
nor U12409 (N_12409,N_5274,N_2020);
nand U12410 (N_12410,N_7450,N_882);
nor U12411 (N_12411,N_8965,N_5957);
or U12412 (N_12412,N_5614,N_1067);
xor U12413 (N_12413,N_8404,N_8554);
xor U12414 (N_12414,N_9107,N_5230);
and U12415 (N_12415,N_674,N_8715);
and U12416 (N_12416,N_9973,N_3757);
or U12417 (N_12417,N_8254,N_3554);
and U12418 (N_12418,N_4715,N_269);
and U12419 (N_12419,N_2395,N_6019);
nor U12420 (N_12420,N_4615,N_2178);
nand U12421 (N_12421,N_7192,N_2971);
and U12422 (N_12422,N_1145,N_5775);
nand U12423 (N_12423,N_7443,N_1552);
nand U12424 (N_12424,N_3284,N_4588);
xnor U12425 (N_12425,N_4985,N_6279);
nand U12426 (N_12426,N_680,N_313);
or U12427 (N_12427,N_2159,N_8451);
and U12428 (N_12428,N_8988,N_5852);
and U12429 (N_12429,N_7800,N_5715);
xor U12430 (N_12430,N_4343,N_3009);
nand U12431 (N_12431,N_6602,N_7226);
xnor U12432 (N_12432,N_354,N_6106);
nor U12433 (N_12433,N_6109,N_1803);
nor U12434 (N_12434,N_4227,N_4395);
and U12435 (N_12435,N_4473,N_2701);
nand U12436 (N_12436,N_1976,N_3769);
nand U12437 (N_12437,N_7791,N_8573);
or U12438 (N_12438,N_7742,N_989);
or U12439 (N_12439,N_6268,N_4183);
nor U12440 (N_12440,N_7119,N_749);
nand U12441 (N_12441,N_9188,N_3305);
or U12442 (N_12442,N_5170,N_6288);
nand U12443 (N_12443,N_4298,N_8043);
nor U12444 (N_12444,N_938,N_249);
nor U12445 (N_12445,N_859,N_4260);
nor U12446 (N_12446,N_6504,N_7011);
nor U12447 (N_12447,N_8468,N_9504);
or U12448 (N_12448,N_4891,N_5416);
nand U12449 (N_12449,N_4241,N_6110);
nand U12450 (N_12450,N_1697,N_1268);
or U12451 (N_12451,N_9120,N_8731);
nor U12452 (N_12452,N_9597,N_3662);
and U12453 (N_12453,N_6045,N_62);
nor U12454 (N_12454,N_2273,N_4180);
nand U12455 (N_12455,N_7669,N_3844);
and U12456 (N_12456,N_7996,N_8236);
and U12457 (N_12457,N_7602,N_329);
nor U12458 (N_12458,N_5313,N_460);
nand U12459 (N_12459,N_2073,N_7392);
nand U12460 (N_12460,N_7736,N_1738);
nand U12461 (N_12461,N_5787,N_763);
or U12462 (N_12462,N_6644,N_3936);
nor U12463 (N_12463,N_4827,N_2201);
or U12464 (N_12464,N_8156,N_2602);
nor U12465 (N_12465,N_6030,N_5737);
nor U12466 (N_12466,N_82,N_5377);
xnor U12467 (N_12467,N_9654,N_9458);
nand U12468 (N_12468,N_1879,N_5115);
and U12469 (N_12469,N_8701,N_4822);
and U12470 (N_12470,N_4101,N_8270);
and U12471 (N_12471,N_8375,N_2449);
xor U12472 (N_12472,N_9125,N_1795);
and U12473 (N_12473,N_8971,N_6325);
or U12474 (N_12474,N_3091,N_2777);
xor U12475 (N_12475,N_9434,N_9555);
or U12476 (N_12476,N_7315,N_1138);
nor U12477 (N_12477,N_8241,N_1043);
nand U12478 (N_12478,N_45,N_9965);
nor U12479 (N_12479,N_5977,N_6223);
nand U12480 (N_12480,N_7599,N_8341);
nand U12481 (N_12481,N_711,N_890);
xor U12482 (N_12482,N_2480,N_635);
or U12483 (N_12483,N_5030,N_9991);
and U12484 (N_12484,N_1704,N_8952);
and U12485 (N_12485,N_9546,N_8296);
xor U12486 (N_12486,N_52,N_9069);
and U12487 (N_12487,N_1008,N_7092);
nor U12488 (N_12488,N_4457,N_1588);
nand U12489 (N_12489,N_4010,N_837);
and U12490 (N_12490,N_8810,N_242);
nand U12491 (N_12491,N_8577,N_3426);
nor U12492 (N_12492,N_8790,N_8622);
nor U12493 (N_12493,N_7047,N_8011);
nand U12494 (N_12494,N_6683,N_9138);
or U12495 (N_12495,N_9964,N_4281);
or U12496 (N_12496,N_8311,N_4254);
and U12497 (N_12497,N_7155,N_7096);
nand U12498 (N_12498,N_8558,N_8247);
or U12499 (N_12499,N_564,N_2572);
or U12500 (N_12500,N_615,N_617);
or U12501 (N_12501,N_1582,N_5895);
and U12502 (N_12502,N_9370,N_5083);
nor U12503 (N_12503,N_9223,N_7772);
nor U12504 (N_12504,N_2057,N_5627);
or U12505 (N_12505,N_1602,N_8946);
nand U12506 (N_12506,N_4255,N_471);
and U12507 (N_12507,N_7078,N_8355);
nand U12508 (N_12508,N_520,N_3022);
and U12509 (N_12509,N_699,N_7607);
or U12510 (N_12510,N_8883,N_3654);
or U12511 (N_12511,N_4628,N_4074);
or U12512 (N_12512,N_1071,N_7390);
and U12513 (N_12513,N_4604,N_8797);
nor U12514 (N_12514,N_8113,N_6895);
and U12515 (N_12515,N_2197,N_7837);
or U12516 (N_12516,N_1336,N_5191);
nor U12517 (N_12517,N_2688,N_1674);
and U12518 (N_12518,N_2309,N_8327);
nor U12519 (N_12519,N_2240,N_8762);
and U12520 (N_12520,N_6884,N_3734);
nor U12521 (N_12521,N_4670,N_5750);
nor U12522 (N_12522,N_5922,N_5121);
nor U12523 (N_12523,N_2549,N_3144);
nand U12524 (N_12524,N_7700,N_2131);
nand U12525 (N_12525,N_9338,N_7723);
and U12526 (N_12526,N_6831,N_2990);
nand U12527 (N_12527,N_8571,N_7644);
nor U12528 (N_12528,N_1964,N_8502);
or U12529 (N_12529,N_7048,N_7017);
and U12530 (N_12530,N_2724,N_8756);
and U12531 (N_12531,N_994,N_606);
and U12532 (N_12532,N_8004,N_2805);
nand U12533 (N_12533,N_5681,N_6950);
or U12534 (N_12534,N_6728,N_2947);
or U12535 (N_12535,N_6810,N_3070);
nor U12536 (N_12536,N_9143,N_8964);
nor U12537 (N_12537,N_8139,N_6138);
and U12538 (N_12538,N_2768,N_7144);
and U12539 (N_12539,N_9187,N_6174);
and U12540 (N_12540,N_3232,N_2626);
and U12541 (N_12541,N_548,N_4816);
nor U12542 (N_12542,N_1468,N_1021);
nand U12543 (N_12543,N_4638,N_6757);
or U12544 (N_12544,N_9236,N_4128);
nand U12545 (N_12545,N_7255,N_6920);
nor U12546 (N_12546,N_8855,N_9714);
nand U12547 (N_12547,N_9859,N_1861);
or U12548 (N_12548,N_6086,N_7501);
and U12549 (N_12549,N_7089,N_6631);
and U12550 (N_12550,N_3648,N_9554);
or U12551 (N_12551,N_9310,N_6061);
and U12552 (N_12552,N_2657,N_1959);
nor U12553 (N_12553,N_6623,N_9592);
or U12554 (N_12554,N_6894,N_6379);
or U12555 (N_12555,N_8921,N_7597);
nand U12556 (N_12556,N_6955,N_3373);
xnor U12557 (N_12557,N_9163,N_8515);
or U12558 (N_12558,N_8399,N_1109);
nor U12559 (N_12559,N_9158,N_4430);
xnor U12560 (N_12560,N_4360,N_7378);
nand U12561 (N_12561,N_5252,N_658);
and U12562 (N_12562,N_4494,N_409);
or U12563 (N_12563,N_5519,N_3311);
or U12564 (N_12564,N_7156,N_4838);
and U12565 (N_12565,N_1204,N_5952);
nor U12566 (N_12566,N_1899,N_4542);
or U12567 (N_12567,N_4251,N_8634);
nand U12568 (N_12568,N_352,N_8092);
and U12569 (N_12569,N_6095,N_102);
nor U12570 (N_12570,N_9046,N_5385);
nor U12571 (N_12571,N_9283,N_3343);
and U12572 (N_12572,N_2910,N_3474);
and U12573 (N_12573,N_6559,N_7261);
nand U12574 (N_12574,N_3132,N_4330);
or U12575 (N_12575,N_1006,N_1346);
nor U12576 (N_12576,N_7006,N_4842);
and U12577 (N_12577,N_4113,N_4197);
and U12578 (N_12578,N_3976,N_9044);
nor U12579 (N_12579,N_7097,N_1007);
xnor U12580 (N_12580,N_9292,N_3631);
and U12581 (N_12581,N_4677,N_6374);
or U12582 (N_12582,N_819,N_9429);
nor U12583 (N_12583,N_4868,N_9427);
nor U12584 (N_12584,N_1205,N_8322);
or U12585 (N_12585,N_7898,N_2412);
nor U12586 (N_12586,N_3367,N_3710);
nand U12587 (N_12587,N_2215,N_8926);
and U12588 (N_12588,N_7300,N_3056);
or U12589 (N_12589,N_5538,N_501);
xnor U12590 (N_12590,N_1396,N_7797);
or U12591 (N_12591,N_7297,N_4919);
and U12592 (N_12592,N_3160,N_6836);
nand U12593 (N_12593,N_2585,N_7319);
and U12594 (N_12594,N_8050,N_5841);
nand U12595 (N_12595,N_3217,N_1221);
and U12596 (N_12596,N_9999,N_4978);
nor U12597 (N_12597,N_8609,N_4652);
xnor U12598 (N_12598,N_2185,N_7882);
nor U12599 (N_12599,N_522,N_7935);
or U12600 (N_12600,N_3142,N_4844);
and U12601 (N_12601,N_1638,N_2834);
or U12602 (N_12602,N_4627,N_2587);
nand U12603 (N_12603,N_1405,N_7036);
nand U12604 (N_12604,N_7449,N_2110);
xor U12605 (N_12605,N_5143,N_1931);
and U12606 (N_12606,N_4688,N_9954);
xor U12607 (N_12607,N_1012,N_1777);
nor U12608 (N_12608,N_9492,N_8910);
or U12609 (N_12609,N_8563,N_4597);
or U12610 (N_12610,N_8697,N_6794);
nor U12611 (N_12611,N_3514,N_3101);
or U12612 (N_12612,N_4366,N_7573);
nor U12613 (N_12613,N_94,N_4116);
nor U12614 (N_12614,N_321,N_2578);
and U12615 (N_12615,N_8180,N_5725);
nand U12616 (N_12616,N_8733,N_8362);
nor U12617 (N_12617,N_1619,N_834);
nor U12618 (N_12618,N_4920,N_282);
nor U12619 (N_12619,N_7232,N_4526);
or U12620 (N_12620,N_7928,N_9583);
xnor U12621 (N_12621,N_6232,N_715);
nor U12622 (N_12622,N_8406,N_3866);
or U12623 (N_12623,N_4322,N_2234);
nor U12624 (N_12624,N_4082,N_5423);
or U12625 (N_12625,N_8229,N_8852);
and U12626 (N_12626,N_9639,N_8217);
or U12627 (N_12627,N_6580,N_6044);
nor U12628 (N_12628,N_5332,N_318);
and U12629 (N_12629,N_8633,N_7593);
xnor U12630 (N_12630,N_3744,N_6322);
nand U12631 (N_12631,N_5980,N_8920);
nand U12632 (N_12632,N_238,N_5637);
and U12633 (N_12633,N_2483,N_4091);
nor U12634 (N_12634,N_9196,N_7526);
and U12635 (N_12635,N_5208,N_2618);
xnor U12636 (N_12636,N_479,N_3380);
nor U12637 (N_12637,N_1219,N_9647);
or U12638 (N_12638,N_8030,N_2379);
xor U12639 (N_12639,N_4477,N_1333);
and U12640 (N_12640,N_7722,N_3711);
and U12641 (N_12641,N_8282,N_5145);
nor U12642 (N_12642,N_4492,N_3139);
nor U12643 (N_12643,N_7065,N_4676);
and U12644 (N_12644,N_6337,N_2706);
nor U12645 (N_12645,N_6305,N_6693);
and U12646 (N_12646,N_5752,N_7105);
and U12647 (N_12647,N_6651,N_2398);
nor U12648 (N_12648,N_9580,N_8618);
nand U12649 (N_12649,N_6,N_4982);
nor U12650 (N_12650,N_3985,N_6521);
or U12651 (N_12651,N_4699,N_2373);
xor U12652 (N_12652,N_4732,N_1747);
nand U12653 (N_12653,N_8767,N_7787);
and U12654 (N_12654,N_2919,N_3350);
and U12655 (N_12655,N_7429,N_8351);
or U12656 (N_12656,N_1930,N_9888);
nand U12657 (N_12657,N_194,N_2046);
nand U12658 (N_12658,N_6100,N_8842);
or U12659 (N_12659,N_7502,N_8808);
nor U12660 (N_12660,N_694,N_7845);
and U12661 (N_12661,N_4419,N_7648);
nand U12662 (N_12662,N_9226,N_1715);
nor U12663 (N_12663,N_1069,N_2441);
nor U12664 (N_12664,N_2327,N_7393);
and U12665 (N_12665,N_5463,N_4882);
or U12666 (N_12666,N_5797,N_4061);
or U12667 (N_12667,N_8714,N_4339);
nand U12668 (N_12668,N_3154,N_254);
and U12669 (N_12669,N_4051,N_340);
or U12670 (N_12670,N_8957,N_175);
or U12671 (N_12671,N_1503,N_6857);
or U12672 (N_12672,N_2363,N_9161);
and U12673 (N_12673,N_1522,N_4024);
nand U12674 (N_12674,N_6500,N_2615);
and U12675 (N_12675,N_7672,N_129);
and U12676 (N_12676,N_4877,N_2295);
nor U12677 (N_12677,N_4523,N_4826);
or U12678 (N_12678,N_5151,N_2269);
nor U12679 (N_12679,N_8437,N_2434);
nand U12680 (N_12680,N_1714,N_1838);
nand U12681 (N_12681,N_9005,N_8074);
or U12682 (N_12682,N_4942,N_7208);
or U12683 (N_12683,N_179,N_8885);
nor U12684 (N_12684,N_8220,N_7026);
nand U12685 (N_12685,N_272,N_5733);
nor U12686 (N_12686,N_2292,N_6398);
or U12687 (N_12687,N_9052,N_5817);
nor U12688 (N_12688,N_5192,N_599);
nand U12689 (N_12689,N_230,N_594);
xor U12690 (N_12690,N_5204,N_3061);
nor U12691 (N_12691,N_9959,N_7153);
nor U12692 (N_12692,N_6236,N_2886);
nor U12693 (N_12693,N_7353,N_3407);
nor U12694 (N_12694,N_9886,N_5558);
nor U12695 (N_12695,N_5163,N_5566);
xor U12696 (N_12696,N_2608,N_5147);
nor U12697 (N_12697,N_3007,N_3527);
xor U12698 (N_12698,N_5945,N_9821);
nand U12699 (N_12699,N_1929,N_5507);
nor U12700 (N_12700,N_5591,N_5838);
nor U12701 (N_12701,N_3729,N_323);
nand U12702 (N_12702,N_583,N_4404);
nand U12703 (N_12703,N_6264,N_8564);
nor U12704 (N_12704,N_2105,N_1856);
and U12705 (N_12705,N_3224,N_6008);
and U12706 (N_12706,N_7242,N_4655);
or U12707 (N_12707,N_9248,N_4038);
xnor U12708 (N_12708,N_5766,N_5008);
or U12709 (N_12709,N_7402,N_6840);
or U12710 (N_12710,N_9133,N_1500);
nor U12711 (N_12711,N_6556,N_7636);
nand U12712 (N_12712,N_8032,N_553);
nor U12713 (N_12713,N_5118,N_2242);
nor U12714 (N_12714,N_536,N_4757);
and U12715 (N_12715,N_5701,N_5586);
and U12716 (N_12716,N_8370,N_4568);
and U12717 (N_12717,N_5250,N_1471);
or U12718 (N_12718,N_9271,N_2279);
or U12719 (N_12719,N_2291,N_897);
and U12720 (N_12720,N_4355,N_8140);
or U12721 (N_12721,N_3356,N_1478);
nor U12722 (N_12722,N_640,N_6593);
nand U12723 (N_12723,N_265,N_7243);
nor U12724 (N_12724,N_8906,N_1988);
nand U12725 (N_12725,N_9000,N_1770);
or U12726 (N_12726,N_1883,N_6830);
nor U12727 (N_12727,N_5139,N_2217);
nor U12728 (N_12728,N_7049,N_4535);
and U12729 (N_12729,N_6970,N_2140);
and U12730 (N_12730,N_2619,N_466);
xnor U12731 (N_12731,N_5571,N_9270);
nand U12732 (N_12732,N_5378,N_5712);
and U12733 (N_12733,N_298,N_1698);
or U12734 (N_12734,N_239,N_1089);
or U12735 (N_12735,N_6344,N_1614);
or U12736 (N_12736,N_6272,N_9866);
and U12737 (N_12737,N_857,N_4252);
xor U12738 (N_12738,N_5906,N_2556);
nor U12739 (N_12739,N_9895,N_3780);
or U12740 (N_12740,N_3810,N_4737);
and U12741 (N_12741,N_9388,N_9102);
nand U12742 (N_12742,N_3772,N_2982);
nand U12743 (N_12743,N_3591,N_3405);
and U12744 (N_12744,N_4901,N_1189);
xnor U12745 (N_12745,N_8953,N_1970);
and U12746 (N_12746,N_3331,N_6171);
nand U12747 (N_12747,N_9266,N_2967);
or U12748 (N_12748,N_5682,N_2262);
and U12749 (N_12749,N_6465,N_3809);
and U12750 (N_12750,N_9170,N_2558);
nand U12751 (N_12751,N_3084,N_4681);
and U12752 (N_12752,N_9070,N_4565);
and U12753 (N_12753,N_8859,N_6183);
or U12754 (N_12754,N_4776,N_6256);
or U12755 (N_12755,N_9298,N_393);
nor U12756 (N_12756,N_4020,N_6584);
and U12757 (N_12757,N_2893,N_7970);
or U12758 (N_12758,N_2774,N_906);
or U12759 (N_12759,N_3961,N_8463);
and U12760 (N_12760,N_2985,N_3255);
and U12761 (N_12761,N_5850,N_9560);
nor U12762 (N_12762,N_360,N_6635);
or U12763 (N_12763,N_81,N_682);
nor U12764 (N_12764,N_2944,N_3685);
and U12765 (N_12765,N_2953,N_7613);
and U12766 (N_12766,N_149,N_5183);
or U12767 (N_12767,N_5452,N_3384);
nand U12768 (N_12768,N_3584,N_3106);
nor U12769 (N_12769,N_3965,N_5928);
nand U12770 (N_12770,N_5031,N_5740);
nor U12771 (N_12771,N_289,N_6755);
or U12772 (N_12772,N_457,N_8948);
nor U12773 (N_12773,N_1542,N_1713);
xor U12774 (N_12774,N_8891,N_3090);
xor U12775 (N_12775,N_1606,N_367);
and U12776 (N_12776,N_3510,N_6445);
nor U12777 (N_12777,N_8872,N_6946);
nand U12778 (N_12778,N_5404,N_6725);
and U12779 (N_12779,N_3834,N_4513);
nor U12780 (N_12780,N_9730,N_1207);
and U12781 (N_12781,N_5226,N_506);
nor U12782 (N_12782,N_2848,N_3151);
and U12783 (N_12783,N_3149,N_9444);
xnor U12784 (N_12784,N_4444,N_9192);
or U12785 (N_12785,N_2336,N_5281);
or U12786 (N_12786,N_2443,N_2883);
xor U12787 (N_12787,N_43,N_8405);
nand U12788 (N_12788,N_2086,N_1448);
nand U12789 (N_12789,N_4459,N_627);
nor U12790 (N_12790,N_3203,N_1630);
nand U12791 (N_12791,N_4516,N_1093);
nand U12792 (N_12792,N_6402,N_3545);
xnor U12793 (N_12793,N_5486,N_3095);
nand U12794 (N_12794,N_6195,N_8187);
xor U12795 (N_12795,N_2403,N_8252);
or U12796 (N_12796,N_4862,N_5016);
nand U12797 (N_12797,N_4057,N_2416);
nand U12798 (N_12798,N_6888,N_4373);
and U12799 (N_12799,N_6663,N_27);
nand U12800 (N_12800,N_9986,N_319);
nand U12801 (N_12801,N_7992,N_8557);
and U12802 (N_12802,N_3141,N_9523);
or U12803 (N_12803,N_2998,N_4712);
nor U12804 (N_12804,N_4717,N_8771);
or U12805 (N_12805,N_809,N_9897);
nand U12806 (N_12806,N_9257,N_3450);
or U12807 (N_12807,N_6994,N_6283);
and U12808 (N_12808,N_3521,N_8427);
or U12809 (N_12809,N_7942,N_5551);
or U12810 (N_12810,N_8249,N_8061);
nand U12811 (N_12811,N_7997,N_1608);
nand U12812 (N_12812,N_9265,N_3509);
or U12813 (N_12813,N_3946,N_3477);
or U12814 (N_12814,N_5268,N_7929);
nor U12815 (N_12815,N_9433,N_7724);
nand U12816 (N_12816,N_9336,N_3901);
nor U12817 (N_12817,N_2435,N_6131);
xor U12818 (N_12818,N_1502,N_2943);
nand U12819 (N_12819,N_9252,N_5547);
nand U12820 (N_12820,N_8789,N_236);
nand U12821 (N_12821,N_122,N_8250);
nor U12822 (N_12822,N_6848,N_9320);
or U12823 (N_12823,N_7986,N_4416);
and U12824 (N_12824,N_8289,N_3964);
xor U12825 (N_12825,N_1317,N_5197);
and U12826 (N_12826,N_6145,N_2356);
nor U12827 (N_12827,N_5685,N_9242);
nor U12828 (N_12828,N_3664,N_8049);
xor U12829 (N_12829,N_9517,N_2345);
nor U12830 (N_12830,N_3158,N_7265);
and U12831 (N_12831,N_4689,N_3318);
nor U12832 (N_12832,N_363,N_41);
nor U12833 (N_12833,N_6231,N_3842);
or U12834 (N_12834,N_6846,N_3119);
and U12835 (N_12835,N_2437,N_5186);
nor U12836 (N_12836,N_9782,N_740);
or U12837 (N_12837,N_7157,N_8420);
nand U12838 (N_12838,N_6698,N_8611);
nor U12839 (N_12839,N_9538,N_914);
and U12840 (N_12840,N_6615,N_7821);
xor U12841 (N_12841,N_5213,N_3865);
nor U12842 (N_12842,N_6139,N_5807);
xnor U12843 (N_12843,N_7673,N_940);
xor U12844 (N_12844,N_9097,N_2569);
and U12845 (N_12845,N_5126,N_7336);
and U12846 (N_12846,N_6772,N_6356);
and U12847 (N_12847,N_7332,N_2095);
or U12848 (N_12848,N_9985,N_3783);
nand U12849 (N_12849,N_8343,N_4031);
nor U12850 (N_12850,N_5360,N_6852);
xnor U12851 (N_12851,N_1260,N_2082);
and U12852 (N_12852,N_5695,N_5825);
and U12853 (N_12853,N_5999,N_333);
nand U12854 (N_12854,N_138,N_6854);
and U12855 (N_12855,N_3750,N_7863);
and U12856 (N_12856,N_3863,N_2548);
xnor U12857 (N_12857,N_7906,N_5658);
nor U12858 (N_12858,N_5693,N_2);
or U12859 (N_12859,N_3105,N_7990);
or U12860 (N_12860,N_7594,N_1998);
nand U12861 (N_12861,N_3361,N_7445);
or U12862 (N_12862,N_6647,N_7073);
and U12863 (N_12863,N_6254,N_8966);
and U12864 (N_12864,N_6941,N_7364);
and U12865 (N_12865,N_6096,N_6054);
xor U12866 (N_12866,N_9282,N_6306);
nand U12867 (N_12867,N_1367,N_3666);
or U12868 (N_12868,N_6332,N_6137);
nor U12869 (N_12869,N_874,N_535);
nand U12870 (N_12870,N_9105,N_3531);
or U12871 (N_12871,N_9942,N_5490);
xnor U12872 (N_12872,N_5890,N_3630);
nand U12873 (N_12873,N_1100,N_5202);
nor U12874 (N_12874,N_810,N_1004);
nor U12875 (N_12875,N_5286,N_1742);
or U12876 (N_12876,N_8022,N_2069);
nand U12877 (N_12877,N_8120,N_8553);
xor U12878 (N_12878,N_5942,N_5124);
and U12879 (N_12879,N_7487,N_5426);
nor U12880 (N_12880,N_8396,N_8612);
or U12881 (N_12881,N_1754,N_6210);
nand U12882 (N_12882,N_5185,N_9198);
nand U12883 (N_12883,N_8619,N_517);
nand U12884 (N_12884,N_8949,N_6097);
nand U12885 (N_12885,N_2979,N_7541);
nand U12886 (N_12886,N_8968,N_7216);
nand U12887 (N_12887,N_3234,N_7745);
or U12888 (N_12888,N_342,N_3944);
xor U12889 (N_12889,N_816,N_8292);
and U12890 (N_12890,N_8549,N_2290);
and U12891 (N_12891,N_4003,N_4356);
and U12892 (N_12892,N_6995,N_7596);
xnor U12893 (N_12893,N_4425,N_4279);
or U12894 (N_12894,N_1064,N_9146);
or U12895 (N_12895,N_7493,N_9903);
nand U12896 (N_12896,N_5408,N_7847);
and U12897 (N_12897,N_8728,N_7975);
xnor U12898 (N_12898,N_4933,N_2051);
or U12899 (N_12899,N_5943,N_5365);
nand U12900 (N_12900,N_6064,N_5529);
and U12901 (N_12901,N_1284,N_9116);
nand U12902 (N_12902,N_5104,N_305);
or U12903 (N_12903,N_6712,N_6579);
or U12904 (N_12904,N_8166,N_6302);
and U12905 (N_12905,N_456,N_8150);
or U12906 (N_12906,N_3722,N_7535);
or U12907 (N_12907,N_9218,N_5088);
and U12908 (N_12908,N_6028,N_7136);
or U12909 (N_12909,N_5992,N_3274);
or U12910 (N_12910,N_8277,N_8664);
nand U12911 (N_12911,N_1447,N_4593);
nor U12912 (N_12912,N_9789,N_7178);
nor U12913 (N_12913,N_9761,N_883);
and U12914 (N_12914,N_8629,N_6779);
or U12915 (N_12915,N_4409,N_1629);
nor U12916 (N_12916,N_4324,N_659);
and U12917 (N_12917,N_4992,N_5348);
and U12918 (N_12918,N_7245,N_2511);
xnor U12919 (N_12919,N_1886,N_5487);
and U12920 (N_12920,N_9796,N_3484);
and U12921 (N_12921,N_1338,N_5813);
nor U12922 (N_12922,N_3990,N_5014);
and U12923 (N_12923,N_4997,N_1372);
nor U12924 (N_12924,N_8053,N_4501);
nand U12925 (N_12925,N_547,N_3288);
nand U12926 (N_12926,N_9073,N_6737);
and U12927 (N_12927,N_4096,N_5209);
or U12928 (N_12928,N_577,N_7270);
nor U12929 (N_12929,N_3168,N_3372);
nand U12930 (N_12930,N_4808,N_9683);
nand U12931 (N_12931,N_3050,N_2522);
nand U12932 (N_12932,N_8318,N_1855);
and U12933 (N_12933,N_6867,N_2039);
xor U12934 (N_12934,N_6730,N_1594);
or U12935 (N_12935,N_4934,N_8324);
nand U12936 (N_12936,N_2212,N_8902);
xnor U12937 (N_12937,N_7367,N_8976);
xor U12938 (N_12938,N_5249,N_6694);
nand U12939 (N_12939,N_6767,N_3053);
nand U12940 (N_12940,N_9274,N_5223);
and U12941 (N_12941,N_6642,N_7063);
nand U12942 (N_12942,N_8963,N_3316);
nor U12943 (N_12943,N_4539,N_2988);
and U12944 (N_12944,N_7828,N_3241);
and U12945 (N_12945,N_8938,N_2603);
nor U12946 (N_12946,N_8225,N_1504);
and U12947 (N_12947,N_8504,N_6471);
nor U12948 (N_12948,N_8800,N_8445);
nor U12949 (N_12949,N_5167,N_896);
nand U12950 (N_12950,N_8023,N_8838);
and U12951 (N_12951,N_5339,N_6277);
nor U12952 (N_12952,N_2079,N_2936);
nand U12953 (N_12953,N_8422,N_8119);
nor U12954 (N_12954,N_6511,N_8261);
or U12955 (N_12955,N_993,N_5382);
nor U12956 (N_12956,N_386,N_1966);
or U12957 (N_12957,N_6263,N_8242);
and U12958 (N_12958,N_3480,N_9479);
nor U12959 (N_12959,N_2426,N_497);
and U12960 (N_12960,N_9563,N_731);
or U12961 (N_12961,N_750,N_5704);
xnor U12962 (N_12962,N_3498,N_4811);
nor U12963 (N_12963,N_9963,N_105);
or U12964 (N_12964,N_1262,N_5691);
and U12965 (N_12965,N_5774,N_4493);
nor U12966 (N_12966,N_2640,N_6524);
or U12967 (N_12967,N_5946,N_7857);
xnor U12968 (N_12968,N_1063,N_451);
or U12969 (N_12969,N_7658,N_3002);
nand U12970 (N_12970,N_1032,N_2466);
and U12971 (N_12971,N_8167,N_1074);
nor U12972 (N_12972,N_353,N_7999);
nand U12973 (N_12973,N_2470,N_1325);
and U12974 (N_12974,N_6359,N_8109);
nand U12975 (N_12975,N_2543,N_1702);
or U12976 (N_12976,N_2544,N_7490);
nor U12977 (N_12977,N_2676,N_7389);
nor U12978 (N_12978,N_1158,N_3942);
or U12979 (N_12979,N_5362,N_8625);
or U12980 (N_12980,N_3803,N_646);
or U12981 (N_12981,N_7705,N_3671);
or U12982 (N_12982,N_6442,N_7670);
or U12983 (N_12983,N_7974,N_6480);
xor U12984 (N_12984,N_9822,N_9111);
and U12985 (N_12985,N_1078,N_3459);
nor U12986 (N_12986,N_6093,N_3708);
and U12987 (N_12987,N_8621,N_7291);
or U12988 (N_12988,N_8995,N_3069);
nor U12989 (N_12989,N_117,N_2228);
and U12990 (N_12990,N_3089,N_5485);
or U12991 (N_12991,N_9207,N_2897);
and U12992 (N_12992,N_7355,N_9749);
or U12993 (N_12993,N_5899,N_4263);
and U12994 (N_12994,N_6124,N_5575);
nand U12995 (N_12995,N_1729,N_8980);
or U12996 (N_12996,N_4810,N_6051);
or U12997 (N_12997,N_5068,N_8230);
nor U12998 (N_12998,N_605,N_4435);
or U12999 (N_12999,N_1688,N_6238);
and U13000 (N_13000,N_286,N_8488);
or U13001 (N_13001,N_4787,N_8550);
or U13002 (N_13002,N_6383,N_2334);
nand U13003 (N_13003,N_4143,N_5631);
nor U13004 (N_13004,N_9705,N_3121);
nor U13005 (N_13005,N_2775,N_4432);
and U13006 (N_13006,N_3301,N_245);
or U13007 (N_13007,N_4305,N_2607);
xnor U13008 (N_13008,N_6612,N_6760);
nand U13009 (N_13009,N_6634,N_1806);
nor U13010 (N_13010,N_1758,N_7522);
nor U13011 (N_13011,N_6491,N_1082);
nor U13012 (N_13012,N_8581,N_6060);
or U13013 (N_13013,N_5853,N_3175);
nor U13014 (N_13014,N_5799,N_9040);
xor U13015 (N_13015,N_6853,N_6369);
or U13016 (N_13016,N_3841,N_8494);
and U13017 (N_13017,N_3635,N_5912);
nand U13018 (N_13018,N_7662,N_2330);
nand U13019 (N_13019,N_5934,N_563);
nand U13020 (N_13020,N_2861,N_3759);
xnor U13021 (N_13021,N_4708,N_4949);
nand U13022 (N_13022,N_1996,N_4256);
and U13023 (N_13023,N_660,N_4333);
nor U13024 (N_13024,N_2170,N_9858);
or U13025 (N_13025,N_2531,N_5392);
or U13026 (N_13026,N_3209,N_8593);
nor U13027 (N_13027,N_8734,N_9319);
nand U13028 (N_13028,N_8329,N_7310);
and U13029 (N_13029,N_4392,N_1439);
or U13030 (N_13030,N_3826,N_669);
and U13031 (N_13031,N_28,N_4935);
nor U13032 (N_13032,N_9732,N_3539);
or U13033 (N_13033,N_4417,N_8857);
nand U13034 (N_13034,N_9602,N_6113);
or U13035 (N_13035,N_2410,N_7598);
nand U13036 (N_13036,N_1267,N_6170);
and U13037 (N_13037,N_7738,N_1476);
nor U13038 (N_13038,N_1402,N_1895);
and U13039 (N_13039,N_6809,N_4309);
and U13040 (N_13040,N_6308,N_2911);
or U13041 (N_13041,N_153,N_8320);
or U13042 (N_13042,N_5412,N_500);
xnor U13043 (N_13043,N_6586,N_1125);
nor U13044 (N_13044,N_9405,N_4337);
nor U13045 (N_13045,N_8716,N_1417);
and U13046 (N_13046,N_2099,N_9001);
nor U13047 (N_13047,N_8689,N_4164);
or U13048 (N_13048,N_988,N_6865);
and U13049 (N_13049,N_5835,N_8025);
or U13050 (N_13050,N_4073,N_9762);
or U13051 (N_13051,N_3903,N_9013);
nand U13052 (N_13052,N_8904,N_4441);
or U13053 (N_13053,N_929,N_6294);
nand U13054 (N_13054,N_58,N_1009);
and U13055 (N_13055,N_2637,N_5786);
or U13056 (N_13056,N_4316,N_8194);
and U13057 (N_13057,N_1139,N_1720);
nand U13058 (N_13058,N_6112,N_5573);
and U13059 (N_13059,N_964,N_9060);
and U13060 (N_13060,N_1884,N_3869);
xnor U13061 (N_13061,N_3443,N_1864);
and U13062 (N_13062,N_7914,N_6167);
and U13063 (N_13063,N_3107,N_6532);
xor U13064 (N_13064,N_8929,N_5436);
and U13065 (N_13065,N_2920,N_5481);
or U13066 (N_13066,N_8671,N_6732);
xnor U13067 (N_13067,N_2375,N_2955);
or U13068 (N_13068,N_1914,N_2554);
xnor U13069 (N_13069,N_7009,N_532);
or U13070 (N_13070,N_8546,N_5696);
and U13071 (N_13071,N_2176,N_9845);
or U13072 (N_13072,N_6321,N_527);
or U13073 (N_13073,N_519,N_5639);
nand U13074 (N_13074,N_6235,N_7807);
nand U13075 (N_13075,N_5652,N_2797);
nor U13076 (N_13076,N_2402,N_6923);
xnor U13077 (N_13077,N_4317,N_8104);
nand U13078 (N_13078,N_5265,N_5150);
nand U13079 (N_13079,N_8284,N_4389);
and U13080 (N_13080,N_4801,N_3738);
nor U13081 (N_13081,N_5846,N_190);
nor U13082 (N_13082,N_2098,N_8637);
nand U13083 (N_13083,N_5876,N_24);
nand U13084 (N_13084,N_9485,N_8537);
and U13085 (N_13085,N_7329,N_4386);
xor U13086 (N_13086,N_8982,N_6804);
nor U13087 (N_13087,N_3145,N_2321);
and U13088 (N_13088,N_3465,N_1299);
nor U13089 (N_13089,N_6601,N_6386);
nor U13090 (N_13090,N_5855,N_6645);
xor U13091 (N_13091,N_2821,N_9630);
or U13092 (N_13092,N_8461,N_9123);
or U13093 (N_13093,N_4540,N_8310);
or U13094 (N_13094,N_523,N_511);
nand U13095 (N_13095,N_7239,N_1844);
nand U13096 (N_13096,N_3934,N_7871);
nor U13097 (N_13097,N_6416,N_7130);
xnor U13098 (N_13098,N_4135,N_5650);
nor U13099 (N_13099,N_1298,N_273);
nor U13100 (N_13100,N_8063,N_4522);
nor U13101 (N_13101,N_955,N_7484);
nor U13102 (N_13102,N_8257,N_1434);
xor U13103 (N_13103,N_2813,N_9431);
and U13104 (N_13104,N_1072,N_2641);
nand U13105 (N_13105,N_374,N_6911);
nand U13106 (N_13106,N_8046,N_1523);
nand U13107 (N_13107,N_2749,N_6324);
nor U13108 (N_13108,N_6062,N_4374);
or U13109 (N_13109,N_1979,N_7981);
nand U13110 (N_13110,N_901,N_3247);
and U13111 (N_13111,N_1610,N_6847);
xnor U13112 (N_13112,N_8402,N_9940);
or U13113 (N_13113,N_951,N_8878);
or U13114 (N_13114,N_5893,N_9211);
or U13115 (N_13115,N_6744,N_8860);
nor U13116 (N_13116,N_1975,N_6569);
and U13117 (N_13117,N_3246,N_926);
xnor U13118 (N_13118,N_6525,N_7578);
nor U13119 (N_13119,N_9567,N_8951);
nor U13120 (N_13120,N_1003,N_3360);
or U13121 (N_13121,N_8015,N_4766);
nand U13122 (N_13122,N_6967,N_1640);
nor U13123 (N_13123,N_8309,N_5405);
xor U13124 (N_13124,N_1557,N_8603);
nor U13125 (N_13125,N_2387,N_1400);
or U13126 (N_13126,N_4957,N_9547);
or U13127 (N_13127,N_2595,N_5749);
xor U13128 (N_13128,N_1271,N_4528);
xor U13129 (N_13129,N_9740,N_8267);
nor U13130 (N_13130,N_9733,N_5110);
nor U13131 (N_13131,N_6039,N_6898);
or U13132 (N_13132,N_1470,N_9171);
and U13133 (N_13133,N_1645,N_8694);
nor U13134 (N_13134,N_4178,N_114);
or U13135 (N_13135,N_7949,N_9363);
and U13136 (N_13136,N_5435,N_3909);
nand U13137 (N_13137,N_292,N_1094);
nor U13138 (N_13138,N_3039,N_1156);
and U13139 (N_13139,N_7860,N_8244);
and U13140 (N_13140,N_5461,N_4352);
nand U13141 (N_13141,N_4654,N_9039);
and U13142 (N_13142,N_3483,N_4853);
nand U13143 (N_13143,N_5949,N_7207);
or U13144 (N_13144,N_8359,N_1053);
and U13145 (N_13145,N_4577,N_9823);
and U13146 (N_13146,N_589,N_8572);
nor U13147 (N_13147,N_8510,N_602);
or U13148 (N_13148,N_7824,N_7612);
and U13149 (N_13149,N_9081,N_7344);
or U13150 (N_13150,N_3319,N_5732);
xnor U13151 (N_13151,N_8495,N_3999);
nor U13152 (N_13152,N_6266,N_8804);
nor U13153 (N_13153,N_2325,N_8522);
nor U13154 (N_13154,N_9432,N_7013);
nor U13155 (N_13155,N_8681,N_7469);
or U13156 (N_13156,N_14,N_7169);
and U13157 (N_13157,N_662,N_2696);
or U13158 (N_13158,N_3340,N_9246);
nor U13159 (N_13159,N_9413,N_3072);
nor U13160 (N_13160,N_6803,N_1495);
or U13161 (N_13161,N_1615,N_5002);
nor U13162 (N_13162,N_1521,N_2623);
nor U13163 (N_13163,N_2539,N_7420);
and U13164 (N_13164,N_8124,N_345);
nor U13165 (N_13165,N_805,N_7964);
or U13166 (N_13166,N_5076,N_4497);
and U13167 (N_13167,N_8969,N_2436);
nand U13168 (N_13168,N_2815,N_6542);
nand U13169 (N_13169,N_1408,N_3836);
nand U13170 (N_13170,N_5210,N_5981);
and U13171 (N_13171,N_2161,N_7842);
nand U13172 (N_13172,N_5039,N_8639);
xor U13173 (N_13173,N_8811,N_858);
and U13174 (N_13174,N_5598,N_9159);
nand U13175 (N_13175,N_2351,N_2071);
or U13176 (N_13176,N_7915,N_2678);
nor U13177 (N_13177,N_5300,N_4754);
nor U13178 (N_13178,N_6978,N_7504);
and U13179 (N_13179,N_3911,N_3475);
nand U13180 (N_13180,N_753,N_3716);
nand U13181 (N_13181,N_1596,N_186);
and U13182 (N_13182,N_4661,N_8730);
and U13183 (N_13183,N_8597,N_2743);
xnor U13184 (N_13184,N_5493,N_1599);
or U13185 (N_13185,N_3478,N_3577);
or U13186 (N_13186,N_9197,N_1216);
nor U13187 (N_13187,N_833,N_3712);
and U13188 (N_13188,N_5656,N_3717);
or U13189 (N_13189,N_5063,N_3449);
nand U13190 (N_13190,N_2828,N_7649);
nor U13191 (N_13191,N_8844,N_5793);
or U13192 (N_13192,N_9425,N_104);
or U13193 (N_13193,N_8213,N_6265);
nand U13194 (N_13194,N_8670,N_7951);
nand U13195 (N_13195,N_1151,N_7307);
and U13196 (N_13196,N_8669,N_2097);
nor U13197 (N_13197,N_4261,N_3887);
or U13198 (N_13198,N_5235,N_7223);
nor U13199 (N_13199,N_5878,N_1554);
or U13200 (N_13200,N_845,N_4450);
xor U13201 (N_13201,N_8014,N_5193);
or U13202 (N_13202,N_8108,N_879);
xnor U13203 (N_13203,N_1240,N_8095);
nor U13204 (N_13204,N_1076,N_4950);
nand U13205 (N_13205,N_7281,N_6071);
xor U13206 (N_13206,N_3163,N_246);
and U13207 (N_13207,N_6983,N_9875);
nand U13208 (N_13208,N_120,N_1700);
and U13209 (N_13209,N_4083,N_5261);
or U13210 (N_13210,N_8978,N_675);
nand U13211 (N_13211,N_6392,N_7171);
and U13212 (N_13212,N_6565,N_3285);
nor U13213 (N_13213,N_2083,N_5844);
nand U13214 (N_13214,N_4621,N_4515);
nand U13215 (N_13215,N_6553,N_3295);
and U13216 (N_13216,N_505,N_1535);
nor U13217 (N_13217,N_4150,N_2106);
and U13218 (N_13218,N_6057,N_6748);
nand U13219 (N_13219,N_452,N_7991);
nand U13220 (N_13220,N_3414,N_8922);
and U13221 (N_13221,N_3689,N_7183);
nand U13222 (N_13222,N_2506,N_5173);
nand U13223 (N_13223,N_5864,N_397);
nor U13224 (N_13224,N_4216,N_3430);
and U13225 (N_13225,N_2419,N_1046);
nand U13226 (N_13226,N_6319,N_2742);
xor U13227 (N_13227,N_4733,N_4029);
nand U13228 (N_13228,N_8693,N_4290);
nand U13229 (N_13229,N_5770,N_7912);
nand U13230 (N_13230,N_3607,N_6415);
or U13231 (N_13231,N_70,N_1195);
nor U13232 (N_13232,N_7399,N_6837);
nand U13233 (N_13233,N_5040,N_4132);
nor U13234 (N_13234,N_922,N_9930);
and U13235 (N_13235,N_9003,N_3977);
xor U13236 (N_13236,N_1973,N_1927);
nand U13237 (N_13237,N_6408,N_9981);
nand U13238 (N_13238,N_6163,N_5138);
nand U13239 (N_13239,N_7762,N_7967);
and U13240 (N_13240,N_7360,N_5806);
nor U13241 (N_13241,N_4698,N_9312);
or U13242 (N_13242,N_2266,N_3741);
nand U13243 (N_13243,N_5882,N_7051);
or U13244 (N_13244,N_5080,N_2183);
nand U13245 (N_13245,N_2127,N_2575);
xor U13246 (N_13246,N_1472,N_7719);
nor U13247 (N_13247,N_3829,N_1381);
and U13248 (N_13248,N_9608,N_5159);
nor U13249 (N_13249,N_6141,N_3254);
and U13250 (N_13250,N_6128,N_317);
nand U13251 (N_13251,N_5113,N_2621);
nand U13252 (N_13252,N_7337,N_1971);
or U13253 (N_13253,N_4072,N_5324);
and U13254 (N_13254,N_1460,N_6357);
nand U13255 (N_13255,N_5731,N_8216);
nor U13256 (N_13256,N_5669,N_4349);
nand U13257 (N_13257,N_891,N_3395);
and U13258 (N_13258,N_3015,N_9484);
and U13259 (N_13259,N_3099,N_6032);
nor U13260 (N_13260,N_7884,N_5334);
and U13261 (N_13261,N_8830,N_8979);
nand U13262 (N_13262,N_2277,N_9926);
nand U13263 (N_13263,N_4126,N_9752);
nand U13264 (N_13264,N_5137,N_3524);
or U13265 (N_13265,N_6701,N_3496);
nor U13266 (N_13266,N_4289,N_6173);
nor U13267 (N_13267,N_9374,N_7110);
xor U13268 (N_13268,N_9328,N_5454);
and U13269 (N_13269,N_9264,N_1968);
or U13270 (N_13270,N_6410,N_9132);
and U13271 (N_13271,N_1834,N_552);
and U13272 (N_13272,N_8312,N_2391);
nor U13273 (N_13273,N_2126,N_9807);
nor U13274 (N_13274,N_8849,N_4491);
xor U13275 (N_13275,N_3458,N_3461);
or U13276 (N_13276,N_8819,N_6081);
or U13277 (N_13277,N_2400,N_4221);
nor U13278 (N_13278,N_3891,N_1214);
and U13279 (N_13279,N_3059,N_7086);
or U13280 (N_13280,N_3735,N_5971);
and U13281 (N_13281,N_2182,N_4345);
nand U13282 (N_13282,N_5154,N_7547);
and U13283 (N_13283,N_9698,N_6221);
xnor U13284 (N_13284,N_6444,N_6792);
or U13285 (N_13285,N_2613,N_3492);
or U13286 (N_13286,N_9543,N_4100);
and U13287 (N_13287,N_4294,N_9380);
and U13288 (N_13288,N_2362,N_9355);
or U13289 (N_13289,N_676,N_6048);
or U13290 (N_13290,N_5778,N_5683);
or U13291 (N_13291,N_6688,N_373);
or U13292 (N_13292,N_3228,N_3534);
or U13293 (N_13293,N_434,N_9737);
xnor U13294 (N_13294,N_6659,N_3075);
or U13295 (N_13295,N_9200,N_852);
or U13296 (N_13296,N_3264,N_7782);
and U13297 (N_13297,N_8440,N_7186);
or U13298 (N_13298,N_5811,N_2484);
nor U13299 (N_13299,N_4039,N_2891);
or U13300 (N_13300,N_2997,N_5429);
and U13301 (N_13301,N_2024,N_9872);
or U13302 (N_13302,N_2404,N_9009);
nand U13303 (N_13303,N_2843,N_6158);
and U13304 (N_13304,N_1200,N_4284);
nand U13305 (N_13305,N_4783,N_1960);
and U13306 (N_13306,N_6022,N_2909);
nand U13307 (N_13307,N_5720,N_2029);
or U13308 (N_13308,N_8737,N_8021);
or U13309 (N_13309,N_913,N_3001);
nand U13310 (N_13310,N_1612,N_7212);
nand U13311 (N_13311,N_4751,N_3174);
nand U13312 (N_13312,N_9285,N_1796);
or U13313 (N_13313,N_9082,N_781);
nor U13314 (N_13314,N_5119,N_2244);
xnor U13315 (N_13315,N_831,N_5938);
xnor U13316 (N_13316,N_1779,N_3064);
and U13317 (N_13317,N_9945,N_6769);
nor U13318 (N_13318,N_1459,N_9758);
and U13319 (N_13319,N_5865,N_143);
and U13320 (N_13320,N_1273,N_5051);
or U13321 (N_13321,N_1319,N_8099);
nand U13322 (N_13322,N_3705,N_5160);
or U13323 (N_13323,N_3567,N_8026);
nor U13324 (N_13324,N_5858,N_4088);
and U13325 (N_13325,N_7124,N_3719);
nor U13326 (N_13326,N_5273,N_4480);
nand U13327 (N_13327,N_9284,N_3728);
nand U13328 (N_13328,N_5936,N_3959);
nand U13329 (N_13329,N_3913,N_9756);
nor U13330 (N_13330,N_3819,N_954);
nand U13331 (N_13331,N_4034,N_8606);
and U13332 (N_13332,N_5777,N_2666);
and U13333 (N_13333,N_4812,N_8854);
xnor U13334 (N_13334,N_4772,N_5920);
xnor U13335 (N_13335,N_2622,N_7711);
nor U13336 (N_13336,N_9549,N_7267);
nor U13337 (N_13337,N_8576,N_1873);
and U13338 (N_13338,N_5711,N_8583);
and U13339 (N_13339,N_1669,N_9404);
xnor U13340 (N_13340,N_270,N_8456);
nand U13341 (N_13341,N_6395,N_283);
nand U13342 (N_13342,N_7544,N_9641);
or U13343 (N_13343,N_7993,N_8516);
or U13344 (N_13344,N_1410,N_3739);
nand U13345 (N_13345,N_7132,N_3533);
and U13346 (N_13346,N_4554,N_8817);
nand U13347 (N_13347,N_8565,N_7041);
and U13348 (N_13348,N_9325,N_493);
nor U13349 (N_13349,N_7140,N_4520);
and U13350 (N_13350,N_3885,N_3843);
nand U13351 (N_13351,N_3770,N_5097);
nor U13352 (N_13352,N_8642,N_2211);
or U13353 (N_13353,N_5482,N_7901);
nand U13354 (N_13354,N_4929,N_5072);
and U13355 (N_13355,N_530,N_9946);
and U13356 (N_13356,N_2283,N_7159);
nand U13357 (N_13357,N_7830,N_61);
xor U13358 (N_13358,N_2235,N_6329);
nand U13359 (N_13359,N_1433,N_3444);
nand U13360 (N_13360,N_1023,N_2163);
nand U13361 (N_13361,N_6479,N_1681);
or U13362 (N_13362,N_7870,N_5200);
nand U13363 (N_13363,N_4380,N_3559);
nand U13364 (N_13364,N_6930,N_314);
or U13365 (N_13365,N_5329,N_2551);
nor U13366 (N_13366,N_7437,N_6682);
nand U13367 (N_13367,N_3472,N_4220);
nor U13368 (N_13368,N_5356,N_4455);
nor U13369 (N_13369,N_9228,N_6362);
nor U13370 (N_13370,N_9900,N_9779);
nand U13371 (N_13371,N_9145,N_3198);
nor U13372 (N_13372,N_1531,N_4557);
and U13373 (N_13373,N_6468,N_3272);
nand U13374 (N_13374,N_1320,N_8772);
and U13375 (N_13375,N_4690,N_4845);
nand U13376 (N_13376,N_1002,N_1652);
and U13377 (N_13377,N_7278,N_3281);
or U13378 (N_13378,N_7189,N_8276);
nor U13379 (N_13379,N_8478,N_9023);
nor U13380 (N_13380,N_848,N_2491);
and U13381 (N_13381,N_5029,N_4669);
and U13382 (N_13382,N_9361,N_4789);
nor U13383 (N_13383,N_6870,N_7492);
and U13384 (N_13384,N_5279,N_7760);
nand U13385 (N_13385,N_2670,N_3327);
or U13386 (N_13386,N_3956,N_8315);
nand U13387 (N_13387,N_6736,N_7634);
nand U13388 (N_13388,N_4311,N_8330);
and U13389 (N_13389,N_4723,N_8107);
and U13390 (N_13390,N_2028,N_1385);
nand U13391 (N_13391,N_7413,N_2133);
or U13392 (N_13392,N_9024,N_9465);
and U13393 (N_13393,N_3540,N_1079);
and U13394 (N_13394,N_8879,N_2816);
nand U13395 (N_13395,N_4157,N_1636);
nor U13396 (N_13396,N_1534,N_6918);
nand U13397 (N_13397,N_6543,N_795);
nor U13398 (N_13398,N_6862,N_3048);
nand U13399 (N_13399,N_3643,N_8548);
or U13400 (N_13400,N_4016,N_2329);
nand U13401 (N_13401,N_1444,N_5212);
or U13402 (N_13402,N_1775,N_7298);
or U13403 (N_13403,N_3817,N_2454);
nand U13404 (N_13404,N_6002,N_7127);
nor U13405 (N_13405,N_1278,N_8248);
or U13406 (N_13406,N_6592,N_8519);
nor U13407 (N_13407,N_863,N_8426);
or U13408 (N_13408,N_1517,N_5881);
or U13409 (N_13409,N_6313,N_4780);
nand U13410 (N_13410,N_1167,N_1509);
nand U13411 (N_13411,N_1830,N_5898);
and U13412 (N_13412,N_6629,N_8163);
or U13413 (N_13413,N_7467,N_5337);
nor U13414 (N_13414,N_9243,N_19);
nand U13415 (N_13415,N_5386,N_2043);
nor U13416 (N_13416,N_7205,N_2899);
xnor U13417 (N_13417,N_5199,N_6815);
nand U13418 (N_13418,N_9460,N_7400);
and U13419 (N_13419,N_7034,N_5527);
nand U13420 (N_13420,N_9628,N_9774);
nor U13421 (N_13421,N_3237,N_264);
nor U13422 (N_13422,N_9324,N_2705);
or U13423 (N_13423,N_267,N_4456);
or U13424 (N_13424,N_3297,N_8627);
or U13425 (N_13425,N_3971,N_3433);
xnor U13426 (N_13426,N_5282,N_3292);
and U13427 (N_13427,N_2063,N_764);
nand U13428 (N_13428,N_2294,N_5278);
nand U13429 (N_13429,N_1936,N_4610);
xnor U13430 (N_13430,N_4198,N_2415);
nor U13431 (N_13431,N_4875,N_2092);
and U13432 (N_13432,N_854,N_6497);
and U13433 (N_13433,N_9879,N_9245);
xnor U13434 (N_13434,N_2050,N_1233);
nor U13435 (N_13435,N_7856,N_8503);
nor U13436 (N_13436,N_3043,N_488);
nor U13437 (N_13437,N_4533,N_1545);
and U13438 (N_13438,N_3725,N_4531);
nand U13439 (N_13439,N_4334,N_1384);
and U13440 (N_13440,N_9969,N_3709);
or U13441 (N_13441,N_9532,N_5654);
nor U13442 (N_13442,N_707,N_7145);
or U13443 (N_13443,N_6204,N_5432);
xor U13444 (N_13444,N_6300,N_5795);
and U13445 (N_13445,N_7945,N_7785);
nand U13446 (N_13446,N_1279,N_1159);
nor U13447 (N_13447,N_3563,N_9332);
or U13448 (N_13448,N_7177,N_8682);
or U13449 (N_13449,N_2592,N_7211);
or U13450 (N_13450,N_2740,N_9988);
nand U13451 (N_13451,N_3409,N_3177);
and U13452 (N_13452,N_8662,N_7376);
or U13453 (N_13453,N_8533,N_2865);
and U13454 (N_13454,N_1616,N_6980);
or U13455 (N_13455,N_294,N_7335);
nor U13456 (N_13456,N_6947,N_5670);
xnor U13457 (N_13457,N_2962,N_191);
nor U13458 (N_13458,N_6245,N_2857);
and U13459 (N_13459,N_5970,N_4582);
nor U13460 (N_13460,N_7494,N_7234);
nand U13461 (N_13461,N_8500,N_7846);
nand U13462 (N_13462,N_8146,N_7276);
nand U13463 (N_13463,N_5383,N_2135);
or U13464 (N_13464,N_941,N_8483);
nor U13465 (N_13465,N_7984,N_4368);
or U13466 (N_13466,N_512,N_7708);
xor U13467 (N_13467,N_2761,N_7911);
and U13468 (N_13468,N_3193,N_9096);
nor U13469 (N_13469,N_2310,N_232);
xor U13470 (N_13470,N_2521,N_1984);
xor U13471 (N_13471,N_1349,N_6509);
xnor U13472 (N_13472,N_1866,N_4897);
and U13473 (N_13473,N_4086,N_5095);
nand U13474 (N_13474,N_724,N_3737);
nor U13475 (N_13475,N_8085,N_6648);
or U13476 (N_13476,N_6187,N_3339);
nand U13477 (N_13477,N_8620,N_1690);
and U13478 (N_13478,N_6985,N_7552);
nor U13479 (N_13479,N_26,N_6669);
nor U13480 (N_13480,N_9667,N_2527);
nand U13481 (N_13481,N_8491,N_8831);
and U13482 (N_13482,N_1249,N_5394);
and U13483 (N_13483,N_8380,N_322);
or U13484 (N_13484,N_1401,N_4602);
or U13485 (N_13485,N_4314,N_1066);
and U13486 (N_13486,N_3908,N_4382);
xor U13487 (N_13487,N_9232,N_241);
or U13488 (N_13488,N_71,N_6202);
and U13489 (N_13489,N_4300,N_4947);
or U13490 (N_13490,N_6849,N_4272);
and U13491 (N_13491,N_1269,N_3018);
xnor U13492 (N_13492,N_4993,N_2458);
and U13493 (N_13493,N_8226,N_790);
or U13494 (N_13494,N_2514,N_6196);
and U13495 (N_13495,N_4267,N_2064);
and U13496 (N_13496,N_8569,N_7524);
nor U13497 (N_13497,N_4738,N_7116);
nor U13498 (N_13498,N_7691,N_2938);
and U13499 (N_13499,N_4498,N_9259);
or U13500 (N_13500,N_9435,N_2831);
and U13501 (N_13501,N_2299,N_9190);
or U13502 (N_13502,N_1263,N_1126);
nor U13503 (N_13503,N_4931,N_327);
and U13504 (N_13504,N_5542,N_3578);
and U13505 (N_13505,N_1764,N_8442);
nor U13506 (N_13506,N_1083,N_8528);
or U13507 (N_13507,N_2247,N_6670);
or U13508 (N_13508,N_2147,N_418);
nand U13509 (N_13509,N_2286,N_8602);
nand U13510 (N_13510,N_9586,N_8698);
and U13511 (N_13511,N_8870,N_5244);
and U13512 (N_13512,N_6244,N_3612);
and U13513 (N_13513,N_4553,N_402);
nand U13514 (N_13514,N_8243,N_4623);
nand U13515 (N_13515,N_8301,N_7904);
nor U13516 (N_13516,N_7334,N_3560);
or U13517 (N_13517,N_5322,N_5497);
nand U13518 (N_13518,N_2809,N_745);
and U13519 (N_13519,N_178,N_237);
nor U13520 (N_13520,N_8786,N_1451);
nand U13521 (N_13521,N_3953,N_3473);
or U13522 (N_13522,N_224,N_3789);
or U13523 (N_13523,N_6454,N_2213);
nand U13524 (N_13524,N_1954,N_6046);
nand U13525 (N_13525,N_4648,N_350);
or U13526 (N_13526,N_843,N_146);
nand U13527 (N_13527,N_4021,N_1575);
or U13528 (N_13528,N_8415,N_7137);
or U13529 (N_13529,N_1603,N_4525);
xor U13530 (N_13530,N_990,N_3507);
or U13531 (N_13531,N_1330,N_717);
or U13532 (N_13532,N_2442,N_9063);
nor U13533 (N_13533,N_3795,N_1234);
xnor U13534 (N_13534,N_4890,N_3775);
nand U13535 (N_13535,N_6118,N_4619);
and U13536 (N_13536,N_7922,N_8290);
and U13537 (N_13537,N_3383,N_5027);
and U13538 (N_13538,N_6877,N_752);
nand U13539 (N_13539,N_4189,N_8752);
xor U13540 (N_13540,N_9615,N_9569);
nand U13541 (N_13541,N_7425,N_8408);
or U13542 (N_13542,N_6973,N_1276);
nor U13543 (N_13543,N_4598,N_2298);
and U13544 (N_13544,N_8794,N_3679);
nor U13545 (N_13545,N_4326,N_5043);
xor U13546 (N_13546,N_8784,N_5061);
or U13547 (N_13547,N_1718,N_1989);
and U13548 (N_13548,N_4788,N_4657);
nand U13549 (N_13549,N_7491,N_3347);
nor U13550 (N_13550,N_1831,N_6735);
or U13551 (N_13551,N_720,N_8003);
nand U13552 (N_13552,N_942,N_2620);
nand U13553 (N_13553,N_4590,N_3325);
and U13554 (N_13554,N_7812,N_6738);
nand U13555 (N_13555,N_799,N_2654);
or U13556 (N_13556,N_1088,N_8338);
nor U13557 (N_13557,N_4023,N_6756);
nor U13558 (N_13558,N_4304,N_7892);
nand U13559 (N_13559,N_1047,N_3923);
and U13560 (N_13560,N_7652,N_8051);
or U13561 (N_13561,N_7147,N_7148);
or U13562 (N_13562,N_147,N_4194);
nand U13563 (N_13563,N_9974,N_8986);
nor U13564 (N_13564,N_8086,N_5744);
and U13565 (N_13565,N_7354,N_9584);
or U13566 (N_13566,N_3205,N_4902);
or U13567 (N_13567,N_2392,N_5052);
nand U13568 (N_13568,N_4486,N_4139);
and U13569 (N_13569,N_1583,N_7375);
nor U13570 (N_13570,N_1836,N_9062);
and U13571 (N_13571,N_6689,N_3984);
and U13572 (N_13572,N_4369,N_1881);
nand U13573 (N_13573,N_792,N_8045);
nand U13574 (N_13574,N_2001,N_5289);
xnor U13575 (N_13575,N_7015,N_6718);
nor U13576 (N_13576,N_7431,N_3969);
and U13577 (N_13577,N_8894,N_3776);
and U13578 (N_13578,N_2610,N_4009);
or U13579 (N_13579,N_4551,N_5338);
and U13580 (N_13580,N_263,N_1555);
nor U13581 (N_13581,N_6370,N_2305);
xor U13582 (N_13582,N_3152,N_5556);
nand U13583 (N_13583,N_9387,N_7350);
and U13584 (N_13584,N_2322,N_8035);
or U13585 (N_13585,N_5094,N_2561);
or U13586 (N_13586,N_5302,N_2718);
and U13587 (N_13587,N_6286,N_7229);
and U13588 (N_13588,N_5054,N_6317);
or U13589 (N_13589,N_8552,N_9022);
nor U13590 (N_13590,N_4472,N_4240);
nand U13591 (N_13591,N_9685,N_974);
nand U13592 (N_13592,N_60,N_7792);
nor U13593 (N_13593,N_6570,N_6561);
nand U13594 (N_13594,N_1465,N_6169);
nor U13595 (N_13595,N_748,N_5311);
nand U13596 (N_13596,N_4438,N_637);
or U13597 (N_13597,N_2565,N_2754);
and U13598 (N_13598,N_7164,N_4506);
or U13599 (N_13599,N_3365,N_900);
nor U13600 (N_13600,N_6275,N_4797);
or U13601 (N_13601,N_2928,N_2062);
nor U13602 (N_13602,N_9505,N_6284);
or U13603 (N_13603,N_3012,N_5294);
or U13604 (N_13604,N_1735,N_424);
and U13605 (N_13605,N_7893,N_3019);
nor U13606 (N_13606,N_921,N_6496);
nand U13607 (N_13607,N_9816,N_2636);
and U13608 (N_13608,N_648,N_5630);
or U13609 (N_13609,N_2941,N_5424);
nor U13610 (N_13610,N_7382,N_8776);
or U13611 (N_13611,N_8526,N_6518);
or U13612 (N_13612,N_1474,N_8101);
or U13613 (N_13613,N_4803,N_550);
nand U13614 (N_13614,N_767,N_4182);
nor U13615 (N_13615,N_3403,N_8007);
xor U13616 (N_13616,N_7623,N_5469);
and U13617 (N_13617,N_5370,N_1292);
nor U13618 (N_13618,N_9788,N_1784);
or U13619 (N_13619,N_9160,N_2677);
and U13620 (N_13620,N_2154,N_8199);
nor U13621 (N_13621,N_9590,N_3346);
and U13622 (N_13622,N_2037,N_5716);
or U13623 (N_13623,N_8258,N_2478);
xnor U13624 (N_13624,N_6673,N_6819);
nor U13625 (N_13625,N_3248,N_1922);
nor U13626 (N_13626,N_6470,N_7976);
nand U13627 (N_13627,N_6455,N_116);
xnor U13628 (N_13628,N_2751,N_4247);
xnor U13629 (N_13629,N_5747,N_9469);
and U13630 (N_13630,N_2271,N_3815);
or U13631 (N_13631,N_1130,N_6821);
and U13632 (N_13632,N_5034,N_2875);
xor U13633 (N_13633,N_3211,N_4692);
nand U13634 (N_13634,N_9121,N_3231);
and U13635 (N_13635,N_9894,N_6835);
nand U13636 (N_13636,N_7989,N_6657);
nor U13637 (N_13637,N_3868,N_127);
nand U13638 (N_13638,N_1274,N_244);
nand U13639 (N_13639,N_7944,N_7697);
xor U13640 (N_13640,N_1841,N_7236);
or U13641 (N_13641,N_9428,N_4687);
and U13642 (N_13642,N_1281,N_8586);
nor U13643 (N_13643,N_4536,N_8350);
or U13644 (N_13644,N_9656,N_6667);
or U13645 (N_13645,N_4040,N_9837);
or U13646 (N_13646,N_4697,N_6188);
nor U13647 (N_13647,N_5690,N_3159);
and U13648 (N_13648,N_5116,N_6519);
and U13649 (N_13649,N_9825,N_5827);
xnor U13650 (N_13650,N_6520,N_5616);
nor U13651 (N_13651,N_3447,N_6934);
nor U13652 (N_13652,N_7373,N_5087);
or U13653 (N_13653,N_103,N_9148);
nor U13654 (N_13654,N_4895,N_346);
nor U13655 (N_13655,N_7396,N_4437);
and U13656 (N_13656,N_6557,N_2474);
xor U13657 (N_13657,N_7941,N_8133);
xnor U13658 (N_13658,N_6091,N_7381);
or U13659 (N_13659,N_6910,N_3504);
and U13660 (N_13660,N_3520,N_1057);
nor U13661 (N_13661,N_2671,N_3771);
or U13662 (N_13662,N_4814,N_4719);
nand U13663 (N_13663,N_9178,N_3434);
or U13664 (N_13664,N_9340,N_712);
nor U13665 (N_13665,N_1731,N_3195);
and U13666 (N_13666,N_6900,N_4018);
xor U13667 (N_13667,N_7667,N_8083);
and U13668 (N_13668,N_9090,N_8721);
and U13669 (N_13669,N_5509,N_6084);
nand U13670 (N_13670,N_6240,N_878);
nand U13671 (N_13671,N_947,N_8031);
or U13672 (N_13672,N_7927,N_9996);
xor U13673 (N_13673,N_3136,N_9544);
nand U13674 (N_13674,N_7054,N_4972);
and U13675 (N_13675,N_5930,N_4614);
or U13676 (N_13676,N_798,N_2697);
nor U13677 (N_13677,N_4532,N_3823);
xor U13678 (N_13678,N_5983,N_576);
or U13679 (N_13679,N_8818,N_4925);
nand U13680 (N_13680,N_9033,N_5672);
and U13681 (N_13681,N_4760,N_6872);
and U13682 (N_13682,N_9185,N_1011);
xor U13683 (N_13683,N_9817,N_5155);
nand U13684 (N_13684,N_8078,N_1091);
or U13685 (N_13685,N_4529,N_5982);
or U13686 (N_13686,N_8774,N_9764);
and U13687 (N_13687,N_9775,N_2946);
nand U13688 (N_13688,N_8903,N_6783);
or U13689 (N_13689,N_1304,N_7516);
nor U13690 (N_13690,N_3471,N_6010);
nand U13691 (N_13691,N_3695,N_6650);
xnor U13692 (N_13692,N_755,N_7180);
nand U13693 (N_13693,N_3611,N_1365);
and U13694 (N_13694,N_3805,N_3410);
and U13695 (N_13695,N_9038,N_4841);
nand U13696 (N_13696,N_4696,N_8009);
xor U13697 (N_13697,N_5130,N_7464);
xor U13698 (N_13698,N_48,N_5905);
nor U13699 (N_13699,N_7536,N_5521);
or U13700 (N_13700,N_4388,N_6786);
nor U13701 (N_13701,N_9244,N_436);
nor U13702 (N_13702,N_7338,N_7654);
and U13703 (N_13703,N_4566,N_507);
or U13704 (N_13704,N_3040,N_7008);
nor U13705 (N_13705,N_6191,N_1734);
nand U13706 (N_13706,N_3382,N_8132);
nand U13707 (N_13707,N_973,N_1654);
nand U13708 (N_13708,N_1529,N_5045);
or U13709 (N_13709,N_6285,N_8317);
and U13710 (N_13710,N_3066,N_830);
and U13711 (N_13711,N_4819,N_7209);
and U13712 (N_13712,N_3859,N_2425);
nand U13713 (N_13713,N_5867,N_6969);
xnor U13714 (N_13714,N_9893,N_6640);
and U13715 (N_13715,N_5028,N_8136);
nand U13716 (N_13716,N_4508,N_6472);
nand U13717 (N_13717,N_8148,N_8130);
or U13718 (N_13718,N_873,N_3150);
or U13719 (N_13719,N_1827,N_3487);
and U13720 (N_13720,N_136,N_7262);
xor U13721 (N_13721,N_7681,N_8834);
xor U13722 (N_13722,N_5089,N_3077);
and U13723 (N_13723,N_5376,N_8617);
or U13724 (N_13724,N_8865,N_5495);
nor U13725 (N_13725,N_645,N_4235);
or U13726 (N_13726,N_9616,N_484);
and U13727 (N_13727,N_7699,N_8768);
nand U13728 (N_13728,N_3042,N_2444);
nor U13729 (N_13729,N_5354,N_2546);
and U13730 (N_13730,N_3880,N_9934);
xnor U13731 (N_13731,N_9606,N_469);
or U13732 (N_13732,N_1527,N_6076);
nor U13733 (N_13733,N_2485,N_4546);
xor U13734 (N_13734,N_7340,N_5788);
nor U13735 (N_13735,N_1551,N_2814);
and U13736 (N_13736,N_5550,N_8524);
nor U13737 (N_13737,N_4983,N_626);
nand U13738 (N_13738,N_5962,N_2825);
and U13739 (N_13739,N_1256,N_8389);
nor U13740 (N_13740,N_8125,N_7256);
or U13741 (N_13741,N_5448,N_8887);
nand U13742 (N_13742,N_817,N_1755);
nand U13743 (N_13743,N_8781,N_2475);
nand U13744 (N_13744,N_734,N_6320);
nor U13745 (N_13745,N_5236,N_9834);
xnor U13746 (N_13746,N_2827,N_3278);
or U13747 (N_13747,N_9810,N_1421);
and U13748 (N_13748,N_8933,N_4647);
or U13749 (N_13749,N_4959,N_3781);
and U13750 (N_13750,N_7461,N_3693);
nand U13751 (N_13751,N_2109,N_9215);
nand U13752 (N_13752,N_7238,N_930);
nand U13753 (N_13753,N_6255,N_6916);
or U13754 (N_13754,N_6678,N_3571);
nor U13755 (N_13755,N_3273,N_6249);
and U13756 (N_13756,N_9947,N_904);
or U13757 (N_13757,N_6652,N_9972);
or U13758 (N_13758,N_3958,N_1096);
nand U13759 (N_13759,N_6921,N_88);
or U13760 (N_13760,N_1655,N_6035);
and U13761 (N_13761,N_4422,N_4108);
or U13762 (N_13762,N_1705,N_419);
nor U13763 (N_13763,N_3103,N_8560);
nand U13764 (N_13764,N_4718,N_5636);
nand U13765 (N_13765,N_8645,N_5959);
and U13766 (N_13766,N_5633,N_3135);
and U13767 (N_13767,N_3651,N_7656);
and U13768 (N_13768,N_3766,N_8840);
nor U13769 (N_13769,N_9717,N_6999);
nor U13770 (N_13770,N_8518,N_1210);
or U13771 (N_13771,N_387,N_9109);
nor U13772 (N_13772,N_1511,N_1569);
nand U13773 (N_13773,N_8749,N_8600);
or U13774 (N_13774,N_3421,N_154);
nand U13775 (N_13775,N_8610,N_6527);
and U13776 (N_13776,N_3169,N_5277);
or U13777 (N_13777,N_6428,N_8880);
and U13778 (N_13778,N_1178,N_3123);
nand U13779 (N_13779,N_9304,N_5870);
nor U13780 (N_13780,N_7059,N_5024);
or U13781 (N_13781,N_3948,N_2794);
nand U13782 (N_13782,N_3031,N_1371);
nor U13783 (N_13783,N_836,N_1466);
xor U13784 (N_13784,N_9938,N_9506);
or U13785 (N_13785,N_1044,N_6225);
or U13786 (N_13786,N_8746,N_2165);
nor U13787 (N_13787,N_5260,N_8833);
and U13788 (N_13788,N_396,N_7710);
nand U13789 (N_13789,N_5837,N_1928);
or U13790 (N_13790,N_2113,N_6573);
nand U13791 (N_13791,N_1693,N_1105);
or U13792 (N_13792,N_8724,N_1154);
and U13793 (N_13793,N_5288,N_3955);
nor U13794 (N_13794,N_2992,N_7052);
nor U13795 (N_13795,N_7196,N_972);
nor U13796 (N_13796,N_4909,N_7184);
or U13797 (N_13797,N_6905,N_7190);
and U13798 (N_13798,N_8984,N_1481);
and U13799 (N_13799,N_1847,N_5333);
or U13800 (N_13800,N_7222,N_9088);
and U13801 (N_13801,N_5327,N_255);
nor U13802 (N_13802,N_6951,N_7576);
nand U13803 (N_13803,N_7357,N_5198);
or U13804 (N_13804,N_1198,N_572);
xor U13805 (N_13805,N_5688,N_3982);
nor U13806 (N_13806,N_8279,N_1173);
nor U13807 (N_13807,N_4851,N_3413);
nor U13808 (N_13808,N_106,N_8893);
nand U13809 (N_13809,N_3324,N_743);
xor U13810 (N_13810,N_8985,N_5555);
xnor U13811 (N_13811,N_5866,N_7587);
nor U13812 (N_13812,N_8950,N_4981);
and U13813 (N_13813,N_531,N_1736);
nand U13814 (N_13814,N_7804,N_4631);
nor U13815 (N_13815,N_9149,N_5168);
or U13816 (N_13816,N_3561,N_5929);
or U13817 (N_13817,N_9960,N_2058);
xor U13818 (N_13818,N_2559,N_903);
or U13819 (N_13819,N_1398,N_1685);
nor U13820 (N_13820,N_1409,N_3688);
and U13821 (N_13821,N_3647,N_4205);
nand U13822 (N_13822,N_4237,N_6796);
or U13823 (N_13823,N_1821,N_9028);
nor U13824 (N_13824,N_9651,N_3068);
xor U13825 (N_13825,N_9490,N_3765);
nand U13826 (N_13826,N_7717,N_3087);
nand U13827 (N_13827,N_4270,N_91);
and U13828 (N_13828,N_4482,N_2463);
nor U13829 (N_13829,N_5298,N_3644);
nor U13830 (N_13830,N_2579,N_189);
and U13831 (N_13831,N_2040,N_4736);
or U13832 (N_13832,N_8679,N_679);
nand U13833 (N_13833,N_5535,N_8153);
nor U13834 (N_13834,N_7042,N_3718);
and U13835 (N_13835,N_7683,N_2250);
and U13836 (N_13836,N_7128,N_3114);
nand U13837 (N_13837,N_3249,N_5205);
nand U13838 (N_13838,N_782,N_2353);
and U13839 (N_13839,N_8143,N_2534);
and U13840 (N_13840,N_32,N_5363);
or U13841 (N_13841,N_2702,N_9739);
or U13842 (N_13842,N_6291,N_6147);
nor U13843 (N_13843,N_2523,N_875);
and U13844 (N_13844,N_802,N_8799);
xor U13845 (N_13845,N_9225,N_5417);
nor U13846 (N_13846,N_4926,N_3212);
or U13847 (N_13847,N_6839,N_4918);
nor U13848 (N_13848,N_5948,N_6791);
and U13849 (N_13849,N_1802,N_8345);
nor U13850 (N_13850,N_64,N_1725);
or U13851 (N_13851,N_6165,N_4365);
nor U13852 (N_13852,N_860,N_714);
nor U13853 (N_13853,N_358,N_9720);
or U13854 (N_13854,N_8735,N_1510);
and U13855 (N_13855,N_7702,N_4722);
nor U13856 (N_13856,N_9443,N_8458);
or U13857 (N_13857,N_5462,N_1712);
or U13858 (N_13858,N_7621,N_7881);
or U13859 (N_13859,N_3186,N_4258);
nand U13860 (N_13860,N_9032,N_2308);
and U13861 (N_13861,N_6182,N_8106);
nand U13862 (N_13862,N_7896,N_8638);
nand U13863 (N_13863,N_1963,N_2926);
and U13864 (N_13864,N_8899,N_6596);
or U13865 (N_13865,N_5964,N_5856);
and U13866 (N_13866,N_9727,N_2732);
nand U13867 (N_13867,N_9794,N_4080);
or U13868 (N_13868,N_6671,N_8741);
or U13869 (N_13869,N_760,N_5152);
or U13870 (N_13870,N_2067,N_7805);
xor U13871 (N_13871,N_7247,N_6754);
nand U13872 (N_13872,N_8240,N_4871);
or U13873 (N_13873,N_5047,N_9079);
or U13874 (N_13874,N_6414,N_1648);
xnor U13875 (N_13875,N_2866,N_5857);
xor U13876 (N_13876,N_9307,N_3073);
nand U13877 (N_13877,N_8897,N_828);
nand U13878 (N_13878,N_6127,N_1366);
xor U13879 (N_13879,N_5900,N_1566);
xnor U13880 (N_13880,N_797,N_4658);
and U13881 (N_13881,N_7299,N_482);
and U13882 (N_13882,N_7940,N_4641);
nor U13883 (N_13883,N_2512,N_7371);
or U13884 (N_13884,N_2080,N_1403);
and U13885 (N_13885,N_2499,N_7947);
or U13886 (N_13886,N_7108,N_9928);
xnor U13887 (N_13887,N_822,N_8821);
xor U13888 (N_13888,N_9975,N_8598);
nor U13889 (N_13889,N_5824,N_2650);
nor U13890 (N_13890,N_2822,N_6841);
and U13891 (N_13891,N_8846,N_4912);
xnor U13892 (N_13892,N_6802,N_5178);
and U13893 (N_13893,N_3606,N_8118);
nor U13894 (N_13894,N_5158,N_7567);
nand U13895 (N_13895,N_8037,N_2386);
nand U13896 (N_13896,N_8624,N_8005);
nor U13897 (N_13897,N_1818,N_1258);
nor U13898 (N_13898,N_3100,N_8378);
nor U13899 (N_13899,N_8650,N_6937);
and U13900 (N_13900,N_3286,N_665);
nand U13901 (N_13901,N_5888,N_6144);
nor U13902 (N_13902,N_1436,N_3201);
or U13903 (N_13903,N_3973,N_7202);
or U13904 (N_13904,N_430,N_769);
xnor U13905 (N_13905,N_5074,N_5989);
nor U13906 (N_13906,N_3625,N_8190);
or U13907 (N_13907,N_4408,N_7620);
nand U13908 (N_13908,N_1773,N_1322);
and U13909 (N_13909,N_8751,N_8745);
and U13910 (N_13910,N_7347,N_4462);
nor U13911 (N_13911,N_1090,N_6340);
nand U13912 (N_13912,N_9748,N_9217);
and U13913 (N_13913,N_4495,N_5057);
xnor U13914 (N_13914,N_341,N_355);
xor U13915 (N_13915,N_1208,N_2863);
nand U13916 (N_13916,N_1227,N_4302);
and U13917 (N_13917,N_2032,N_7795);
nor U13918 (N_13918,N_2942,N_647);
xor U13919 (N_13919,N_596,N_3788);
nand U13920 (N_13920,N_7657,N_4986);
nand U13921 (N_13921,N_3294,N_9746);
and U13922 (N_13922,N_2500,N_8585);
nor U13923 (N_13923,N_7304,N_2770);
or U13924 (N_13924,N_3393,N_3881);
and U13925 (N_13925,N_480,N_4144);
or U13926 (N_13926,N_6687,N_5181);
nand U13927 (N_13927,N_7895,N_8006);
xnor U13928 (N_13928,N_8898,N_4075);
nor U13929 (N_13929,N_9655,N_5760);
and U13930 (N_13930,N_3787,N_1706);
nor U13931 (N_13931,N_4340,N_3455);
xor U13932 (N_13932,N_8959,N_1639);
nor U13933 (N_13933,N_4589,N_1118);
or U13934 (N_13934,N_5066,N_7377);
or U13935 (N_13935,N_5875,N_6012);
nand U13936 (N_13936,N_8732,N_8814);
or U13937 (N_13937,N_3466,N_1898);
nand U13938 (N_13938,N_1241,N_8358);
or U13939 (N_13939,N_9152,N_6246);
nand U13940 (N_13940,N_7465,N_1683);
nand U13941 (N_13941,N_3223,N_8251);
and U13942 (N_13942,N_3599,N_306);
and U13943 (N_13943,N_8690,N_4412);
or U13944 (N_13944,N_4958,N_7018);
xor U13945 (N_13945,N_4607,N_2054);
and U13946 (N_13946,N_7855,N_2424);
or U13947 (N_13947,N_1383,N_8255);
nand U13948 (N_13948,N_7316,N_44);
or U13949 (N_13949,N_3847,N_2937);
or U13950 (N_13950,N_3354,N_7561);
nand U13951 (N_13951,N_1815,N_3604);
nand U13952 (N_13952,N_4351,N_3603);
nand U13953 (N_13953,N_3300,N_3926);
nand U13954 (N_13954,N_5179,N_8486);
or U13955 (N_13955,N_6546,N_6197);
nor U13956 (N_13956,N_2588,N_9478);
nand U13957 (N_13957,N_1165,N_6250);
nand U13958 (N_13958,N_7012,N_3269);
and U13959 (N_13959,N_1446,N_6564);
or U13960 (N_13960,N_4071,N_5474);
or U13961 (N_13961,N_9610,N_9707);
nand U13962 (N_13962,N_4118,N_7653);
and U13963 (N_13963,N_3851,N_5730);
nand U13964 (N_13964,N_9983,N_1604);
and U13965 (N_13965,N_6797,N_9333);
and U13966 (N_13966,N_5842,N_4802);
nand U13967 (N_13967,N_1485,N_757);
or U13968 (N_13968,N_1562,N_7266);
or U13969 (N_13969,N_6429,N_5442);
or U13970 (N_13970,N_1170,N_2864);
nor U13971 (N_13971,N_5464,N_6675);
nand U13972 (N_13972,N_3856,N_3147);
nand U13973 (N_13973,N_3293,N_9297);
nand U13974 (N_13974,N_4965,N_4793);
xnor U13975 (N_13975,N_4815,N_5789);
nand U13976 (N_13976,N_1892,N_4050);
and U13977 (N_13977,N_1058,N_3855);
or U13978 (N_13978,N_4307,N_4721);
or U13979 (N_13979,N_3794,N_3930);
nor U13980 (N_13980,N_3879,N_9659);
xor U13981 (N_13981,N_4407,N_1580);
and U13982 (N_13982,N_5401,N_8431);
or U13983 (N_13983,N_3515,N_2008);
nand U13984 (N_13984,N_8680,N_6721);
nand U13985 (N_13985,N_9352,N_5389);
and U13986 (N_13986,N_3493,N_9681);
nand U13987 (N_13987,N_399,N_2233);
or U13988 (N_13988,N_4036,N_3076);
and U13989 (N_13989,N_5102,N_3753);
nor U13990 (N_13990,N_2367,N_7909);
nor U13991 (N_13991,N_8530,N_1507);
nor U13992 (N_13992,N_2003,N_6771);
nor U13993 (N_13993,N_1247,N_6152);
nand U13994 (N_13994,N_4202,N_8806);
or U13995 (N_13995,N_1196,N_1907);
nand U13996 (N_13996,N_1741,N_8089);
nor U13997 (N_13997,N_4467,N_5745);
and U13998 (N_13998,N_3330,N_5742);
or U13999 (N_13999,N_2152,N_9778);
nand U14000 (N_14000,N_6957,N_1176);
xor U14001 (N_14001,N_6493,N_9317);
xor U14002 (N_14002,N_7551,N_4618);
and U14003 (N_14003,N_9348,N_2074);
and U14004 (N_14004,N_5257,N_6892);
nor U14005 (N_14005,N_7690,N_7325);
nor U14006 (N_14006,N_7601,N_7517);
nand U14007 (N_14007,N_5123,N_3058);
nor U14008 (N_14008,N_6101,N_1851);
or U14009 (N_14009,N_1946,N_4056);
and U14010 (N_14010,N_7135,N_5105);
and U14011 (N_14011,N_6462,N_9167);
or U14012 (N_14012,N_701,N_1380);
xor U14013 (N_14013,N_7826,N_6469);
nor U14014 (N_14014,N_8847,N_8367);
nor U14015 (N_14015,N_7874,N_9445);
nand U14016 (N_14016,N_301,N_789);
nand U14017 (N_14017,N_6806,N_5395);
nand U14018 (N_14018,N_3970,N_8054);
nor U14019 (N_14019,N_3886,N_3253);
nand U14020 (N_14020,N_4832,N_4773);
and U14021 (N_14021,N_3939,N_1708);
nand U14022 (N_14022,N_9695,N_6711);
nor U14023 (N_14023,N_8644,N_6216);
nor U14024 (N_14024,N_6406,N_1586);
nor U14025 (N_14025,N_991,N_8316);
or U14026 (N_14026,N_9556,N_842);
xnor U14027 (N_14027,N_7133,N_4341);
nor U14028 (N_14028,N_673,N_5427);
nand U14029 (N_14029,N_6976,N_5590);
or U14030 (N_14030,N_7244,N_6707);
nor U14031 (N_14031,N_9393,N_1452);
nand U14032 (N_14032,N_7321,N_6874);
and U14033 (N_14033,N_279,N_9978);
nand U14034 (N_14034,N_8168,N_7283);
nand U14035 (N_14035,N_1703,N_176);
nand U14036 (N_14036,N_8556,N_5973);
or U14037 (N_14037,N_2186,N_4866);
or U14038 (N_14038,N_823,N_4828);
and U14039 (N_14039,N_5292,N_7765);
and U14040 (N_14040,N_9692,N_2076);
and U14041 (N_14041,N_9258,N_7479);
and U14042 (N_14042,N_4608,N_4651);
nand U14043 (N_14043,N_207,N_174);
nor U14044 (N_14044,N_4741,N_5746);
nor U14045 (N_14045,N_3041,N_1027);
xor U14046 (N_14046,N_6089,N_6530);
and U14047 (N_14047,N_2012,N_5993);
nor U14048 (N_14048,N_9383,N_2431);
and U14049 (N_14049,N_1664,N_2917);
nand U14050 (N_14050,N_2642,N_5156);
and U14051 (N_14051,N_7839,N_6387);
and U14052 (N_14052,N_6407,N_7823);
or U14053 (N_14053,N_8874,N_6176);
nor U14054 (N_14054,N_4883,N_2342);
or U14055 (N_14055,N_6897,N_9818);
nand U14056 (N_14056,N_5444,N_6271);
nand U14057 (N_14057,N_1166,N_5000);
and U14058 (N_14058,N_74,N_8820);
or U14059 (N_14059,N_4666,N_3037);
or U14060 (N_14060,N_3677,N_9617);
nor U14061 (N_14061,N_3026,N_7240);
nand U14062 (N_14062,N_3835,N_1416);
xor U14063 (N_14063,N_6492,N_4564);
xor U14064 (N_14064,N_7796,N_25);
nand U14065 (N_14065,N_2175,N_2407);
nand U14066 (N_14066,N_4939,N_5879);
nor U14067 (N_14067,N_5768,N_556);
nor U14068 (N_14068,N_8770,N_365);
nor U14069 (N_14069,N_6773,N_2346);
or U14070 (N_14070,N_7085,N_6156);
nand U14071 (N_14071,N_9227,N_7579);
nor U14072 (N_14072,N_9057,N_3456);
nand U14073 (N_14073,N_7626,N_5894);
or U14074 (N_14074,N_6720,N_1750);
or U14075 (N_14075,N_2128,N_5415);
xor U14076 (N_14076,N_401,N_6979);
nor U14077 (N_14077,N_6537,N_5531);
or U14078 (N_14078,N_5344,N_5915);
and U14079 (N_14079,N_3595,N_1231);
nor U14080 (N_14080,N_8356,N_3754);
or U14081 (N_14081,N_5149,N_4821);
nand U14082 (N_14082,N_7053,N_6199);
xnor U14083 (N_14083,N_542,N_2157);
or U14084 (N_14084,N_4226,N_7696);
or U14085 (N_14085,N_6293,N_7410);
nand U14086 (N_14086,N_5563,N_8308);
nor U14087 (N_14087,N_3553,N_8659);
nand U14088 (N_14088,N_6807,N_4560);
and U14089 (N_14089,N_1691,N_4049);
nand U14090 (N_14090,N_6949,N_5466);
nand U14091 (N_14091,N_4656,N_3745);
and U14092 (N_14092,N_9637,N_4236);
nand U14093 (N_14093,N_3342,N_9411);
and U14094 (N_14094,N_8209,N_257);
nor U14095 (N_14095,N_2072,N_1490);
xor U14096 (N_14096,N_761,N_467);
or U14097 (N_14097,N_8545,N_3277);
nand U14098 (N_14098,N_9129,N_5818);
nor U14099 (N_14099,N_5036,N_7463);
nand U14100 (N_14100,N_1005,N_5937);
nor U14101 (N_14101,N_864,N_2869);
nand U14102 (N_14102,N_4673,N_6948);
xor U14103 (N_14103,N_6954,N_5494);
and U14104 (N_14104,N_4353,N_6134);
nand U14105 (N_14105,N_5552,N_150);
and U14106 (N_14106,N_1136,N_3730);
or U14107 (N_14107,N_7397,N_442);
and U14108 (N_14108,N_2557,N_2081);
and U14109 (N_14109,N_2335,N_1293);
nor U14110 (N_14110,N_6582,N_7165);
nand U14111 (N_14111,N_2728,N_4282);
xnor U14112 (N_14112,N_7685,N_5947);
or U14113 (N_14113,N_6315,N_3134);
nand U14114 (N_14114,N_2606,N_1202);
or U14115 (N_14115,N_6526,N_1212);
and U14116 (N_14116,N_9291,N_6654);
or U14117 (N_14117,N_9454,N_4794);
or U14118 (N_14118,N_5909,N_5790);
nor U14119 (N_14119,N_773,N_5743);
and U14120 (N_14120,N_525,N_3943);
xor U14121 (N_14121,N_8531,N_5926);
nor U14122 (N_14122,N_3250,N_6993);
or U14123 (N_14123,N_93,N_9943);
or U14124 (N_14124,N_6352,N_9329);
and U14125 (N_14125,N_8211,N_8115);
nor U14126 (N_14126,N_9423,N_12);
and U14127 (N_14127,N_7,N_8073);
or U14128 (N_14128,N_351,N_2450);
and U14129 (N_14129,N_7924,N_4155);
xnor U14130 (N_14130,N_5647,N_4583);
nand U14131 (N_14131,N_6610,N_4596);
nand U14132 (N_14132,N_8016,N_9334);
nand U14133 (N_14133,N_8851,N_641);
and U14134 (N_14134,N_4259,N_3335);
and U14135 (N_14135,N_8839,N_5184);
or U14136 (N_14136,N_6456,N_7023);
xnor U14137 (N_14137,N_2975,N_4725);
nand U14138 (N_14138,N_8970,N_1978);
nor U14139 (N_14139,N_1042,N_5889);
or U14140 (N_14140,N_54,N_384);
xor U14141 (N_14141,N_7521,N_6925);
xor U14142 (N_14142,N_7185,N_4834);
nor U14143 (N_14143,N_1430,N_7611);
nor U14144 (N_14144,N_7067,N_1728);
and U14145 (N_14145,N_8916,N_6820);
or U14146 (N_14146,N_9545,N_4095);
and U14147 (N_14147,N_8975,N_1671);
xor U14148 (N_14148,N_5851,N_2177);
and U14149 (N_14149,N_5956,N_3489);
or U14150 (N_14150,N_9493,N_4612);
or U14151 (N_14151,N_4937,N_1453);
and U14152 (N_14152,N_600,N_5919);
nand U14153 (N_14153,N_3130,N_7663);
and U14154 (N_14154,N_2272,N_3659);
and U14155 (N_14155,N_5661,N_2107);
nand U14156 (N_14156,N_1155,N_8170);
xor U14157 (N_14157,N_9220,N_3242);
nand U14158 (N_14158,N_7113,N_9302);
or U14159 (N_14159,N_8117,N_1727);
nand U14160 (N_14160,N_7886,N_9633);
or U14161 (N_14161,N_1311,N_8773);
nand U14162 (N_14162,N_6333,N_7057);
nand U14163 (N_14163,N_6180,N_8000);
nor U14164 (N_14164,N_3876,N_6397);
or U14165 (N_14165,N_9416,N_8476);
or U14166 (N_14166,N_5058,N_9982);
nor U14167 (N_14167,N_6529,N_5082);
nand U14168 (N_14168,N_9477,N_4269);
nor U14169 (N_14169,N_6539,N_4537);
and U14170 (N_14170,N_1637,N_2945);
xor U14171 (N_14171,N_1826,N_8691);
and U14172 (N_14172,N_2232,N_7070);
nand U14173 (N_14173,N_961,N_8480);
xor U14174 (N_14174,N_290,N_454);
nand U14175 (N_14175,N_8337,N_5642);
and U14176 (N_14176,N_8630,N_7025);
or U14177 (N_14177,N_288,N_5511);
nor U14178 (N_14178,N_4809,N_5443);
nor U14179 (N_14179,N_7902,N_5548);
or U14180 (N_14180,N_6226,N_6094);
or U14181 (N_14181,N_6040,N_3724);
and U14182 (N_14182,N_3673,N_5738);
and U14183 (N_14183,N_5012,N_6832);
or U14184 (N_14184,N_7715,N_2867);
xor U14185 (N_14185,N_1916,N_9670);
nand U14186 (N_14186,N_4079,N_1462);
nor U14187 (N_14187,N_6741,N_113);
and U14188 (N_14188,N_1108,N_4347);
xnor U14189 (N_14189,N_1823,N_9041);
or U14190 (N_14190,N_2358,N_2995);
xor U14191 (N_14191,N_7966,N_2752);
and U14192 (N_14192,N_1553,N_4076);
nand U14193 (N_14193,N_9708,N_9233);
nand U14194 (N_14194,N_3854,N_9518);
or U14195 (N_14195,N_8561,N_7194);
and U14196 (N_14196,N_925,N_7549);
nor U14197 (N_14197,N_9854,N_5907);
nor U14198 (N_14198,N_6882,N_3057);
or U14199 (N_14199,N_2653,N_4674);
nor U14200 (N_14200,N_5653,N_8605);
and U14201 (N_14201,N_1574,N_9351);
and U14202 (N_14202,N_5270,N_5599);
or U14203 (N_14203,N_3723,N_2720);
nand U14204 (N_14204,N_7172,N_8080);
and U14205 (N_14205,N_6512,N_2218);
and U14206 (N_14206,N_6653,N_8967);
nand U14207 (N_14207,N_2101,N_2760);
nand U14208 (N_14208,N_325,N_9091);
xor U14209 (N_14209,N_8183,N_956);
nand U14210 (N_14210,N_1295,N_8739);
and U14211 (N_14211,N_3871,N_4701);
nor U14212 (N_14212,N_1549,N_3334);
nand U14213 (N_14213,N_1180,N_7624);
nand U14214 (N_14214,N_2370,N_4605);
nand U14215 (N_14215,N_8253,N_9058);
xor U14216 (N_14216,N_7004,N_9801);
xnor U14217 (N_14217,N_5903,N_2710);
nor U14218 (N_14218,N_9571,N_9496);
xnor U14219 (N_14219,N_7258,N_9564);
nor U14220 (N_14220,N_7118,N_7799);
nand U14221 (N_14221,N_9525,N_4678);
nor U14222 (N_14222,N_3921,N_1340);
or U14223 (N_14223,N_9014,N_7701);
and U14224 (N_14224,N_8041,N_76);
or U14225 (N_14225,N_4988,N_4332);
nor U14226 (N_14226,N_4257,N_5620);
and U14227 (N_14227,N_7313,N_7474);
nor U14228 (N_14228,N_1387,N_2376);
nor U14229 (N_14229,N_8262,N_3230);
xor U14230 (N_14230,N_9293,N_3011);
xnor U14231 (N_14231,N_2555,N_5668);
and U14232 (N_14232,N_7139,N_4045);
xor U14233 (N_14233,N_9933,N_5505);
nand U14234 (N_14234,N_2993,N_9176);
and U14235 (N_14235,N_7031,N_8227);
nor U14236 (N_14236,N_9004,N_3446);
nand U14237 (N_14237,N_5358,N_5251);
nor U14238 (N_14238,N_7349,N_3476);
or U14239 (N_14239,N_5923,N_611);
nand U14240 (N_14240,N_5331,N_8841);
nor U14241 (N_14241,N_6859,N_7758);
nor U14242 (N_14242,N_5953,N_9962);
nor U14243 (N_14243,N_2203,N_7608);
or U14244 (N_14244,N_2456,N_6390);
nand U14245 (N_14245,N_4511,N_4541);
nand U14246 (N_14246,N_4371,N_3629);
and U14247 (N_14247,N_5972,N_5413);
nor U14248 (N_14248,N_5296,N_6793);
xor U14249 (N_14249,N_4154,N_3890);
or U14250 (N_14250,N_2429,N_5927);
nand U14251 (N_14251,N_2876,N_6467);
and U14252 (N_14252,N_15,N_8325);
nor U14253 (N_14253,N_5258,N_5540);
xnor U14254 (N_14254,N_8763,N_8535);
nor U14255 (N_14255,N_7028,N_3564);
nor U14256 (N_14256,N_1532,N_9669);
nand U14257 (N_14257,N_2394,N_9447);
or U14258 (N_14258,N_3715,N_328);
xnor U14259 (N_14259,N_6639,N_9719);
xnor U14260 (N_14260,N_6148,N_4168);
and U14261 (N_14261,N_4423,N_2530);
or U14262 (N_14262,N_6871,N_616);
nor U14263 (N_14263,N_7024,N_2904);
xnor U14264 (N_14264,N_3494,N_8816);
and U14265 (N_14265,N_2047,N_2231);
nand U14266 (N_14266,N_1957,N_1761);
and U14267 (N_14267,N_6295,N_2341);
xnor U14268 (N_14268,N_4782,N_5955);
nor U14269 (N_14269,N_6724,N_2108);
and U14270 (N_14270,N_8149,N_6104);
or U14271 (N_14271,N_2791,N_8100);
nor U14272 (N_14272,N_7641,N_9562);
or U14273 (N_14273,N_7913,N_5536);
or U14274 (N_14274,N_9902,N_4584);
and U14275 (N_14275,N_4055,N_9124);
or U14276 (N_14276,N_3637,N_7622);
nand U14277 (N_14277,N_1024,N_5176);
nor U14278 (N_14278,N_7260,N_3646);
nor U14279 (N_14279,N_8785,N_7292);
or U14280 (N_14280,N_1699,N_1880);
or U14281 (N_14281,N_9944,N_2508);
nand U14282 (N_14282,N_6929,N_3532);
nor U14283 (N_14283,N_6105,N_1701);
nor U14284 (N_14284,N_9919,N_3499);
and U14285 (N_14285,N_5411,N_6902);
nor U14286 (N_14286,N_1544,N_2388);
and U14287 (N_14287,N_9135,N_3464);
or U14288 (N_14288,N_8205,N_5755);
and U14289 (N_14289,N_3381,N_7749);
nor U14290 (N_14290,N_9871,N_3721);
and U14291 (N_14291,N_8298,N_7233);
and U14292 (N_14292,N_4990,N_8900);
and U14293 (N_14293,N_432,N_228);
and U14294 (N_14294,N_5804,N_3676);
nand U14295 (N_14295,N_5133,N_2142);
nor U14296 (N_14296,N_3102,N_5589);
nand U14297 (N_14297,N_4008,N_4856);
nor U14298 (N_14298,N_5659,N_4030);
or U14299 (N_14299,N_3761,N_3402);
and U14300 (N_14300,N_7220,N_4622);
nor U14301 (N_14301,N_3375,N_5217);
xor U14302 (N_14302,N_5979,N_5196);
or U14303 (N_14303,N_3398,N_1059);
or U14304 (N_14304,N_9395,N_7001);
and U14305 (N_14305,N_8940,N_812);
xnor U14306 (N_14306,N_4869,N_8237);
or U14307 (N_14307,N_6508,N_1776);
or U14308 (N_14308,N_2806,N_6723);
xnor U14309 (N_14309,N_2593,N_3187);
nand U14310 (N_14310,N_840,N_6088);
and U14311 (N_14311,N_9997,N_4650);
xor U14312 (N_14312,N_2368,N_9486);
and U14313 (N_14313,N_6620,N_4672);
or U14314 (N_14314,N_5613,N_5692);
nor U14315 (N_14315,N_8412,N_700);
or U14316 (N_14316,N_3621,N_3898);
nor U14317 (N_14317,N_6660,N_9873);
nand U14318 (N_14318,N_6365,N_1235);
nor U14319 (N_14319,N_2600,N_8873);
and U14320 (N_14320,N_2352,N_7318);
and U14321 (N_14321,N_4876,N_7214);
nand U14322 (N_14322,N_7030,N_6795);
and U14323 (N_14323,N_4767,N_1528);
or U14324 (N_14324,N_3322,N_1739);
or U14325 (N_14325,N_6956,N_2258);
and U14326 (N_14326,N_6143,N_8397);
and U14327 (N_14327,N_6475,N_1499);
or U14328 (N_14328,N_6598,N_7277);
nand U14329 (N_14329,N_3995,N_4805);
nor U14330 (N_14330,N_9061,N_6193);
or U14331 (N_14331,N_2830,N_8407);
or U14332 (N_14332,N_1062,N_1197);
nor U14333 (N_14333,N_3900,N_5643);
and U14334 (N_14334,N_5129,N_9256);
nor U14335 (N_14335,N_2652,N_7938);
or U14336 (N_14336,N_4140,N_829);
nor U14337 (N_14337,N_2807,N_7588);
nor U14338 (N_14338,N_3861,N_1121);
or U14339 (N_14339,N_8044,N_9927);
nand U14340 (N_14340,N_7069,N_8266);
and U14341 (N_14341,N_7455,N_3435);
nand U14342 (N_14342,N_9327,N_166);
and U14343 (N_14343,N_8281,N_1314);
nand U14344 (N_14344,N_4044,N_8845);
and U14345 (N_14345,N_3261,N_8525);
xnor U14346 (N_14346,N_908,N_6207);
and U14347 (N_14347,N_4479,N_4724);
or U14348 (N_14348,N_6099,N_3547);
nor U14349 (N_14349,N_2698,N_7462);
xnor U14350 (N_14350,N_3016,N_3658);
or U14351 (N_14351,N_5600,N_8764);
or U14352 (N_14352,N_1337,N_5299);
or U14353 (N_14353,N_303,N_192);
or U14354 (N_14354,N_1492,N_2493);
or U14355 (N_14355,N_1857,N_6079);
nand U14356 (N_14356,N_2278,N_2031);
nand U14357 (N_14357,N_7731,N_2924);
and U14358 (N_14358,N_5434,N_8460);
or U14359 (N_14359,N_5819,N_6014);
nand U14360 (N_14360,N_7322,N_7252);
nor U14361 (N_14361,N_5524,N_6625);
nor U14362 (N_14362,N_7950,N_4855);
and U14363 (N_14363,N_9672,N_7889);
or U14364 (N_14364,N_6125,N_1050);
or U14365 (N_14365,N_5635,N_9743);
nor U14366 (N_14366,N_1839,N_5518);
and U14367 (N_14367,N_4310,N_4956);
or U14368 (N_14368,N_7446,N_4538);
or U14369 (N_14369,N_3080,N_5148);
nand U14370 (N_14370,N_5287,N_16);
nor U14371 (N_14371,N_6364,N_3008);
or U14372 (N_14372,N_9826,N_8383);
xor U14373 (N_14373,N_3364,N_5697);
or U14374 (N_14374,N_1868,N_2948);
nor U14375 (N_14375,N_5508,N_4475);
or U14376 (N_14376,N_5144,N_4971);
and U14377 (N_14377,N_3748,N_2708);
or U14378 (N_14378,N_4000,N_7112);
nor U14379 (N_14379,N_4510,N_7825);
or U14380 (N_14380,N_8179,N_7910);
or U14381 (N_14381,N_6733,N_8918);
and U14382 (N_14382,N_5860,N_6851);
and U14383 (N_14383,N_5078,N_3156);
and U14384 (N_14384,N_1300,N_6697);
nand U14385 (N_14385,N_400,N_8722);
nand U14386 (N_14386,N_4271,N_3184);
nor U14387 (N_14387,N_6856,N_7246);
or U14388 (N_14388,N_1303,N_7546);
and U14389 (N_14389,N_8783,N_5756);
and U14390 (N_14390,N_1129,N_6339);
nand U14391 (N_14391,N_3674,N_9912);
nor U14392 (N_14392,N_4854,N_3226);
nand U14393 (N_14393,N_5336,N_4756);
nor U14394 (N_14394,N_9130,N_2750);
nor U14395 (N_14395,N_3569,N_5932);
nand U14396 (N_14396,N_1150,N_7750);
or U14397 (N_14397,N_6372,N_1972);
or U14398 (N_14398,N_9635,N_2026);
or U14399 (N_14399,N_7687,N_4691);
nand U14400 (N_14400,N_4980,N_4273);
or U14401 (N_14401,N_8013,N_2417);
and U14402 (N_14402,N_3208,N_7045);
nor U14403 (N_14403,N_3394,N_9750);
and U14404 (N_14404,N_7495,N_8592);
nor U14405 (N_14405,N_9269,N_4449);
and U14406 (N_14406,N_5638,N_4707);
or U14407 (N_14407,N_5419,N_123);
nor U14408 (N_14408,N_4364,N_7342);
and U14409 (N_14409,N_651,N_3233);
nand U14410 (N_14410,N_3438,N_9330);
nand U14411 (N_14411,N_8429,N_5726);
or U14412 (N_14412,N_7565,N_8219);
nor U14413 (N_14413,N_3949,N_8036);
nand U14414 (N_14414,N_124,N_9205);
and U14415 (N_14415,N_2459,N_3323);
or U14416 (N_14416,N_591,N_6185);
or U14417 (N_14417,N_9305,N_9844);
nor U14418 (N_14418,N_6550,N_8836);
xnor U14419 (N_14419,N_2994,N_4277);
nor U14420 (N_14420,N_4763,N_9408);
or U14421 (N_14421,N_3321,N_5352);
xnor U14422 (N_14422,N_364,N_2716);
or U14423 (N_14423,N_3329,N_4534);
and U14424 (N_14424,N_3502,N_6400);
nand U14425 (N_14425,N_8188,N_4181);
xnor U14426 (N_14426,N_1350,N_2574);
and U14427 (N_14427,N_2528,N_1188);
nor U14428 (N_14428,N_7529,N_920);
and U14429 (N_14429,N_8994,N_2581);
nand U14430 (N_14430,N_2802,N_73);
xnor U14431 (N_14431,N_3638,N_6162);
nand U14432 (N_14432,N_2219,N_3283);
and U14433 (N_14433,N_6189,N_8661);
or U14434 (N_14434,N_5228,N_5624);
and U14435 (N_14435,N_9450,N_9745);
xor U14436 (N_14436,N_6710,N_8379);
nand U14437 (N_14437,N_5785,N_6457);
xor U14438 (N_14438,N_8945,N_3060);
and U14439 (N_14439,N_9147,N_8514);
nor U14440 (N_14440,N_6619,N_441);
and U14441 (N_14441,N_9861,N_7037);
nand U14442 (N_14442,N_9646,N_2497);
or U14443 (N_14443,N_9557,N_3083);
or U14444 (N_14444,N_2304,N_6403);
nor U14445 (N_14445,N_4436,N_1000);
nand U14446 (N_14446,N_4274,N_9718);
or U14447 (N_14447,N_3074,N_1901);
and U14448 (N_14448,N_5801,N_6547);
nand U14449 (N_14449,N_2560,N_78);
or U14450 (N_14450,N_824,N_8866);
nor U14451 (N_14451,N_2880,N_426);
xnor U14452 (N_14452,N_7444,N_5645);
nand U14453 (N_14453,N_8711,N_3773);
or U14454 (N_14454,N_5025,N_3179);
or U14455 (N_14455,N_6763,N_9313);
nor U14456 (N_14456,N_6155,N_4191);
nand U14457 (N_14457,N_8366,N_4714);
xor U14458 (N_14458,N_1789,N_9209);
nor U14459 (N_14459,N_9103,N_6435);
nor U14460 (N_14460,N_9860,N_7751);
nand U14461 (N_14461,N_2601,N_4609);
nand U14462 (N_14462,N_9238,N_7789);
and U14463 (N_14463,N_8176,N_2439);
nor U14464 (N_14464,N_7346,N_9604);
nand U14465 (N_14465,N_5001,N_6513);
or U14466 (N_14466,N_6376,N_6597);
or U14467 (N_14467,N_38,N_6412);
and U14468 (N_14468,N_1199,N_8069);
and U14469 (N_14469,N_2584,N_6997);
nand U14470 (N_14470,N_3420,N_5056);
and U14471 (N_14471,N_7548,N_8395);
or U14472 (N_14472,N_2281,N_1694);
nor U14473 (N_14473,N_297,N_1623);
nor U14474 (N_14474,N_2344,N_8678);
nand U14475 (N_14475,N_2725,N_1312);
nor U14476 (N_14476,N_5722,N_8273);
and U14477 (N_14477,N_4874,N_1853);
xor U14478 (N_14478,N_7272,N_476);
nor U14479 (N_14479,N_6533,N_2311);
nand U14480 (N_14480,N_7411,N_1538);
and U14481 (N_14481,N_4915,N_5754);
or U14482 (N_14482,N_2744,N_5297);
or U14483 (N_14483,N_3,N_7497);
nor U14484 (N_14484,N_8939,N_20);
nor U14485 (N_14485,N_447,N_4233);
nand U14486 (N_14486,N_1646,N_2090);
and U14487 (N_14487,N_656,N_2790);
nor U14488 (N_14488,N_821,N_948);
or U14489 (N_14489,N_8365,N_8435);
or U14490 (N_14490,N_133,N_4114);
nor U14491 (N_14491,N_6998,N_4070);
nor U14492 (N_14492,N_2892,N_8040);
nand U14493 (N_14493,N_2462,N_8815);
nor U14494 (N_14494,N_912,N_5723);
nor U14495 (N_14495,N_4403,N_783);
xnor U14496 (N_14496,N_2005,N_6585);
xor U14497 (N_14497,N_2986,N_4504);
nand U14498 (N_14498,N_754,N_1323);
and U14499 (N_14499,N_6378,N_8738);
nand U14500 (N_14500,N_3351,N_1526);
and U14501 (N_14501,N_3219,N_4790);
or U14502 (N_14502,N_158,N_3980);
nand U14503 (N_14503,N_6677,N_3997);
nor U14504 (N_14504,N_2787,N_2789);
and U14505 (N_14505,N_6972,N_2195);
nor U14506 (N_14506,N_3751,N_3337);
and U14507 (N_14507,N_139,N_1095);
nand U14508 (N_14508,N_2687,N_7415);
nand U14509 (N_14509,N_3482,N_8323);
and U14510 (N_14510,N_6349,N_6549);
nor U14511 (N_14511,N_9201,N_962);
or U14512 (N_14512,N_5602,N_9189);
or U14513 (N_14513,N_3215,N_7668);
nor U14514 (N_14514,N_9036,N_8116);
or U14515 (N_14515,N_7475,N_5532);
xor U14516 (N_14516,N_4572,N_49);
nor U14517 (N_14517,N_1254,N_1277);
nand U14518 (N_14518,N_6742,N_6419);
xnor U14519 (N_14519,N_8283,N_2405);
nand U14520 (N_14520,N_5169,N_59);
and U14521 (N_14521,N_1893,N_7575);
or U14522 (N_14522,N_4161,N_112);
nor U14523 (N_14523,N_9112,N_5700);
nand U14524 (N_14524,N_6121,N_5628);
nor U14525 (N_14525,N_5053,N_4580);
nor U14526 (N_14526,N_558,N_7442);
and U14527 (N_14527,N_1991,N_4424);
nand U14528 (N_14528,N_4312,N_8779);
xnor U14529 (N_14529,N_910,N_8727);
nor U14530 (N_14530,N_9527,N_4033);
xnor U14531 (N_14531,N_7370,N_9624);
nor U14532 (N_14532,N_7538,N_4894);
and U14533 (N_14533,N_3178,N_6843);
or U14534 (N_14534,N_8263,N_6267);
or U14535 (N_14535,N_8706,N_7131);
and U14536 (N_14536,N_4527,N_8594);
or U14537 (N_14537,N_8596,N_5776);
nor U14538 (N_14538,N_7958,N_8935);
nor U14539 (N_14539,N_6307,N_1687);
nor U14540 (N_14540,N_4636,N_3720);
nor U14541 (N_14541,N_388,N_4567);
and U14542 (N_14542,N_5460,N_2061);
or U14543 (N_14543,N_461,N_5729);
or U14544 (N_14544,N_4067,N_7282);
xnor U14545 (N_14545,N_7427,N_5784);
nand U14546 (N_14546,N_6316,N_2795);
or U14547 (N_14547,N_613,N_1556);
and U14548 (N_14548,N_1106,N_7916);
or U14549 (N_14549,N_2378,N_7339);
or U14550 (N_14550,N_3200,N_4887);
or U14551 (N_14551,N_5393,N_1506);
or U14552 (N_14552,N_141,N_3792);
and U14553 (N_14553,N_4649,N_9108);
xor U14554 (N_14554,N_2236,N_4124);
or U14555 (N_14555,N_5272,N_9760);
or U14556 (N_14556,N_932,N_1117);
or U14557 (N_14557,N_3258,N_992);
nor U14558 (N_14558,N_6115,N_5449);
and U14559 (N_14559,N_4229,N_3094);
or U14560 (N_14560,N_9468,N_1848);
and U14561 (N_14561,N_8717,N_3029);
and U14562 (N_14562,N_4946,N_8513);
or U14563 (N_14563,N_4671,N_7783);
or U14564 (N_14564,N_2248,N_7317);
nor U14565 (N_14565,N_4133,N_1624);
and U14566 (N_14566,N_1084,N_9295);
and U14567 (N_14567,N_4060,N_8506);
nand U14568 (N_14568,N_6604,N_7798);
or U14569 (N_14569,N_8555,N_7730);
xor U14570 (N_14570,N_9303,N_999);
nor U14571 (N_14571,N_3839,N_3778);
and U14572 (N_14572,N_9916,N_8570);
or U14573 (N_14573,N_9508,N_730);
and U14574 (N_14574,N_9573,N_5491);
and U14575 (N_14575,N_3508,N_2878);
nand U14576 (N_14576,N_5112,N_3467);
nand U14577 (N_14577,N_1358,N_7580);
and U14578 (N_14578,N_4359,N_5409);
xor U14579 (N_14579,N_4089,N_5323);
nand U14580 (N_14580,N_8575,N_8332);
nor U14581 (N_14581,N_3883,N_6458);
and U14582 (N_14582,N_8538,N_5640);
or U14583 (N_14583,N_2285,N_5271);
and U14584 (N_14584,N_4328,N_6761);
or U14585 (N_14585,N_5771,N_3374);
nand U14586 (N_14586,N_1891,N_5621);
nand U14587 (N_14587,N_8212,N_6845);
nor U14588 (N_14588,N_7383,N_3691);
nand U14589 (N_14589,N_3706,N_9401);
nor U14590 (N_14590,N_6133,N_2758);
and U14591 (N_14591,N_7629,N_3138);
or U14592 (N_14592,N_8233,N_1787);
nand U14593 (N_14593,N_4276,N_5275);
nor U14594 (N_14594,N_5224,N_703);
or U14595 (N_14595,N_5107,N_2532);
nor U14596 (N_14596,N_6988,N_7134);
nor U14597 (N_14597,N_2571,N_8579);
nor U14598 (N_14598,N_5800,N_6154);
nor U14599 (N_14599,N_3632,N_6257);
or U14600 (N_14600,N_5753,N_2873);
or U14601 (N_14601,N_9281,N_5869);
or U14602 (N_14602,N_2189,N_9418);
nand U14603 (N_14603,N_5091,N_877);
nand U14604 (N_14604,N_4433,N_464);
nand U14605 (N_14605,N_7686,N_1958);
and U14606 (N_14606,N_3425,N_9710);
or U14607 (N_14607,N_3166,N_3479);
nand U14608 (N_14608,N_3370,N_206);
nand U14609 (N_14609,N_657,N_4250);
and U14610 (N_14610,N_2681,N_7505);
and U14611 (N_14611,N_1817,N_468);
nand U14612 (N_14612,N_6774,N_4109);
or U14613 (N_14613,N_4964,N_2122);
xor U14614 (N_14614,N_7204,N_2205);
nor U14615 (N_14615,N_8287,N_8760);
or U14616 (N_14616,N_2264,N_8665);
and U14617 (N_14617,N_7016,N_9932);
xor U14618 (N_14618,N_3582,N_4704);
or U14619 (N_14619,N_5984,N_4217);
nand U14620 (N_14620,N_8775,N_359);
nand U14621 (N_14621,N_4469,N_1440);
nand U14622 (N_14622,N_1266,N_390);
and U14623 (N_14623,N_8019,N_4575);
or U14624 (N_14624,N_9214,N_7210);
and U14625 (N_14625,N_5679,N_1965);
nor U14626 (N_14626,N_1252,N_937);
nor U14627 (N_14627,N_6021,N_5335);
and U14628 (N_14628,N_6627,N_9809);
or U14629 (N_14629,N_9937,N_7046);
xnor U14630 (N_14630,N_5916,N_9728);
and U14631 (N_14631,N_5615,N_4514);
and U14632 (N_14632,N_299,N_3390);
nor U14633 (N_14633,N_6026,N_9280);
or U14634 (N_14634,N_4640,N_9877);
nand U14635 (N_14635,N_5418,N_2612);
nor U14636 (N_14636,N_939,N_198);
and U14637 (N_14637,N_7228,N_6992);
nand U14638 (N_14638,N_7257,N_7835);
nor U14639 (N_14639,N_1567,N_9093);
or U14640 (N_14640,N_4552,N_7388);
xor U14641 (N_14641,N_723,N_8409);
and U14642 (N_14642,N_3282,N_4363);
nand U14643 (N_14643,N_9155,N_1375);
nand U14644 (N_14644,N_6816,N_6577);
nand U14645 (N_14645,N_9054,N_3358);
and U14646 (N_14646,N_6608,N_9755);
nor U14647 (N_14647,N_7254,N_39);
or U14648 (N_14648,N_9769,N_8517);
xor U14649 (N_14649,N_7918,N_1620);
nand U14650 (N_14650,N_6962,N_7301);
nand U14651 (N_14651,N_6368,N_1668);
and U14652 (N_14652,N_1876,N_248);
nand U14653 (N_14653,N_7693,N_1766);
nor U14654 (N_14654,N_9658,N_8280);
nand U14655 (N_14655,N_3522,N_252);
xor U14656 (N_14656,N_9693,N_3790);
nand U14657 (N_14657,N_9992,N_89);
or U14658 (N_14658,N_945,N_643);
and U14659 (N_14659,N_5675,N_7403);
nand U14660 (N_14660,N_9803,N_5567);
and U14661 (N_14661,N_5032,N_8084);
or U14662 (N_14662,N_4225,N_6025);
and U14663 (N_14663,N_5471,N_1497);
or U14664 (N_14664,N_413,N_8400);
xnor U14665 (N_14665,N_5504,N_6587);
nor U14666 (N_14666,N_3238,N_9905);
nor U14667 (N_14667,N_4642,N_361);
nand U14668 (N_14668,N_3743,N_6709);
nor U14669 (N_14669,N_201,N_9398);
nor U14670 (N_14670,N_8314,N_5489);
nor U14671 (N_14671,N_33,N_7815);
or U14672 (N_14672,N_6000,N_5751);
nor U14673 (N_14673,N_8649,N_9977);
nand U14674 (N_14674,N_6276,N_253);
nand U14675 (N_14675,N_6875,N_1232);
nand U14676 (N_14676,N_6868,N_4011);
xor U14677 (N_14677,N_3697,N_7977);
or U14678 (N_14678,N_5396,N_7138);
and U14679 (N_14679,N_7584,N_3027);
or U14680 (N_14680,N_446,N_5761);
xnor U14681 (N_14681,N_6588,N_538);
nor U14682 (N_14682,N_9237,N_6423);
nand U14683 (N_14683,N_5913,N_1940);
and U14684 (N_14684,N_312,N_8223);
nor U14685 (N_14685,N_8454,N_9051);
and U14686 (N_14686,N_8890,N_6705);
and U14687 (N_14687,N_6209,N_2014);
nand U14688 (N_14688,N_3945,N_975);
or U14689 (N_14689,N_4755,N_516);
xnor U14690 (N_14690,N_391,N_5055);
and U14691 (N_14691,N_6568,N_7532);
and U14692 (N_14692,N_7115,N_6380);
or U14693 (N_14693,N_2779,N_8719);
or U14694 (N_14694,N_1316,N_8861);
nand U14695 (N_14695,N_1378,N_6702);
nor U14696 (N_14696,N_9747,N_8464);
or U14697 (N_14697,N_22,N_557);
or U14698 (N_14698,N_4131,N_5308);
nand U14699 (N_14699,N_2820,N_1967);
or U14700 (N_14700,N_1187,N_8192);
or U14701 (N_14701,N_6404,N_7814);
nand U14702 (N_14702,N_9579,N_9680);
nor U14703 (N_14703,N_6981,N_4786);
or U14704 (N_14704,N_1745,N_1805);
and U14705 (N_14705,N_6975,N_5164);
nor U14706 (N_14706,N_1565,N_9578);
nand U14707 (N_14707,N_7459,N_6991);
or U14708 (N_14708,N_9948,N_4481);
nor U14709 (N_14709,N_1399,N_2366);
nand U14710 (N_14710,N_8126,N_1239);
nor U14711 (N_14711,N_2148,N_2490);
nor U14712 (N_14712,N_5975,N_4836);
and U14713 (N_14713,N_5510,N_3317);
nand U14714 (N_14714,N_5781,N_2507);
nor U14715 (N_14715,N_5686,N_1835);
nand U14716 (N_14716,N_2847,N_2100);
or U14717 (N_14717,N_4296,N_6024);
nor U14718 (N_14718,N_5724,N_6684);
and U14719 (N_14719,N_3035,N_1662);
nor U14720 (N_14720,N_5897,N_6798);
nor U14721 (N_14721,N_4004,N_6059);
nor U14722 (N_14722,N_1001,N_7520);
or U14723 (N_14723,N_9898,N_5871);
xnor U14724 (N_14724,N_8489,N_3684);
nor U14725 (N_14725,N_3796,N_485);
nand U14726 (N_14726,N_6149,N_7939);
and U14727 (N_14727,N_6330,N_8246);
or U14728 (N_14728,N_251,N_2859);
xor U14729 (N_14729,N_2550,N_7809);
nor U14730 (N_14730,N_3546,N_1820);
nand U14731 (N_14731,N_6787,N_2380);
and U14732 (N_14732,N_9626,N_5433);
and U14733 (N_14733,N_8088,N_3652);
or U14734 (N_14734,N_8540,N_8792);
xor U14735 (N_14735,N_7527,N_9095);
or U14736 (N_14736,N_5263,N_2785);
or U14737 (N_14737,N_9157,N_2536);
xnor U14738 (N_14738,N_4046,N_5374);
nor U14739 (N_14739,N_449,N_6164);
xor U14740 (N_14740,N_6194,N_9627);
nand U14741 (N_14741,N_7763,N_6114);
or U14742 (N_14742,N_378,N_608);
nor U14743 (N_14743,N_4019,N_7640);
and U14744 (N_14744,N_8128,N_3468);
or U14745 (N_14745,N_3023,N_5611);
or U14746 (N_14746,N_2978,N_1035);
nor U14747 (N_14747,N_8881,N_6259);
xnor U14748 (N_14748,N_704,N_7170);
nor U14749 (N_14749,N_2989,N_5122);
nand U14750 (N_14750,N_7936,N_7903);
nor U14751 (N_14751,N_7533,N_3259);
or U14752 (N_14752,N_8384,N_3580);
xor U14753 (N_14753,N_7759,N_9613);
xor U14754 (N_14754,N_1131,N_2693);
and U14755 (N_14755,N_226,N_8414);
nand U14756 (N_14756,N_5349,N_2137);
nor U14757 (N_14757,N_5702,N_6206);
nand U14758 (N_14758,N_7507,N_3543);
xnor U14759 (N_14759,N_1558,N_9889);
xor U14760 (N_14760,N_4466,N_3442);
and U14761 (N_14761,N_800,N_2721);
nor U14762 (N_14762,N_8471,N_4346);
nor U14763 (N_14763,N_5539,N_3093);
and U14764 (N_14764,N_4768,N_3592);
nand U14765 (N_14765,N_7095,N_3853);
and U14766 (N_14766,N_3086,N_219);
and U14767 (N_14767,N_892,N_5305);
nor U14768 (N_14768,N_6896,N_3460);
nor U14769 (N_14769,N_4850,N_9343);
and U14770 (N_14770,N_6522,N_1845);
nor U14771 (N_14771,N_4865,N_9210);
and U14772 (N_14772,N_1206,N_8539);
xor U14773 (N_14773,N_7352,N_4174);
and U14774 (N_14774,N_5839,N_905);
and U14775 (N_14775,N_4861,N_3256);
nand U14776 (N_14776,N_8521,N_2526);
or U14777 (N_14777,N_966,N_9910);
and U14778 (N_14778,N_4362,N_6488);
nor U14779 (N_14779,N_3512,N_2686);
or U14780 (N_14780,N_7288,N_5439);
nand U14781 (N_14781,N_2870,N_5085);
or U14782 (N_14782,N_6248,N_739);
or U14783 (N_14783,N_2576,N_8832);
xor U14784 (N_14784,N_4881,N_5484);
nand U14785 (N_14785,N_811,N_7684);
and U14786 (N_14786,N_3265,N_7706);
and U14787 (N_14787,N_2447,N_6355);
nor U14788 (N_14788,N_6665,N_3601);
xnor U14789 (N_14789,N_4451,N_3746);
nand U14790 (N_14790,N_2517,N_8993);
and U14791 (N_14791,N_4613,N_7473);
and U14792 (N_14792,N_9904,N_1537);
and U14793 (N_14793,N_2158,N_6943);
or U14794 (N_14794,N_8684,N_6326);
nor U14795 (N_14795,N_3914,N_7853);
and U14796 (N_14796,N_4458,N_1191);
nor U14797 (N_14797,N_8934,N_3801);
nor U14798 (N_14798,N_2088,N_9402);
or U14799 (N_14799,N_2384,N_3377);
nor U14800 (N_14800,N_9367,N_5307);
xnor U14801 (N_14801,N_1846,N_7647);
nand U14802 (N_14802,N_381,N_7080);
nand U14803 (N_14803,N_3501,N_4173);
and U14804 (N_14804,N_8632,N_450);
or U14805 (N_14805,N_4928,N_8470);
or U14806 (N_14806,N_697,N_3302);
or U14807 (N_14807,N_3197,N_8131);
nand U14808 (N_14808,N_7241,N_1793);
nand U14809 (N_14809,N_3755,N_7694);
xor U14810 (N_14810,N_2139,N_1933);
nor U14811 (N_14811,N_8511,N_3593);
or U14812 (N_14812,N_2823,N_8418);
nand U14813 (N_14813,N_965,N_6828);
or U14814 (N_14814,N_9565,N_3115);
or U14815 (N_14815,N_4585,N_7510);
nor U14816 (N_14816,N_4924,N_8342);
and U14817 (N_14817,N_7534,N_1228);
nand U14818 (N_14818,N_7275,N_654);
nor U14819 (N_14819,N_7582,N_7542);
xor U14820 (N_14820,N_1144,N_4421);
nand U14821 (N_14821,N_5968,N_1160);
nand U14822 (N_14822,N_445,N_9083);
and U14823 (N_14823,N_6622,N_3206);
or U14824 (N_14824,N_376,N_6986);
or U14825 (N_14825,N_8648,N_6788);
nand U14826 (N_14826,N_1479,N_8932);
xnor U14827 (N_14827,N_2817,N_5207);
nand U14828 (N_14828,N_6578,N_8747);
nor U14829 (N_14829,N_8759,N_3146);
nand U14830 (N_14830,N_5081,N_5958);
and U14831 (N_14831,N_6290,N_6917);
nor U14832 (N_14832,N_6800,N_8191);
and U14833 (N_14833,N_1923,N_50);
or U14834 (N_14834,N_6939,N_5861);
or U14835 (N_14835,N_8882,N_8765);
xnor U14836 (N_14836,N_6287,N_6371);
or U14837 (N_14837,N_4084,N_2427);
or U14838 (N_14838,N_3155,N_8755);
xnor U14839 (N_14839,N_2668,N_8428);
nor U14840 (N_14840,N_431,N_9221);
nor U14841 (N_14841,N_8905,N_3941);
nor U14842 (N_14842,N_8867,N_9174);
or U14843 (N_14843,N_5985,N_5234);
and U14844 (N_14844,N_2268,N_5646);
or U14845 (N_14845,N_1428,N_1355);
nor U14846 (N_14846,N_7191,N_9862);
and U14847 (N_14847,N_1051,N_7850);
nand U14848 (N_14848,N_3633,N_9476);
nor U14849 (N_14849,N_6068,N_7218);
nor U14850 (N_14850,N_5387,N_6234);
or U14851 (N_14851,N_8306,N_8354);
or U14852 (N_14852,N_6662,N_7819);
or U14853 (N_14853,N_8919,N_3749);
and U14854 (N_14854,N_3804,N_9531);
nand U14855 (N_14855,N_2858,N_3454);
nand U14856 (N_14856,N_5153,N_8626);
nor U14857 (N_14857,N_8038,N_2661);
or U14858 (N_14858,N_4081,N_1220);
nand U14859 (N_14859,N_6903,N_4218);
nand U14860 (N_14860,N_1217,N_5648);
nor U14861 (N_14861,N_8791,N_2089);
nor U14862 (N_14862,N_1161,N_4686);
nor U14863 (N_14863,N_5255,N_5231);
or U14864 (N_14864,N_281,N_6334);
nand U14865 (N_14865,N_9856,N_1407);
xor U14866 (N_14866,N_2119,N_5222);
or U14867 (N_14867,N_2723,N_1874);
and U14868 (N_14868,N_8411,N_7827);
nand U14869 (N_14869,N_3661,N_2343);
nand U14870 (N_14870,N_7060,N_1915);
nor U14871 (N_14871,N_475,N_1294);
nor U14872 (N_14872,N_7908,N_2041);
nor U14873 (N_14873,N_4727,N_8487);
nor U14874 (N_14874,N_1419,N_2369);
nand U14875 (N_14875,N_4028,N_42);
and U14876 (N_14876,N_9240,N_66);
and U14877 (N_14877,N_1486,N_813);
nor U14878 (N_14878,N_250,N_2393);
nor U14879 (N_14879,N_3369,N_4739);
nand U14880 (N_14880,N_348,N_8264);
or U14881 (N_14881,N_8374,N_3986);
nand U14882 (N_14882,N_689,N_6431);
and U14883 (N_14883,N_3006,N_7107);
or U14884 (N_14884,N_7972,N_1458);
nor U14885 (N_14885,N_1438,N_6037);
xor U14886 (N_14886,N_6751,N_6426);
or U14887 (N_14887,N_804,N_8614);
nand U14888 (N_14888,N_696,N_8065);
nand U14889 (N_14889,N_2206,N_4555);
nor U14890 (N_14890,N_5976,N_1015);
nand U14891 (N_14891,N_2598,N_5215);
nor U14892 (N_14892,N_574,N_729);
or U14893 (N_14893,N_9802,N_2259);
nor U14894 (N_14894,N_5005,N_5399);
and U14895 (N_14895,N_9715,N_6448);
nor U14896 (N_14896,N_3332,N_9066);
or U14897 (N_14897,N_4989,N_196);
nor U14898 (N_14898,N_6420,N_90);
or U14899 (N_14899,N_9168,N_9634);
nand U14900 (N_14900,N_6422,N_1887);
or U14901 (N_14901,N_3878,N_1153);
xnor U14902 (N_14902,N_9186,N_7151);
nand U14903 (N_14903,N_7934,N_8992);
xnor U14904 (N_14904,N_4798,N_8924);
and U14905 (N_14905,N_2599,N_7822);
or U14906 (N_14906,N_9618,N_7500);
nand U14907 (N_14907,N_3588,N_4752);
and U14908 (N_14908,N_6643,N_223);
nand U14909 (N_14909,N_1048,N_4911);
and U14910 (N_14910,N_7988,N_1122);
nand U14911 (N_14911,N_9711,N_8566);
and U14912 (N_14912,N_9392,N_9503);
and U14913 (N_14913,N_2800,N_5901);
xnor U14914 (N_14914,N_8347,N_9574);
nor U14915 (N_14915,N_1484,N_2838);
and U14916 (N_14916,N_741,N_2180);
and U14917 (N_14917,N_4396,N_3758);
and U14918 (N_14918,N_9386,N_9216);
or U14919 (N_14919,N_4860,N_6050);
nor U14920 (N_14920,N_1885,N_9629);
and U14921 (N_14921,N_6960,N_7564);
xor U14922 (N_14922,N_2465,N_7447);
or U14923 (N_14923,N_7725,N_7488);
and U14924 (N_14924,N_3033,N_8954);
nor U14925 (N_14925,N_1068,N_2973);
and U14926 (N_14926,N_8368,N_3098);
nor U14927 (N_14927,N_7408,N_5931);
nand U14928 (N_14928,N_8937,N_8393);
and U14929 (N_14929,N_2239,N_6680);
nor U14930 (N_14930,N_7087,N_2428);
xor U14931 (N_14931,N_9831,N_1751);
nor U14932 (N_14932,N_3062,N_4447);
nand U14933 (N_14933,N_3153,N_7810);
nand U14934 (N_14934,N_5468,N_2096);
and U14935 (N_14935,N_7703,N_1877);
and U14936 (N_14936,N_9795,N_473);
nor U14937 (N_14937,N_3870,N_463);
or U14938 (N_14938,N_5676,N_425);
or U14939 (N_14939,N_7959,N_3998);
and U14940 (N_14940,N_2649,N_9162);
and U14941 (N_14941,N_170,N_9169);
xor U14942 (N_14942,N_1242,N_9321);
xor U14943 (N_14943,N_725,N_2181);
nor U14944 (N_14944,N_1904,N_9953);
nand U14945 (N_14945,N_1123,N_1875);
or U14946 (N_14946,N_4434,N_8692);
nand U14947 (N_14947,N_326,N_3181);
nor U14948 (N_14948,N_6439,N_2207);
and U14949 (N_14949,N_3875,N_1116);
and U14950 (N_14950,N_8801,N_6523);
nand U14951 (N_14951,N_2348,N_5227);
nor U14952 (N_14952,N_4559,N_6036);
and U14953 (N_14953,N_5940,N_2390);
xnor U14954 (N_14954,N_2594,N_6215);
or U14955 (N_14955,N_4068,N_6440);
and U14956 (N_14956,N_6540,N_2015);
or U14957 (N_14957,N_5810,N_2469);
or U14958 (N_14958,N_3814,N_7033);
xnor U14959 (N_14959,N_4778,N_4548);
xor U14960 (N_14960,N_5887,N_3620);
nand U14961 (N_14961,N_3171,N_1379);
and U14962 (N_14962,N_3873,N_2819);
nand U14963 (N_14963,N_5037,N_3014);
and U14964 (N_14964,N_2567,N_6538);
nor U14965 (N_14965,N_3882,N_7581);
xor U14966 (N_14966,N_4795,N_2323);
nand U14967 (N_14967,N_9591,N_1104);
xnor U14968 (N_14968,N_6434,N_7746);
nand U14969 (N_14969,N_8245,N_7600);
xor U14970 (N_14970,N_6729,N_3656);
or U14971 (N_14971,N_5816,N_9621);
xor U14972 (N_14972,N_8232,N_3005);
nand U14973 (N_14973,N_9971,N_4204);
nand U14974 (N_14974,N_3832,N_4485);
nand U14975 (N_14975,N_9906,N_9379);
nor U14976 (N_14976,N_4344,N_561);
nor U14977 (N_14977,N_4001,N_8465);
nand U14978 (N_14978,N_7326,N_5303);
nand U14979 (N_14979,N_4047,N_7754);
nor U14980 (N_14980,N_6367,N_4974);
nor U14981 (N_14981,N_661,N_4952);
nand U14982 (N_14982,N_9098,N_7563);
nand U14983 (N_14983,N_3116,N_6805);
or U14984 (N_14984,N_4234,N_4390);
and U14985 (N_14985,N_3055,N_1348);
and U14986 (N_14986,N_815,N_3404);
or U14987 (N_14987,N_7558,N_1236);
xnor U14988 (N_14988,N_7498,N_7293);
and U14989 (N_14989,N_477,N_4910);
nand U14990 (N_14990,N_7351,N_8239);
or U14991 (N_14991,N_4606,N_950);
or U14992 (N_14992,N_632,N_5364);
and U14993 (N_14993,N_3243,N_4224);
nor U14994 (N_14994,N_9451,N_4549);
nor U14995 (N_14995,N_3893,N_7550);
or U14996 (N_14996,N_4863,N_1756);
nand U14997 (N_14997,N_2553,N_2987);
nor U14998 (N_14998,N_6844,N_4152);
or U14999 (N_14999,N_4119,N_7286);
nor U15000 (N_15000,N_1885,N_5240);
and U15001 (N_15001,N_4566,N_3017);
or U15002 (N_15002,N_2580,N_9079);
nand U15003 (N_15003,N_2918,N_89);
and U15004 (N_15004,N_8476,N_9175);
and U15005 (N_15005,N_2572,N_4096);
xnor U15006 (N_15006,N_2288,N_3017);
xnor U15007 (N_15007,N_1029,N_8942);
and U15008 (N_15008,N_4384,N_3433);
nor U15009 (N_15009,N_2337,N_5308);
and U15010 (N_15010,N_1329,N_4912);
nand U15011 (N_15011,N_2121,N_4328);
or U15012 (N_15012,N_6743,N_5113);
xor U15013 (N_15013,N_7890,N_7869);
or U15014 (N_15014,N_5727,N_4899);
nand U15015 (N_15015,N_4613,N_284);
xor U15016 (N_15016,N_5615,N_83);
nand U15017 (N_15017,N_8110,N_810);
nor U15018 (N_15018,N_7612,N_5953);
nor U15019 (N_15019,N_3910,N_4342);
nor U15020 (N_15020,N_3524,N_4006);
nand U15021 (N_15021,N_4634,N_5001);
nor U15022 (N_15022,N_4647,N_8917);
and U15023 (N_15023,N_6492,N_6053);
nand U15024 (N_15024,N_9262,N_9336);
xnor U15025 (N_15025,N_3609,N_22);
nand U15026 (N_15026,N_4670,N_7369);
or U15027 (N_15027,N_5338,N_223);
or U15028 (N_15028,N_8732,N_663);
nor U15029 (N_15029,N_2516,N_3238);
xor U15030 (N_15030,N_258,N_7395);
and U15031 (N_15031,N_5239,N_7301);
and U15032 (N_15032,N_4538,N_459);
nand U15033 (N_15033,N_2062,N_5166);
nand U15034 (N_15034,N_4885,N_1201);
nor U15035 (N_15035,N_4242,N_1506);
and U15036 (N_15036,N_6009,N_4341);
or U15037 (N_15037,N_1752,N_5288);
xnor U15038 (N_15038,N_7641,N_7299);
and U15039 (N_15039,N_7552,N_5222);
nor U15040 (N_15040,N_6903,N_4252);
or U15041 (N_15041,N_247,N_1352);
or U15042 (N_15042,N_7783,N_6130);
and U15043 (N_15043,N_5997,N_8738);
nand U15044 (N_15044,N_1208,N_3374);
or U15045 (N_15045,N_2686,N_8894);
nor U15046 (N_15046,N_1845,N_2091);
nor U15047 (N_15047,N_7542,N_4576);
and U15048 (N_15048,N_5643,N_753);
nand U15049 (N_15049,N_1876,N_5326);
xnor U15050 (N_15050,N_5135,N_7262);
and U15051 (N_15051,N_1355,N_7595);
nor U15052 (N_15052,N_5903,N_4322);
or U15053 (N_15053,N_3081,N_7649);
nand U15054 (N_15054,N_6359,N_7483);
or U15055 (N_15055,N_2619,N_1875);
or U15056 (N_15056,N_3710,N_8782);
nor U15057 (N_15057,N_1078,N_9413);
or U15058 (N_15058,N_6981,N_5286);
and U15059 (N_15059,N_7720,N_5132);
or U15060 (N_15060,N_7137,N_6938);
nand U15061 (N_15061,N_5704,N_7509);
and U15062 (N_15062,N_4663,N_863);
nand U15063 (N_15063,N_2565,N_8406);
or U15064 (N_15064,N_6083,N_9946);
or U15065 (N_15065,N_9703,N_3753);
and U15066 (N_15066,N_4300,N_8312);
nand U15067 (N_15067,N_5099,N_4763);
nand U15068 (N_15068,N_3095,N_8043);
xnor U15069 (N_15069,N_6532,N_5508);
and U15070 (N_15070,N_7046,N_5920);
nand U15071 (N_15071,N_3442,N_4885);
nor U15072 (N_15072,N_45,N_1476);
and U15073 (N_15073,N_2514,N_21);
and U15074 (N_15074,N_6956,N_1533);
nor U15075 (N_15075,N_6421,N_7502);
nor U15076 (N_15076,N_9848,N_869);
nor U15077 (N_15077,N_5577,N_9612);
nor U15078 (N_15078,N_1538,N_6845);
nor U15079 (N_15079,N_7100,N_3274);
nand U15080 (N_15080,N_8214,N_2622);
and U15081 (N_15081,N_4920,N_6296);
nor U15082 (N_15082,N_7526,N_4463);
or U15083 (N_15083,N_6596,N_6289);
xor U15084 (N_15084,N_2724,N_2699);
nor U15085 (N_15085,N_1548,N_8609);
nor U15086 (N_15086,N_2120,N_6567);
and U15087 (N_15087,N_1265,N_1370);
nor U15088 (N_15088,N_4466,N_7187);
and U15089 (N_15089,N_4683,N_5741);
and U15090 (N_15090,N_4411,N_8959);
nor U15091 (N_15091,N_6367,N_3078);
xor U15092 (N_15092,N_4991,N_8497);
or U15093 (N_15093,N_1606,N_8816);
nor U15094 (N_15094,N_6687,N_7192);
or U15095 (N_15095,N_65,N_1340);
or U15096 (N_15096,N_9521,N_8285);
nand U15097 (N_15097,N_9178,N_8873);
nand U15098 (N_15098,N_5819,N_5705);
and U15099 (N_15099,N_267,N_276);
and U15100 (N_15100,N_1472,N_3179);
xor U15101 (N_15101,N_1247,N_9281);
or U15102 (N_15102,N_9185,N_6696);
or U15103 (N_15103,N_2068,N_5323);
nand U15104 (N_15104,N_3324,N_3984);
and U15105 (N_15105,N_6447,N_6369);
xnor U15106 (N_15106,N_4570,N_6320);
xor U15107 (N_15107,N_1007,N_1939);
or U15108 (N_15108,N_7836,N_5485);
nand U15109 (N_15109,N_2640,N_1031);
or U15110 (N_15110,N_3159,N_7129);
or U15111 (N_15111,N_1602,N_8226);
xnor U15112 (N_15112,N_1289,N_3338);
xnor U15113 (N_15113,N_455,N_5479);
and U15114 (N_15114,N_3920,N_9067);
nand U15115 (N_15115,N_9993,N_2741);
nor U15116 (N_15116,N_2632,N_6763);
nand U15117 (N_15117,N_4182,N_3841);
or U15118 (N_15118,N_9014,N_5269);
nand U15119 (N_15119,N_6517,N_7829);
nand U15120 (N_15120,N_9386,N_362);
or U15121 (N_15121,N_3684,N_2004);
nor U15122 (N_15122,N_4030,N_3644);
nor U15123 (N_15123,N_5525,N_2052);
or U15124 (N_15124,N_9555,N_3614);
nor U15125 (N_15125,N_6010,N_2079);
nand U15126 (N_15126,N_1990,N_5139);
nor U15127 (N_15127,N_1810,N_2686);
and U15128 (N_15128,N_5520,N_7595);
nor U15129 (N_15129,N_7789,N_7490);
nand U15130 (N_15130,N_9621,N_5213);
xnor U15131 (N_15131,N_2591,N_752);
xnor U15132 (N_15132,N_3398,N_9471);
nor U15133 (N_15133,N_3357,N_3783);
and U15134 (N_15134,N_4808,N_5858);
or U15135 (N_15135,N_364,N_4901);
or U15136 (N_15136,N_9266,N_238);
nor U15137 (N_15137,N_7445,N_4200);
xor U15138 (N_15138,N_1048,N_1450);
nor U15139 (N_15139,N_9971,N_6981);
nor U15140 (N_15140,N_9368,N_8853);
xnor U15141 (N_15141,N_1015,N_1361);
xor U15142 (N_15142,N_7696,N_3447);
or U15143 (N_15143,N_3327,N_8015);
nand U15144 (N_15144,N_543,N_2945);
and U15145 (N_15145,N_704,N_3237);
xnor U15146 (N_15146,N_3668,N_4306);
and U15147 (N_15147,N_3878,N_6942);
nor U15148 (N_15148,N_4658,N_1820);
and U15149 (N_15149,N_5444,N_124);
nor U15150 (N_15150,N_7123,N_7997);
and U15151 (N_15151,N_9120,N_1474);
nor U15152 (N_15152,N_478,N_5428);
nor U15153 (N_15153,N_8455,N_2049);
or U15154 (N_15154,N_1144,N_6698);
nor U15155 (N_15155,N_3307,N_6387);
nand U15156 (N_15156,N_9222,N_2885);
and U15157 (N_15157,N_58,N_2207);
or U15158 (N_15158,N_2220,N_5807);
xnor U15159 (N_15159,N_8001,N_1313);
nand U15160 (N_15160,N_1502,N_5088);
nor U15161 (N_15161,N_974,N_83);
nand U15162 (N_15162,N_3753,N_5347);
and U15163 (N_15163,N_7601,N_6594);
nand U15164 (N_15164,N_3939,N_3098);
nand U15165 (N_15165,N_1758,N_6834);
or U15166 (N_15166,N_6259,N_9334);
and U15167 (N_15167,N_1441,N_5783);
nand U15168 (N_15168,N_3356,N_1625);
xor U15169 (N_15169,N_1479,N_8387);
nor U15170 (N_15170,N_3892,N_7839);
nor U15171 (N_15171,N_4955,N_1858);
nor U15172 (N_15172,N_8013,N_6283);
nand U15173 (N_15173,N_6653,N_575);
and U15174 (N_15174,N_6987,N_3029);
or U15175 (N_15175,N_1196,N_3822);
and U15176 (N_15176,N_3766,N_7115);
nand U15177 (N_15177,N_3983,N_2029);
nor U15178 (N_15178,N_3489,N_8074);
and U15179 (N_15179,N_2766,N_841);
nand U15180 (N_15180,N_3899,N_326);
or U15181 (N_15181,N_1423,N_5716);
nand U15182 (N_15182,N_3200,N_2132);
and U15183 (N_15183,N_5205,N_460);
or U15184 (N_15184,N_9394,N_3414);
nor U15185 (N_15185,N_7165,N_9655);
and U15186 (N_15186,N_5416,N_3713);
xor U15187 (N_15187,N_2791,N_3697);
and U15188 (N_15188,N_8585,N_4921);
or U15189 (N_15189,N_3562,N_2222);
nor U15190 (N_15190,N_3392,N_4279);
nor U15191 (N_15191,N_7429,N_7967);
xnor U15192 (N_15192,N_3157,N_1564);
nand U15193 (N_15193,N_6233,N_152);
and U15194 (N_15194,N_4325,N_4803);
nand U15195 (N_15195,N_6071,N_2608);
and U15196 (N_15196,N_8208,N_780);
or U15197 (N_15197,N_5425,N_6981);
nor U15198 (N_15198,N_8334,N_2459);
and U15199 (N_15199,N_2302,N_9274);
nand U15200 (N_15200,N_1035,N_7458);
nor U15201 (N_15201,N_4669,N_499);
and U15202 (N_15202,N_7123,N_7910);
and U15203 (N_15203,N_4311,N_3968);
and U15204 (N_15204,N_5330,N_6039);
or U15205 (N_15205,N_1857,N_6184);
nand U15206 (N_15206,N_5814,N_3132);
or U15207 (N_15207,N_7320,N_8917);
xnor U15208 (N_15208,N_2960,N_2503);
nor U15209 (N_15209,N_3456,N_9985);
xor U15210 (N_15210,N_9864,N_4751);
nand U15211 (N_15211,N_1907,N_5775);
or U15212 (N_15212,N_7830,N_2150);
or U15213 (N_15213,N_8857,N_6661);
or U15214 (N_15214,N_6165,N_8851);
nand U15215 (N_15215,N_7626,N_5669);
nor U15216 (N_15216,N_3515,N_7518);
nand U15217 (N_15217,N_4901,N_6177);
nor U15218 (N_15218,N_634,N_6031);
xnor U15219 (N_15219,N_5034,N_4172);
xnor U15220 (N_15220,N_4137,N_3230);
and U15221 (N_15221,N_7383,N_2403);
nand U15222 (N_15222,N_2291,N_177);
nor U15223 (N_15223,N_9201,N_5650);
nor U15224 (N_15224,N_1966,N_7990);
or U15225 (N_15225,N_8343,N_388);
nand U15226 (N_15226,N_3629,N_6179);
and U15227 (N_15227,N_6400,N_8919);
or U15228 (N_15228,N_9577,N_8343);
and U15229 (N_15229,N_5577,N_9348);
nand U15230 (N_15230,N_5295,N_4188);
or U15231 (N_15231,N_9841,N_2013);
nand U15232 (N_15232,N_5631,N_2573);
and U15233 (N_15233,N_7338,N_2598);
nor U15234 (N_15234,N_3255,N_5672);
nor U15235 (N_15235,N_6537,N_817);
or U15236 (N_15236,N_9517,N_4428);
nor U15237 (N_15237,N_8298,N_2311);
xnor U15238 (N_15238,N_6232,N_8773);
xor U15239 (N_15239,N_3017,N_8941);
and U15240 (N_15240,N_4353,N_3001);
or U15241 (N_15241,N_678,N_7097);
or U15242 (N_15242,N_7408,N_9688);
or U15243 (N_15243,N_6805,N_3383);
or U15244 (N_15244,N_1839,N_404);
or U15245 (N_15245,N_5431,N_9771);
and U15246 (N_15246,N_1799,N_1);
or U15247 (N_15247,N_3184,N_2628);
or U15248 (N_15248,N_1437,N_9255);
nand U15249 (N_15249,N_4492,N_741);
and U15250 (N_15250,N_4436,N_6825);
and U15251 (N_15251,N_1475,N_6752);
and U15252 (N_15252,N_7260,N_9188);
nor U15253 (N_15253,N_4782,N_694);
and U15254 (N_15254,N_4976,N_848);
nor U15255 (N_15255,N_8997,N_9536);
nor U15256 (N_15256,N_6415,N_8439);
or U15257 (N_15257,N_31,N_2640);
or U15258 (N_15258,N_2173,N_5721);
and U15259 (N_15259,N_6360,N_8123);
xor U15260 (N_15260,N_246,N_6639);
and U15261 (N_15261,N_44,N_8820);
or U15262 (N_15262,N_7485,N_4100);
and U15263 (N_15263,N_1705,N_4361);
nor U15264 (N_15264,N_4575,N_3779);
xor U15265 (N_15265,N_1714,N_1265);
nor U15266 (N_15266,N_9051,N_9825);
nor U15267 (N_15267,N_3005,N_6789);
or U15268 (N_15268,N_9769,N_6699);
nor U15269 (N_15269,N_4370,N_5040);
and U15270 (N_15270,N_6005,N_9117);
nand U15271 (N_15271,N_5411,N_5797);
nand U15272 (N_15272,N_3069,N_2887);
and U15273 (N_15273,N_9979,N_5434);
and U15274 (N_15274,N_4089,N_4553);
or U15275 (N_15275,N_8303,N_1676);
or U15276 (N_15276,N_4085,N_6113);
nand U15277 (N_15277,N_1290,N_7986);
or U15278 (N_15278,N_5736,N_8730);
or U15279 (N_15279,N_6252,N_3806);
or U15280 (N_15280,N_2169,N_2186);
nand U15281 (N_15281,N_283,N_7748);
or U15282 (N_15282,N_8978,N_7895);
nor U15283 (N_15283,N_7803,N_7943);
or U15284 (N_15284,N_3099,N_6133);
nor U15285 (N_15285,N_3410,N_1794);
xor U15286 (N_15286,N_562,N_4383);
and U15287 (N_15287,N_9549,N_2795);
nor U15288 (N_15288,N_3426,N_6025);
nand U15289 (N_15289,N_7720,N_233);
nand U15290 (N_15290,N_7589,N_1800);
nand U15291 (N_15291,N_1867,N_9639);
and U15292 (N_15292,N_1636,N_6578);
and U15293 (N_15293,N_3020,N_4051);
nor U15294 (N_15294,N_8678,N_7270);
nor U15295 (N_15295,N_2472,N_9012);
nor U15296 (N_15296,N_2880,N_7141);
xor U15297 (N_15297,N_351,N_8695);
or U15298 (N_15298,N_9703,N_4376);
nand U15299 (N_15299,N_1515,N_2302);
or U15300 (N_15300,N_9144,N_8144);
or U15301 (N_15301,N_240,N_5311);
nand U15302 (N_15302,N_876,N_9138);
xor U15303 (N_15303,N_6071,N_8149);
xor U15304 (N_15304,N_8946,N_5932);
nor U15305 (N_15305,N_7664,N_1551);
or U15306 (N_15306,N_9858,N_4759);
nand U15307 (N_15307,N_3820,N_3032);
or U15308 (N_15308,N_63,N_7326);
nor U15309 (N_15309,N_5562,N_8051);
nor U15310 (N_15310,N_8481,N_7618);
and U15311 (N_15311,N_7306,N_9689);
or U15312 (N_15312,N_1049,N_2466);
nand U15313 (N_15313,N_6211,N_4685);
nand U15314 (N_15314,N_6126,N_763);
and U15315 (N_15315,N_9259,N_1804);
or U15316 (N_15316,N_7302,N_5594);
nor U15317 (N_15317,N_8079,N_1454);
and U15318 (N_15318,N_4572,N_7419);
xor U15319 (N_15319,N_5425,N_1514);
and U15320 (N_15320,N_6578,N_422);
nor U15321 (N_15321,N_8709,N_9812);
and U15322 (N_15322,N_5197,N_8427);
nor U15323 (N_15323,N_2657,N_1529);
xnor U15324 (N_15324,N_3702,N_5967);
and U15325 (N_15325,N_8171,N_1082);
or U15326 (N_15326,N_7202,N_3815);
and U15327 (N_15327,N_7818,N_6596);
and U15328 (N_15328,N_9787,N_3663);
and U15329 (N_15329,N_6645,N_6063);
and U15330 (N_15330,N_5406,N_8364);
nand U15331 (N_15331,N_8699,N_3916);
nor U15332 (N_15332,N_3999,N_8730);
nand U15333 (N_15333,N_8918,N_171);
or U15334 (N_15334,N_3450,N_4227);
nor U15335 (N_15335,N_1970,N_6126);
and U15336 (N_15336,N_6108,N_8807);
xor U15337 (N_15337,N_8739,N_3524);
nor U15338 (N_15338,N_7716,N_1158);
xor U15339 (N_15339,N_4150,N_8541);
nor U15340 (N_15340,N_5013,N_8696);
xnor U15341 (N_15341,N_1926,N_3444);
or U15342 (N_15342,N_806,N_8309);
and U15343 (N_15343,N_4954,N_9910);
or U15344 (N_15344,N_4109,N_2377);
or U15345 (N_15345,N_9015,N_1384);
nand U15346 (N_15346,N_5734,N_6454);
and U15347 (N_15347,N_775,N_9933);
or U15348 (N_15348,N_6043,N_880);
nor U15349 (N_15349,N_7445,N_1591);
nor U15350 (N_15350,N_7696,N_6598);
and U15351 (N_15351,N_6622,N_4581);
or U15352 (N_15352,N_8233,N_7014);
nand U15353 (N_15353,N_5798,N_5035);
nor U15354 (N_15354,N_5,N_4407);
xor U15355 (N_15355,N_1593,N_2309);
and U15356 (N_15356,N_2473,N_5220);
nand U15357 (N_15357,N_856,N_8471);
and U15358 (N_15358,N_2838,N_5387);
or U15359 (N_15359,N_8612,N_4153);
and U15360 (N_15360,N_1819,N_1212);
nor U15361 (N_15361,N_4629,N_512);
or U15362 (N_15362,N_4718,N_9607);
and U15363 (N_15363,N_7281,N_1887);
nand U15364 (N_15364,N_2570,N_4536);
nor U15365 (N_15365,N_2386,N_4038);
or U15366 (N_15366,N_3954,N_2029);
xnor U15367 (N_15367,N_7723,N_7310);
or U15368 (N_15368,N_4066,N_5334);
nand U15369 (N_15369,N_7094,N_9454);
and U15370 (N_15370,N_9688,N_1771);
nor U15371 (N_15371,N_6579,N_7290);
nand U15372 (N_15372,N_6760,N_4491);
and U15373 (N_15373,N_8719,N_1764);
and U15374 (N_15374,N_4862,N_3410);
nand U15375 (N_15375,N_2782,N_1872);
nand U15376 (N_15376,N_7857,N_4620);
and U15377 (N_15377,N_4780,N_5475);
and U15378 (N_15378,N_5472,N_1283);
nor U15379 (N_15379,N_7514,N_4490);
nand U15380 (N_15380,N_9613,N_9435);
nand U15381 (N_15381,N_6036,N_6311);
xnor U15382 (N_15382,N_5716,N_6767);
or U15383 (N_15383,N_5219,N_624);
nand U15384 (N_15384,N_355,N_9550);
or U15385 (N_15385,N_9066,N_3807);
nor U15386 (N_15386,N_3941,N_696);
or U15387 (N_15387,N_4079,N_2337);
xor U15388 (N_15388,N_6450,N_4191);
and U15389 (N_15389,N_6132,N_62);
nor U15390 (N_15390,N_7585,N_6587);
nor U15391 (N_15391,N_4891,N_7083);
nand U15392 (N_15392,N_6453,N_248);
nor U15393 (N_15393,N_3164,N_8470);
or U15394 (N_15394,N_1266,N_5814);
and U15395 (N_15395,N_6731,N_5686);
or U15396 (N_15396,N_5980,N_8919);
nor U15397 (N_15397,N_1228,N_9259);
nand U15398 (N_15398,N_6949,N_9342);
nand U15399 (N_15399,N_2439,N_2657);
or U15400 (N_15400,N_7454,N_6717);
or U15401 (N_15401,N_4809,N_7444);
nand U15402 (N_15402,N_4537,N_5102);
and U15403 (N_15403,N_2949,N_658);
nor U15404 (N_15404,N_506,N_2465);
nor U15405 (N_15405,N_4588,N_2662);
and U15406 (N_15406,N_9700,N_928);
and U15407 (N_15407,N_9678,N_7230);
or U15408 (N_15408,N_5993,N_2565);
or U15409 (N_15409,N_1968,N_5031);
nor U15410 (N_15410,N_1582,N_773);
xnor U15411 (N_15411,N_2879,N_1209);
or U15412 (N_15412,N_680,N_9696);
or U15413 (N_15413,N_1549,N_7039);
and U15414 (N_15414,N_7073,N_5760);
nor U15415 (N_15415,N_2659,N_1315);
nor U15416 (N_15416,N_4720,N_347);
and U15417 (N_15417,N_4295,N_1560);
nand U15418 (N_15418,N_2139,N_7601);
nand U15419 (N_15419,N_7459,N_1901);
xnor U15420 (N_15420,N_6533,N_1965);
and U15421 (N_15421,N_4981,N_1146);
or U15422 (N_15422,N_1645,N_7634);
nor U15423 (N_15423,N_881,N_5161);
and U15424 (N_15424,N_7337,N_662);
nand U15425 (N_15425,N_6597,N_1056);
or U15426 (N_15426,N_234,N_9509);
or U15427 (N_15427,N_7833,N_7362);
nor U15428 (N_15428,N_7043,N_8156);
or U15429 (N_15429,N_7425,N_2296);
nand U15430 (N_15430,N_9349,N_2383);
or U15431 (N_15431,N_1724,N_1861);
xor U15432 (N_15432,N_8982,N_5209);
xnor U15433 (N_15433,N_17,N_3770);
and U15434 (N_15434,N_9483,N_7735);
nand U15435 (N_15435,N_6181,N_184);
or U15436 (N_15436,N_4681,N_636);
and U15437 (N_15437,N_4127,N_9596);
nand U15438 (N_15438,N_445,N_2337);
or U15439 (N_15439,N_7313,N_411);
xnor U15440 (N_15440,N_8036,N_7801);
or U15441 (N_15441,N_8463,N_640);
nand U15442 (N_15442,N_5643,N_9931);
nor U15443 (N_15443,N_4149,N_2204);
or U15444 (N_15444,N_1775,N_8854);
and U15445 (N_15445,N_833,N_5854);
nand U15446 (N_15446,N_824,N_5670);
nor U15447 (N_15447,N_2068,N_3692);
xnor U15448 (N_15448,N_2706,N_9231);
nor U15449 (N_15449,N_9482,N_1690);
nand U15450 (N_15450,N_1013,N_9351);
nand U15451 (N_15451,N_3620,N_7670);
and U15452 (N_15452,N_167,N_8886);
nor U15453 (N_15453,N_3867,N_2040);
nor U15454 (N_15454,N_6474,N_8295);
and U15455 (N_15455,N_3058,N_561);
nand U15456 (N_15456,N_5996,N_2220);
and U15457 (N_15457,N_6599,N_1289);
nand U15458 (N_15458,N_6386,N_6592);
or U15459 (N_15459,N_8616,N_1471);
and U15460 (N_15460,N_9010,N_8352);
nor U15461 (N_15461,N_903,N_417);
nand U15462 (N_15462,N_2260,N_4240);
or U15463 (N_15463,N_7655,N_3341);
nand U15464 (N_15464,N_2935,N_3711);
nor U15465 (N_15465,N_7050,N_3995);
nor U15466 (N_15466,N_4749,N_3687);
or U15467 (N_15467,N_4699,N_651);
nand U15468 (N_15468,N_318,N_6370);
xor U15469 (N_15469,N_618,N_8286);
xor U15470 (N_15470,N_1890,N_9305);
and U15471 (N_15471,N_4914,N_2144);
or U15472 (N_15472,N_3344,N_9299);
nand U15473 (N_15473,N_3656,N_6379);
and U15474 (N_15474,N_6090,N_2826);
and U15475 (N_15475,N_8575,N_7765);
nor U15476 (N_15476,N_1074,N_4359);
xnor U15477 (N_15477,N_5206,N_9335);
nand U15478 (N_15478,N_3275,N_4875);
and U15479 (N_15479,N_4828,N_9878);
or U15480 (N_15480,N_304,N_5609);
or U15481 (N_15481,N_1578,N_4136);
nand U15482 (N_15482,N_8264,N_6504);
and U15483 (N_15483,N_6269,N_3422);
or U15484 (N_15484,N_1192,N_2636);
nand U15485 (N_15485,N_7761,N_3013);
nand U15486 (N_15486,N_1783,N_9153);
nor U15487 (N_15487,N_6440,N_5962);
and U15488 (N_15488,N_5828,N_2981);
and U15489 (N_15489,N_9443,N_7629);
and U15490 (N_15490,N_826,N_4802);
nor U15491 (N_15491,N_3502,N_7814);
nand U15492 (N_15492,N_6521,N_4935);
nand U15493 (N_15493,N_4356,N_4268);
nor U15494 (N_15494,N_514,N_1394);
or U15495 (N_15495,N_5686,N_5205);
and U15496 (N_15496,N_5809,N_6259);
and U15497 (N_15497,N_2842,N_2419);
or U15498 (N_15498,N_7319,N_6117);
or U15499 (N_15499,N_5843,N_9282);
or U15500 (N_15500,N_981,N_7040);
or U15501 (N_15501,N_9229,N_2395);
xor U15502 (N_15502,N_6683,N_5475);
nand U15503 (N_15503,N_338,N_6551);
nor U15504 (N_15504,N_1403,N_8774);
nand U15505 (N_15505,N_4771,N_229);
and U15506 (N_15506,N_9477,N_4355);
and U15507 (N_15507,N_8475,N_9172);
xnor U15508 (N_15508,N_5261,N_3479);
nor U15509 (N_15509,N_8302,N_1432);
nand U15510 (N_15510,N_599,N_3526);
or U15511 (N_15511,N_1964,N_865);
nor U15512 (N_15512,N_8519,N_1154);
and U15513 (N_15513,N_6220,N_7586);
and U15514 (N_15514,N_2357,N_4557);
and U15515 (N_15515,N_6961,N_1290);
and U15516 (N_15516,N_5090,N_9697);
and U15517 (N_15517,N_7226,N_4994);
and U15518 (N_15518,N_8621,N_2008);
nand U15519 (N_15519,N_5461,N_2637);
and U15520 (N_15520,N_8351,N_6780);
or U15521 (N_15521,N_9811,N_821);
nand U15522 (N_15522,N_3488,N_36);
and U15523 (N_15523,N_4188,N_8778);
nand U15524 (N_15524,N_9225,N_6691);
nor U15525 (N_15525,N_391,N_3769);
nor U15526 (N_15526,N_6652,N_4694);
or U15527 (N_15527,N_3647,N_9486);
or U15528 (N_15528,N_1036,N_8470);
nand U15529 (N_15529,N_4044,N_1455);
nand U15530 (N_15530,N_6463,N_7041);
nor U15531 (N_15531,N_4310,N_7829);
xnor U15532 (N_15532,N_9079,N_8862);
or U15533 (N_15533,N_8411,N_6870);
or U15534 (N_15534,N_5444,N_5073);
nand U15535 (N_15535,N_2002,N_8116);
or U15536 (N_15536,N_251,N_4572);
or U15537 (N_15537,N_9690,N_2846);
or U15538 (N_15538,N_1523,N_4973);
or U15539 (N_15539,N_8369,N_2118);
or U15540 (N_15540,N_2410,N_7433);
or U15541 (N_15541,N_9175,N_4082);
nand U15542 (N_15542,N_3092,N_9781);
or U15543 (N_15543,N_4548,N_5583);
nor U15544 (N_15544,N_3310,N_8090);
nand U15545 (N_15545,N_7761,N_9858);
nor U15546 (N_15546,N_6927,N_9753);
and U15547 (N_15547,N_8267,N_3684);
and U15548 (N_15548,N_2960,N_3091);
xnor U15549 (N_15549,N_7032,N_3230);
or U15550 (N_15550,N_9083,N_642);
nor U15551 (N_15551,N_2350,N_1682);
nor U15552 (N_15552,N_3572,N_3123);
or U15553 (N_15553,N_7954,N_6942);
or U15554 (N_15554,N_8174,N_4945);
nor U15555 (N_15555,N_8751,N_2425);
nor U15556 (N_15556,N_3735,N_2505);
or U15557 (N_15557,N_1195,N_2695);
nand U15558 (N_15558,N_5065,N_9069);
or U15559 (N_15559,N_7453,N_1663);
and U15560 (N_15560,N_8081,N_1727);
nor U15561 (N_15561,N_1169,N_7048);
nand U15562 (N_15562,N_6287,N_8941);
nor U15563 (N_15563,N_7599,N_2448);
nor U15564 (N_15564,N_1210,N_4086);
nand U15565 (N_15565,N_6715,N_4412);
nor U15566 (N_15566,N_1011,N_4928);
nand U15567 (N_15567,N_3446,N_3514);
and U15568 (N_15568,N_317,N_8793);
nand U15569 (N_15569,N_4945,N_8415);
nand U15570 (N_15570,N_7992,N_9903);
or U15571 (N_15571,N_4262,N_7542);
or U15572 (N_15572,N_4164,N_8696);
and U15573 (N_15573,N_4767,N_243);
nor U15574 (N_15574,N_4163,N_336);
nor U15575 (N_15575,N_6165,N_4500);
nand U15576 (N_15576,N_1120,N_8925);
nand U15577 (N_15577,N_300,N_1800);
or U15578 (N_15578,N_4818,N_8741);
xnor U15579 (N_15579,N_3943,N_1196);
or U15580 (N_15580,N_2545,N_379);
nand U15581 (N_15581,N_1366,N_5339);
xor U15582 (N_15582,N_6461,N_859);
or U15583 (N_15583,N_4716,N_5550);
or U15584 (N_15584,N_4391,N_5528);
nand U15585 (N_15585,N_1881,N_5230);
nor U15586 (N_15586,N_7509,N_3503);
nand U15587 (N_15587,N_2490,N_3056);
or U15588 (N_15588,N_2283,N_8356);
and U15589 (N_15589,N_1190,N_9018);
xor U15590 (N_15590,N_9902,N_5329);
nor U15591 (N_15591,N_7412,N_3918);
xor U15592 (N_15592,N_4444,N_346);
xor U15593 (N_15593,N_2060,N_9254);
nand U15594 (N_15594,N_5976,N_5281);
or U15595 (N_15595,N_6879,N_4342);
nor U15596 (N_15596,N_4050,N_6569);
nand U15597 (N_15597,N_5195,N_6912);
nand U15598 (N_15598,N_9460,N_9949);
nand U15599 (N_15599,N_5292,N_2409);
nand U15600 (N_15600,N_2917,N_2638);
or U15601 (N_15601,N_252,N_4224);
xor U15602 (N_15602,N_8398,N_9689);
nand U15603 (N_15603,N_7519,N_9387);
nor U15604 (N_15604,N_653,N_7572);
nand U15605 (N_15605,N_8419,N_7039);
and U15606 (N_15606,N_8812,N_6849);
xor U15607 (N_15607,N_9799,N_43);
nor U15608 (N_15608,N_8242,N_7763);
and U15609 (N_15609,N_8824,N_9445);
nand U15610 (N_15610,N_9707,N_1760);
nor U15611 (N_15611,N_465,N_7948);
nor U15612 (N_15612,N_6164,N_3318);
and U15613 (N_15613,N_7820,N_6925);
and U15614 (N_15614,N_1864,N_2861);
nor U15615 (N_15615,N_7317,N_6293);
xnor U15616 (N_15616,N_5478,N_9814);
nand U15617 (N_15617,N_2789,N_6259);
nor U15618 (N_15618,N_1582,N_525);
nand U15619 (N_15619,N_4124,N_625);
nand U15620 (N_15620,N_397,N_6786);
and U15621 (N_15621,N_1004,N_1811);
and U15622 (N_15622,N_5812,N_6357);
nand U15623 (N_15623,N_9854,N_1873);
nand U15624 (N_15624,N_6930,N_2511);
and U15625 (N_15625,N_7748,N_4934);
and U15626 (N_15626,N_376,N_3256);
xor U15627 (N_15627,N_9654,N_9431);
nand U15628 (N_15628,N_1209,N_8884);
nor U15629 (N_15629,N_8275,N_3144);
nand U15630 (N_15630,N_5577,N_3821);
nor U15631 (N_15631,N_7639,N_9480);
nor U15632 (N_15632,N_4473,N_4647);
nor U15633 (N_15633,N_4809,N_9199);
nand U15634 (N_15634,N_9973,N_1148);
and U15635 (N_15635,N_9937,N_6212);
or U15636 (N_15636,N_3654,N_2356);
and U15637 (N_15637,N_5081,N_4856);
or U15638 (N_15638,N_9203,N_717);
nand U15639 (N_15639,N_9298,N_5527);
or U15640 (N_15640,N_4518,N_8146);
nor U15641 (N_15641,N_3958,N_4583);
nand U15642 (N_15642,N_5768,N_5039);
nand U15643 (N_15643,N_6021,N_1160);
and U15644 (N_15644,N_9320,N_969);
nand U15645 (N_15645,N_7591,N_9553);
xor U15646 (N_15646,N_5525,N_3665);
nand U15647 (N_15647,N_1632,N_333);
and U15648 (N_15648,N_6607,N_3194);
xor U15649 (N_15649,N_7616,N_688);
nor U15650 (N_15650,N_7399,N_9742);
nand U15651 (N_15651,N_7643,N_6473);
or U15652 (N_15652,N_8834,N_1788);
and U15653 (N_15653,N_440,N_8317);
nand U15654 (N_15654,N_3270,N_9774);
nor U15655 (N_15655,N_5929,N_999);
or U15656 (N_15656,N_7342,N_1951);
nor U15657 (N_15657,N_1259,N_7863);
or U15658 (N_15658,N_8520,N_1056);
or U15659 (N_15659,N_2406,N_8643);
xor U15660 (N_15660,N_7966,N_4450);
or U15661 (N_15661,N_2255,N_681);
nor U15662 (N_15662,N_8146,N_8737);
nor U15663 (N_15663,N_5270,N_2124);
nor U15664 (N_15664,N_2191,N_4351);
or U15665 (N_15665,N_6255,N_2497);
or U15666 (N_15666,N_488,N_2674);
and U15667 (N_15667,N_3485,N_4215);
and U15668 (N_15668,N_4467,N_6091);
and U15669 (N_15669,N_9354,N_2008);
and U15670 (N_15670,N_3335,N_9445);
nand U15671 (N_15671,N_4695,N_7452);
nand U15672 (N_15672,N_8516,N_122);
nor U15673 (N_15673,N_6919,N_8523);
and U15674 (N_15674,N_7335,N_1570);
nand U15675 (N_15675,N_6552,N_3673);
nor U15676 (N_15676,N_5502,N_3250);
and U15677 (N_15677,N_9472,N_7885);
nand U15678 (N_15678,N_1154,N_1390);
or U15679 (N_15679,N_6174,N_6789);
nand U15680 (N_15680,N_247,N_8066);
nand U15681 (N_15681,N_2340,N_341);
or U15682 (N_15682,N_8814,N_3221);
nor U15683 (N_15683,N_9681,N_8904);
or U15684 (N_15684,N_6914,N_4222);
and U15685 (N_15685,N_6814,N_9264);
and U15686 (N_15686,N_7546,N_7263);
and U15687 (N_15687,N_8011,N_798);
nor U15688 (N_15688,N_1918,N_9968);
or U15689 (N_15689,N_3671,N_6285);
and U15690 (N_15690,N_2339,N_9161);
nor U15691 (N_15691,N_213,N_2063);
nor U15692 (N_15692,N_2873,N_503);
and U15693 (N_15693,N_4659,N_8165);
nand U15694 (N_15694,N_1646,N_7709);
nor U15695 (N_15695,N_4776,N_6629);
nand U15696 (N_15696,N_9712,N_3667);
nand U15697 (N_15697,N_2791,N_2886);
nand U15698 (N_15698,N_5194,N_731);
or U15699 (N_15699,N_9263,N_4179);
and U15700 (N_15700,N_8845,N_349);
nor U15701 (N_15701,N_1698,N_534);
and U15702 (N_15702,N_2654,N_168);
and U15703 (N_15703,N_5729,N_61);
and U15704 (N_15704,N_3589,N_9031);
nor U15705 (N_15705,N_783,N_9680);
nand U15706 (N_15706,N_6973,N_9555);
and U15707 (N_15707,N_9,N_5842);
or U15708 (N_15708,N_3054,N_3092);
nand U15709 (N_15709,N_1353,N_4550);
nand U15710 (N_15710,N_3518,N_857);
nand U15711 (N_15711,N_4641,N_8810);
nor U15712 (N_15712,N_7246,N_5777);
nor U15713 (N_15713,N_2661,N_4068);
or U15714 (N_15714,N_7095,N_7472);
nand U15715 (N_15715,N_6419,N_681);
xor U15716 (N_15716,N_9531,N_2188);
or U15717 (N_15717,N_5429,N_4866);
or U15718 (N_15718,N_6212,N_524);
and U15719 (N_15719,N_3183,N_6074);
nor U15720 (N_15720,N_7864,N_4056);
nand U15721 (N_15721,N_657,N_4126);
or U15722 (N_15722,N_3688,N_7406);
or U15723 (N_15723,N_4653,N_4962);
or U15724 (N_15724,N_7189,N_8956);
and U15725 (N_15725,N_2915,N_8271);
nand U15726 (N_15726,N_4534,N_6650);
or U15727 (N_15727,N_1990,N_5234);
nor U15728 (N_15728,N_8546,N_6626);
nand U15729 (N_15729,N_2260,N_3615);
or U15730 (N_15730,N_1252,N_9442);
xor U15731 (N_15731,N_2765,N_2264);
nand U15732 (N_15732,N_9297,N_7138);
or U15733 (N_15733,N_2720,N_2366);
nand U15734 (N_15734,N_1889,N_5127);
nand U15735 (N_15735,N_5426,N_7502);
and U15736 (N_15736,N_3367,N_5487);
xnor U15737 (N_15737,N_8562,N_609);
nand U15738 (N_15738,N_7198,N_6931);
nor U15739 (N_15739,N_9185,N_9644);
and U15740 (N_15740,N_9157,N_1680);
and U15741 (N_15741,N_2720,N_6197);
nand U15742 (N_15742,N_2643,N_4222);
nor U15743 (N_15743,N_9446,N_1766);
nor U15744 (N_15744,N_7596,N_5126);
or U15745 (N_15745,N_636,N_3288);
nor U15746 (N_15746,N_8134,N_7068);
and U15747 (N_15747,N_5280,N_562);
and U15748 (N_15748,N_7103,N_3307);
nor U15749 (N_15749,N_2450,N_3027);
nor U15750 (N_15750,N_3667,N_7536);
or U15751 (N_15751,N_4474,N_133);
nor U15752 (N_15752,N_6206,N_8402);
and U15753 (N_15753,N_1160,N_2692);
and U15754 (N_15754,N_3120,N_235);
or U15755 (N_15755,N_5089,N_8142);
xor U15756 (N_15756,N_2610,N_1931);
and U15757 (N_15757,N_1465,N_7775);
and U15758 (N_15758,N_4446,N_7402);
nor U15759 (N_15759,N_4850,N_466);
nand U15760 (N_15760,N_347,N_4725);
nor U15761 (N_15761,N_9159,N_4816);
xnor U15762 (N_15762,N_8133,N_2819);
nor U15763 (N_15763,N_1659,N_3919);
or U15764 (N_15764,N_8868,N_2575);
nand U15765 (N_15765,N_2116,N_8066);
and U15766 (N_15766,N_6856,N_2518);
nor U15767 (N_15767,N_8689,N_7074);
or U15768 (N_15768,N_5267,N_4540);
and U15769 (N_15769,N_7935,N_6589);
xor U15770 (N_15770,N_1495,N_4147);
nand U15771 (N_15771,N_5910,N_619);
xor U15772 (N_15772,N_4279,N_9813);
nor U15773 (N_15773,N_6638,N_5538);
xor U15774 (N_15774,N_1224,N_9275);
nor U15775 (N_15775,N_6632,N_5109);
or U15776 (N_15776,N_2305,N_8458);
or U15777 (N_15777,N_375,N_8924);
xnor U15778 (N_15778,N_5386,N_6320);
nor U15779 (N_15779,N_7784,N_1856);
nand U15780 (N_15780,N_5752,N_1264);
or U15781 (N_15781,N_4907,N_290);
nor U15782 (N_15782,N_4362,N_2538);
nand U15783 (N_15783,N_3600,N_3342);
nand U15784 (N_15784,N_2771,N_2445);
nor U15785 (N_15785,N_8986,N_2836);
or U15786 (N_15786,N_1953,N_2671);
and U15787 (N_15787,N_724,N_5947);
nor U15788 (N_15788,N_6556,N_4760);
nand U15789 (N_15789,N_8302,N_7601);
nor U15790 (N_15790,N_2846,N_7417);
or U15791 (N_15791,N_8185,N_9372);
or U15792 (N_15792,N_7058,N_5518);
or U15793 (N_15793,N_4972,N_5102);
or U15794 (N_15794,N_4969,N_3141);
nor U15795 (N_15795,N_9726,N_2474);
nand U15796 (N_15796,N_6472,N_882);
nor U15797 (N_15797,N_4321,N_9573);
and U15798 (N_15798,N_1962,N_3871);
or U15799 (N_15799,N_3546,N_4034);
and U15800 (N_15800,N_2258,N_9816);
or U15801 (N_15801,N_688,N_1872);
nand U15802 (N_15802,N_3460,N_3342);
or U15803 (N_15803,N_5788,N_9110);
or U15804 (N_15804,N_840,N_7416);
or U15805 (N_15805,N_3149,N_8485);
xnor U15806 (N_15806,N_5832,N_4493);
and U15807 (N_15807,N_6234,N_1807);
or U15808 (N_15808,N_7414,N_8378);
nor U15809 (N_15809,N_7152,N_2716);
nor U15810 (N_15810,N_519,N_5499);
or U15811 (N_15811,N_7707,N_6003);
nor U15812 (N_15812,N_5665,N_5641);
nor U15813 (N_15813,N_3043,N_4508);
and U15814 (N_15814,N_2400,N_8999);
nand U15815 (N_15815,N_1430,N_5462);
nor U15816 (N_15816,N_8190,N_6893);
or U15817 (N_15817,N_8830,N_8267);
or U15818 (N_15818,N_5326,N_4881);
xnor U15819 (N_15819,N_5708,N_9816);
or U15820 (N_15820,N_3921,N_4021);
nand U15821 (N_15821,N_4108,N_7244);
nor U15822 (N_15822,N_2138,N_8827);
and U15823 (N_15823,N_6089,N_4198);
nor U15824 (N_15824,N_1753,N_9205);
nor U15825 (N_15825,N_6180,N_8005);
nor U15826 (N_15826,N_6841,N_9638);
nand U15827 (N_15827,N_8375,N_2972);
xnor U15828 (N_15828,N_4295,N_7860);
nand U15829 (N_15829,N_5684,N_1998);
and U15830 (N_15830,N_2249,N_4738);
and U15831 (N_15831,N_4236,N_3382);
nor U15832 (N_15832,N_7608,N_7374);
and U15833 (N_15833,N_7878,N_998);
nor U15834 (N_15834,N_6611,N_5727);
and U15835 (N_15835,N_2279,N_5);
nor U15836 (N_15836,N_963,N_6964);
and U15837 (N_15837,N_3479,N_5821);
nor U15838 (N_15838,N_5073,N_5750);
nor U15839 (N_15839,N_7027,N_7640);
nand U15840 (N_15840,N_3622,N_5723);
and U15841 (N_15841,N_3084,N_865);
or U15842 (N_15842,N_249,N_6936);
nand U15843 (N_15843,N_4841,N_4187);
nand U15844 (N_15844,N_694,N_1072);
nand U15845 (N_15845,N_1642,N_552);
xnor U15846 (N_15846,N_3516,N_7813);
nor U15847 (N_15847,N_1072,N_1939);
nor U15848 (N_15848,N_2644,N_1169);
or U15849 (N_15849,N_4976,N_7657);
nor U15850 (N_15850,N_8692,N_4193);
nand U15851 (N_15851,N_8586,N_8869);
and U15852 (N_15852,N_5732,N_8446);
nand U15853 (N_15853,N_6391,N_2689);
or U15854 (N_15854,N_330,N_5938);
nand U15855 (N_15855,N_784,N_3675);
and U15856 (N_15856,N_690,N_3526);
xor U15857 (N_15857,N_1307,N_1752);
or U15858 (N_15858,N_7884,N_9648);
nor U15859 (N_15859,N_5808,N_3881);
nand U15860 (N_15860,N_4996,N_4026);
or U15861 (N_15861,N_8461,N_1270);
nor U15862 (N_15862,N_8243,N_6212);
nand U15863 (N_15863,N_0,N_2822);
or U15864 (N_15864,N_2110,N_1368);
nor U15865 (N_15865,N_7001,N_6841);
and U15866 (N_15866,N_9444,N_7373);
or U15867 (N_15867,N_5446,N_822);
nand U15868 (N_15868,N_5157,N_255);
and U15869 (N_15869,N_2262,N_9751);
nor U15870 (N_15870,N_7788,N_7266);
or U15871 (N_15871,N_8315,N_444);
nand U15872 (N_15872,N_1622,N_2964);
nand U15873 (N_15873,N_4220,N_6843);
nand U15874 (N_15874,N_721,N_2221);
nor U15875 (N_15875,N_1553,N_7806);
nand U15876 (N_15876,N_3980,N_823);
nor U15877 (N_15877,N_9626,N_1895);
or U15878 (N_15878,N_9856,N_3961);
or U15879 (N_15879,N_8329,N_1308);
nand U15880 (N_15880,N_2435,N_6374);
nand U15881 (N_15881,N_97,N_5938);
nand U15882 (N_15882,N_5680,N_3027);
nand U15883 (N_15883,N_9738,N_3134);
xor U15884 (N_15884,N_2316,N_7586);
nand U15885 (N_15885,N_4115,N_7686);
or U15886 (N_15886,N_2199,N_6177);
nand U15887 (N_15887,N_6009,N_4376);
and U15888 (N_15888,N_6822,N_6903);
nor U15889 (N_15889,N_5978,N_3223);
or U15890 (N_15890,N_2266,N_1369);
nand U15891 (N_15891,N_5716,N_5681);
and U15892 (N_15892,N_7227,N_4981);
xnor U15893 (N_15893,N_1562,N_4472);
and U15894 (N_15894,N_6387,N_200);
nor U15895 (N_15895,N_554,N_6388);
or U15896 (N_15896,N_7063,N_6073);
and U15897 (N_15897,N_6880,N_8376);
nor U15898 (N_15898,N_3898,N_8746);
nor U15899 (N_15899,N_9908,N_9480);
nor U15900 (N_15900,N_1925,N_7555);
or U15901 (N_15901,N_7507,N_9863);
or U15902 (N_15902,N_654,N_9805);
xnor U15903 (N_15903,N_5827,N_4347);
or U15904 (N_15904,N_7137,N_8623);
nor U15905 (N_15905,N_4193,N_5509);
nor U15906 (N_15906,N_451,N_6238);
or U15907 (N_15907,N_7196,N_7571);
and U15908 (N_15908,N_6454,N_8005);
nand U15909 (N_15909,N_1981,N_2869);
nor U15910 (N_15910,N_5536,N_8679);
nand U15911 (N_15911,N_6270,N_1191);
nor U15912 (N_15912,N_2984,N_101);
and U15913 (N_15913,N_3368,N_6001);
and U15914 (N_15914,N_4663,N_4673);
xnor U15915 (N_15915,N_5526,N_4409);
and U15916 (N_15916,N_745,N_1746);
nand U15917 (N_15917,N_6493,N_9728);
nand U15918 (N_15918,N_2143,N_5943);
or U15919 (N_15919,N_5458,N_4006);
and U15920 (N_15920,N_8785,N_7811);
nor U15921 (N_15921,N_9502,N_8192);
xor U15922 (N_15922,N_9624,N_6902);
nand U15923 (N_15923,N_7705,N_9888);
nand U15924 (N_15924,N_2089,N_4119);
nand U15925 (N_15925,N_1362,N_7340);
and U15926 (N_15926,N_9955,N_7809);
nand U15927 (N_15927,N_4011,N_4416);
nor U15928 (N_15928,N_6418,N_3673);
nand U15929 (N_15929,N_9672,N_6298);
or U15930 (N_15930,N_8413,N_6625);
nand U15931 (N_15931,N_1053,N_8384);
nand U15932 (N_15932,N_6413,N_7884);
xnor U15933 (N_15933,N_267,N_268);
and U15934 (N_15934,N_9567,N_7749);
and U15935 (N_15935,N_7365,N_4509);
nand U15936 (N_15936,N_1852,N_2586);
and U15937 (N_15937,N_6513,N_6783);
nand U15938 (N_15938,N_7649,N_5362);
nor U15939 (N_15939,N_1792,N_652);
or U15940 (N_15940,N_3892,N_5132);
nor U15941 (N_15941,N_9769,N_6225);
nor U15942 (N_15942,N_9554,N_2136);
xor U15943 (N_15943,N_795,N_5469);
or U15944 (N_15944,N_8369,N_7694);
nor U15945 (N_15945,N_7081,N_3486);
or U15946 (N_15946,N_4504,N_6844);
and U15947 (N_15947,N_9237,N_5373);
and U15948 (N_15948,N_8314,N_7929);
xor U15949 (N_15949,N_5519,N_6465);
and U15950 (N_15950,N_9415,N_1618);
nand U15951 (N_15951,N_8054,N_4960);
xnor U15952 (N_15952,N_2261,N_7275);
nor U15953 (N_15953,N_8661,N_598);
nor U15954 (N_15954,N_7013,N_2889);
nor U15955 (N_15955,N_2072,N_451);
or U15956 (N_15956,N_7188,N_836);
nor U15957 (N_15957,N_3570,N_143);
or U15958 (N_15958,N_2224,N_8913);
nand U15959 (N_15959,N_110,N_2244);
nand U15960 (N_15960,N_2857,N_2686);
and U15961 (N_15961,N_3215,N_7273);
nor U15962 (N_15962,N_2490,N_9181);
or U15963 (N_15963,N_6816,N_5831);
xnor U15964 (N_15964,N_6996,N_1636);
xor U15965 (N_15965,N_2992,N_1030);
nor U15966 (N_15966,N_7082,N_362);
nor U15967 (N_15967,N_5130,N_4811);
nand U15968 (N_15968,N_2588,N_2086);
or U15969 (N_15969,N_5341,N_4619);
or U15970 (N_15970,N_42,N_6150);
or U15971 (N_15971,N_2905,N_3916);
or U15972 (N_15972,N_9250,N_9755);
xor U15973 (N_15973,N_7595,N_620);
and U15974 (N_15974,N_2649,N_1493);
and U15975 (N_15975,N_6961,N_439);
nand U15976 (N_15976,N_8064,N_6991);
nand U15977 (N_15977,N_5070,N_1214);
and U15978 (N_15978,N_4887,N_7238);
nor U15979 (N_15979,N_645,N_2054);
nor U15980 (N_15980,N_8182,N_9674);
or U15981 (N_15981,N_3631,N_8770);
nand U15982 (N_15982,N_2729,N_1679);
nor U15983 (N_15983,N_187,N_340);
and U15984 (N_15984,N_3989,N_7870);
or U15985 (N_15985,N_386,N_2696);
or U15986 (N_15986,N_8903,N_9916);
and U15987 (N_15987,N_4329,N_8191);
and U15988 (N_15988,N_3830,N_2597);
nand U15989 (N_15989,N_7905,N_6485);
nor U15990 (N_15990,N_9323,N_3194);
or U15991 (N_15991,N_9028,N_3282);
and U15992 (N_15992,N_9370,N_4635);
nor U15993 (N_15993,N_1027,N_1231);
nand U15994 (N_15994,N_1872,N_117);
and U15995 (N_15995,N_6146,N_8061);
nand U15996 (N_15996,N_7514,N_2116);
nand U15997 (N_15997,N_7080,N_4417);
nor U15998 (N_15998,N_7554,N_1223);
nand U15999 (N_15999,N_5166,N_6836);
and U16000 (N_16000,N_2986,N_9538);
and U16001 (N_16001,N_5207,N_1682);
and U16002 (N_16002,N_4020,N_8324);
and U16003 (N_16003,N_7596,N_7103);
and U16004 (N_16004,N_5673,N_3612);
or U16005 (N_16005,N_4977,N_7219);
or U16006 (N_16006,N_1311,N_8451);
nor U16007 (N_16007,N_5913,N_2296);
nand U16008 (N_16008,N_2097,N_5932);
or U16009 (N_16009,N_206,N_6457);
nand U16010 (N_16010,N_7065,N_6227);
and U16011 (N_16011,N_308,N_8168);
nor U16012 (N_16012,N_5942,N_8423);
nor U16013 (N_16013,N_6965,N_2972);
and U16014 (N_16014,N_7313,N_531);
nor U16015 (N_16015,N_8035,N_236);
nor U16016 (N_16016,N_3519,N_6408);
nor U16017 (N_16017,N_7595,N_9650);
and U16018 (N_16018,N_8946,N_8902);
nand U16019 (N_16019,N_4535,N_3856);
nor U16020 (N_16020,N_8296,N_6149);
and U16021 (N_16021,N_7163,N_23);
and U16022 (N_16022,N_3654,N_9120);
and U16023 (N_16023,N_6443,N_7567);
and U16024 (N_16024,N_4238,N_1800);
or U16025 (N_16025,N_8750,N_8054);
nand U16026 (N_16026,N_7415,N_7766);
and U16027 (N_16027,N_2758,N_1822);
and U16028 (N_16028,N_7242,N_2489);
nor U16029 (N_16029,N_6110,N_1055);
and U16030 (N_16030,N_7348,N_5208);
and U16031 (N_16031,N_4437,N_5838);
and U16032 (N_16032,N_3544,N_2400);
xnor U16033 (N_16033,N_7612,N_8311);
and U16034 (N_16034,N_3794,N_7143);
nor U16035 (N_16035,N_763,N_1933);
nand U16036 (N_16036,N_1571,N_7131);
or U16037 (N_16037,N_4506,N_5627);
nand U16038 (N_16038,N_736,N_6917);
and U16039 (N_16039,N_5828,N_9232);
nor U16040 (N_16040,N_1477,N_1500);
nand U16041 (N_16041,N_79,N_7751);
and U16042 (N_16042,N_5196,N_642);
nor U16043 (N_16043,N_3607,N_9365);
or U16044 (N_16044,N_7404,N_1711);
nand U16045 (N_16045,N_2872,N_7623);
nor U16046 (N_16046,N_2545,N_9688);
xor U16047 (N_16047,N_8592,N_579);
nand U16048 (N_16048,N_9478,N_7645);
and U16049 (N_16049,N_3780,N_6374);
or U16050 (N_16050,N_9528,N_9368);
and U16051 (N_16051,N_3200,N_3715);
or U16052 (N_16052,N_9493,N_1784);
nor U16053 (N_16053,N_567,N_5226);
and U16054 (N_16054,N_455,N_6725);
nand U16055 (N_16055,N_7733,N_194);
nand U16056 (N_16056,N_1280,N_9909);
nor U16057 (N_16057,N_372,N_9163);
nor U16058 (N_16058,N_3519,N_8385);
and U16059 (N_16059,N_5158,N_8849);
nand U16060 (N_16060,N_7908,N_9036);
and U16061 (N_16061,N_7373,N_8392);
xnor U16062 (N_16062,N_5309,N_5825);
or U16063 (N_16063,N_69,N_5534);
xor U16064 (N_16064,N_8850,N_5905);
xnor U16065 (N_16065,N_5142,N_8162);
and U16066 (N_16066,N_6637,N_3617);
or U16067 (N_16067,N_5441,N_1515);
nand U16068 (N_16068,N_1493,N_1666);
nor U16069 (N_16069,N_2582,N_8026);
and U16070 (N_16070,N_4686,N_6698);
or U16071 (N_16071,N_4773,N_7499);
nor U16072 (N_16072,N_9991,N_2420);
nand U16073 (N_16073,N_662,N_1103);
nand U16074 (N_16074,N_5434,N_696);
nor U16075 (N_16075,N_9583,N_5690);
and U16076 (N_16076,N_8541,N_4596);
or U16077 (N_16077,N_40,N_6461);
and U16078 (N_16078,N_1755,N_734);
or U16079 (N_16079,N_1660,N_6064);
xnor U16080 (N_16080,N_8229,N_9243);
nor U16081 (N_16081,N_7646,N_3319);
nor U16082 (N_16082,N_3196,N_3508);
and U16083 (N_16083,N_6663,N_3069);
and U16084 (N_16084,N_5362,N_5430);
and U16085 (N_16085,N_7509,N_2611);
or U16086 (N_16086,N_6163,N_7749);
nand U16087 (N_16087,N_9846,N_9184);
or U16088 (N_16088,N_5605,N_8688);
or U16089 (N_16089,N_2770,N_2628);
and U16090 (N_16090,N_210,N_5049);
or U16091 (N_16091,N_7314,N_6209);
and U16092 (N_16092,N_9798,N_1191);
and U16093 (N_16093,N_4558,N_1290);
and U16094 (N_16094,N_5560,N_3974);
or U16095 (N_16095,N_186,N_8143);
and U16096 (N_16096,N_6991,N_5930);
nand U16097 (N_16097,N_9242,N_942);
nor U16098 (N_16098,N_8151,N_4107);
or U16099 (N_16099,N_5320,N_4612);
and U16100 (N_16100,N_4667,N_2221);
and U16101 (N_16101,N_2651,N_1054);
nand U16102 (N_16102,N_9386,N_4403);
and U16103 (N_16103,N_6139,N_4423);
nand U16104 (N_16104,N_9645,N_860);
nor U16105 (N_16105,N_1121,N_1714);
or U16106 (N_16106,N_340,N_331);
or U16107 (N_16107,N_9994,N_7426);
nand U16108 (N_16108,N_2317,N_3467);
and U16109 (N_16109,N_3715,N_1279);
or U16110 (N_16110,N_4721,N_9435);
nand U16111 (N_16111,N_6577,N_939);
nand U16112 (N_16112,N_8773,N_645);
or U16113 (N_16113,N_7973,N_132);
and U16114 (N_16114,N_3238,N_6360);
nand U16115 (N_16115,N_4928,N_413);
nor U16116 (N_16116,N_2814,N_7193);
nand U16117 (N_16117,N_4926,N_4116);
nor U16118 (N_16118,N_3915,N_897);
nand U16119 (N_16119,N_164,N_9619);
nor U16120 (N_16120,N_7169,N_101);
nor U16121 (N_16121,N_8217,N_4611);
or U16122 (N_16122,N_5382,N_5351);
xnor U16123 (N_16123,N_9423,N_8193);
nor U16124 (N_16124,N_621,N_9069);
xnor U16125 (N_16125,N_1634,N_8971);
xnor U16126 (N_16126,N_6918,N_336);
xor U16127 (N_16127,N_45,N_2509);
or U16128 (N_16128,N_3443,N_3447);
xnor U16129 (N_16129,N_8853,N_2851);
nand U16130 (N_16130,N_4451,N_6161);
nand U16131 (N_16131,N_9858,N_7792);
nor U16132 (N_16132,N_2161,N_9682);
nand U16133 (N_16133,N_6654,N_1173);
nand U16134 (N_16134,N_9969,N_4905);
xnor U16135 (N_16135,N_6013,N_8207);
nor U16136 (N_16136,N_2704,N_217);
nand U16137 (N_16137,N_2592,N_6406);
nand U16138 (N_16138,N_8422,N_7583);
nand U16139 (N_16139,N_8903,N_2399);
or U16140 (N_16140,N_7614,N_9297);
and U16141 (N_16141,N_7027,N_1809);
nor U16142 (N_16142,N_485,N_360);
or U16143 (N_16143,N_6182,N_9277);
nor U16144 (N_16144,N_4920,N_362);
nand U16145 (N_16145,N_2553,N_6242);
or U16146 (N_16146,N_5016,N_6672);
nand U16147 (N_16147,N_9979,N_7794);
xnor U16148 (N_16148,N_2463,N_1210);
and U16149 (N_16149,N_8629,N_1062);
and U16150 (N_16150,N_5640,N_6491);
or U16151 (N_16151,N_1368,N_4042);
and U16152 (N_16152,N_6701,N_8024);
and U16153 (N_16153,N_9571,N_6201);
nor U16154 (N_16154,N_509,N_6316);
or U16155 (N_16155,N_8028,N_517);
or U16156 (N_16156,N_120,N_5987);
nor U16157 (N_16157,N_5216,N_317);
and U16158 (N_16158,N_512,N_800);
nand U16159 (N_16159,N_9167,N_2544);
and U16160 (N_16160,N_3945,N_2556);
nor U16161 (N_16161,N_8592,N_224);
nand U16162 (N_16162,N_9876,N_1238);
xor U16163 (N_16163,N_3120,N_8946);
nand U16164 (N_16164,N_9435,N_653);
and U16165 (N_16165,N_7530,N_941);
or U16166 (N_16166,N_7979,N_120);
nor U16167 (N_16167,N_4035,N_7069);
nor U16168 (N_16168,N_6516,N_8127);
nand U16169 (N_16169,N_3384,N_1465);
xnor U16170 (N_16170,N_9153,N_8634);
nor U16171 (N_16171,N_328,N_6508);
or U16172 (N_16172,N_5430,N_7712);
and U16173 (N_16173,N_1797,N_9324);
nand U16174 (N_16174,N_7358,N_5991);
xnor U16175 (N_16175,N_9087,N_6840);
xor U16176 (N_16176,N_953,N_7170);
nand U16177 (N_16177,N_5769,N_7628);
nand U16178 (N_16178,N_7797,N_2589);
or U16179 (N_16179,N_1351,N_3742);
or U16180 (N_16180,N_4964,N_1134);
nand U16181 (N_16181,N_4278,N_233);
nor U16182 (N_16182,N_2600,N_6908);
or U16183 (N_16183,N_8810,N_4299);
nor U16184 (N_16184,N_9435,N_5470);
nand U16185 (N_16185,N_7025,N_311);
or U16186 (N_16186,N_4027,N_904);
or U16187 (N_16187,N_5648,N_306);
nor U16188 (N_16188,N_1907,N_4644);
or U16189 (N_16189,N_8718,N_6683);
nand U16190 (N_16190,N_3555,N_8898);
or U16191 (N_16191,N_4257,N_8848);
nand U16192 (N_16192,N_5721,N_7709);
and U16193 (N_16193,N_8144,N_6958);
nor U16194 (N_16194,N_4428,N_4509);
nand U16195 (N_16195,N_3435,N_8607);
and U16196 (N_16196,N_6189,N_1307);
and U16197 (N_16197,N_9222,N_5651);
and U16198 (N_16198,N_9350,N_7744);
nand U16199 (N_16199,N_3966,N_7401);
nand U16200 (N_16200,N_9665,N_996);
nor U16201 (N_16201,N_3578,N_9577);
xnor U16202 (N_16202,N_7067,N_8470);
nor U16203 (N_16203,N_9862,N_9738);
or U16204 (N_16204,N_4956,N_7235);
nand U16205 (N_16205,N_4731,N_962);
or U16206 (N_16206,N_1482,N_2108);
nand U16207 (N_16207,N_8772,N_7402);
nand U16208 (N_16208,N_1052,N_7620);
nand U16209 (N_16209,N_4743,N_7963);
and U16210 (N_16210,N_2883,N_2282);
or U16211 (N_16211,N_5361,N_7813);
nand U16212 (N_16212,N_1597,N_4140);
nor U16213 (N_16213,N_8228,N_1626);
nor U16214 (N_16214,N_8579,N_9782);
and U16215 (N_16215,N_9868,N_9083);
and U16216 (N_16216,N_4073,N_1266);
and U16217 (N_16217,N_6602,N_9110);
and U16218 (N_16218,N_6896,N_7664);
xnor U16219 (N_16219,N_2161,N_4167);
or U16220 (N_16220,N_5810,N_3210);
and U16221 (N_16221,N_3859,N_837);
or U16222 (N_16222,N_8425,N_8713);
nor U16223 (N_16223,N_7835,N_896);
xnor U16224 (N_16224,N_3165,N_1963);
nor U16225 (N_16225,N_2551,N_3669);
nand U16226 (N_16226,N_3904,N_4304);
xor U16227 (N_16227,N_638,N_9763);
nand U16228 (N_16228,N_7424,N_7494);
nor U16229 (N_16229,N_1202,N_8801);
nor U16230 (N_16230,N_5052,N_7528);
nor U16231 (N_16231,N_1397,N_8853);
nand U16232 (N_16232,N_9853,N_9871);
and U16233 (N_16233,N_7445,N_524);
nor U16234 (N_16234,N_8089,N_1267);
and U16235 (N_16235,N_8037,N_8306);
nor U16236 (N_16236,N_779,N_1751);
or U16237 (N_16237,N_7132,N_8562);
nand U16238 (N_16238,N_2815,N_4801);
nor U16239 (N_16239,N_5873,N_7972);
xnor U16240 (N_16240,N_861,N_3786);
nor U16241 (N_16241,N_2738,N_231);
and U16242 (N_16242,N_102,N_3601);
and U16243 (N_16243,N_7469,N_7750);
nand U16244 (N_16244,N_928,N_5080);
or U16245 (N_16245,N_1487,N_4005);
and U16246 (N_16246,N_2313,N_1690);
nor U16247 (N_16247,N_3166,N_2975);
nand U16248 (N_16248,N_2588,N_668);
nor U16249 (N_16249,N_1039,N_5868);
nor U16250 (N_16250,N_9392,N_3445);
or U16251 (N_16251,N_8335,N_807);
and U16252 (N_16252,N_856,N_2098);
xor U16253 (N_16253,N_7452,N_311);
xor U16254 (N_16254,N_7890,N_5260);
nand U16255 (N_16255,N_3651,N_4687);
or U16256 (N_16256,N_1648,N_2554);
nand U16257 (N_16257,N_7865,N_352);
and U16258 (N_16258,N_6885,N_9004);
nand U16259 (N_16259,N_1268,N_1574);
nand U16260 (N_16260,N_6416,N_564);
nand U16261 (N_16261,N_2600,N_7363);
or U16262 (N_16262,N_2363,N_499);
xor U16263 (N_16263,N_4088,N_7742);
xnor U16264 (N_16264,N_1999,N_1392);
nand U16265 (N_16265,N_9338,N_7731);
nor U16266 (N_16266,N_5366,N_4389);
nor U16267 (N_16267,N_4938,N_7641);
nor U16268 (N_16268,N_2073,N_3112);
or U16269 (N_16269,N_7121,N_650);
nor U16270 (N_16270,N_1781,N_5370);
and U16271 (N_16271,N_9111,N_8395);
or U16272 (N_16272,N_4782,N_2000);
and U16273 (N_16273,N_908,N_3700);
xor U16274 (N_16274,N_453,N_953);
xor U16275 (N_16275,N_2509,N_751);
xor U16276 (N_16276,N_1798,N_6760);
nor U16277 (N_16277,N_142,N_5783);
or U16278 (N_16278,N_3658,N_820);
and U16279 (N_16279,N_5297,N_9379);
or U16280 (N_16280,N_5651,N_7895);
or U16281 (N_16281,N_6223,N_2223);
and U16282 (N_16282,N_9512,N_3932);
nor U16283 (N_16283,N_4612,N_9499);
nor U16284 (N_16284,N_1703,N_9907);
nand U16285 (N_16285,N_9894,N_8832);
nor U16286 (N_16286,N_8858,N_1048);
nand U16287 (N_16287,N_2553,N_4555);
nand U16288 (N_16288,N_3156,N_9302);
nand U16289 (N_16289,N_7287,N_6514);
nor U16290 (N_16290,N_9989,N_8115);
or U16291 (N_16291,N_7930,N_1831);
nand U16292 (N_16292,N_4607,N_9641);
nor U16293 (N_16293,N_2139,N_9876);
nand U16294 (N_16294,N_4154,N_5814);
and U16295 (N_16295,N_9190,N_9026);
or U16296 (N_16296,N_3806,N_2129);
or U16297 (N_16297,N_8345,N_7104);
xor U16298 (N_16298,N_3370,N_2947);
or U16299 (N_16299,N_1754,N_8596);
nor U16300 (N_16300,N_4247,N_8300);
and U16301 (N_16301,N_4497,N_4768);
xnor U16302 (N_16302,N_2106,N_4783);
nor U16303 (N_16303,N_5644,N_7338);
xor U16304 (N_16304,N_5287,N_7504);
and U16305 (N_16305,N_1140,N_4135);
xnor U16306 (N_16306,N_4942,N_9388);
nor U16307 (N_16307,N_1367,N_3609);
nor U16308 (N_16308,N_5319,N_1486);
or U16309 (N_16309,N_1152,N_5280);
or U16310 (N_16310,N_6962,N_9187);
xnor U16311 (N_16311,N_4413,N_2122);
nand U16312 (N_16312,N_2818,N_3151);
and U16313 (N_16313,N_6035,N_3573);
nand U16314 (N_16314,N_9287,N_4865);
or U16315 (N_16315,N_310,N_3853);
or U16316 (N_16316,N_9804,N_9240);
or U16317 (N_16317,N_4025,N_2460);
xnor U16318 (N_16318,N_7958,N_3556);
nor U16319 (N_16319,N_5270,N_544);
nand U16320 (N_16320,N_6907,N_1913);
nor U16321 (N_16321,N_510,N_8251);
or U16322 (N_16322,N_3530,N_5586);
and U16323 (N_16323,N_2745,N_7522);
nand U16324 (N_16324,N_9413,N_7648);
nand U16325 (N_16325,N_8493,N_6496);
nor U16326 (N_16326,N_806,N_1191);
nor U16327 (N_16327,N_5067,N_9427);
or U16328 (N_16328,N_6247,N_9064);
nor U16329 (N_16329,N_9339,N_5630);
or U16330 (N_16330,N_9092,N_2987);
and U16331 (N_16331,N_357,N_3012);
nor U16332 (N_16332,N_5057,N_1944);
xnor U16333 (N_16333,N_3962,N_6809);
or U16334 (N_16334,N_50,N_8077);
nand U16335 (N_16335,N_3002,N_3680);
or U16336 (N_16336,N_5015,N_2592);
and U16337 (N_16337,N_5538,N_755);
and U16338 (N_16338,N_4705,N_9501);
or U16339 (N_16339,N_5493,N_979);
and U16340 (N_16340,N_2946,N_5701);
or U16341 (N_16341,N_8291,N_4931);
nor U16342 (N_16342,N_4959,N_4970);
or U16343 (N_16343,N_1836,N_7111);
nor U16344 (N_16344,N_3277,N_5234);
and U16345 (N_16345,N_6929,N_1028);
nand U16346 (N_16346,N_6777,N_4391);
or U16347 (N_16347,N_6495,N_5744);
and U16348 (N_16348,N_525,N_680);
or U16349 (N_16349,N_2749,N_6899);
xnor U16350 (N_16350,N_8745,N_9312);
or U16351 (N_16351,N_2536,N_1912);
nand U16352 (N_16352,N_2834,N_460);
and U16353 (N_16353,N_2200,N_4164);
nand U16354 (N_16354,N_7902,N_6759);
or U16355 (N_16355,N_516,N_7640);
or U16356 (N_16356,N_4865,N_2493);
nand U16357 (N_16357,N_9247,N_3474);
and U16358 (N_16358,N_724,N_2974);
nor U16359 (N_16359,N_2834,N_9923);
and U16360 (N_16360,N_7950,N_4387);
and U16361 (N_16361,N_7918,N_8407);
nor U16362 (N_16362,N_3898,N_7454);
xor U16363 (N_16363,N_6036,N_7126);
nand U16364 (N_16364,N_2807,N_879);
nand U16365 (N_16365,N_3190,N_9256);
or U16366 (N_16366,N_5378,N_7861);
nor U16367 (N_16367,N_3212,N_31);
and U16368 (N_16368,N_4899,N_1130);
and U16369 (N_16369,N_7454,N_4135);
or U16370 (N_16370,N_5084,N_2849);
nand U16371 (N_16371,N_2609,N_8359);
nand U16372 (N_16372,N_9904,N_2101);
nor U16373 (N_16373,N_350,N_3931);
and U16374 (N_16374,N_9420,N_1754);
or U16375 (N_16375,N_8910,N_8306);
nand U16376 (N_16376,N_1385,N_9136);
or U16377 (N_16377,N_8830,N_5482);
or U16378 (N_16378,N_7125,N_9036);
nor U16379 (N_16379,N_8822,N_5428);
and U16380 (N_16380,N_3109,N_7856);
nor U16381 (N_16381,N_3971,N_5802);
nand U16382 (N_16382,N_438,N_3023);
nor U16383 (N_16383,N_7486,N_8513);
nand U16384 (N_16384,N_9802,N_840);
nor U16385 (N_16385,N_1509,N_3127);
nor U16386 (N_16386,N_8482,N_6250);
nor U16387 (N_16387,N_3640,N_3839);
or U16388 (N_16388,N_9731,N_5449);
or U16389 (N_16389,N_370,N_4024);
and U16390 (N_16390,N_2467,N_8653);
nand U16391 (N_16391,N_1084,N_3362);
and U16392 (N_16392,N_2563,N_4550);
nor U16393 (N_16393,N_3333,N_6233);
nor U16394 (N_16394,N_3538,N_4248);
xnor U16395 (N_16395,N_8029,N_3989);
nand U16396 (N_16396,N_831,N_9160);
nand U16397 (N_16397,N_1120,N_2106);
or U16398 (N_16398,N_2050,N_7883);
or U16399 (N_16399,N_4691,N_2226);
nor U16400 (N_16400,N_7927,N_1230);
nor U16401 (N_16401,N_9887,N_6019);
or U16402 (N_16402,N_6852,N_6083);
nor U16403 (N_16403,N_9353,N_9583);
and U16404 (N_16404,N_2926,N_1525);
nor U16405 (N_16405,N_5270,N_209);
nor U16406 (N_16406,N_6171,N_3247);
nor U16407 (N_16407,N_4935,N_9248);
and U16408 (N_16408,N_863,N_7298);
nor U16409 (N_16409,N_1232,N_1572);
nor U16410 (N_16410,N_2442,N_641);
or U16411 (N_16411,N_7899,N_4772);
nand U16412 (N_16412,N_9796,N_4347);
and U16413 (N_16413,N_8577,N_1803);
or U16414 (N_16414,N_4601,N_6403);
nand U16415 (N_16415,N_1801,N_1887);
or U16416 (N_16416,N_5221,N_7535);
xor U16417 (N_16417,N_2326,N_8639);
nand U16418 (N_16418,N_9956,N_1167);
nor U16419 (N_16419,N_2198,N_3789);
and U16420 (N_16420,N_3713,N_5801);
and U16421 (N_16421,N_7007,N_2631);
and U16422 (N_16422,N_7011,N_630);
and U16423 (N_16423,N_889,N_2819);
nand U16424 (N_16424,N_132,N_1346);
or U16425 (N_16425,N_9651,N_2453);
xnor U16426 (N_16426,N_4834,N_2017);
nor U16427 (N_16427,N_2609,N_5549);
or U16428 (N_16428,N_9382,N_1181);
nand U16429 (N_16429,N_5981,N_197);
and U16430 (N_16430,N_3787,N_3696);
nor U16431 (N_16431,N_3415,N_6012);
xnor U16432 (N_16432,N_7300,N_3602);
or U16433 (N_16433,N_3871,N_165);
and U16434 (N_16434,N_8507,N_3536);
xor U16435 (N_16435,N_1283,N_2262);
or U16436 (N_16436,N_6349,N_5242);
nor U16437 (N_16437,N_7077,N_4172);
or U16438 (N_16438,N_5933,N_7758);
nor U16439 (N_16439,N_890,N_442);
nor U16440 (N_16440,N_9731,N_2424);
nand U16441 (N_16441,N_1177,N_4746);
and U16442 (N_16442,N_8736,N_1908);
and U16443 (N_16443,N_2563,N_7816);
xor U16444 (N_16444,N_6892,N_7510);
nand U16445 (N_16445,N_6924,N_1505);
or U16446 (N_16446,N_1054,N_9296);
or U16447 (N_16447,N_961,N_7449);
or U16448 (N_16448,N_8949,N_2119);
nand U16449 (N_16449,N_1917,N_6035);
xor U16450 (N_16450,N_4510,N_2612);
nand U16451 (N_16451,N_4616,N_1707);
xnor U16452 (N_16452,N_6431,N_1663);
and U16453 (N_16453,N_1090,N_3463);
and U16454 (N_16454,N_4731,N_5010);
or U16455 (N_16455,N_8381,N_2107);
xnor U16456 (N_16456,N_974,N_4382);
nand U16457 (N_16457,N_6546,N_6344);
xor U16458 (N_16458,N_8152,N_5281);
nand U16459 (N_16459,N_8326,N_4965);
or U16460 (N_16460,N_6476,N_8475);
nor U16461 (N_16461,N_7079,N_6672);
and U16462 (N_16462,N_4175,N_9417);
nand U16463 (N_16463,N_4000,N_2672);
and U16464 (N_16464,N_3320,N_6858);
nor U16465 (N_16465,N_6322,N_9502);
nor U16466 (N_16466,N_6135,N_9926);
xnor U16467 (N_16467,N_6707,N_7727);
and U16468 (N_16468,N_8068,N_5700);
nor U16469 (N_16469,N_8649,N_4337);
or U16470 (N_16470,N_3829,N_8280);
nand U16471 (N_16471,N_8069,N_6337);
or U16472 (N_16472,N_1340,N_321);
or U16473 (N_16473,N_8758,N_2755);
and U16474 (N_16474,N_455,N_9802);
nand U16475 (N_16475,N_5011,N_7336);
or U16476 (N_16476,N_5786,N_9147);
nand U16477 (N_16477,N_6276,N_8871);
or U16478 (N_16478,N_8766,N_8314);
xor U16479 (N_16479,N_5736,N_4883);
or U16480 (N_16480,N_9992,N_2699);
xor U16481 (N_16481,N_6248,N_3994);
nor U16482 (N_16482,N_3237,N_6476);
or U16483 (N_16483,N_969,N_9091);
and U16484 (N_16484,N_8941,N_8358);
and U16485 (N_16485,N_8649,N_1255);
and U16486 (N_16486,N_5739,N_6527);
and U16487 (N_16487,N_1613,N_1845);
or U16488 (N_16488,N_8389,N_4219);
and U16489 (N_16489,N_801,N_9191);
nand U16490 (N_16490,N_8058,N_1819);
and U16491 (N_16491,N_6821,N_238);
and U16492 (N_16492,N_2064,N_570);
and U16493 (N_16493,N_3577,N_8385);
and U16494 (N_16494,N_6834,N_6646);
nand U16495 (N_16495,N_5032,N_5234);
nor U16496 (N_16496,N_3328,N_3886);
xnor U16497 (N_16497,N_8491,N_4944);
nor U16498 (N_16498,N_3119,N_6887);
and U16499 (N_16499,N_2151,N_7889);
nor U16500 (N_16500,N_2887,N_9099);
nor U16501 (N_16501,N_180,N_945);
nor U16502 (N_16502,N_9675,N_7001);
nor U16503 (N_16503,N_2756,N_1912);
and U16504 (N_16504,N_7340,N_9889);
and U16505 (N_16505,N_5516,N_1737);
and U16506 (N_16506,N_7032,N_4665);
and U16507 (N_16507,N_6742,N_1874);
or U16508 (N_16508,N_8684,N_3267);
or U16509 (N_16509,N_3684,N_517);
and U16510 (N_16510,N_4215,N_4295);
and U16511 (N_16511,N_977,N_8180);
and U16512 (N_16512,N_4975,N_2530);
or U16513 (N_16513,N_1694,N_4555);
or U16514 (N_16514,N_1164,N_7420);
nand U16515 (N_16515,N_3027,N_9314);
nand U16516 (N_16516,N_7911,N_3412);
nand U16517 (N_16517,N_2276,N_655);
nor U16518 (N_16518,N_8235,N_691);
or U16519 (N_16519,N_6140,N_754);
nand U16520 (N_16520,N_9304,N_5687);
or U16521 (N_16521,N_6071,N_1395);
nand U16522 (N_16522,N_5931,N_9037);
and U16523 (N_16523,N_9865,N_9267);
nor U16524 (N_16524,N_401,N_3494);
and U16525 (N_16525,N_1280,N_6962);
nor U16526 (N_16526,N_4415,N_7089);
and U16527 (N_16527,N_6256,N_3447);
xnor U16528 (N_16528,N_7853,N_8136);
nor U16529 (N_16529,N_6174,N_7786);
or U16530 (N_16530,N_8340,N_4179);
nand U16531 (N_16531,N_6906,N_9692);
xnor U16532 (N_16532,N_9811,N_5492);
or U16533 (N_16533,N_2661,N_2513);
nand U16534 (N_16534,N_9453,N_4213);
xor U16535 (N_16535,N_2668,N_6232);
nand U16536 (N_16536,N_8850,N_292);
and U16537 (N_16537,N_8814,N_3283);
nand U16538 (N_16538,N_4043,N_3112);
nand U16539 (N_16539,N_8160,N_2907);
nand U16540 (N_16540,N_1613,N_355);
nand U16541 (N_16541,N_2501,N_987);
and U16542 (N_16542,N_2363,N_8413);
nand U16543 (N_16543,N_350,N_5230);
and U16544 (N_16544,N_2177,N_9211);
or U16545 (N_16545,N_2301,N_1861);
xnor U16546 (N_16546,N_1070,N_542);
xnor U16547 (N_16547,N_3275,N_1513);
nor U16548 (N_16548,N_9809,N_7495);
or U16549 (N_16549,N_4460,N_8254);
and U16550 (N_16550,N_4025,N_5438);
nor U16551 (N_16551,N_9631,N_9206);
nor U16552 (N_16552,N_1654,N_2042);
and U16553 (N_16553,N_1973,N_1378);
or U16554 (N_16554,N_3704,N_1873);
nand U16555 (N_16555,N_6528,N_1278);
or U16556 (N_16556,N_7216,N_5809);
nand U16557 (N_16557,N_8831,N_9177);
and U16558 (N_16558,N_6226,N_1833);
xor U16559 (N_16559,N_2245,N_1822);
nor U16560 (N_16560,N_6340,N_9925);
or U16561 (N_16561,N_1973,N_9236);
nand U16562 (N_16562,N_7687,N_37);
nand U16563 (N_16563,N_6930,N_9589);
and U16564 (N_16564,N_4185,N_4160);
nand U16565 (N_16565,N_5584,N_8179);
nor U16566 (N_16566,N_9368,N_5703);
and U16567 (N_16567,N_5969,N_7978);
or U16568 (N_16568,N_5309,N_9759);
xor U16569 (N_16569,N_2659,N_3885);
nand U16570 (N_16570,N_2352,N_3853);
and U16571 (N_16571,N_4428,N_1479);
nor U16572 (N_16572,N_5868,N_3399);
nor U16573 (N_16573,N_7921,N_8526);
or U16574 (N_16574,N_4571,N_1619);
nor U16575 (N_16575,N_9478,N_0);
or U16576 (N_16576,N_7150,N_1715);
xnor U16577 (N_16577,N_651,N_8736);
nor U16578 (N_16578,N_5218,N_4784);
nor U16579 (N_16579,N_3298,N_3367);
or U16580 (N_16580,N_8302,N_5642);
or U16581 (N_16581,N_9235,N_7909);
xor U16582 (N_16582,N_5186,N_6092);
xnor U16583 (N_16583,N_1709,N_2180);
nor U16584 (N_16584,N_1659,N_6929);
nand U16585 (N_16585,N_9331,N_2714);
or U16586 (N_16586,N_6767,N_5002);
and U16587 (N_16587,N_5729,N_3010);
nor U16588 (N_16588,N_2887,N_1132);
nand U16589 (N_16589,N_6149,N_1271);
nand U16590 (N_16590,N_5712,N_1869);
nor U16591 (N_16591,N_2937,N_7913);
xor U16592 (N_16592,N_3959,N_2380);
or U16593 (N_16593,N_4760,N_5429);
or U16594 (N_16594,N_3380,N_6616);
nand U16595 (N_16595,N_8436,N_5621);
nor U16596 (N_16596,N_460,N_5025);
or U16597 (N_16597,N_5882,N_8549);
or U16598 (N_16598,N_5009,N_5188);
xnor U16599 (N_16599,N_2365,N_2530);
or U16600 (N_16600,N_2489,N_7144);
nor U16601 (N_16601,N_7946,N_9263);
nor U16602 (N_16602,N_2378,N_9023);
or U16603 (N_16603,N_482,N_3524);
nand U16604 (N_16604,N_455,N_6277);
and U16605 (N_16605,N_8863,N_1411);
or U16606 (N_16606,N_2370,N_3102);
nor U16607 (N_16607,N_8088,N_2148);
or U16608 (N_16608,N_7192,N_9312);
nor U16609 (N_16609,N_1319,N_2897);
and U16610 (N_16610,N_6266,N_7234);
and U16611 (N_16611,N_1461,N_2718);
or U16612 (N_16612,N_2260,N_5473);
or U16613 (N_16613,N_6212,N_2160);
and U16614 (N_16614,N_2546,N_9102);
nor U16615 (N_16615,N_6167,N_4432);
nand U16616 (N_16616,N_6487,N_7857);
nand U16617 (N_16617,N_4255,N_5695);
or U16618 (N_16618,N_8950,N_6632);
and U16619 (N_16619,N_7240,N_3075);
or U16620 (N_16620,N_8525,N_4863);
nor U16621 (N_16621,N_7854,N_5756);
and U16622 (N_16622,N_5740,N_3202);
nor U16623 (N_16623,N_2421,N_5863);
nor U16624 (N_16624,N_14,N_8057);
and U16625 (N_16625,N_9256,N_5596);
xor U16626 (N_16626,N_1827,N_97);
or U16627 (N_16627,N_8926,N_9587);
and U16628 (N_16628,N_7522,N_104);
and U16629 (N_16629,N_6686,N_9676);
nor U16630 (N_16630,N_145,N_1689);
and U16631 (N_16631,N_9817,N_2003);
nand U16632 (N_16632,N_2435,N_78);
and U16633 (N_16633,N_3025,N_8403);
or U16634 (N_16634,N_3216,N_307);
or U16635 (N_16635,N_8777,N_8897);
or U16636 (N_16636,N_8112,N_2461);
nor U16637 (N_16637,N_5765,N_1410);
nor U16638 (N_16638,N_2612,N_5171);
nand U16639 (N_16639,N_8523,N_6741);
and U16640 (N_16640,N_3030,N_4972);
or U16641 (N_16641,N_5700,N_8820);
nand U16642 (N_16642,N_3887,N_6534);
or U16643 (N_16643,N_1700,N_3744);
or U16644 (N_16644,N_764,N_4263);
nor U16645 (N_16645,N_6953,N_9211);
nor U16646 (N_16646,N_9509,N_5536);
nor U16647 (N_16647,N_313,N_3484);
xor U16648 (N_16648,N_4240,N_8881);
or U16649 (N_16649,N_7509,N_1723);
nand U16650 (N_16650,N_7650,N_3918);
nor U16651 (N_16651,N_2926,N_6037);
nor U16652 (N_16652,N_2138,N_1013);
and U16653 (N_16653,N_7921,N_6205);
and U16654 (N_16654,N_377,N_5170);
nor U16655 (N_16655,N_737,N_3814);
or U16656 (N_16656,N_8533,N_5465);
nand U16657 (N_16657,N_2154,N_6987);
and U16658 (N_16658,N_1898,N_6823);
nor U16659 (N_16659,N_1995,N_6061);
or U16660 (N_16660,N_273,N_1095);
nor U16661 (N_16661,N_6186,N_6880);
nand U16662 (N_16662,N_897,N_7811);
and U16663 (N_16663,N_9544,N_9494);
and U16664 (N_16664,N_2206,N_3023);
nand U16665 (N_16665,N_2141,N_797);
and U16666 (N_16666,N_9461,N_8761);
nand U16667 (N_16667,N_8544,N_9967);
xnor U16668 (N_16668,N_6391,N_2353);
or U16669 (N_16669,N_1602,N_5901);
xor U16670 (N_16670,N_1124,N_7103);
or U16671 (N_16671,N_1582,N_4667);
or U16672 (N_16672,N_6967,N_5429);
nand U16673 (N_16673,N_8313,N_8365);
or U16674 (N_16674,N_6231,N_434);
nand U16675 (N_16675,N_7989,N_5772);
nor U16676 (N_16676,N_9318,N_9390);
nand U16677 (N_16677,N_6772,N_3905);
or U16678 (N_16678,N_4398,N_2090);
nand U16679 (N_16679,N_5452,N_7625);
and U16680 (N_16680,N_1503,N_2955);
and U16681 (N_16681,N_9370,N_8932);
nand U16682 (N_16682,N_980,N_3764);
nor U16683 (N_16683,N_7491,N_9707);
nor U16684 (N_16684,N_8467,N_2517);
nand U16685 (N_16685,N_6556,N_2377);
nand U16686 (N_16686,N_9742,N_8366);
and U16687 (N_16687,N_1001,N_7833);
nand U16688 (N_16688,N_5189,N_6281);
xor U16689 (N_16689,N_7682,N_8062);
and U16690 (N_16690,N_8208,N_144);
or U16691 (N_16691,N_5461,N_2587);
xnor U16692 (N_16692,N_1781,N_2217);
nand U16693 (N_16693,N_5271,N_9823);
xor U16694 (N_16694,N_1341,N_9183);
nor U16695 (N_16695,N_5549,N_90);
and U16696 (N_16696,N_6987,N_8365);
and U16697 (N_16697,N_5893,N_6590);
nor U16698 (N_16698,N_5111,N_1569);
xnor U16699 (N_16699,N_6408,N_5258);
or U16700 (N_16700,N_6448,N_6845);
or U16701 (N_16701,N_7436,N_4114);
nor U16702 (N_16702,N_4207,N_2509);
and U16703 (N_16703,N_2498,N_3242);
or U16704 (N_16704,N_7457,N_2614);
nand U16705 (N_16705,N_4011,N_6262);
nand U16706 (N_16706,N_3942,N_7436);
nor U16707 (N_16707,N_4656,N_5590);
nor U16708 (N_16708,N_9206,N_6774);
nand U16709 (N_16709,N_8450,N_6591);
nor U16710 (N_16710,N_1876,N_860);
nand U16711 (N_16711,N_3179,N_6613);
nor U16712 (N_16712,N_7538,N_8824);
and U16713 (N_16713,N_7874,N_8959);
and U16714 (N_16714,N_5758,N_1358);
nor U16715 (N_16715,N_8160,N_9646);
nor U16716 (N_16716,N_4382,N_4659);
nand U16717 (N_16717,N_3918,N_8855);
and U16718 (N_16718,N_3206,N_4667);
nand U16719 (N_16719,N_4849,N_994);
nand U16720 (N_16720,N_7014,N_9040);
nor U16721 (N_16721,N_88,N_3265);
or U16722 (N_16722,N_3957,N_8825);
nand U16723 (N_16723,N_410,N_8963);
xor U16724 (N_16724,N_9248,N_3451);
nand U16725 (N_16725,N_8183,N_1011);
nor U16726 (N_16726,N_6389,N_2071);
or U16727 (N_16727,N_9023,N_597);
nand U16728 (N_16728,N_7021,N_6868);
nor U16729 (N_16729,N_327,N_5659);
nor U16730 (N_16730,N_4370,N_2358);
nor U16731 (N_16731,N_8087,N_3689);
and U16732 (N_16732,N_1364,N_2132);
nand U16733 (N_16733,N_2820,N_7998);
xor U16734 (N_16734,N_8749,N_4619);
and U16735 (N_16735,N_1081,N_1026);
nand U16736 (N_16736,N_1747,N_6705);
nand U16737 (N_16737,N_6174,N_886);
nor U16738 (N_16738,N_8596,N_9714);
and U16739 (N_16739,N_6607,N_3552);
nor U16740 (N_16740,N_9992,N_3291);
nor U16741 (N_16741,N_8924,N_807);
nor U16742 (N_16742,N_8523,N_8396);
or U16743 (N_16743,N_3363,N_7397);
nor U16744 (N_16744,N_8530,N_912);
nor U16745 (N_16745,N_6553,N_8611);
nor U16746 (N_16746,N_976,N_5917);
nor U16747 (N_16747,N_9592,N_6092);
or U16748 (N_16748,N_1177,N_3381);
and U16749 (N_16749,N_4875,N_7068);
nor U16750 (N_16750,N_2238,N_7423);
nor U16751 (N_16751,N_5834,N_2970);
nor U16752 (N_16752,N_6745,N_2702);
and U16753 (N_16753,N_4893,N_5482);
or U16754 (N_16754,N_1895,N_1400);
xnor U16755 (N_16755,N_8794,N_9171);
and U16756 (N_16756,N_1155,N_1706);
and U16757 (N_16757,N_6990,N_3012);
xor U16758 (N_16758,N_9315,N_8271);
nand U16759 (N_16759,N_8533,N_5615);
or U16760 (N_16760,N_1577,N_3321);
nand U16761 (N_16761,N_9453,N_1439);
or U16762 (N_16762,N_5780,N_4065);
or U16763 (N_16763,N_6578,N_4561);
nand U16764 (N_16764,N_9230,N_7920);
or U16765 (N_16765,N_7435,N_5443);
nor U16766 (N_16766,N_9734,N_7053);
nand U16767 (N_16767,N_6921,N_9398);
or U16768 (N_16768,N_7641,N_4526);
and U16769 (N_16769,N_373,N_3130);
or U16770 (N_16770,N_6283,N_1611);
and U16771 (N_16771,N_9618,N_7129);
or U16772 (N_16772,N_1752,N_8360);
or U16773 (N_16773,N_776,N_6997);
or U16774 (N_16774,N_1107,N_7693);
nand U16775 (N_16775,N_7318,N_9597);
or U16776 (N_16776,N_5923,N_476);
or U16777 (N_16777,N_2528,N_6949);
nand U16778 (N_16778,N_5054,N_2294);
nor U16779 (N_16779,N_6949,N_3323);
xor U16780 (N_16780,N_3476,N_8617);
nor U16781 (N_16781,N_9058,N_4580);
nand U16782 (N_16782,N_4819,N_2016);
nor U16783 (N_16783,N_5660,N_1141);
or U16784 (N_16784,N_3968,N_1349);
nor U16785 (N_16785,N_1888,N_3662);
and U16786 (N_16786,N_5562,N_3861);
and U16787 (N_16787,N_3939,N_7000);
nand U16788 (N_16788,N_1365,N_8974);
and U16789 (N_16789,N_7253,N_3253);
nor U16790 (N_16790,N_68,N_1408);
and U16791 (N_16791,N_2473,N_1772);
nor U16792 (N_16792,N_6155,N_7041);
and U16793 (N_16793,N_8705,N_7306);
nand U16794 (N_16794,N_2830,N_513);
nor U16795 (N_16795,N_9815,N_9248);
nand U16796 (N_16796,N_2732,N_5557);
nor U16797 (N_16797,N_2793,N_4894);
nor U16798 (N_16798,N_3390,N_9168);
xnor U16799 (N_16799,N_5644,N_8579);
nor U16800 (N_16800,N_4636,N_9355);
nand U16801 (N_16801,N_6638,N_2791);
nor U16802 (N_16802,N_6452,N_8022);
or U16803 (N_16803,N_9042,N_8231);
nor U16804 (N_16804,N_3914,N_3447);
or U16805 (N_16805,N_5126,N_4777);
nor U16806 (N_16806,N_118,N_5832);
and U16807 (N_16807,N_1495,N_7587);
nor U16808 (N_16808,N_4073,N_3936);
nand U16809 (N_16809,N_3759,N_6572);
nor U16810 (N_16810,N_4175,N_1554);
nand U16811 (N_16811,N_8449,N_2207);
nor U16812 (N_16812,N_1286,N_1650);
nor U16813 (N_16813,N_7518,N_6185);
and U16814 (N_16814,N_983,N_813);
or U16815 (N_16815,N_3181,N_2020);
and U16816 (N_16816,N_477,N_3335);
and U16817 (N_16817,N_6432,N_8616);
nor U16818 (N_16818,N_3831,N_1753);
nand U16819 (N_16819,N_1662,N_8838);
or U16820 (N_16820,N_3287,N_3614);
and U16821 (N_16821,N_3220,N_3427);
nor U16822 (N_16822,N_8370,N_3379);
or U16823 (N_16823,N_1736,N_6738);
xor U16824 (N_16824,N_9296,N_4738);
nand U16825 (N_16825,N_2279,N_9111);
nor U16826 (N_16826,N_7727,N_4654);
nor U16827 (N_16827,N_2652,N_1348);
xor U16828 (N_16828,N_5370,N_7296);
or U16829 (N_16829,N_7717,N_4926);
nand U16830 (N_16830,N_4592,N_1224);
nand U16831 (N_16831,N_4101,N_1619);
nand U16832 (N_16832,N_3156,N_4574);
nor U16833 (N_16833,N_7532,N_1397);
nor U16834 (N_16834,N_4998,N_8865);
or U16835 (N_16835,N_9434,N_9815);
and U16836 (N_16836,N_532,N_5490);
and U16837 (N_16837,N_9920,N_5040);
or U16838 (N_16838,N_716,N_8367);
and U16839 (N_16839,N_7363,N_6992);
and U16840 (N_16840,N_5526,N_6626);
nand U16841 (N_16841,N_5165,N_7980);
nor U16842 (N_16842,N_6042,N_374);
and U16843 (N_16843,N_1487,N_8839);
or U16844 (N_16844,N_9787,N_5114);
nand U16845 (N_16845,N_3084,N_3916);
or U16846 (N_16846,N_747,N_7358);
and U16847 (N_16847,N_3949,N_1972);
nor U16848 (N_16848,N_4144,N_664);
and U16849 (N_16849,N_8289,N_1755);
nand U16850 (N_16850,N_6837,N_2333);
and U16851 (N_16851,N_4602,N_1841);
or U16852 (N_16852,N_1624,N_2147);
nor U16853 (N_16853,N_8336,N_715);
nor U16854 (N_16854,N_6849,N_5892);
or U16855 (N_16855,N_3734,N_8397);
and U16856 (N_16856,N_9071,N_7564);
and U16857 (N_16857,N_8542,N_1686);
or U16858 (N_16858,N_2768,N_1721);
or U16859 (N_16859,N_9411,N_7457);
and U16860 (N_16860,N_6185,N_7895);
or U16861 (N_16861,N_6711,N_9369);
or U16862 (N_16862,N_5325,N_5025);
and U16863 (N_16863,N_9460,N_3024);
nor U16864 (N_16864,N_8733,N_8791);
nor U16865 (N_16865,N_9053,N_8339);
nand U16866 (N_16866,N_7457,N_4009);
and U16867 (N_16867,N_809,N_3915);
nand U16868 (N_16868,N_1652,N_5759);
or U16869 (N_16869,N_9910,N_142);
nand U16870 (N_16870,N_66,N_7774);
nand U16871 (N_16871,N_4921,N_5441);
and U16872 (N_16872,N_4322,N_978);
nor U16873 (N_16873,N_6901,N_2939);
nand U16874 (N_16874,N_8125,N_5843);
and U16875 (N_16875,N_2052,N_6335);
nand U16876 (N_16876,N_7152,N_1360);
nor U16877 (N_16877,N_6873,N_3513);
nor U16878 (N_16878,N_8619,N_388);
or U16879 (N_16879,N_3017,N_9197);
nor U16880 (N_16880,N_6702,N_6090);
or U16881 (N_16881,N_3704,N_5582);
nand U16882 (N_16882,N_4196,N_8476);
and U16883 (N_16883,N_7663,N_5838);
xnor U16884 (N_16884,N_3466,N_8206);
nand U16885 (N_16885,N_2804,N_6975);
or U16886 (N_16886,N_5444,N_8783);
or U16887 (N_16887,N_4601,N_9297);
nand U16888 (N_16888,N_2607,N_5798);
or U16889 (N_16889,N_7674,N_1667);
nor U16890 (N_16890,N_9534,N_1236);
nor U16891 (N_16891,N_821,N_1964);
and U16892 (N_16892,N_3104,N_8688);
xor U16893 (N_16893,N_4229,N_5734);
nor U16894 (N_16894,N_2864,N_4534);
nor U16895 (N_16895,N_4980,N_6562);
or U16896 (N_16896,N_8989,N_5893);
nand U16897 (N_16897,N_7637,N_2613);
and U16898 (N_16898,N_9391,N_9509);
and U16899 (N_16899,N_8468,N_7790);
and U16900 (N_16900,N_4277,N_2092);
or U16901 (N_16901,N_8454,N_8382);
nand U16902 (N_16902,N_572,N_6546);
nand U16903 (N_16903,N_3094,N_8240);
nand U16904 (N_16904,N_1247,N_5925);
and U16905 (N_16905,N_4373,N_6052);
xor U16906 (N_16906,N_5652,N_9039);
and U16907 (N_16907,N_4206,N_4848);
and U16908 (N_16908,N_6986,N_1138);
nor U16909 (N_16909,N_2108,N_2890);
nor U16910 (N_16910,N_2461,N_8713);
and U16911 (N_16911,N_7791,N_95);
or U16912 (N_16912,N_6114,N_4875);
and U16913 (N_16913,N_1475,N_4242);
or U16914 (N_16914,N_3306,N_7419);
or U16915 (N_16915,N_9356,N_3446);
and U16916 (N_16916,N_2952,N_4463);
nor U16917 (N_16917,N_4653,N_2426);
xnor U16918 (N_16918,N_6172,N_847);
nor U16919 (N_16919,N_5959,N_3772);
and U16920 (N_16920,N_7037,N_1497);
nor U16921 (N_16921,N_6721,N_143);
nand U16922 (N_16922,N_3702,N_7359);
and U16923 (N_16923,N_9033,N_7912);
nor U16924 (N_16924,N_5985,N_5718);
nand U16925 (N_16925,N_3965,N_2972);
and U16926 (N_16926,N_691,N_4574);
and U16927 (N_16927,N_3382,N_8646);
nand U16928 (N_16928,N_2314,N_6174);
xnor U16929 (N_16929,N_8105,N_6847);
nand U16930 (N_16930,N_1022,N_8603);
and U16931 (N_16931,N_4600,N_2814);
nor U16932 (N_16932,N_6820,N_9118);
xor U16933 (N_16933,N_4468,N_7730);
and U16934 (N_16934,N_2253,N_6467);
and U16935 (N_16935,N_8850,N_6678);
or U16936 (N_16936,N_7338,N_9264);
and U16937 (N_16937,N_7881,N_5833);
nand U16938 (N_16938,N_2917,N_3426);
or U16939 (N_16939,N_1397,N_9269);
xnor U16940 (N_16940,N_3194,N_6313);
nand U16941 (N_16941,N_9170,N_6789);
or U16942 (N_16942,N_9201,N_5226);
or U16943 (N_16943,N_6539,N_3176);
or U16944 (N_16944,N_694,N_9277);
nand U16945 (N_16945,N_9414,N_4834);
nand U16946 (N_16946,N_2306,N_2131);
nand U16947 (N_16947,N_1457,N_6102);
and U16948 (N_16948,N_4782,N_3543);
nand U16949 (N_16949,N_56,N_84);
and U16950 (N_16950,N_5745,N_8447);
or U16951 (N_16951,N_4190,N_1375);
nand U16952 (N_16952,N_4435,N_8726);
or U16953 (N_16953,N_8686,N_9185);
or U16954 (N_16954,N_8194,N_6372);
and U16955 (N_16955,N_3392,N_1917);
nor U16956 (N_16956,N_1719,N_6161);
xnor U16957 (N_16957,N_4279,N_5394);
and U16958 (N_16958,N_3009,N_5497);
and U16959 (N_16959,N_7594,N_4524);
nand U16960 (N_16960,N_896,N_7157);
nand U16961 (N_16961,N_2091,N_5000);
or U16962 (N_16962,N_784,N_5224);
or U16963 (N_16963,N_5436,N_5240);
or U16964 (N_16964,N_8441,N_2063);
nand U16965 (N_16965,N_9976,N_5871);
nor U16966 (N_16966,N_3047,N_7836);
and U16967 (N_16967,N_7044,N_2216);
or U16968 (N_16968,N_7946,N_1203);
nand U16969 (N_16969,N_7336,N_7518);
nand U16970 (N_16970,N_7841,N_2850);
nor U16971 (N_16971,N_7353,N_5581);
or U16972 (N_16972,N_2639,N_5682);
and U16973 (N_16973,N_374,N_127);
nand U16974 (N_16974,N_7716,N_5338);
or U16975 (N_16975,N_1661,N_9957);
nor U16976 (N_16976,N_5240,N_507);
xor U16977 (N_16977,N_6644,N_6769);
nand U16978 (N_16978,N_9061,N_9523);
nor U16979 (N_16979,N_6518,N_2825);
or U16980 (N_16980,N_212,N_8108);
nand U16981 (N_16981,N_3205,N_7448);
or U16982 (N_16982,N_8119,N_6729);
nand U16983 (N_16983,N_5061,N_8510);
and U16984 (N_16984,N_4846,N_4028);
and U16985 (N_16985,N_3401,N_1153);
nor U16986 (N_16986,N_6984,N_4369);
nor U16987 (N_16987,N_3244,N_8386);
and U16988 (N_16988,N_2230,N_8091);
nor U16989 (N_16989,N_2296,N_4029);
or U16990 (N_16990,N_6683,N_2534);
and U16991 (N_16991,N_8351,N_2734);
nor U16992 (N_16992,N_1726,N_2606);
nor U16993 (N_16993,N_5022,N_4881);
and U16994 (N_16994,N_1120,N_1100);
xor U16995 (N_16995,N_1809,N_817);
nand U16996 (N_16996,N_2414,N_1599);
or U16997 (N_16997,N_8686,N_4810);
nand U16998 (N_16998,N_6749,N_8399);
or U16999 (N_16999,N_6376,N_7646);
and U17000 (N_17000,N_1757,N_1677);
nand U17001 (N_17001,N_1182,N_2191);
nor U17002 (N_17002,N_1916,N_1012);
or U17003 (N_17003,N_3035,N_9895);
xnor U17004 (N_17004,N_5167,N_5714);
and U17005 (N_17005,N_761,N_7481);
nand U17006 (N_17006,N_3925,N_2156);
nand U17007 (N_17007,N_1859,N_1342);
nand U17008 (N_17008,N_2383,N_6907);
nand U17009 (N_17009,N_5334,N_182);
nor U17010 (N_17010,N_9116,N_6541);
nand U17011 (N_17011,N_8738,N_475);
and U17012 (N_17012,N_8515,N_9954);
xor U17013 (N_17013,N_5861,N_9910);
xnor U17014 (N_17014,N_3222,N_8943);
nand U17015 (N_17015,N_2708,N_5580);
nor U17016 (N_17016,N_9892,N_261);
nand U17017 (N_17017,N_8505,N_6826);
or U17018 (N_17018,N_6359,N_4836);
nor U17019 (N_17019,N_9405,N_1945);
or U17020 (N_17020,N_5087,N_804);
and U17021 (N_17021,N_8811,N_6249);
and U17022 (N_17022,N_416,N_6292);
nand U17023 (N_17023,N_5979,N_1318);
nand U17024 (N_17024,N_3184,N_6838);
nand U17025 (N_17025,N_6538,N_4932);
nor U17026 (N_17026,N_4128,N_7821);
or U17027 (N_17027,N_8242,N_3944);
or U17028 (N_17028,N_1220,N_4163);
nand U17029 (N_17029,N_6551,N_8591);
and U17030 (N_17030,N_6169,N_7146);
xnor U17031 (N_17031,N_5777,N_2396);
nor U17032 (N_17032,N_914,N_7259);
or U17033 (N_17033,N_1104,N_9914);
or U17034 (N_17034,N_4270,N_9191);
nor U17035 (N_17035,N_8522,N_6130);
and U17036 (N_17036,N_8086,N_2515);
nor U17037 (N_17037,N_6117,N_7087);
xnor U17038 (N_17038,N_1222,N_4052);
and U17039 (N_17039,N_1687,N_6018);
xnor U17040 (N_17040,N_9192,N_6783);
nor U17041 (N_17041,N_5443,N_6605);
nor U17042 (N_17042,N_2546,N_1582);
nor U17043 (N_17043,N_8826,N_3952);
and U17044 (N_17044,N_7845,N_674);
nand U17045 (N_17045,N_3279,N_4625);
nand U17046 (N_17046,N_3977,N_7382);
and U17047 (N_17047,N_7201,N_6349);
or U17048 (N_17048,N_3567,N_652);
nor U17049 (N_17049,N_4419,N_4997);
nor U17050 (N_17050,N_4144,N_3680);
nor U17051 (N_17051,N_8364,N_3286);
nor U17052 (N_17052,N_2621,N_8347);
or U17053 (N_17053,N_8624,N_102);
nor U17054 (N_17054,N_449,N_5868);
or U17055 (N_17055,N_2723,N_6760);
and U17056 (N_17056,N_8879,N_1941);
and U17057 (N_17057,N_1055,N_9964);
and U17058 (N_17058,N_7644,N_2166);
nand U17059 (N_17059,N_9570,N_4347);
nor U17060 (N_17060,N_7821,N_3975);
xor U17061 (N_17061,N_2029,N_5736);
or U17062 (N_17062,N_8120,N_4605);
nand U17063 (N_17063,N_1229,N_4665);
or U17064 (N_17064,N_4130,N_5448);
nand U17065 (N_17065,N_5552,N_2757);
and U17066 (N_17066,N_6141,N_7935);
xor U17067 (N_17067,N_6649,N_7051);
nor U17068 (N_17068,N_6550,N_5560);
nand U17069 (N_17069,N_4151,N_7357);
and U17070 (N_17070,N_7341,N_9613);
and U17071 (N_17071,N_5269,N_7603);
nor U17072 (N_17072,N_7421,N_7548);
xor U17073 (N_17073,N_2992,N_657);
nor U17074 (N_17074,N_2952,N_5237);
nand U17075 (N_17075,N_2325,N_3030);
xor U17076 (N_17076,N_863,N_7529);
and U17077 (N_17077,N_6189,N_6272);
nor U17078 (N_17078,N_7583,N_2027);
or U17079 (N_17079,N_6690,N_3052);
and U17080 (N_17080,N_2822,N_8328);
nor U17081 (N_17081,N_2666,N_7085);
nor U17082 (N_17082,N_1795,N_2680);
or U17083 (N_17083,N_6643,N_6915);
or U17084 (N_17084,N_8729,N_5180);
and U17085 (N_17085,N_3853,N_2927);
and U17086 (N_17086,N_3217,N_8507);
or U17087 (N_17087,N_7083,N_3664);
or U17088 (N_17088,N_4877,N_1405);
and U17089 (N_17089,N_7765,N_4668);
xnor U17090 (N_17090,N_4419,N_5696);
nor U17091 (N_17091,N_6288,N_7887);
nand U17092 (N_17092,N_1039,N_4716);
nor U17093 (N_17093,N_8876,N_9440);
or U17094 (N_17094,N_8881,N_8473);
xnor U17095 (N_17095,N_1788,N_6547);
and U17096 (N_17096,N_4738,N_762);
or U17097 (N_17097,N_2258,N_5791);
and U17098 (N_17098,N_5622,N_4459);
or U17099 (N_17099,N_2666,N_5979);
or U17100 (N_17100,N_4987,N_2515);
or U17101 (N_17101,N_3610,N_6825);
or U17102 (N_17102,N_2405,N_4803);
nand U17103 (N_17103,N_5750,N_2450);
and U17104 (N_17104,N_3276,N_3942);
nor U17105 (N_17105,N_4810,N_1054);
nand U17106 (N_17106,N_9593,N_1338);
and U17107 (N_17107,N_6021,N_6969);
nor U17108 (N_17108,N_5795,N_8451);
nor U17109 (N_17109,N_548,N_7890);
or U17110 (N_17110,N_3348,N_1044);
nand U17111 (N_17111,N_868,N_2179);
nor U17112 (N_17112,N_5071,N_2070);
nand U17113 (N_17113,N_888,N_2127);
or U17114 (N_17114,N_1364,N_8498);
or U17115 (N_17115,N_792,N_4723);
and U17116 (N_17116,N_7266,N_2745);
and U17117 (N_17117,N_7011,N_9909);
and U17118 (N_17118,N_3728,N_8297);
nor U17119 (N_17119,N_5829,N_2495);
nand U17120 (N_17120,N_6151,N_6908);
nand U17121 (N_17121,N_99,N_1107);
or U17122 (N_17122,N_9324,N_9071);
and U17123 (N_17123,N_5348,N_6312);
nand U17124 (N_17124,N_5604,N_7317);
or U17125 (N_17125,N_8033,N_4968);
and U17126 (N_17126,N_8617,N_5850);
and U17127 (N_17127,N_1763,N_3062);
nand U17128 (N_17128,N_5209,N_5651);
nor U17129 (N_17129,N_7672,N_6750);
nand U17130 (N_17130,N_2164,N_8711);
and U17131 (N_17131,N_1832,N_3719);
nand U17132 (N_17132,N_1172,N_1313);
nor U17133 (N_17133,N_1118,N_8102);
nand U17134 (N_17134,N_9132,N_8859);
nand U17135 (N_17135,N_3663,N_3001);
nand U17136 (N_17136,N_2594,N_2674);
nor U17137 (N_17137,N_3612,N_6416);
nand U17138 (N_17138,N_7883,N_579);
or U17139 (N_17139,N_550,N_7391);
nor U17140 (N_17140,N_8788,N_7547);
and U17141 (N_17141,N_2288,N_7755);
xnor U17142 (N_17142,N_3326,N_3341);
nor U17143 (N_17143,N_9707,N_333);
or U17144 (N_17144,N_147,N_5089);
and U17145 (N_17145,N_4356,N_4166);
nor U17146 (N_17146,N_7490,N_9668);
nand U17147 (N_17147,N_142,N_5128);
nor U17148 (N_17148,N_6394,N_191);
xnor U17149 (N_17149,N_1388,N_1139);
or U17150 (N_17150,N_1577,N_3260);
xnor U17151 (N_17151,N_9375,N_9337);
nor U17152 (N_17152,N_5283,N_4049);
nor U17153 (N_17153,N_6727,N_5986);
xor U17154 (N_17154,N_3468,N_671);
xor U17155 (N_17155,N_3925,N_1457);
nand U17156 (N_17156,N_8977,N_5917);
xnor U17157 (N_17157,N_7238,N_3070);
nand U17158 (N_17158,N_4893,N_7700);
and U17159 (N_17159,N_9069,N_535);
nor U17160 (N_17160,N_2463,N_2682);
nand U17161 (N_17161,N_5184,N_6745);
nand U17162 (N_17162,N_138,N_2176);
and U17163 (N_17163,N_8221,N_2727);
and U17164 (N_17164,N_4795,N_1685);
nand U17165 (N_17165,N_8942,N_4282);
and U17166 (N_17166,N_3962,N_8198);
nand U17167 (N_17167,N_3917,N_8980);
and U17168 (N_17168,N_2806,N_4460);
nand U17169 (N_17169,N_3802,N_3601);
xor U17170 (N_17170,N_7682,N_5284);
nand U17171 (N_17171,N_8091,N_8880);
and U17172 (N_17172,N_9608,N_7652);
nor U17173 (N_17173,N_2184,N_340);
and U17174 (N_17174,N_6571,N_6643);
nor U17175 (N_17175,N_8221,N_4785);
nand U17176 (N_17176,N_6728,N_9598);
nor U17177 (N_17177,N_5344,N_3502);
nand U17178 (N_17178,N_891,N_4219);
nand U17179 (N_17179,N_4159,N_8362);
xnor U17180 (N_17180,N_5804,N_6957);
and U17181 (N_17181,N_9596,N_1870);
nand U17182 (N_17182,N_3090,N_3552);
and U17183 (N_17183,N_9527,N_6064);
or U17184 (N_17184,N_6497,N_6642);
nand U17185 (N_17185,N_1032,N_1490);
or U17186 (N_17186,N_4438,N_5788);
and U17187 (N_17187,N_5995,N_7708);
and U17188 (N_17188,N_9261,N_9710);
and U17189 (N_17189,N_4615,N_968);
nand U17190 (N_17190,N_2405,N_5308);
xnor U17191 (N_17191,N_3932,N_5228);
nor U17192 (N_17192,N_3164,N_8551);
nand U17193 (N_17193,N_2432,N_9684);
or U17194 (N_17194,N_6700,N_6820);
nor U17195 (N_17195,N_7347,N_1091);
and U17196 (N_17196,N_2887,N_7371);
nor U17197 (N_17197,N_5004,N_4310);
nor U17198 (N_17198,N_7322,N_287);
and U17199 (N_17199,N_9859,N_6582);
nor U17200 (N_17200,N_3716,N_983);
xnor U17201 (N_17201,N_6691,N_2735);
nand U17202 (N_17202,N_795,N_7129);
or U17203 (N_17203,N_6245,N_6304);
xnor U17204 (N_17204,N_8323,N_2312);
nand U17205 (N_17205,N_2802,N_3559);
and U17206 (N_17206,N_1472,N_5270);
xor U17207 (N_17207,N_1906,N_8110);
nor U17208 (N_17208,N_464,N_9299);
or U17209 (N_17209,N_2595,N_1051);
or U17210 (N_17210,N_5066,N_718);
xnor U17211 (N_17211,N_1872,N_8567);
nand U17212 (N_17212,N_9831,N_9828);
nor U17213 (N_17213,N_4802,N_1676);
nand U17214 (N_17214,N_3644,N_9001);
and U17215 (N_17215,N_5603,N_7391);
and U17216 (N_17216,N_2041,N_6457);
and U17217 (N_17217,N_4135,N_7491);
nor U17218 (N_17218,N_5193,N_4150);
nor U17219 (N_17219,N_4834,N_4285);
nand U17220 (N_17220,N_2803,N_2048);
and U17221 (N_17221,N_5167,N_8730);
nand U17222 (N_17222,N_3587,N_2843);
nor U17223 (N_17223,N_7488,N_7277);
xnor U17224 (N_17224,N_3808,N_8445);
nor U17225 (N_17225,N_6430,N_9157);
and U17226 (N_17226,N_9642,N_1343);
xnor U17227 (N_17227,N_5434,N_2501);
and U17228 (N_17228,N_5948,N_397);
or U17229 (N_17229,N_2065,N_8722);
nor U17230 (N_17230,N_2052,N_5311);
or U17231 (N_17231,N_3458,N_1922);
and U17232 (N_17232,N_9372,N_6834);
nand U17233 (N_17233,N_4560,N_8708);
or U17234 (N_17234,N_9725,N_528);
or U17235 (N_17235,N_6635,N_9114);
or U17236 (N_17236,N_3719,N_8351);
nand U17237 (N_17237,N_3850,N_6595);
xnor U17238 (N_17238,N_9917,N_8754);
nand U17239 (N_17239,N_7575,N_2495);
nor U17240 (N_17240,N_2338,N_464);
and U17241 (N_17241,N_4570,N_9136);
and U17242 (N_17242,N_1565,N_8763);
or U17243 (N_17243,N_3485,N_8426);
and U17244 (N_17244,N_9541,N_531);
nand U17245 (N_17245,N_7401,N_6248);
nand U17246 (N_17246,N_6391,N_9786);
or U17247 (N_17247,N_9256,N_6209);
nand U17248 (N_17248,N_4707,N_4904);
nor U17249 (N_17249,N_1335,N_1388);
xor U17250 (N_17250,N_7527,N_1307);
nand U17251 (N_17251,N_4825,N_1304);
or U17252 (N_17252,N_7960,N_190);
nand U17253 (N_17253,N_3148,N_4015);
and U17254 (N_17254,N_6611,N_8768);
nor U17255 (N_17255,N_3413,N_7485);
xnor U17256 (N_17256,N_170,N_7358);
or U17257 (N_17257,N_9910,N_6865);
and U17258 (N_17258,N_4558,N_6237);
xnor U17259 (N_17259,N_2650,N_6175);
or U17260 (N_17260,N_1103,N_941);
and U17261 (N_17261,N_7062,N_5606);
nand U17262 (N_17262,N_3685,N_1763);
nor U17263 (N_17263,N_7686,N_2276);
and U17264 (N_17264,N_634,N_330);
nor U17265 (N_17265,N_1152,N_4189);
nand U17266 (N_17266,N_3202,N_8345);
or U17267 (N_17267,N_6320,N_5039);
and U17268 (N_17268,N_915,N_3858);
nand U17269 (N_17269,N_5650,N_6345);
and U17270 (N_17270,N_7108,N_3254);
nand U17271 (N_17271,N_495,N_2409);
and U17272 (N_17272,N_7418,N_7976);
or U17273 (N_17273,N_6752,N_2829);
nor U17274 (N_17274,N_4454,N_4834);
nor U17275 (N_17275,N_9958,N_5461);
nand U17276 (N_17276,N_7086,N_9527);
nor U17277 (N_17277,N_7262,N_8305);
nand U17278 (N_17278,N_3167,N_9234);
nor U17279 (N_17279,N_5276,N_2098);
xor U17280 (N_17280,N_4579,N_218);
or U17281 (N_17281,N_3989,N_6588);
nand U17282 (N_17282,N_6725,N_9489);
or U17283 (N_17283,N_981,N_6062);
nor U17284 (N_17284,N_4639,N_1227);
nor U17285 (N_17285,N_7030,N_3746);
or U17286 (N_17286,N_5181,N_2045);
and U17287 (N_17287,N_543,N_9504);
and U17288 (N_17288,N_8413,N_4587);
nor U17289 (N_17289,N_7155,N_2609);
or U17290 (N_17290,N_4110,N_6607);
or U17291 (N_17291,N_8487,N_5402);
nand U17292 (N_17292,N_4392,N_5923);
and U17293 (N_17293,N_8617,N_6777);
nand U17294 (N_17294,N_762,N_2904);
nor U17295 (N_17295,N_5804,N_4209);
and U17296 (N_17296,N_7087,N_3689);
and U17297 (N_17297,N_1303,N_5900);
and U17298 (N_17298,N_2109,N_7130);
nand U17299 (N_17299,N_3630,N_1005);
or U17300 (N_17300,N_711,N_3496);
nor U17301 (N_17301,N_8315,N_5838);
nand U17302 (N_17302,N_2854,N_7082);
nor U17303 (N_17303,N_3696,N_4510);
and U17304 (N_17304,N_3922,N_8098);
nor U17305 (N_17305,N_3602,N_7672);
and U17306 (N_17306,N_9709,N_2784);
and U17307 (N_17307,N_1997,N_7580);
nor U17308 (N_17308,N_4051,N_3311);
or U17309 (N_17309,N_7892,N_9906);
and U17310 (N_17310,N_8451,N_7051);
nor U17311 (N_17311,N_9551,N_5179);
or U17312 (N_17312,N_9856,N_1216);
nor U17313 (N_17313,N_9542,N_9459);
or U17314 (N_17314,N_7737,N_6991);
xnor U17315 (N_17315,N_2448,N_8309);
and U17316 (N_17316,N_7168,N_7669);
and U17317 (N_17317,N_9370,N_133);
nor U17318 (N_17318,N_3881,N_4310);
or U17319 (N_17319,N_9476,N_760);
nand U17320 (N_17320,N_9184,N_207);
or U17321 (N_17321,N_9020,N_8684);
and U17322 (N_17322,N_6358,N_9646);
nor U17323 (N_17323,N_2068,N_5815);
nor U17324 (N_17324,N_5712,N_8099);
or U17325 (N_17325,N_5390,N_7595);
nand U17326 (N_17326,N_5522,N_4921);
xnor U17327 (N_17327,N_5872,N_5758);
and U17328 (N_17328,N_791,N_817);
nor U17329 (N_17329,N_8154,N_673);
nand U17330 (N_17330,N_4426,N_1027);
and U17331 (N_17331,N_5585,N_5547);
nand U17332 (N_17332,N_5366,N_3781);
nand U17333 (N_17333,N_4271,N_5290);
nor U17334 (N_17334,N_6763,N_3820);
nor U17335 (N_17335,N_3693,N_4343);
nand U17336 (N_17336,N_7540,N_276);
nor U17337 (N_17337,N_5579,N_8471);
or U17338 (N_17338,N_8341,N_1046);
and U17339 (N_17339,N_8113,N_9922);
and U17340 (N_17340,N_2945,N_4354);
nor U17341 (N_17341,N_7362,N_6173);
xnor U17342 (N_17342,N_9659,N_5123);
nand U17343 (N_17343,N_4570,N_2164);
nor U17344 (N_17344,N_143,N_18);
nand U17345 (N_17345,N_1015,N_8786);
nor U17346 (N_17346,N_7024,N_962);
nand U17347 (N_17347,N_563,N_4925);
and U17348 (N_17348,N_7038,N_458);
nor U17349 (N_17349,N_9342,N_4010);
or U17350 (N_17350,N_9904,N_6102);
nor U17351 (N_17351,N_1280,N_5289);
nor U17352 (N_17352,N_6648,N_438);
or U17353 (N_17353,N_3485,N_7454);
nor U17354 (N_17354,N_2744,N_7724);
or U17355 (N_17355,N_5530,N_7633);
xor U17356 (N_17356,N_5529,N_1625);
or U17357 (N_17357,N_4716,N_3003);
nand U17358 (N_17358,N_3586,N_451);
and U17359 (N_17359,N_4177,N_6468);
or U17360 (N_17360,N_4018,N_6211);
and U17361 (N_17361,N_8982,N_5846);
or U17362 (N_17362,N_9712,N_7381);
and U17363 (N_17363,N_5550,N_921);
xor U17364 (N_17364,N_991,N_9747);
nor U17365 (N_17365,N_5817,N_3918);
or U17366 (N_17366,N_4623,N_4243);
nand U17367 (N_17367,N_6602,N_2067);
and U17368 (N_17368,N_6155,N_5374);
xor U17369 (N_17369,N_3890,N_9206);
nand U17370 (N_17370,N_9496,N_5378);
or U17371 (N_17371,N_7377,N_9322);
or U17372 (N_17372,N_5213,N_3030);
nand U17373 (N_17373,N_7595,N_6436);
or U17374 (N_17374,N_3811,N_649);
and U17375 (N_17375,N_7292,N_9694);
xor U17376 (N_17376,N_4632,N_5945);
nor U17377 (N_17377,N_7251,N_5144);
nor U17378 (N_17378,N_1635,N_4162);
nor U17379 (N_17379,N_115,N_6609);
nor U17380 (N_17380,N_8704,N_7770);
or U17381 (N_17381,N_3329,N_8253);
and U17382 (N_17382,N_8009,N_1436);
xor U17383 (N_17383,N_6841,N_8036);
and U17384 (N_17384,N_1468,N_8107);
and U17385 (N_17385,N_7787,N_9638);
and U17386 (N_17386,N_7804,N_2752);
xor U17387 (N_17387,N_9526,N_817);
or U17388 (N_17388,N_5156,N_4306);
xnor U17389 (N_17389,N_9008,N_8862);
nand U17390 (N_17390,N_9243,N_5331);
and U17391 (N_17391,N_2552,N_4399);
and U17392 (N_17392,N_2542,N_6370);
nand U17393 (N_17393,N_5394,N_4339);
or U17394 (N_17394,N_4688,N_532);
and U17395 (N_17395,N_1930,N_8096);
or U17396 (N_17396,N_9124,N_1351);
nor U17397 (N_17397,N_4373,N_3218);
or U17398 (N_17398,N_150,N_506);
or U17399 (N_17399,N_8053,N_5296);
nor U17400 (N_17400,N_1694,N_2661);
and U17401 (N_17401,N_4121,N_8152);
nor U17402 (N_17402,N_7769,N_368);
nand U17403 (N_17403,N_5103,N_1643);
xnor U17404 (N_17404,N_9212,N_1683);
nand U17405 (N_17405,N_5835,N_3568);
nand U17406 (N_17406,N_1472,N_1240);
xnor U17407 (N_17407,N_4143,N_5910);
xnor U17408 (N_17408,N_3578,N_5603);
xor U17409 (N_17409,N_5856,N_8275);
nor U17410 (N_17410,N_4873,N_6152);
and U17411 (N_17411,N_4813,N_348);
nand U17412 (N_17412,N_2125,N_4420);
and U17413 (N_17413,N_9667,N_526);
and U17414 (N_17414,N_8554,N_6441);
and U17415 (N_17415,N_2249,N_9930);
or U17416 (N_17416,N_6926,N_4910);
nand U17417 (N_17417,N_8551,N_7257);
and U17418 (N_17418,N_617,N_4424);
or U17419 (N_17419,N_5917,N_3422);
nand U17420 (N_17420,N_3415,N_2755);
and U17421 (N_17421,N_4745,N_9476);
or U17422 (N_17422,N_1038,N_3343);
xnor U17423 (N_17423,N_6733,N_7312);
and U17424 (N_17424,N_7442,N_452);
nor U17425 (N_17425,N_1634,N_3251);
xnor U17426 (N_17426,N_3244,N_7710);
nor U17427 (N_17427,N_1123,N_2343);
nand U17428 (N_17428,N_9496,N_8228);
nand U17429 (N_17429,N_418,N_5404);
nand U17430 (N_17430,N_7295,N_7688);
and U17431 (N_17431,N_8731,N_7811);
or U17432 (N_17432,N_5582,N_5228);
or U17433 (N_17433,N_4087,N_8252);
nand U17434 (N_17434,N_4955,N_7898);
and U17435 (N_17435,N_5036,N_1717);
or U17436 (N_17436,N_2929,N_908);
or U17437 (N_17437,N_5275,N_9157);
nor U17438 (N_17438,N_8854,N_1223);
and U17439 (N_17439,N_2796,N_248);
nor U17440 (N_17440,N_5694,N_1932);
nand U17441 (N_17441,N_2519,N_4526);
nand U17442 (N_17442,N_7175,N_9409);
nand U17443 (N_17443,N_8270,N_2790);
nand U17444 (N_17444,N_2819,N_9005);
nand U17445 (N_17445,N_1168,N_548);
nand U17446 (N_17446,N_5793,N_5182);
nor U17447 (N_17447,N_9157,N_7602);
or U17448 (N_17448,N_7304,N_2600);
or U17449 (N_17449,N_3831,N_4511);
xnor U17450 (N_17450,N_6159,N_3641);
and U17451 (N_17451,N_8884,N_363);
or U17452 (N_17452,N_6413,N_3478);
and U17453 (N_17453,N_707,N_5014);
or U17454 (N_17454,N_8110,N_9258);
nand U17455 (N_17455,N_571,N_8136);
or U17456 (N_17456,N_9586,N_1503);
nor U17457 (N_17457,N_7147,N_6365);
or U17458 (N_17458,N_8341,N_2658);
nor U17459 (N_17459,N_1615,N_1781);
nand U17460 (N_17460,N_813,N_6967);
and U17461 (N_17461,N_4901,N_6791);
and U17462 (N_17462,N_259,N_8739);
and U17463 (N_17463,N_2228,N_5483);
nand U17464 (N_17464,N_5324,N_1802);
or U17465 (N_17465,N_8770,N_7759);
nand U17466 (N_17466,N_5221,N_4250);
and U17467 (N_17467,N_322,N_1020);
nand U17468 (N_17468,N_7446,N_969);
nand U17469 (N_17469,N_1457,N_6460);
or U17470 (N_17470,N_7584,N_1186);
nor U17471 (N_17471,N_7990,N_5565);
xnor U17472 (N_17472,N_9758,N_6197);
and U17473 (N_17473,N_7331,N_3526);
or U17474 (N_17474,N_1121,N_7581);
nand U17475 (N_17475,N_6504,N_4533);
and U17476 (N_17476,N_2053,N_9140);
nor U17477 (N_17477,N_8179,N_5103);
and U17478 (N_17478,N_3855,N_9761);
nand U17479 (N_17479,N_3884,N_6472);
nor U17480 (N_17480,N_5645,N_6077);
or U17481 (N_17481,N_4197,N_8715);
nand U17482 (N_17482,N_3795,N_5883);
or U17483 (N_17483,N_8301,N_8947);
nand U17484 (N_17484,N_794,N_9352);
nand U17485 (N_17485,N_5972,N_1781);
nor U17486 (N_17486,N_6966,N_7317);
xor U17487 (N_17487,N_9990,N_1983);
and U17488 (N_17488,N_7882,N_4507);
and U17489 (N_17489,N_8904,N_7811);
nand U17490 (N_17490,N_6005,N_1069);
or U17491 (N_17491,N_4012,N_6855);
nor U17492 (N_17492,N_2221,N_6161);
nand U17493 (N_17493,N_4378,N_1848);
nand U17494 (N_17494,N_1069,N_384);
or U17495 (N_17495,N_6010,N_6811);
or U17496 (N_17496,N_9534,N_7742);
nand U17497 (N_17497,N_1512,N_4213);
or U17498 (N_17498,N_6578,N_3779);
xnor U17499 (N_17499,N_7011,N_2082);
nor U17500 (N_17500,N_2470,N_2065);
nor U17501 (N_17501,N_1619,N_2991);
xor U17502 (N_17502,N_7763,N_2115);
nand U17503 (N_17503,N_5383,N_9442);
xnor U17504 (N_17504,N_8480,N_2255);
and U17505 (N_17505,N_7062,N_5322);
and U17506 (N_17506,N_4296,N_3334);
nor U17507 (N_17507,N_4852,N_4179);
xor U17508 (N_17508,N_6805,N_9934);
and U17509 (N_17509,N_2091,N_5155);
nor U17510 (N_17510,N_2807,N_632);
and U17511 (N_17511,N_751,N_4713);
and U17512 (N_17512,N_1411,N_3385);
or U17513 (N_17513,N_6315,N_3577);
nand U17514 (N_17514,N_5521,N_6220);
nand U17515 (N_17515,N_2511,N_5703);
nand U17516 (N_17516,N_7937,N_4812);
and U17517 (N_17517,N_3061,N_4869);
and U17518 (N_17518,N_9895,N_5368);
nor U17519 (N_17519,N_8743,N_9424);
nor U17520 (N_17520,N_9467,N_3960);
and U17521 (N_17521,N_9445,N_540);
nor U17522 (N_17522,N_9291,N_8907);
xor U17523 (N_17523,N_9767,N_4513);
and U17524 (N_17524,N_7525,N_2491);
nor U17525 (N_17525,N_3548,N_6629);
nor U17526 (N_17526,N_715,N_2015);
nor U17527 (N_17527,N_7320,N_1788);
nor U17528 (N_17528,N_400,N_2354);
nand U17529 (N_17529,N_4810,N_6892);
and U17530 (N_17530,N_3498,N_4887);
xnor U17531 (N_17531,N_6620,N_4205);
and U17532 (N_17532,N_3876,N_6568);
nand U17533 (N_17533,N_8879,N_9644);
or U17534 (N_17534,N_1098,N_3342);
nand U17535 (N_17535,N_980,N_1226);
or U17536 (N_17536,N_8148,N_2086);
nand U17537 (N_17537,N_2025,N_3679);
xnor U17538 (N_17538,N_4332,N_6707);
nor U17539 (N_17539,N_2857,N_8056);
or U17540 (N_17540,N_8710,N_5215);
or U17541 (N_17541,N_4256,N_171);
nor U17542 (N_17542,N_59,N_4725);
xnor U17543 (N_17543,N_3157,N_4556);
nand U17544 (N_17544,N_1614,N_103);
nor U17545 (N_17545,N_7310,N_2968);
and U17546 (N_17546,N_5405,N_6772);
and U17547 (N_17547,N_2838,N_5510);
nand U17548 (N_17548,N_9291,N_2036);
or U17549 (N_17549,N_8280,N_1142);
and U17550 (N_17550,N_9183,N_6590);
xor U17551 (N_17551,N_5773,N_5323);
nand U17552 (N_17552,N_5393,N_2784);
nand U17553 (N_17553,N_9892,N_9713);
nand U17554 (N_17554,N_6504,N_2010);
nor U17555 (N_17555,N_4304,N_4204);
and U17556 (N_17556,N_6804,N_5094);
or U17557 (N_17557,N_7714,N_5111);
and U17558 (N_17558,N_7272,N_239);
or U17559 (N_17559,N_4326,N_447);
nand U17560 (N_17560,N_5075,N_4559);
nand U17561 (N_17561,N_975,N_2080);
nor U17562 (N_17562,N_3389,N_8803);
and U17563 (N_17563,N_5411,N_9919);
nand U17564 (N_17564,N_8685,N_8716);
nor U17565 (N_17565,N_4231,N_4787);
xor U17566 (N_17566,N_2525,N_2724);
nand U17567 (N_17567,N_2711,N_637);
nor U17568 (N_17568,N_5040,N_6747);
nand U17569 (N_17569,N_7477,N_1972);
and U17570 (N_17570,N_1545,N_6523);
and U17571 (N_17571,N_9411,N_4276);
nor U17572 (N_17572,N_7721,N_5154);
or U17573 (N_17573,N_4276,N_4825);
or U17574 (N_17574,N_3513,N_3950);
or U17575 (N_17575,N_1162,N_5870);
nor U17576 (N_17576,N_995,N_4181);
and U17577 (N_17577,N_9419,N_5460);
nand U17578 (N_17578,N_1147,N_9142);
nor U17579 (N_17579,N_5674,N_1220);
and U17580 (N_17580,N_8041,N_8478);
nand U17581 (N_17581,N_3789,N_1963);
nand U17582 (N_17582,N_9588,N_8916);
nor U17583 (N_17583,N_1109,N_9632);
and U17584 (N_17584,N_140,N_5284);
or U17585 (N_17585,N_1558,N_6049);
nor U17586 (N_17586,N_6176,N_8919);
nor U17587 (N_17587,N_9152,N_3217);
xor U17588 (N_17588,N_7686,N_8662);
or U17589 (N_17589,N_5153,N_5740);
nand U17590 (N_17590,N_9440,N_8898);
nand U17591 (N_17591,N_7359,N_8232);
and U17592 (N_17592,N_7108,N_7663);
nand U17593 (N_17593,N_7018,N_3827);
nand U17594 (N_17594,N_1488,N_402);
nand U17595 (N_17595,N_3413,N_2838);
and U17596 (N_17596,N_3610,N_9037);
nor U17597 (N_17597,N_1251,N_7020);
nand U17598 (N_17598,N_4188,N_4976);
and U17599 (N_17599,N_6291,N_8797);
or U17600 (N_17600,N_4810,N_2831);
and U17601 (N_17601,N_4385,N_8941);
nand U17602 (N_17602,N_2895,N_1588);
nor U17603 (N_17603,N_8643,N_1004);
or U17604 (N_17604,N_3918,N_4934);
nor U17605 (N_17605,N_4137,N_5645);
nor U17606 (N_17606,N_7808,N_5324);
xnor U17607 (N_17607,N_3541,N_2880);
and U17608 (N_17608,N_2495,N_2218);
xor U17609 (N_17609,N_482,N_4483);
nand U17610 (N_17610,N_2465,N_6371);
nand U17611 (N_17611,N_1644,N_5012);
or U17612 (N_17612,N_7814,N_6536);
or U17613 (N_17613,N_1617,N_2784);
or U17614 (N_17614,N_5148,N_8095);
nor U17615 (N_17615,N_2393,N_8307);
or U17616 (N_17616,N_9277,N_3828);
and U17617 (N_17617,N_1222,N_3895);
nor U17618 (N_17618,N_9610,N_3386);
nor U17619 (N_17619,N_3460,N_7828);
and U17620 (N_17620,N_1788,N_9655);
xnor U17621 (N_17621,N_364,N_1554);
nor U17622 (N_17622,N_8658,N_9578);
and U17623 (N_17623,N_1448,N_4369);
nand U17624 (N_17624,N_8396,N_4691);
nor U17625 (N_17625,N_8785,N_3276);
and U17626 (N_17626,N_2514,N_9759);
or U17627 (N_17627,N_9182,N_2984);
nand U17628 (N_17628,N_7128,N_9977);
or U17629 (N_17629,N_1610,N_209);
or U17630 (N_17630,N_4341,N_1302);
xnor U17631 (N_17631,N_8393,N_1808);
or U17632 (N_17632,N_5716,N_7188);
nor U17633 (N_17633,N_9983,N_5023);
nand U17634 (N_17634,N_553,N_6038);
nand U17635 (N_17635,N_4246,N_4730);
or U17636 (N_17636,N_8321,N_5348);
nand U17637 (N_17637,N_2639,N_3446);
and U17638 (N_17638,N_4035,N_2072);
or U17639 (N_17639,N_9690,N_4786);
xor U17640 (N_17640,N_4288,N_6857);
nor U17641 (N_17641,N_1307,N_6875);
or U17642 (N_17642,N_9927,N_9011);
nand U17643 (N_17643,N_8628,N_8435);
and U17644 (N_17644,N_9347,N_9448);
nor U17645 (N_17645,N_4835,N_4315);
nor U17646 (N_17646,N_9949,N_921);
nor U17647 (N_17647,N_2256,N_7779);
nor U17648 (N_17648,N_1085,N_5766);
nand U17649 (N_17649,N_9926,N_6773);
nor U17650 (N_17650,N_3985,N_9235);
nand U17651 (N_17651,N_4680,N_445);
nor U17652 (N_17652,N_731,N_8489);
nor U17653 (N_17653,N_2364,N_813);
and U17654 (N_17654,N_9358,N_9239);
nor U17655 (N_17655,N_7887,N_8174);
nand U17656 (N_17656,N_1054,N_5804);
nor U17657 (N_17657,N_8134,N_9713);
nand U17658 (N_17658,N_9838,N_5328);
nand U17659 (N_17659,N_5302,N_5152);
nand U17660 (N_17660,N_9168,N_6460);
or U17661 (N_17661,N_4002,N_9767);
or U17662 (N_17662,N_6460,N_1334);
nor U17663 (N_17663,N_4249,N_4514);
nor U17664 (N_17664,N_551,N_9444);
nor U17665 (N_17665,N_4409,N_225);
or U17666 (N_17666,N_6264,N_5245);
or U17667 (N_17667,N_4980,N_9770);
or U17668 (N_17668,N_768,N_5730);
nand U17669 (N_17669,N_561,N_4394);
nand U17670 (N_17670,N_9866,N_8572);
nand U17671 (N_17671,N_1412,N_6023);
and U17672 (N_17672,N_722,N_2711);
xor U17673 (N_17673,N_4739,N_9760);
nand U17674 (N_17674,N_473,N_8513);
xnor U17675 (N_17675,N_6219,N_6063);
xor U17676 (N_17676,N_2998,N_5042);
and U17677 (N_17677,N_1840,N_8802);
or U17678 (N_17678,N_3135,N_9460);
nor U17679 (N_17679,N_3284,N_8572);
and U17680 (N_17680,N_1011,N_6912);
or U17681 (N_17681,N_873,N_1434);
nor U17682 (N_17682,N_625,N_5034);
and U17683 (N_17683,N_2445,N_2665);
or U17684 (N_17684,N_6561,N_1487);
and U17685 (N_17685,N_2629,N_2218);
and U17686 (N_17686,N_8908,N_7198);
or U17687 (N_17687,N_6279,N_4143);
and U17688 (N_17688,N_7473,N_4872);
nand U17689 (N_17689,N_1534,N_5470);
and U17690 (N_17690,N_3441,N_9576);
nand U17691 (N_17691,N_540,N_4175);
and U17692 (N_17692,N_3639,N_3847);
or U17693 (N_17693,N_2096,N_3627);
nand U17694 (N_17694,N_4193,N_7611);
nor U17695 (N_17695,N_1697,N_7825);
and U17696 (N_17696,N_4439,N_7363);
and U17697 (N_17697,N_9664,N_3486);
xnor U17698 (N_17698,N_1963,N_302);
or U17699 (N_17699,N_1329,N_8188);
or U17700 (N_17700,N_1939,N_2803);
nor U17701 (N_17701,N_6654,N_652);
nor U17702 (N_17702,N_4461,N_5989);
nor U17703 (N_17703,N_8184,N_8335);
nor U17704 (N_17704,N_4652,N_9539);
and U17705 (N_17705,N_6574,N_5190);
nand U17706 (N_17706,N_6488,N_233);
and U17707 (N_17707,N_8019,N_6093);
nor U17708 (N_17708,N_2473,N_101);
nor U17709 (N_17709,N_8138,N_7601);
or U17710 (N_17710,N_6279,N_8868);
and U17711 (N_17711,N_1030,N_3977);
and U17712 (N_17712,N_5184,N_4473);
xor U17713 (N_17713,N_1616,N_5730);
nor U17714 (N_17714,N_2027,N_3981);
nand U17715 (N_17715,N_838,N_6043);
nand U17716 (N_17716,N_6396,N_1399);
nor U17717 (N_17717,N_1003,N_5300);
or U17718 (N_17718,N_6888,N_6747);
nor U17719 (N_17719,N_8103,N_5088);
nand U17720 (N_17720,N_1601,N_8663);
and U17721 (N_17721,N_3958,N_1862);
or U17722 (N_17722,N_869,N_3759);
and U17723 (N_17723,N_2144,N_944);
nand U17724 (N_17724,N_482,N_4712);
and U17725 (N_17725,N_6449,N_5402);
nand U17726 (N_17726,N_4272,N_4325);
and U17727 (N_17727,N_4117,N_5799);
nand U17728 (N_17728,N_8988,N_6646);
nand U17729 (N_17729,N_8662,N_8937);
and U17730 (N_17730,N_5454,N_3855);
nor U17731 (N_17731,N_5449,N_6286);
or U17732 (N_17732,N_7645,N_7979);
nor U17733 (N_17733,N_2878,N_2897);
and U17734 (N_17734,N_9025,N_5745);
nand U17735 (N_17735,N_1027,N_5777);
and U17736 (N_17736,N_8774,N_6591);
nand U17737 (N_17737,N_2468,N_17);
or U17738 (N_17738,N_9591,N_5075);
nand U17739 (N_17739,N_3259,N_4494);
xnor U17740 (N_17740,N_3700,N_9340);
and U17741 (N_17741,N_601,N_576);
and U17742 (N_17742,N_8871,N_6057);
nor U17743 (N_17743,N_8944,N_5175);
nand U17744 (N_17744,N_8112,N_3494);
nand U17745 (N_17745,N_3591,N_8912);
nor U17746 (N_17746,N_4844,N_5075);
nor U17747 (N_17747,N_3829,N_9062);
or U17748 (N_17748,N_94,N_4621);
and U17749 (N_17749,N_3657,N_4346);
and U17750 (N_17750,N_1503,N_4616);
xor U17751 (N_17751,N_26,N_6835);
nand U17752 (N_17752,N_5784,N_2211);
xor U17753 (N_17753,N_2817,N_3700);
and U17754 (N_17754,N_8380,N_5663);
and U17755 (N_17755,N_1049,N_8158);
xnor U17756 (N_17756,N_244,N_9757);
and U17757 (N_17757,N_3378,N_7610);
and U17758 (N_17758,N_2872,N_6863);
nand U17759 (N_17759,N_954,N_5939);
nand U17760 (N_17760,N_7285,N_3760);
nand U17761 (N_17761,N_1903,N_5229);
nor U17762 (N_17762,N_2463,N_594);
or U17763 (N_17763,N_4250,N_997);
and U17764 (N_17764,N_4570,N_3846);
nand U17765 (N_17765,N_5628,N_8473);
nand U17766 (N_17766,N_9617,N_7146);
or U17767 (N_17767,N_9899,N_5988);
or U17768 (N_17768,N_4498,N_975);
nor U17769 (N_17769,N_7379,N_4020);
nor U17770 (N_17770,N_5102,N_1940);
and U17771 (N_17771,N_1590,N_1383);
and U17772 (N_17772,N_1403,N_7061);
and U17773 (N_17773,N_5972,N_4946);
nand U17774 (N_17774,N_1,N_3976);
and U17775 (N_17775,N_1182,N_4773);
or U17776 (N_17776,N_4022,N_5452);
nand U17777 (N_17777,N_1071,N_9730);
nand U17778 (N_17778,N_7399,N_2061);
nand U17779 (N_17779,N_5747,N_4170);
and U17780 (N_17780,N_8975,N_8300);
and U17781 (N_17781,N_1123,N_4150);
nor U17782 (N_17782,N_6772,N_4170);
and U17783 (N_17783,N_6020,N_8545);
nor U17784 (N_17784,N_4794,N_9923);
nor U17785 (N_17785,N_9852,N_5365);
and U17786 (N_17786,N_6474,N_678);
nor U17787 (N_17787,N_844,N_2177);
nor U17788 (N_17788,N_5673,N_6190);
and U17789 (N_17789,N_8874,N_9149);
nor U17790 (N_17790,N_9250,N_3855);
or U17791 (N_17791,N_8819,N_7929);
and U17792 (N_17792,N_711,N_5639);
or U17793 (N_17793,N_4464,N_7632);
nand U17794 (N_17794,N_1893,N_2985);
or U17795 (N_17795,N_4213,N_2500);
nor U17796 (N_17796,N_1001,N_114);
nor U17797 (N_17797,N_2687,N_5758);
and U17798 (N_17798,N_206,N_1125);
nand U17799 (N_17799,N_7721,N_6046);
or U17800 (N_17800,N_5403,N_3225);
nor U17801 (N_17801,N_9869,N_2666);
or U17802 (N_17802,N_147,N_2995);
nand U17803 (N_17803,N_4507,N_2532);
and U17804 (N_17804,N_3893,N_6439);
or U17805 (N_17805,N_8597,N_7457);
and U17806 (N_17806,N_3130,N_1828);
or U17807 (N_17807,N_4322,N_7916);
nand U17808 (N_17808,N_5751,N_7895);
nor U17809 (N_17809,N_9937,N_6902);
nand U17810 (N_17810,N_575,N_5616);
xor U17811 (N_17811,N_9028,N_1050);
and U17812 (N_17812,N_4965,N_7795);
nor U17813 (N_17813,N_109,N_2051);
nor U17814 (N_17814,N_8138,N_6894);
and U17815 (N_17815,N_2196,N_1152);
or U17816 (N_17816,N_6211,N_2659);
or U17817 (N_17817,N_289,N_7201);
or U17818 (N_17818,N_8152,N_2460);
and U17819 (N_17819,N_8342,N_6219);
xor U17820 (N_17820,N_3650,N_1092);
or U17821 (N_17821,N_5016,N_1960);
and U17822 (N_17822,N_4781,N_1044);
or U17823 (N_17823,N_5322,N_7836);
and U17824 (N_17824,N_2685,N_5674);
nand U17825 (N_17825,N_4402,N_238);
or U17826 (N_17826,N_8190,N_2365);
nand U17827 (N_17827,N_2917,N_5225);
nand U17828 (N_17828,N_7358,N_366);
nor U17829 (N_17829,N_7170,N_9323);
nand U17830 (N_17830,N_1946,N_3743);
and U17831 (N_17831,N_8729,N_1364);
nor U17832 (N_17832,N_1955,N_676);
or U17833 (N_17833,N_1157,N_6834);
nor U17834 (N_17834,N_6566,N_7483);
and U17835 (N_17835,N_2053,N_4013);
nand U17836 (N_17836,N_6629,N_7018);
or U17837 (N_17837,N_8607,N_4019);
nor U17838 (N_17838,N_1819,N_2382);
xnor U17839 (N_17839,N_6613,N_9223);
nor U17840 (N_17840,N_4782,N_3601);
nand U17841 (N_17841,N_7168,N_1040);
nand U17842 (N_17842,N_8423,N_8611);
nand U17843 (N_17843,N_8836,N_7701);
or U17844 (N_17844,N_5482,N_5773);
nor U17845 (N_17845,N_5306,N_5008);
nor U17846 (N_17846,N_9516,N_3253);
nor U17847 (N_17847,N_519,N_331);
nand U17848 (N_17848,N_6790,N_3137);
nand U17849 (N_17849,N_293,N_1998);
nor U17850 (N_17850,N_9323,N_2434);
nand U17851 (N_17851,N_2568,N_2794);
nor U17852 (N_17852,N_1874,N_6677);
nand U17853 (N_17853,N_743,N_8450);
and U17854 (N_17854,N_7467,N_5376);
or U17855 (N_17855,N_8387,N_3084);
or U17856 (N_17856,N_7677,N_3562);
nor U17857 (N_17857,N_202,N_199);
and U17858 (N_17858,N_1148,N_8778);
and U17859 (N_17859,N_7731,N_8040);
or U17860 (N_17860,N_139,N_1294);
nand U17861 (N_17861,N_8410,N_8343);
and U17862 (N_17862,N_5179,N_7562);
nand U17863 (N_17863,N_7368,N_9578);
or U17864 (N_17864,N_6712,N_8807);
or U17865 (N_17865,N_1907,N_617);
and U17866 (N_17866,N_8042,N_1986);
nand U17867 (N_17867,N_3676,N_9933);
nor U17868 (N_17868,N_1282,N_851);
nand U17869 (N_17869,N_7355,N_4051);
nor U17870 (N_17870,N_5715,N_4616);
xor U17871 (N_17871,N_6827,N_2766);
nand U17872 (N_17872,N_793,N_1160);
nor U17873 (N_17873,N_354,N_6627);
and U17874 (N_17874,N_4947,N_5677);
xnor U17875 (N_17875,N_6591,N_8559);
and U17876 (N_17876,N_7485,N_2356);
and U17877 (N_17877,N_9502,N_5387);
or U17878 (N_17878,N_9848,N_2781);
and U17879 (N_17879,N_5161,N_611);
nand U17880 (N_17880,N_1379,N_124);
and U17881 (N_17881,N_8220,N_153);
nand U17882 (N_17882,N_7457,N_900);
nand U17883 (N_17883,N_3310,N_5814);
or U17884 (N_17884,N_1342,N_7486);
and U17885 (N_17885,N_7132,N_5899);
nor U17886 (N_17886,N_484,N_3468);
nor U17887 (N_17887,N_4809,N_5344);
nor U17888 (N_17888,N_5745,N_6037);
nand U17889 (N_17889,N_595,N_1561);
xor U17890 (N_17890,N_6803,N_4461);
nand U17891 (N_17891,N_7943,N_2446);
or U17892 (N_17892,N_8117,N_8242);
or U17893 (N_17893,N_846,N_8186);
and U17894 (N_17894,N_7897,N_2629);
and U17895 (N_17895,N_7280,N_1612);
or U17896 (N_17896,N_7895,N_1352);
nand U17897 (N_17897,N_731,N_7501);
nand U17898 (N_17898,N_5806,N_6435);
nand U17899 (N_17899,N_1111,N_7769);
nand U17900 (N_17900,N_8201,N_421);
and U17901 (N_17901,N_7276,N_9483);
and U17902 (N_17902,N_4253,N_3092);
nand U17903 (N_17903,N_7750,N_4393);
nor U17904 (N_17904,N_6245,N_1326);
xor U17905 (N_17905,N_7654,N_7318);
nand U17906 (N_17906,N_4365,N_861);
or U17907 (N_17907,N_8016,N_7029);
and U17908 (N_17908,N_9208,N_2548);
and U17909 (N_17909,N_7212,N_3941);
nand U17910 (N_17910,N_1743,N_5008);
nand U17911 (N_17911,N_2267,N_1035);
or U17912 (N_17912,N_772,N_6681);
nand U17913 (N_17913,N_2869,N_4034);
nand U17914 (N_17914,N_280,N_4670);
xor U17915 (N_17915,N_4669,N_3624);
or U17916 (N_17916,N_565,N_6269);
and U17917 (N_17917,N_8309,N_6117);
nor U17918 (N_17918,N_6927,N_5200);
xor U17919 (N_17919,N_1443,N_6050);
nand U17920 (N_17920,N_8013,N_4746);
nor U17921 (N_17921,N_8419,N_4380);
nor U17922 (N_17922,N_8952,N_7511);
or U17923 (N_17923,N_3048,N_7338);
xor U17924 (N_17924,N_6515,N_931);
and U17925 (N_17925,N_4550,N_7245);
xnor U17926 (N_17926,N_697,N_140);
and U17927 (N_17927,N_182,N_1925);
and U17928 (N_17928,N_4392,N_3237);
nor U17929 (N_17929,N_7958,N_1948);
nand U17930 (N_17930,N_471,N_3209);
nand U17931 (N_17931,N_2313,N_720);
and U17932 (N_17932,N_7911,N_6962);
and U17933 (N_17933,N_6870,N_8999);
and U17934 (N_17934,N_2999,N_2732);
xnor U17935 (N_17935,N_5845,N_7412);
or U17936 (N_17936,N_2691,N_356);
nand U17937 (N_17937,N_7405,N_4683);
nand U17938 (N_17938,N_2902,N_8341);
and U17939 (N_17939,N_9041,N_130);
nor U17940 (N_17940,N_5589,N_5345);
nor U17941 (N_17941,N_6899,N_9963);
or U17942 (N_17942,N_9551,N_7141);
nand U17943 (N_17943,N_288,N_891);
nand U17944 (N_17944,N_1618,N_5605);
nand U17945 (N_17945,N_1422,N_8822);
nand U17946 (N_17946,N_5785,N_907);
or U17947 (N_17947,N_2858,N_1644);
nor U17948 (N_17948,N_2946,N_6127);
nand U17949 (N_17949,N_7103,N_5882);
xnor U17950 (N_17950,N_4578,N_4288);
and U17951 (N_17951,N_425,N_5275);
nor U17952 (N_17952,N_6601,N_4111);
nand U17953 (N_17953,N_1666,N_3892);
or U17954 (N_17954,N_8939,N_8592);
xnor U17955 (N_17955,N_3250,N_2442);
or U17956 (N_17956,N_5770,N_2710);
or U17957 (N_17957,N_5653,N_1860);
or U17958 (N_17958,N_3223,N_1433);
and U17959 (N_17959,N_5553,N_6259);
nand U17960 (N_17960,N_4015,N_8878);
nand U17961 (N_17961,N_8633,N_5596);
nand U17962 (N_17962,N_7752,N_1937);
nand U17963 (N_17963,N_153,N_6679);
xor U17964 (N_17964,N_6921,N_8881);
nor U17965 (N_17965,N_1358,N_1922);
nand U17966 (N_17966,N_9676,N_842);
nor U17967 (N_17967,N_6174,N_972);
and U17968 (N_17968,N_8396,N_8057);
nor U17969 (N_17969,N_3600,N_3295);
and U17970 (N_17970,N_9560,N_6542);
nand U17971 (N_17971,N_6298,N_4954);
or U17972 (N_17972,N_9173,N_2818);
or U17973 (N_17973,N_3077,N_321);
nor U17974 (N_17974,N_4051,N_2579);
nor U17975 (N_17975,N_2492,N_8899);
nand U17976 (N_17976,N_993,N_2023);
nor U17977 (N_17977,N_3754,N_546);
nor U17978 (N_17978,N_6671,N_3451);
nand U17979 (N_17979,N_5386,N_9966);
nand U17980 (N_17980,N_51,N_1118);
nor U17981 (N_17981,N_9719,N_9285);
nor U17982 (N_17982,N_3341,N_5690);
xnor U17983 (N_17983,N_199,N_6556);
and U17984 (N_17984,N_1451,N_3470);
and U17985 (N_17985,N_6495,N_4224);
nor U17986 (N_17986,N_447,N_6752);
or U17987 (N_17987,N_3706,N_2302);
and U17988 (N_17988,N_6311,N_3982);
and U17989 (N_17989,N_7734,N_6064);
nand U17990 (N_17990,N_1827,N_6809);
and U17991 (N_17991,N_170,N_5061);
or U17992 (N_17992,N_9808,N_7806);
nand U17993 (N_17993,N_2661,N_8344);
nand U17994 (N_17994,N_7204,N_1928);
nor U17995 (N_17995,N_4199,N_5700);
nor U17996 (N_17996,N_3945,N_8697);
and U17997 (N_17997,N_6885,N_8265);
xor U17998 (N_17998,N_2580,N_1687);
xnor U17999 (N_17999,N_2680,N_4901);
nand U18000 (N_18000,N_8126,N_4938);
nor U18001 (N_18001,N_5131,N_3462);
or U18002 (N_18002,N_7208,N_7680);
nand U18003 (N_18003,N_8775,N_5668);
nand U18004 (N_18004,N_5840,N_3614);
or U18005 (N_18005,N_9289,N_4313);
nor U18006 (N_18006,N_5730,N_6960);
xnor U18007 (N_18007,N_2675,N_1323);
or U18008 (N_18008,N_6107,N_4730);
and U18009 (N_18009,N_8265,N_680);
xor U18010 (N_18010,N_9413,N_6447);
or U18011 (N_18011,N_8835,N_5377);
nor U18012 (N_18012,N_1327,N_7916);
nor U18013 (N_18013,N_8386,N_9247);
xor U18014 (N_18014,N_8225,N_9584);
nor U18015 (N_18015,N_6318,N_1165);
nand U18016 (N_18016,N_8552,N_5406);
nor U18017 (N_18017,N_8691,N_1225);
and U18018 (N_18018,N_3168,N_3187);
and U18019 (N_18019,N_4315,N_5972);
and U18020 (N_18020,N_1456,N_8765);
nor U18021 (N_18021,N_5086,N_124);
and U18022 (N_18022,N_8281,N_8520);
xor U18023 (N_18023,N_6069,N_5823);
nand U18024 (N_18024,N_7211,N_6205);
and U18025 (N_18025,N_8211,N_3349);
or U18026 (N_18026,N_559,N_7579);
or U18027 (N_18027,N_4203,N_4501);
or U18028 (N_18028,N_331,N_3234);
or U18029 (N_18029,N_8293,N_5789);
nand U18030 (N_18030,N_3200,N_4273);
and U18031 (N_18031,N_5545,N_7494);
nand U18032 (N_18032,N_3039,N_2976);
or U18033 (N_18033,N_9344,N_5165);
nor U18034 (N_18034,N_5608,N_658);
nand U18035 (N_18035,N_6174,N_4385);
nand U18036 (N_18036,N_2747,N_2808);
xnor U18037 (N_18037,N_2095,N_3551);
xor U18038 (N_18038,N_2603,N_1401);
nor U18039 (N_18039,N_3112,N_9916);
nand U18040 (N_18040,N_4965,N_2140);
or U18041 (N_18041,N_8463,N_1971);
nor U18042 (N_18042,N_5032,N_5118);
nand U18043 (N_18043,N_4480,N_33);
or U18044 (N_18044,N_5466,N_8979);
xor U18045 (N_18045,N_1205,N_7106);
xnor U18046 (N_18046,N_9747,N_824);
or U18047 (N_18047,N_8292,N_4512);
nand U18048 (N_18048,N_9871,N_8826);
and U18049 (N_18049,N_2083,N_629);
or U18050 (N_18050,N_2247,N_7216);
xnor U18051 (N_18051,N_9312,N_7577);
nor U18052 (N_18052,N_4036,N_9894);
nand U18053 (N_18053,N_5227,N_8723);
nand U18054 (N_18054,N_4591,N_7300);
nor U18055 (N_18055,N_6795,N_6776);
nand U18056 (N_18056,N_7742,N_850);
xnor U18057 (N_18057,N_2356,N_7854);
or U18058 (N_18058,N_6967,N_9981);
nand U18059 (N_18059,N_2371,N_5343);
and U18060 (N_18060,N_1184,N_2951);
nor U18061 (N_18061,N_1602,N_2944);
nand U18062 (N_18062,N_4661,N_2248);
or U18063 (N_18063,N_9533,N_1675);
and U18064 (N_18064,N_6884,N_8217);
or U18065 (N_18065,N_4077,N_8826);
or U18066 (N_18066,N_9946,N_9211);
nand U18067 (N_18067,N_6770,N_9047);
xnor U18068 (N_18068,N_838,N_9211);
nor U18069 (N_18069,N_1361,N_1493);
nand U18070 (N_18070,N_95,N_2033);
nand U18071 (N_18071,N_863,N_9302);
and U18072 (N_18072,N_736,N_9615);
or U18073 (N_18073,N_188,N_2398);
and U18074 (N_18074,N_2997,N_5487);
nor U18075 (N_18075,N_5101,N_8237);
nand U18076 (N_18076,N_1781,N_4645);
nor U18077 (N_18077,N_1685,N_3925);
nand U18078 (N_18078,N_4943,N_1438);
nor U18079 (N_18079,N_1332,N_654);
nand U18080 (N_18080,N_5564,N_3565);
nor U18081 (N_18081,N_1377,N_9077);
nor U18082 (N_18082,N_2681,N_4276);
nor U18083 (N_18083,N_6344,N_1637);
and U18084 (N_18084,N_6122,N_4235);
nor U18085 (N_18085,N_7176,N_9167);
or U18086 (N_18086,N_8756,N_3973);
or U18087 (N_18087,N_808,N_8331);
nand U18088 (N_18088,N_6304,N_4038);
and U18089 (N_18089,N_6805,N_8600);
nor U18090 (N_18090,N_4046,N_4777);
nand U18091 (N_18091,N_5959,N_8752);
nand U18092 (N_18092,N_8515,N_6918);
nor U18093 (N_18093,N_773,N_75);
nor U18094 (N_18094,N_6559,N_4974);
and U18095 (N_18095,N_3262,N_3753);
nand U18096 (N_18096,N_2369,N_4799);
or U18097 (N_18097,N_6342,N_4777);
or U18098 (N_18098,N_526,N_9943);
nand U18099 (N_18099,N_4955,N_3142);
xor U18100 (N_18100,N_5205,N_1969);
xnor U18101 (N_18101,N_2804,N_2705);
or U18102 (N_18102,N_8833,N_2075);
and U18103 (N_18103,N_4123,N_7365);
nor U18104 (N_18104,N_9256,N_7779);
nand U18105 (N_18105,N_202,N_6012);
nand U18106 (N_18106,N_6501,N_8366);
nand U18107 (N_18107,N_3499,N_8898);
nand U18108 (N_18108,N_2621,N_7029);
and U18109 (N_18109,N_3277,N_3498);
or U18110 (N_18110,N_6513,N_7962);
and U18111 (N_18111,N_7984,N_7735);
or U18112 (N_18112,N_1357,N_757);
and U18113 (N_18113,N_6977,N_9862);
nand U18114 (N_18114,N_8915,N_8692);
or U18115 (N_18115,N_9961,N_3218);
nor U18116 (N_18116,N_2344,N_191);
or U18117 (N_18117,N_316,N_6042);
nor U18118 (N_18118,N_4343,N_8986);
nor U18119 (N_18119,N_8067,N_9068);
or U18120 (N_18120,N_6321,N_8305);
nor U18121 (N_18121,N_9762,N_9837);
or U18122 (N_18122,N_4924,N_4532);
or U18123 (N_18123,N_2789,N_6242);
nand U18124 (N_18124,N_9172,N_2559);
nor U18125 (N_18125,N_6039,N_4589);
or U18126 (N_18126,N_6378,N_2053);
or U18127 (N_18127,N_8577,N_7212);
xor U18128 (N_18128,N_371,N_6795);
and U18129 (N_18129,N_760,N_3118);
xor U18130 (N_18130,N_7855,N_4450);
or U18131 (N_18131,N_7254,N_3905);
or U18132 (N_18132,N_1297,N_7619);
and U18133 (N_18133,N_8451,N_967);
xor U18134 (N_18134,N_4105,N_9682);
nor U18135 (N_18135,N_7824,N_2299);
and U18136 (N_18136,N_2198,N_1955);
and U18137 (N_18137,N_7305,N_7831);
and U18138 (N_18138,N_9165,N_3947);
nand U18139 (N_18139,N_6577,N_9322);
nand U18140 (N_18140,N_2201,N_5479);
nand U18141 (N_18141,N_9183,N_7906);
or U18142 (N_18142,N_8825,N_8634);
xnor U18143 (N_18143,N_8539,N_8730);
and U18144 (N_18144,N_4215,N_8771);
and U18145 (N_18145,N_8256,N_9461);
xnor U18146 (N_18146,N_5388,N_3315);
and U18147 (N_18147,N_8627,N_6497);
and U18148 (N_18148,N_8921,N_5803);
nand U18149 (N_18149,N_2601,N_7865);
or U18150 (N_18150,N_1626,N_6551);
and U18151 (N_18151,N_3577,N_3623);
nand U18152 (N_18152,N_7731,N_1262);
or U18153 (N_18153,N_5079,N_6929);
or U18154 (N_18154,N_4130,N_4941);
nand U18155 (N_18155,N_938,N_9826);
or U18156 (N_18156,N_5880,N_8914);
nand U18157 (N_18157,N_9476,N_2078);
nor U18158 (N_18158,N_316,N_4064);
or U18159 (N_18159,N_4184,N_40);
xor U18160 (N_18160,N_1123,N_5075);
and U18161 (N_18161,N_544,N_9370);
and U18162 (N_18162,N_1756,N_4815);
nor U18163 (N_18163,N_3929,N_6900);
and U18164 (N_18164,N_4253,N_2116);
and U18165 (N_18165,N_9976,N_2534);
or U18166 (N_18166,N_5134,N_6443);
nor U18167 (N_18167,N_5327,N_5979);
nor U18168 (N_18168,N_459,N_8180);
and U18169 (N_18169,N_2574,N_8973);
nand U18170 (N_18170,N_3435,N_850);
nor U18171 (N_18171,N_6538,N_4224);
xor U18172 (N_18172,N_564,N_5817);
and U18173 (N_18173,N_9829,N_1643);
xor U18174 (N_18174,N_3605,N_9571);
nor U18175 (N_18175,N_1058,N_9484);
nand U18176 (N_18176,N_5104,N_48);
and U18177 (N_18177,N_1262,N_5214);
and U18178 (N_18178,N_3130,N_1424);
and U18179 (N_18179,N_9474,N_6854);
and U18180 (N_18180,N_9792,N_1174);
or U18181 (N_18181,N_9420,N_8850);
nor U18182 (N_18182,N_2525,N_9350);
nor U18183 (N_18183,N_9067,N_1866);
nand U18184 (N_18184,N_8910,N_8678);
nand U18185 (N_18185,N_3680,N_1698);
or U18186 (N_18186,N_1320,N_2328);
nand U18187 (N_18187,N_9210,N_7465);
nor U18188 (N_18188,N_9403,N_2893);
nor U18189 (N_18189,N_2603,N_6090);
or U18190 (N_18190,N_7599,N_9471);
nor U18191 (N_18191,N_2823,N_8310);
or U18192 (N_18192,N_9671,N_5877);
nor U18193 (N_18193,N_2155,N_9859);
nor U18194 (N_18194,N_5041,N_928);
or U18195 (N_18195,N_1710,N_7388);
and U18196 (N_18196,N_2781,N_1379);
or U18197 (N_18197,N_5711,N_3213);
or U18198 (N_18198,N_8313,N_3533);
xor U18199 (N_18199,N_6963,N_3100);
and U18200 (N_18200,N_7456,N_4986);
or U18201 (N_18201,N_9204,N_9447);
or U18202 (N_18202,N_4365,N_5171);
and U18203 (N_18203,N_6657,N_5238);
or U18204 (N_18204,N_1933,N_772);
nor U18205 (N_18205,N_9384,N_7041);
or U18206 (N_18206,N_2384,N_7527);
or U18207 (N_18207,N_5795,N_5298);
and U18208 (N_18208,N_7442,N_6343);
nand U18209 (N_18209,N_52,N_8945);
or U18210 (N_18210,N_9753,N_8812);
nand U18211 (N_18211,N_5510,N_186);
nand U18212 (N_18212,N_1076,N_6498);
nor U18213 (N_18213,N_6551,N_4970);
nand U18214 (N_18214,N_6549,N_5554);
or U18215 (N_18215,N_3447,N_3408);
xor U18216 (N_18216,N_160,N_4385);
nor U18217 (N_18217,N_3699,N_2868);
nand U18218 (N_18218,N_3898,N_8280);
and U18219 (N_18219,N_9974,N_501);
and U18220 (N_18220,N_6278,N_4559);
or U18221 (N_18221,N_3265,N_5321);
nand U18222 (N_18222,N_9245,N_7905);
or U18223 (N_18223,N_6227,N_3202);
nand U18224 (N_18224,N_2843,N_5258);
nor U18225 (N_18225,N_6617,N_5976);
or U18226 (N_18226,N_2146,N_1399);
nand U18227 (N_18227,N_4848,N_5081);
nor U18228 (N_18228,N_3316,N_7462);
or U18229 (N_18229,N_2899,N_6839);
xor U18230 (N_18230,N_2900,N_4052);
nor U18231 (N_18231,N_7971,N_383);
nand U18232 (N_18232,N_3541,N_3605);
nor U18233 (N_18233,N_3950,N_4212);
or U18234 (N_18234,N_6170,N_1928);
nand U18235 (N_18235,N_2339,N_7532);
nand U18236 (N_18236,N_7415,N_1527);
nor U18237 (N_18237,N_1026,N_6731);
or U18238 (N_18238,N_2914,N_2740);
or U18239 (N_18239,N_6925,N_6176);
nand U18240 (N_18240,N_4757,N_990);
or U18241 (N_18241,N_1533,N_8191);
xor U18242 (N_18242,N_3680,N_9198);
and U18243 (N_18243,N_7521,N_3631);
or U18244 (N_18244,N_143,N_9491);
nand U18245 (N_18245,N_2692,N_5436);
nand U18246 (N_18246,N_1640,N_7711);
or U18247 (N_18247,N_7700,N_1396);
nor U18248 (N_18248,N_3732,N_1024);
or U18249 (N_18249,N_3158,N_7348);
nor U18250 (N_18250,N_60,N_3714);
and U18251 (N_18251,N_8210,N_4466);
nand U18252 (N_18252,N_105,N_5176);
and U18253 (N_18253,N_802,N_9422);
and U18254 (N_18254,N_308,N_7140);
xnor U18255 (N_18255,N_8508,N_5058);
or U18256 (N_18256,N_4985,N_9938);
and U18257 (N_18257,N_956,N_8550);
nand U18258 (N_18258,N_4153,N_3251);
nor U18259 (N_18259,N_1752,N_5839);
xnor U18260 (N_18260,N_4366,N_1051);
or U18261 (N_18261,N_9450,N_8546);
nor U18262 (N_18262,N_1331,N_6321);
or U18263 (N_18263,N_4277,N_9330);
xnor U18264 (N_18264,N_4285,N_2512);
xor U18265 (N_18265,N_2062,N_3033);
or U18266 (N_18266,N_7615,N_4458);
nand U18267 (N_18267,N_1982,N_1638);
nand U18268 (N_18268,N_8135,N_253);
or U18269 (N_18269,N_3375,N_4222);
and U18270 (N_18270,N_505,N_5957);
and U18271 (N_18271,N_8099,N_5037);
nor U18272 (N_18272,N_7517,N_293);
nor U18273 (N_18273,N_6824,N_6955);
or U18274 (N_18274,N_6743,N_401);
xnor U18275 (N_18275,N_245,N_1626);
and U18276 (N_18276,N_9887,N_6140);
or U18277 (N_18277,N_8496,N_4226);
nand U18278 (N_18278,N_1124,N_2931);
and U18279 (N_18279,N_7346,N_7673);
and U18280 (N_18280,N_8643,N_6312);
nand U18281 (N_18281,N_8455,N_3725);
or U18282 (N_18282,N_3615,N_6231);
or U18283 (N_18283,N_9725,N_2287);
nor U18284 (N_18284,N_728,N_5053);
nor U18285 (N_18285,N_2781,N_3454);
nor U18286 (N_18286,N_4949,N_2726);
or U18287 (N_18287,N_6010,N_5401);
or U18288 (N_18288,N_736,N_2763);
and U18289 (N_18289,N_1179,N_204);
or U18290 (N_18290,N_2247,N_4636);
and U18291 (N_18291,N_2654,N_3441);
or U18292 (N_18292,N_2807,N_9929);
nor U18293 (N_18293,N_4277,N_4865);
nand U18294 (N_18294,N_7463,N_1771);
or U18295 (N_18295,N_5979,N_9918);
xnor U18296 (N_18296,N_7968,N_6732);
nor U18297 (N_18297,N_2299,N_6488);
and U18298 (N_18298,N_2706,N_8766);
or U18299 (N_18299,N_3909,N_3722);
or U18300 (N_18300,N_9521,N_5936);
and U18301 (N_18301,N_7837,N_8117);
and U18302 (N_18302,N_4631,N_4798);
xor U18303 (N_18303,N_441,N_1168);
and U18304 (N_18304,N_6655,N_291);
and U18305 (N_18305,N_2397,N_3354);
and U18306 (N_18306,N_1244,N_600);
or U18307 (N_18307,N_4245,N_5744);
and U18308 (N_18308,N_7515,N_6770);
xnor U18309 (N_18309,N_7551,N_2093);
nand U18310 (N_18310,N_8732,N_1940);
xnor U18311 (N_18311,N_7266,N_7348);
or U18312 (N_18312,N_2614,N_1382);
or U18313 (N_18313,N_1950,N_7760);
or U18314 (N_18314,N_8879,N_9237);
nand U18315 (N_18315,N_8363,N_480);
nor U18316 (N_18316,N_6519,N_2177);
nor U18317 (N_18317,N_6234,N_6433);
nor U18318 (N_18318,N_4031,N_4880);
nor U18319 (N_18319,N_1526,N_2217);
and U18320 (N_18320,N_6242,N_8768);
or U18321 (N_18321,N_6839,N_2696);
nand U18322 (N_18322,N_7340,N_2382);
nor U18323 (N_18323,N_6540,N_7110);
and U18324 (N_18324,N_3210,N_2021);
nand U18325 (N_18325,N_2596,N_4484);
or U18326 (N_18326,N_626,N_7014);
and U18327 (N_18327,N_8134,N_2632);
or U18328 (N_18328,N_3125,N_8061);
nor U18329 (N_18329,N_2794,N_6263);
or U18330 (N_18330,N_8725,N_3488);
nand U18331 (N_18331,N_6955,N_3713);
and U18332 (N_18332,N_5778,N_1732);
nor U18333 (N_18333,N_4777,N_2378);
nor U18334 (N_18334,N_2485,N_7668);
nor U18335 (N_18335,N_9897,N_9963);
or U18336 (N_18336,N_9510,N_2252);
nor U18337 (N_18337,N_3643,N_2843);
nand U18338 (N_18338,N_2331,N_6372);
and U18339 (N_18339,N_5745,N_3988);
nand U18340 (N_18340,N_1221,N_5221);
nand U18341 (N_18341,N_1139,N_3791);
nand U18342 (N_18342,N_1319,N_6540);
nor U18343 (N_18343,N_1108,N_9779);
nand U18344 (N_18344,N_3963,N_3996);
and U18345 (N_18345,N_3460,N_1861);
nand U18346 (N_18346,N_5620,N_3607);
and U18347 (N_18347,N_1154,N_3749);
and U18348 (N_18348,N_8909,N_7130);
nand U18349 (N_18349,N_8343,N_1600);
and U18350 (N_18350,N_9906,N_7004);
xor U18351 (N_18351,N_528,N_1061);
nand U18352 (N_18352,N_3416,N_5534);
xor U18353 (N_18353,N_7499,N_8332);
nor U18354 (N_18354,N_7023,N_1099);
and U18355 (N_18355,N_7291,N_6886);
or U18356 (N_18356,N_988,N_8011);
nor U18357 (N_18357,N_9676,N_2853);
or U18358 (N_18358,N_5468,N_6811);
nor U18359 (N_18359,N_6271,N_9402);
and U18360 (N_18360,N_1888,N_6154);
or U18361 (N_18361,N_5588,N_6774);
nor U18362 (N_18362,N_9834,N_9973);
and U18363 (N_18363,N_7358,N_2315);
or U18364 (N_18364,N_1291,N_3405);
and U18365 (N_18365,N_9869,N_8214);
nor U18366 (N_18366,N_7901,N_4093);
nor U18367 (N_18367,N_515,N_4374);
nand U18368 (N_18368,N_6505,N_1387);
and U18369 (N_18369,N_7595,N_6280);
nand U18370 (N_18370,N_9497,N_3929);
and U18371 (N_18371,N_3034,N_3666);
nand U18372 (N_18372,N_3604,N_1488);
nor U18373 (N_18373,N_2107,N_4659);
or U18374 (N_18374,N_3180,N_4044);
xor U18375 (N_18375,N_317,N_3164);
nor U18376 (N_18376,N_7315,N_756);
nand U18377 (N_18377,N_8653,N_6699);
nor U18378 (N_18378,N_9363,N_4524);
nand U18379 (N_18379,N_9644,N_19);
nand U18380 (N_18380,N_3938,N_3109);
or U18381 (N_18381,N_3594,N_4497);
nor U18382 (N_18382,N_2051,N_2153);
nand U18383 (N_18383,N_8034,N_6107);
or U18384 (N_18384,N_9053,N_5285);
xor U18385 (N_18385,N_7484,N_852);
nand U18386 (N_18386,N_709,N_2956);
nor U18387 (N_18387,N_1932,N_3515);
xor U18388 (N_18388,N_2268,N_6719);
nand U18389 (N_18389,N_7937,N_4147);
xor U18390 (N_18390,N_2083,N_3189);
or U18391 (N_18391,N_8325,N_7151);
nand U18392 (N_18392,N_6999,N_9652);
nand U18393 (N_18393,N_408,N_7980);
and U18394 (N_18394,N_7179,N_1933);
nand U18395 (N_18395,N_936,N_465);
or U18396 (N_18396,N_7441,N_6225);
nor U18397 (N_18397,N_4165,N_557);
nand U18398 (N_18398,N_7108,N_6811);
and U18399 (N_18399,N_1803,N_4151);
nand U18400 (N_18400,N_7645,N_6155);
and U18401 (N_18401,N_6792,N_4280);
and U18402 (N_18402,N_2119,N_6131);
or U18403 (N_18403,N_7017,N_3359);
or U18404 (N_18404,N_2459,N_903);
nand U18405 (N_18405,N_1818,N_1514);
nor U18406 (N_18406,N_476,N_3954);
nand U18407 (N_18407,N_714,N_7439);
nor U18408 (N_18408,N_3042,N_100);
xor U18409 (N_18409,N_7861,N_6028);
and U18410 (N_18410,N_449,N_2697);
nand U18411 (N_18411,N_9397,N_3154);
or U18412 (N_18412,N_7267,N_8962);
and U18413 (N_18413,N_2615,N_5119);
and U18414 (N_18414,N_5398,N_3927);
nor U18415 (N_18415,N_368,N_5879);
nand U18416 (N_18416,N_646,N_2915);
xor U18417 (N_18417,N_2397,N_9758);
nor U18418 (N_18418,N_6374,N_9033);
nor U18419 (N_18419,N_9012,N_336);
nand U18420 (N_18420,N_903,N_1838);
nand U18421 (N_18421,N_951,N_7448);
nand U18422 (N_18422,N_8656,N_4313);
nand U18423 (N_18423,N_1516,N_6302);
and U18424 (N_18424,N_3634,N_1219);
and U18425 (N_18425,N_6082,N_8199);
nand U18426 (N_18426,N_278,N_4636);
nand U18427 (N_18427,N_7844,N_4924);
nand U18428 (N_18428,N_2769,N_4282);
nand U18429 (N_18429,N_3473,N_4240);
and U18430 (N_18430,N_7221,N_3317);
and U18431 (N_18431,N_7685,N_5598);
or U18432 (N_18432,N_7468,N_6998);
nor U18433 (N_18433,N_3208,N_5305);
xnor U18434 (N_18434,N_4478,N_7720);
nand U18435 (N_18435,N_2464,N_7933);
or U18436 (N_18436,N_7318,N_8894);
or U18437 (N_18437,N_34,N_8681);
nor U18438 (N_18438,N_9212,N_5706);
or U18439 (N_18439,N_2723,N_974);
and U18440 (N_18440,N_2552,N_5327);
nand U18441 (N_18441,N_8642,N_3704);
nand U18442 (N_18442,N_1934,N_3826);
nor U18443 (N_18443,N_5370,N_3473);
nand U18444 (N_18444,N_8058,N_2654);
xor U18445 (N_18445,N_1563,N_8663);
xnor U18446 (N_18446,N_1259,N_806);
or U18447 (N_18447,N_5855,N_1431);
or U18448 (N_18448,N_241,N_4533);
and U18449 (N_18449,N_4321,N_9119);
and U18450 (N_18450,N_9252,N_1664);
or U18451 (N_18451,N_6145,N_2568);
nor U18452 (N_18452,N_7241,N_7234);
nor U18453 (N_18453,N_3658,N_2346);
or U18454 (N_18454,N_2004,N_5529);
or U18455 (N_18455,N_4523,N_7157);
nor U18456 (N_18456,N_1196,N_1531);
nand U18457 (N_18457,N_6536,N_4205);
nor U18458 (N_18458,N_6232,N_2250);
nor U18459 (N_18459,N_1554,N_7254);
xnor U18460 (N_18460,N_9575,N_8702);
and U18461 (N_18461,N_2874,N_5841);
and U18462 (N_18462,N_9849,N_3254);
or U18463 (N_18463,N_8419,N_7541);
nand U18464 (N_18464,N_8317,N_7814);
nor U18465 (N_18465,N_5940,N_3709);
nor U18466 (N_18466,N_4073,N_7007);
nor U18467 (N_18467,N_9247,N_305);
nand U18468 (N_18468,N_559,N_2298);
or U18469 (N_18469,N_6867,N_2482);
nor U18470 (N_18470,N_4972,N_1058);
nand U18471 (N_18471,N_3159,N_6375);
xnor U18472 (N_18472,N_9203,N_2135);
xnor U18473 (N_18473,N_7169,N_8627);
or U18474 (N_18474,N_7308,N_4316);
or U18475 (N_18475,N_973,N_7287);
or U18476 (N_18476,N_6153,N_4148);
and U18477 (N_18477,N_7295,N_5076);
or U18478 (N_18478,N_5188,N_6227);
or U18479 (N_18479,N_8666,N_6420);
and U18480 (N_18480,N_8706,N_5576);
or U18481 (N_18481,N_8988,N_3572);
nand U18482 (N_18482,N_3873,N_7449);
nand U18483 (N_18483,N_5878,N_7415);
or U18484 (N_18484,N_1488,N_2661);
nor U18485 (N_18485,N_5522,N_2873);
nand U18486 (N_18486,N_7110,N_27);
nand U18487 (N_18487,N_676,N_3036);
and U18488 (N_18488,N_6125,N_4858);
nor U18489 (N_18489,N_5713,N_7329);
or U18490 (N_18490,N_8263,N_2273);
nand U18491 (N_18491,N_588,N_5702);
and U18492 (N_18492,N_6464,N_2723);
or U18493 (N_18493,N_3164,N_5410);
nor U18494 (N_18494,N_2781,N_767);
nor U18495 (N_18495,N_3319,N_2296);
and U18496 (N_18496,N_1977,N_2595);
and U18497 (N_18497,N_5750,N_4083);
nor U18498 (N_18498,N_4372,N_1894);
nor U18499 (N_18499,N_6171,N_9623);
or U18500 (N_18500,N_5070,N_1267);
and U18501 (N_18501,N_6190,N_561);
xnor U18502 (N_18502,N_8611,N_4100);
and U18503 (N_18503,N_6715,N_6575);
nor U18504 (N_18504,N_6806,N_5311);
and U18505 (N_18505,N_3026,N_4378);
and U18506 (N_18506,N_9878,N_8260);
xnor U18507 (N_18507,N_3804,N_758);
xor U18508 (N_18508,N_649,N_8885);
nand U18509 (N_18509,N_5912,N_8151);
xor U18510 (N_18510,N_3449,N_4546);
and U18511 (N_18511,N_5775,N_6628);
or U18512 (N_18512,N_2126,N_6804);
or U18513 (N_18513,N_1741,N_8094);
xor U18514 (N_18514,N_40,N_8500);
nand U18515 (N_18515,N_7473,N_8584);
or U18516 (N_18516,N_3376,N_7010);
xor U18517 (N_18517,N_8286,N_2827);
xnor U18518 (N_18518,N_3527,N_8562);
or U18519 (N_18519,N_496,N_9289);
nor U18520 (N_18520,N_5520,N_1668);
and U18521 (N_18521,N_2476,N_8986);
nand U18522 (N_18522,N_8385,N_9159);
and U18523 (N_18523,N_7565,N_9702);
nand U18524 (N_18524,N_7816,N_4187);
and U18525 (N_18525,N_1952,N_5220);
or U18526 (N_18526,N_5672,N_3217);
and U18527 (N_18527,N_2312,N_6703);
nor U18528 (N_18528,N_7093,N_6350);
or U18529 (N_18529,N_1712,N_8590);
nor U18530 (N_18530,N_1216,N_6234);
nor U18531 (N_18531,N_4424,N_4870);
and U18532 (N_18532,N_1196,N_144);
or U18533 (N_18533,N_1707,N_5597);
and U18534 (N_18534,N_2984,N_6659);
and U18535 (N_18535,N_1192,N_9581);
or U18536 (N_18536,N_9825,N_9019);
nand U18537 (N_18537,N_2675,N_893);
xnor U18538 (N_18538,N_1467,N_7733);
xnor U18539 (N_18539,N_9448,N_2594);
and U18540 (N_18540,N_763,N_5846);
or U18541 (N_18541,N_2167,N_9507);
nand U18542 (N_18542,N_2018,N_5227);
or U18543 (N_18543,N_9786,N_2628);
or U18544 (N_18544,N_2047,N_6467);
and U18545 (N_18545,N_6960,N_8316);
nor U18546 (N_18546,N_9091,N_3027);
and U18547 (N_18547,N_1454,N_8638);
and U18548 (N_18548,N_51,N_8263);
nor U18549 (N_18549,N_5755,N_325);
nor U18550 (N_18550,N_2751,N_4638);
nand U18551 (N_18551,N_1333,N_3802);
and U18552 (N_18552,N_7033,N_5670);
nor U18553 (N_18553,N_8618,N_3303);
or U18554 (N_18554,N_9794,N_8534);
nand U18555 (N_18555,N_8696,N_2690);
nand U18556 (N_18556,N_2993,N_980);
or U18557 (N_18557,N_6928,N_4094);
or U18558 (N_18558,N_2610,N_4736);
and U18559 (N_18559,N_7460,N_2626);
and U18560 (N_18560,N_1850,N_5894);
xnor U18561 (N_18561,N_8072,N_5054);
nor U18562 (N_18562,N_8210,N_6397);
nor U18563 (N_18563,N_9957,N_4419);
or U18564 (N_18564,N_6914,N_428);
nor U18565 (N_18565,N_6074,N_9299);
and U18566 (N_18566,N_7374,N_2868);
xnor U18567 (N_18567,N_605,N_4107);
or U18568 (N_18568,N_4216,N_4706);
xor U18569 (N_18569,N_2796,N_3659);
nor U18570 (N_18570,N_1928,N_8378);
xnor U18571 (N_18571,N_7286,N_9223);
nor U18572 (N_18572,N_9620,N_7727);
nor U18573 (N_18573,N_9148,N_1602);
nand U18574 (N_18574,N_5403,N_7035);
nor U18575 (N_18575,N_7777,N_2337);
and U18576 (N_18576,N_2495,N_1002);
nand U18577 (N_18577,N_2903,N_3070);
nand U18578 (N_18578,N_4314,N_5175);
or U18579 (N_18579,N_5415,N_1463);
nand U18580 (N_18580,N_8751,N_875);
nor U18581 (N_18581,N_6036,N_9425);
nor U18582 (N_18582,N_5971,N_2761);
xor U18583 (N_18583,N_2616,N_922);
or U18584 (N_18584,N_4070,N_9134);
xor U18585 (N_18585,N_7124,N_2828);
nor U18586 (N_18586,N_2460,N_6325);
and U18587 (N_18587,N_1352,N_1420);
xor U18588 (N_18588,N_7403,N_820);
or U18589 (N_18589,N_7788,N_312);
nand U18590 (N_18590,N_275,N_644);
or U18591 (N_18591,N_5794,N_2378);
nor U18592 (N_18592,N_6441,N_9610);
or U18593 (N_18593,N_2522,N_7655);
xnor U18594 (N_18594,N_6181,N_2686);
nor U18595 (N_18595,N_4366,N_7200);
and U18596 (N_18596,N_3257,N_4859);
or U18597 (N_18597,N_4501,N_3056);
nor U18598 (N_18598,N_9679,N_9631);
or U18599 (N_18599,N_8840,N_269);
nor U18600 (N_18600,N_2828,N_7877);
or U18601 (N_18601,N_3337,N_1691);
and U18602 (N_18602,N_1820,N_1364);
or U18603 (N_18603,N_6871,N_8553);
and U18604 (N_18604,N_1148,N_3914);
nand U18605 (N_18605,N_4105,N_831);
nor U18606 (N_18606,N_2164,N_2648);
xnor U18607 (N_18607,N_7278,N_8778);
nand U18608 (N_18608,N_5449,N_8494);
and U18609 (N_18609,N_9028,N_6664);
and U18610 (N_18610,N_9187,N_5162);
nand U18611 (N_18611,N_5357,N_6605);
or U18612 (N_18612,N_736,N_6683);
or U18613 (N_18613,N_4350,N_2936);
or U18614 (N_18614,N_2559,N_660);
xor U18615 (N_18615,N_5299,N_1017);
or U18616 (N_18616,N_729,N_8066);
or U18617 (N_18617,N_9507,N_666);
or U18618 (N_18618,N_3986,N_7403);
and U18619 (N_18619,N_8082,N_7906);
nor U18620 (N_18620,N_7081,N_2342);
xnor U18621 (N_18621,N_348,N_9204);
or U18622 (N_18622,N_2702,N_669);
or U18623 (N_18623,N_2108,N_5213);
nor U18624 (N_18624,N_4519,N_1023);
nand U18625 (N_18625,N_8277,N_3769);
nor U18626 (N_18626,N_6894,N_6610);
and U18627 (N_18627,N_8418,N_9333);
and U18628 (N_18628,N_5926,N_9066);
nand U18629 (N_18629,N_5094,N_6753);
nand U18630 (N_18630,N_4246,N_6657);
nor U18631 (N_18631,N_2768,N_4781);
or U18632 (N_18632,N_1124,N_6109);
or U18633 (N_18633,N_4957,N_9499);
or U18634 (N_18634,N_8825,N_5412);
or U18635 (N_18635,N_9371,N_7052);
nor U18636 (N_18636,N_4646,N_5771);
nor U18637 (N_18637,N_2773,N_7793);
nor U18638 (N_18638,N_7457,N_7941);
nand U18639 (N_18639,N_4604,N_3972);
nor U18640 (N_18640,N_2737,N_6067);
nand U18641 (N_18641,N_3457,N_9751);
nor U18642 (N_18642,N_1956,N_7751);
and U18643 (N_18643,N_4845,N_2417);
or U18644 (N_18644,N_6782,N_8458);
and U18645 (N_18645,N_8522,N_8239);
and U18646 (N_18646,N_2363,N_2329);
nand U18647 (N_18647,N_1601,N_6137);
and U18648 (N_18648,N_5217,N_6912);
nand U18649 (N_18649,N_2773,N_9528);
or U18650 (N_18650,N_2102,N_5179);
nand U18651 (N_18651,N_227,N_735);
xnor U18652 (N_18652,N_1768,N_3041);
nand U18653 (N_18653,N_6108,N_3908);
or U18654 (N_18654,N_7265,N_8314);
and U18655 (N_18655,N_7590,N_9524);
or U18656 (N_18656,N_1369,N_4394);
nor U18657 (N_18657,N_2277,N_9334);
nand U18658 (N_18658,N_1535,N_602);
nor U18659 (N_18659,N_8700,N_9029);
xnor U18660 (N_18660,N_1205,N_7607);
or U18661 (N_18661,N_6576,N_724);
and U18662 (N_18662,N_3682,N_2198);
nand U18663 (N_18663,N_8174,N_4628);
or U18664 (N_18664,N_2134,N_3958);
and U18665 (N_18665,N_57,N_8351);
nand U18666 (N_18666,N_8326,N_3934);
nor U18667 (N_18667,N_3515,N_5631);
nor U18668 (N_18668,N_9769,N_7532);
nor U18669 (N_18669,N_3947,N_8917);
or U18670 (N_18670,N_6282,N_7628);
nor U18671 (N_18671,N_4225,N_8016);
xor U18672 (N_18672,N_7165,N_1585);
xnor U18673 (N_18673,N_9053,N_2606);
nand U18674 (N_18674,N_1246,N_7150);
or U18675 (N_18675,N_3501,N_2754);
and U18676 (N_18676,N_2254,N_9832);
or U18677 (N_18677,N_1953,N_3366);
or U18678 (N_18678,N_4190,N_5112);
or U18679 (N_18679,N_4651,N_2139);
or U18680 (N_18680,N_5143,N_8386);
or U18681 (N_18681,N_9270,N_8212);
nand U18682 (N_18682,N_1952,N_2911);
or U18683 (N_18683,N_1757,N_5602);
xnor U18684 (N_18684,N_1292,N_2196);
or U18685 (N_18685,N_5937,N_2331);
nor U18686 (N_18686,N_5890,N_6867);
and U18687 (N_18687,N_7491,N_2387);
nor U18688 (N_18688,N_6443,N_2447);
nor U18689 (N_18689,N_421,N_1853);
nand U18690 (N_18690,N_3869,N_2218);
nand U18691 (N_18691,N_974,N_1856);
or U18692 (N_18692,N_5948,N_1337);
nand U18693 (N_18693,N_7415,N_1240);
and U18694 (N_18694,N_1163,N_8905);
or U18695 (N_18695,N_9654,N_7175);
or U18696 (N_18696,N_3372,N_8858);
nor U18697 (N_18697,N_1217,N_4605);
nand U18698 (N_18698,N_9649,N_7561);
nand U18699 (N_18699,N_7601,N_1395);
nor U18700 (N_18700,N_5844,N_1138);
and U18701 (N_18701,N_4711,N_3921);
or U18702 (N_18702,N_1050,N_8029);
xor U18703 (N_18703,N_9349,N_6562);
and U18704 (N_18704,N_6723,N_7532);
and U18705 (N_18705,N_3230,N_4588);
and U18706 (N_18706,N_8537,N_6137);
nand U18707 (N_18707,N_8367,N_3391);
and U18708 (N_18708,N_3055,N_8026);
nor U18709 (N_18709,N_9374,N_2807);
or U18710 (N_18710,N_5191,N_415);
or U18711 (N_18711,N_1094,N_9925);
nor U18712 (N_18712,N_9545,N_6746);
and U18713 (N_18713,N_2654,N_2608);
nor U18714 (N_18714,N_8314,N_2393);
or U18715 (N_18715,N_9131,N_1216);
nand U18716 (N_18716,N_3459,N_6005);
nor U18717 (N_18717,N_6307,N_1976);
or U18718 (N_18718,N_6886,N_6896);
and U18719 (N_18719,N_1085,N_2793);
nor U18720 (N_18720,N_9144,N_4242);
nor U18721 (N_18721,N_1013,N_7683);
nand U18722 (N_18722,N_9780,N_3613);
or U18723 (N_18723,N_9369,N_8382);
nor U18724 (N_18724,N_4088,N_7719);
and U18725 (N_18725,N_956,N_6081);
nand U18726 (N_18726,N_8129,N_6650);
nor U18727 (N_18727,N_2099,N_7908);
and U18728 (N_18728,N_3403,N_4133);
nand U18729 (N_18729,N_605,N_9738);
nor U18730 (N_18730,N_1282,N_9137);
nand U18731 (N_18731,N_9314,N_4912);
nand U18732 (N_18732,N_1743,N_4341);
and U18733 (N_18733,N_7085,N_1663);
and U18734 (N_18734,N_4770,N_9959);
or U18735 (N_18735,N_4924,N_3549);
or U18736 (N_18736,N_340,N_5271);
and U18737 (N_18737,N_5745,N_2348);
nor U18738 (N_18738,N_4496,N_5796);
nor U18739 (N_18739,N_6648,N_5204);
xor U18740 (N_18740,N_4166,N_3069);
xor U18741 (N_18741,N_7173,N_4570);
nor U18742 (N_18742,N_5908,N_9320);
and U18743 (N_18743,N_464,N_2636);
or U18744 (N_18744,N_816,N_1032);
and U18745 (N_18745,N_6415,N_2375);
and U18746 (N_18746,N_1065,N_5961);
nand U18747 (N_18747,N_9962,N_2769);
nand U18748 (N_18748,N_8452,N_6468);
and U18749 (N_18749,N_3784,N_7465);
or U18750 (N_18750,N_448,N_6810);
xnor U18751 (N_18751,N_6352,N_3227);
nor U18752 (N_18752,N_1583,N_3984);
or U18753 (N_18753,N_4883,N_2057);
or U18754 (N_18754,N_2030,N_9732);
and U18755 (N_18755,N_3477,N_7504);
nand U18756 (N_18756,N_2961,N_9783);
xnor U18757 (N_18757,N_100,N_8725);
and U18758 (N_18758,N_958,N_5301);
nor U18759 (N_18759,N_1040,N_1120);
or U18760 (N_18760,N_5330,N_4387);
and U18761 (N_18761,N_634,N_3208);
and U18762 (N_18762,N_5699,N_8079);
or U18763 (N_18763,N_3504,N_3475);
and U18764 (N_18764,N_3961,N_2660);
nand U18765 (N_18765,N_1820,N_2195);
and U18766 (N_18766,N_2033,N_8887);
xor U18767 (N_18767,N_2745,N_2123);
nor U18768 (N_18768,N_35,N_1644);
and U18769 (N_18769,N_2529,N_4572);
and U18770 (N_18770,N_6664,N_1998);
nand U18771 (N_18771,N_9027,N_5836);
xor U18772 (N_18772,N_7630,N_743);
xnor U18773 (N_18773,N_3174,N_2128);
xnor U18774 (N_18774,N_8649,N_8479);
or U18775 (N_18775,N_650,N_2631);
xor U18776 (N_18776,N_3968,N_5603);
or U18777 (N_18777,N_1168,N_431);
xor U18778 (N_18778,N_7913,N_9492);
or U18779 (N_18779,N_5231,N_1131);
and U18780 (N_18780,N_1658,N_3197);
xor U18781 (N_18781,N_8353,N_7786);
xnor U18782 (N_18782,N_5479,N_2165);
nand U18783 (N_18783,N_8991,N_5019);
and U18784 (N_18784,N_249,N_5674);
nand U18785 (N_18785,N_9572,N_4990);
and U18786 (N_18786,N_5881,N_9636);
and U18787 (N_18787,N_8164,N_9995);
nand U18788 (N_18788,N_8492,N_4029);
nand U18789 (N_18789,N_6929,N_254);
or U18790 (N_18790,N_4449,N_1514);
nor U18791 (N_18791,N_9682,N_5037);
or U18792 (N_18792,N_7403,N_477);
and U18793 (N_18793,N_6160,N_2719);
nand U18794 (N_18794,N_4816,N_249);
and U18795 (N_18795,N_7405,N_239);
xor U18796 (N_18796,N_5508,N_8660);
xnor U18797 (N_18797,N_9666,N_6441);
nor U18798 (N_18798,N_1,N_5237);
nand U18799 (N_18799,N_7376,N_2464);
nor U18800 (N_18800,N_7364,N_621);
nor U18801 (N_18801,N_1427,N_4171);
or U18802 (N_18802,N_4029,N_8511);
and U18803 (N_18803,N_9217,N_6109);
and U18804 (N_18804,N_3000,N_4085);
and U18805 (N_18805,N_621,N_1607);
or U18806 (N_18806,N_4966,N_7731);
nand U18807 (N_18807,N_7273,N_1320);
nor U18808 (N_18808,N_5047,N_7470);
xnor U18809 (N_18809,N_8364,N_5640);
and U18810 (N_18810,N_8787,N_3521);
or U18811 (N_18811,N_4161,N_6244);
or U18812 (N_18812,N_4478,N_1942);
nor U18813 (N_18813,N_9303,N_834);
nor U18814 (N_18814,N_698,N_809);
or U18815 (N_18815,N_6237,N_109);
or U18816 (N_18816,N_1956,N_7972);
or U18817 (N_18817,N_4832,N_5821);
and U18818 (N_18818,N_8482,N_4133);
and U18819 (N_18819,N_5982,N_7606);
or U18820 (N_18820,N_3257,N_8792);
or U18821 (N_18821,N_8687,N_7283);
or U18822 (N_18822,N_115,N_8154);
or U18823 (N_18823,N_2158,N_1347);
nand U18824 (N_18824,N_8480,N_9159);
or U18825 (N_18825,N_5981,N_3793);
or U18826 (N_18826,N_8098,N_5236);
nor U18827 (N_18827,N_4629,N_5766);
and U18828 (N_18828,N_6363,N_862);
nor U18829 (N_18829,N_9,N_6185);
and U18830 (N_18830,N_7154,N_6288);
or U18831 (N_18831,N_6689,N_5690);
or U18832 (N_18832,N_707,N_8154);
xnor U18833 (N_18833,N_8406,N_1721);
nor U18834 (N_18834,N_8024,N_6769);
xor U18835 (N_18835,N_7086,N_2240);
xor U18836 (N_18836,N_579,N_3402);
xor U18837 (N_18837,N_1236,N_8438);
and U18838 (N_18838,N_5362,N_8623);
nand U18839 (N_18839,N_5030,N_3258);
nand U18840 (N_18840,N_7313,N_3818);
nor U18841 (N_18841,N_7716,N_3243);
and U18842 (N_18842,N_436,N_7620);
and U18843 (N_18843,N_7751,N_8462);
nand U18844 (N_18844,N_8264,N_5466);
or U18845 (N_18845,N_2360,N_8897);
or U18846 (N_18846,N_6949,N_6116);
nand U18847 (N_18847,N_503,N_3883);
xor U18848 (N_18848,N_6125,N_8983);
nor U18849 (N_18849,N_5443,N_7762);
nand U18850 (N_18850,N_2811,N_7958);
or U18851 (N_18851,N_9991,N_2368);
nand U18852 (N_18852,N_8893,N_1497);
and U18853 (N_18853,N_1436,N_821);
nor U18854 (N_18854,N_4660,N_2424);
nor U18855 (N_18855,N_5900,N_3120);
nor U18856 (N_18856,N_6522,N_3423);
xor U18857 (N_18857,N_3928,N_1493);
and U18858 (N_18858,N_7031,N_3913);
nor U18859 (N_18859,N_1353,N_7452);
nand U18860 (N_18860,N_1038,N_2472);
nand U18861 (N_18861,N_6318,N_4748);
nor U18862 (N_18862,N_9054,N_2572);
nor U18863 (N_18863,N_4072,N_5902);
nor U18864 (N_18864,N_8199,N_3034);
xnor U18865 (N_18865,N_3977,N_5413);
xnor U18866 (N_18866,N_6170,N_5745);
or U18867 (N_18867,N_3450,N_2403);
xnor U18868 (N_18868,N_5644,N_4814);
or U18869 (N_18869,N_4920,N_6980);
nor U18870 (N_18870,N_3964,N_7793);
nor U18871 (N_18871,N_4518,N_856);
nor U18872 (N_18872,N_1478,N_111);
nor U18873 (N_18873,N_906,N_4213);
or U18874 (N_18874,N_7608,N_9513);
xnor U18875 (N_18875,N_6124,N_66);
nand U18876 (N_18876,N_2573,N_5516);
or U18877 (N_18877,N_4211,N_1080);
and U18878 (N_18878,N_3605,N_400);
or U18879 (N_18879,N_4,N_3402);
nor U18880 (N_18880,N_6469,N_9614);
nor U18881 (N_18881,N_9190,N_7827);
nand U18882 (N_18882,N_190,N_1405);
and U18883 (N_18883,N_1327,N_3615);
and U18884 (N_18884,N_6220,N_4187);
or U18885 (N_18885,N_8471,N_4786);
nor U18886 (N_18886,N_3967,N_8227);
or U18887 (N_18887,N_3554,N_6829);
nor U18888 (N_18888,N_88,N_3169);
nor U18889 (N_18889,N_4540,N_259);
or U18890 (N_18890,N_5831,N_8191);
and U18891 (N_18891,N_6019,N_3997);
and U18892 (N_18892,N_4241,N_6572);
nand U18893 (N_18893,N_6396,N_9034);
nor U18894 (N_18894,N_9484,N_6856);
xnor U18895 (N_18895,N_4312,N_7829);
and U18896 (N_18896,N_5285,N_8408);
nor U18897 (N_18897,N_6649,N_1880);
or U18898 (N_18898,N_57,N_7036);
xor U18899 (N_18899,N_3168,N_9392);
and U18900 (N_18900,N_1225,N_4798);
xor U18901 (N_18901,N_4322,N_3596);
or U18902 (N_18902,N_6673,N_6777);
nor U18903 (N_18903,N_2722,N_9893);
and U18904 (N_18904,N_7132,N_465);
xor U18905 (N_18905,N_7166,N_3885);
or U18906 (N_18906,N_1884,N_8540);
nor U18907 (N_18907,N_2056,N_838);
and U18908 (N_18908,N_8782,N_381);
nand U18909 (N_18909,N_7139,N_5624);
and U18910 (N_18910,N_4519,N_8852);
xnor U18911 (N_18911,N_5570,N_1103);
nand U18912 (N_18912,N_7970,N_69);
and U18913 (N_18913,N_9908,N_5354);
nor U18914 (N_18914,N_9218,N_9046);
and U18915 (N_18915,N_5306,N_9734);
xnor U18916 (N_18916,N_6867,N_1749);
nand U18917 (N_18917,N_3202,N_2593);
nor U18918 (N_18918,N_4227,N_6214);
and U18919 (N_18919,N_1039,N_9898);
nand U18920 (N_18920,N_7535,N_8752);
and U18921 (N_18921,N_5720,N_9604);
nor U18922 (N_18922,N_2488,N_3519);
and U18923 (N_18923,N_9633,N_9308);
or U18924 (N_18924,N_7995,N_1848);
nand U18925 (N_18925,N_998,N_8847);
and U18926 (N_18926,N_8525,N_4589);
xnor U18927 (N_18927,N_9378,N_6067);
nor U18928 (N_18928,N_9667,N_8228);
or U18929 (N_18929,N_5797,N_5264);
nor U18930 (N_18930,N_6709,N_1184);
nor U18931 (N_18931,N_5983,N_4705);
or U18932 (N_18932,N_4092,N_1130);
and U18933 (N_18933,N_7835,N_5821);
nor U18934 (N_18934,N_3764,N_2539);
or U18935 (N_18935,N_7760,N_9344);
nor U18936 (N_18936,N_6728,N_6426);
xor U18937 (N_18937,N_7707,N_5726);
nor U18938 (N_18938,N_3486,N_6078);
nor U18939 (N_18939,N_6004,N_2909);
nand U18940 (N_18940,N_3464,N_5133);
nor U18941 (N_18941,N_9071,N_789);
and U18942 (N_18942,N_5345,N_1459);
xor U18943 (N_18943,N_4636,N_9242);
nand U18944 (N_18944,N_2827,N_5445);
nor U18945 (N_18945,N_6842,N_7091);
nor U18946 (N_18946,N_8867,N_5182);
xnor U18947 (N_18947,N_9475,N_4380);
nand U18948 (N_18948,N_6350,N_598);
nor U18949 (N_18949,N_9252,N_6492);
nand U18950 (N_18950,N_5872,N_8237);
xnor U18951 (N_18951,N_5757,N_1952);
and U18952 (N_18952,N_2010,N_6873);
nor U18953 (N_18953,N_878,N_7704);
and U18954 (N_18954,N_6867,N_1671);
or U18955 (N_18955,N_4283,N_8806);
or U18956 (N_18956,N_9811,N_2574);
or U18957 (N_18957,N_9713,N_1170);
and U18958 (N_18958,N_5656,N_5723);
nor U18959 (N_18959,N_5861,N_6447);
nand U18960 (N_18960,N_5203,N_1113);
nand U18961 (N_18961,N_4742,N_2317);
nand U18962 (N_18962,N_8017,N_9372);
nor U18963 (N_18963,N_3062,N_753);
and U18964 (N_18964,N_6708,N_4707);
nand U18965 (N_18965,N_1988,N_3255);
and U18966 (N_18966,N_37,N_2778);
or U18967 (N_18967,N_6089,N_3284);
and U18968 (N_18968,N_2138,N_9288);
nand U18969 (N_18969,N_8150,N_6509);
and U18970 (N_18970,N_1408,N_2262);
nand U18971 (N_18971,N_5994,N_6135);
and U18972 (N_18972,N_5762,N_7644);
nor U18973 (N_18973,N_1710,N_3755);
and U18974 (N_18974,N_8649,N_4376);
nand U18975 (N_18975,N_6481,N_28);
nor U18976 (N_18976,N_4606,N_9289);
or U18977 (N_18977,N_1661,N_8456);
nand U18978 (N_18978,N_948,N_8217);
nand U18979 (N_18979,N_8006,N_7166);
and U18980 (N_18980,N_5436,N_257);
and U18981 (N_18981,N_645,N_9814);
nor U18982 (N_18982,N_9090,N_3521);
nand U18983 (N_18983,N_761,N_2937);
nand U18984 (N_18984,N_9220,N_8162);
or U18985 (N_18985,N_5885,N_5169);
or U18986 (N_18986,N_6604,N_4977);
and U18987 (N_18987,N_7769,N_4681);
nand U18988 (N_18988,N_475,N_495);
nor U18989 (N_18989,N_168,N_1420);
nor U18990 (N_18990,N_354,N_4015);
xor U18991 (N_18991,N_3040,N_2253);
or U18992 (N_18992,N_2017,N_354);
nand U18993 (N_18993,N_7805,N_6116);
nor U18994 (N_18994,N_6682,N_6151);
xnor U18995 (N_18995,N_6015,N_9593);
nand U18996 (N_18996,N_6010,N_9583);
or U18997 (N_18997,N_3500,N_3699);
and U18998 (N_18998,N_6981,N_6195);
nor U18999 (N_18999,N_3141,N_2745);
nand U19000 (N_19000,N_8552,N_9729);
and U19001 (N_19001,N_8835,N_6074);
and U19002 (N_19002,N_4972,N_7945);
or U19003 (N_19003,N_8924,N_655);
or U19004 (N_19004,N_8428,N_5601);
and U19005 (N_19005,N_6298,N_2780);
and U19006 (N_19006,N_6041,N_7240);
or U19007 (N_19007,N_8811,N_9897);
nor U19008 (N_19008,N_8877,N_1613);
and U19009 (N_19009,N_2776,N_723);
nand U19010 (N_19010,N_2140,N_210);
nand U19011 (N_19011,N_7040,N_1040);
nor U19012 (N_19012,N_8620,N_7773);
nor U19013 (N_19013,N_3962,N_3596);
or U19014 (N_19014,N_8675,N_3361);
and U19015 (N_19015,N_2966,N_9588);
and U19016 (N_19016,N_8385,N_4762);
nand U19017 (N_19017,N_492,N_8177);
and U19018 (N_19018,N_6667,N_5662);
nor U19019 (N_19019,N_8168,N_9354);
nor U19020 (N_19020,N_4480,N_5628);
or U19021 (N_19021,N_8492,N_7374);
and U19022 (N_19022,N_3012,N_7429);
and U19023 (N_19023,N_3549,N_2061);
nand U19024 (N_19024,N_4692,N_8293);
or U19025 (N_19025,N_94,N_6641);
nand U19026 (N_19026,N_6696,N_9690);
or U19027 (N_19027,N_7839,N_6668);
nand U19028 (N_19028,N_5229,N_1738);
nand U19029 (N_19029,N_2490,N_6129);
nand U19030 (N_19030,N_1313,N_3342);
xor U19031 (N_19031,N_7328,N_2615);
or U19032 (N_19032,N_378,N_5201);
and U19033 (N_19033,N_4347,N_7936);
and U19034 (N_19034,N_9050,N_8268);
xnor U19035 (N_19035,N_5727,N_6103);
nor U19036 (N_19036,N_8946,N_170);
and U19037 (N_19037,N_1852,N_9390);
nor U19038 (N_19038,N_2079,N_1469);
nor U19039 (N_19039,N_8951,N_3443);
nand U19040 (N_19040,N_1775,N_8909);
and U19041 (N_19041,N_1908,N_8567);
and U19042 (N_19042,N_7689,N_4509);
or U19043 (N_19043,N_770,N_7076);
nor U19044 (N_19044,N_2079,N_6316);
nand U19045 (N_19045,N_1533,N_1262);
xor U19046 (N_19046,N_9551,N_2727);
or U19047 (N_19047,N_133,N_9623);
or U19048 (N_19048,N_6805,N_3766);
nand U19049 (N_19049,N_6999,N_8525);
nor U19050 (N_19050,N_8911,N_344);
or U19051 (N_19051,N_7785,N_1848);
xnor U19052 (N_19052,N_6760,N_28);
nand U19053 (N_19053,N_67,N_3556);
or U19054 (N_19054,N_2260,N_9808);
and U19055 (N_19055,N_5052,N_1247);
nor U19056 (N_19056,N_6381,N_9390);
nor U19057 (N_19057,N_911,N_3029);
or U19058 (N_19058,N_4140,N_3713);
or U19059 (N_19059,N_7341,N_4134);
nor U19060 (N_19060,N_4342,N_2603);
and U19061 (N_19061,N_3138,N_2203);
or U19062 (N_19062,N_2517,N_5789);
nor U19063 (N_19063,N_6811,N_9118);
nand U19064 (N_19064,N_5830,N_9631);
nor U19065 (N_19065,N_6023,N_748);
or U19066 (N_19066,N_7615,N_2373);
or U19067 (N_19067,N_2132,N_9925);
or U19068 (N_19068,N_6570,N_8752);
nand U19069 (N_19069,N_3266,N_3066);
nand U19070 (N_19070,N_6843,N_4500);
nand U19071 (N_19071,N_2391,N_9272);
or U19072 (N_19072,N_4352,N_1635);
nor U19073 (N_19073,N_3307,N_6187);
xnor U19074 (N_19074,N_9031,N_5052);
or U19075 (N_19075,N_3897,N_2725);
nor U19076 (N_19076,N_7431,N_49);
nand U19077 (N_19077,N_1996,N_5942);
or U19078 (N_19078,N_9218,N_2338);
and U19079 (N_19079,N_4916,N_9804);
nor U19080 (N_19080,N_1277,N_4708);
and U19081 (N_19081,N_39,N_7748);
and U19082 (N_19082,N_7023,N_1017);
and U19083 (N_19083,N_3651,N_2764);
nor U19084 (N_19084,N_1545,N_9965);
nor U19085 (N_19085,N_9026,N_1280);
and U19086 (N_19086,N_8953,N_1137);
nand U19087 (N_19087,N_2356,N_412);
and U19088 (N_19088,N_7883,N_4280);
nand U19089 (N_19089,N_5386,N_1881);
nand U19090 (N_19090,N_3287,N_4323);
xor U19091 (N_19091,N_6108,N_6566);
and U19092 (N_19092,N_7414,N_5812);
nand U19093 (N_19093,N_7148,N_3054);
nor U19094 (N_19094,N_2120,N_3860);
and U19095 (N_19095,N_349,N_9531);
xnor U19096 (N_19096,N_4337,N_7836);
and U19097 (N_19097,N_9327,N_262);
or U19098 (N_19098,N_7179,N_3838);
nand U19099 (N_19099,N_5713,N_477);
nor U19100 (N_19100,N_8334,N_5891);
and U19101 (N_19101,N_3270,N_1475);
nor U19102 (N_19102,N_3401,N_7536);
xnor U19103 (N_19103,N_8977,N_1681);
nor U19104 (N_19104,N_7613,N_4911);
or U19105 (N_19105,N_2252,N_7829);
nor U19106 (N_19106,N_1843,N_3247);
nand U19107 (N_19107,N_6574,N_2487);
or U19108 (N_19108,N_4508,N_9111);
xor U19109 (N_19109,N_1914,N_1891);
and U19110 (N_19110,N_5406,N_3711);
and U19111 (N_19111,N_7882,N_9538);
and U19112 (N_19112,N_7361,N_2123);
nor U19113 (N_19113,N_4511,N_2929);
and U19114 (N_19114,N_2850,N_2163);
xor U19115 (N_19115,N_1468,N_8832);
nand U19116 (N_19116,N_8896,N_7153);
and U19117 (N_19117,N_5678,N_8526);
nor U19118 (N_19118,N_5500,N_8534);
xor U19119 (N_19119,N_4535,N_8343);
nand U19120 (N_19120,N_1257,N_9316);
and U19121 (N_19121,N_2892,N_9150);
nand U19122 (N_19122,N_8143,N_708);
nand U19123 (N_19123,N_9035,N_19);
xor U19124 (N_19124,N_6953,N_8164);
xor U19125 (N_19125,N_5150,N_7776);
nor U19126 (N_19126,N_5070,N_6312);
nor U19127 (N_19127,N_4128,N_8954);
or U19128 (N_19128,N_7017,N_5687);
nor U19129 (N_19129,N_3545,N_9503);
and U19130 (N_19130,N_1825,N_7696);
and U19131 (N_19131,N_7389,N_9042);
nor U19132 (N_19132,N_9431,N_3778);
nand U19133 (N_19133,N_6091,N_561);
or U19134 (N_19134,N_8595,N_3160);
and U19135 (N_19135,N_5409,N_8826);
and U19136 (N_19136,N_4631,N_4582);
and U19137 (N_19137,N_2674,N_6777);
and U19138 (N_19138,N_8646,N_3396);
nor U19139 (N_19139,N_2742,N_9881);
nand U19140 (N_19140,N_8061,N_5162);
nand U19141 (N_19141,N_5996,N_5011);
or U19142 (N_19142,N_8343,N_6437);
or U19143 (N_19143,N_508,N_7091);
nor U19144 (N_19144,N_8545,N_9916);
nor U19145 (N_19145,N_2474,N_243);
or U19146 (N_19146,N_5558,N_5811);
and U19147 (N_19147,N_2666,N_1985);
nor U19148 (N_19148,N_5183,N_7363);
or U19149 (N_19149,N_436,N_9178);
or U19150 (N_19150,N_1482,N_2384);
or U19151 (N_19151,N_7968,N_3689);
nor U19152 (N_19152,N_5598,N_8872);
nor U19153 (N_19153,N_6647,N_8135);
nor U19154 (N_19154,N_8643,N_6808);
and U19155 (N_19155,N_2391,N_3191);
nand U19156 (N_19156,N_954,N_2912);
and U19157 (N_19157,N_8768,N_4710);
or U19158 (N_19158,N_6109,N_8086);
nand U19159 (N_19159,N_3405,N_8132);
xnor U19160 (N_19160,N_6344,N_8686);
xnor U19161 (N_19161,N_868,N_6004);
nor U19162 (N_19162,N_3567,N_9502);
and U19163 (N_19163,N_7638,N_5151);
xnor U19164 (N_19164,N_8021,N_8729);
or U19165 (N_19165,N_7080,N_6611);
xnor U19166 (N_19166,N_4300,N_7852);
nand U19167 (N_19167,N_7872,N_4502);
nand U19168 (N_19168,N_4240,N_9721);
or U19169 (N_19169,N_5581,N_3794);
xnor U19170 (N_19170,N_7266,N_9261);
nor U19171 (N_19171,N_7850,N_1743);
and U19172 (N_19172,N_397,N_7951);
xor U19173 (N_19173,N_6957,N_3481);
and U19174 (N_19174,N_4005,N_1997);
nor U19175 (N_19175,N_6597,N_2272);
xnor U19176 (N_19176,N_1606,N_9428);
nor U19177 (N_19177,N_5797,N_8327);
xnor U19178 (N_19178,N_5332,N_1074);
xnor U19179 (N_19179,N_8324,N_4175);
or U19180 (N_19180,N_4488,N_1038);
nand U19181 (N_19181,N_6831,N_3353);
nand U19182 (N_19182,N_4180,N_4824);
nor U19183 (N_19183,N_1065,N_3731);
or U19184 (N_19184,N_5878,N_999);
nor U19185 (N_19185,N_436,N_6201);
or U19186 (N_19186,N_4357,N_3761);
xor U19187 (N_19187,N_7806,N_4451);
nor U19188 (N_19188,N_1681,N_1926);
xnor U19189 (N_19189,N_4531,N_9300);
nand U19190 (N_19190,N_1741,N_736);
or U19191 (N_19191,N_7462,N_7833);
and U19192 (N_19192,N_592,N_8630);
nand U19193 (N_19193,N_5282,N_7670);
and U19194 (N_19194,N_6901,N_4703);
and U19195 (N_19195,N_3664,N_5410);
or U19196 (N_19196,N_1195,N_2391);
nor U19197 (N_19197,N_3691,N_4348);
nor U19198 (N_19198,N_8184,N_6821);
and U19199 (N_19199,N_1227,N_7969);
or U19200 (N_19200,N_7004,N_6792);
and U19201 (N_19201,N_1203,N_5433);
xnor U19202 (N_19202,N_5545,N_557);
xnor U19203 (N_19203,N_164,N_6081);
nor U19204 (N_19204,N_3884,N_3144);
nor U19205 (N_19205,N_67,N_1895);
nor U19206 (N_19206,N_7025,N_753);
and U19207 (N_19207,N_5101,N_2444);
nor U19208 (N_19208,N_5698,N_4961);
nor U19209 (N_19209,N_5859,N_7788);
and U19210 (N_19210,N_23,N_4884);
and U19211 (N_19211,N_9159,N_9483);
and U19212 (N_19212,N_3462,N_615);
and U19213 (N_19213,N_6620,N_2839);
and U19214 (N_19214,N_8630,N_9003);
nor U19215 (N_19215,N_7502,N_1323);
or U19216 (N_19216,N_2663,N_6723);
nand U19217 (N_19217,N_1644,N_3613);
nor U19218 (N_19218,N_5737,N_4585);
nor U19219 (N_19219,N_8707,N_1118);
xnor U19220 (N_19220,N_8932,N_1903);
and U19221 (N_19221,N_918,N_9864);
xnor U19222 (N_19222,N_5295,N_4355);
nand U19223 (N_19223,N_8957,N_2634);
xnor U19224 (N_19224,N_3983,N_840);
and U19225 (N_19225,N_670,N_6350);
nor U19226 (N_19226,N_1260,N_7509);
and U19227 (N_19227,N_1385,N_8435);
xnor U19228 (N_19228,N_8087,N_8624);
or U19229 (N_19229,N_843,N_9536);
or U19230 (N_19230,N_8232,N_5505);
nand U19231 (N_19231,N_7995,N_8368);
nand U19232 (N_19232,N_867,N_2660);
and U19233 (N_19233,N_1042,N_6949);
and U19234 (N_19234,N_6379,N_9720);
or U19235 (N_19235,N_4339,N_4041);
nand U19236 (N_19236,N_436,N_9285);
nor U19237 (N_19237,N_3055,N_9181);
nor U19238 (N_19238,N_86,N_4596);
or U19239 (N_19239,N_6740,N_2722);
xnor U19240 (N_19240,N_8492,N_5326);
and U19241 (N_19241,N_8386,N_9151);
xor U19242 (N_19242,N_6690,N_5427);
nand U19243 (N_19243,N_5407,N_3043);
xnor U19244 (N_19244,N_264,N_6134);
nand U19245 (N_19245,N_4428,N_57);
xnor U19246 (N_19246,N_1568,N_9986);
or U19247 (N_19247,N_7489,N_7535);
nand U19248 (N_19248,N_3152,N_6891);
and U19249 (N_19249,N_2290,N_3535);
nand U19250 (N_19250,N_5790,N_610);
or U19251 (N_19251,N_9432,N_437);
nor U19252 (N_19252,N_2040,N_4872);
nand U19253 (N_19253,N_4010,N_7893);
nand U19254 (N_19254,N_5347,N_3954);
nand U19255 (N_19255,N_229,N_4977);
and U19256 (N_19256,N_7895,N_9857);
or U19257 (N_19257,N_6042,N_6848);
or U19258 (N_19258,N_7841,N_6409);
or U19259 (N_19259,N_554,N_7454);
or U19260 (N_19260,N_923,N_5126);
xor U19261 (N_19261,N_2070,N_6845);
or U19262 (N_19262,N_9567,N_1113);
and U19263 (N_19263,N_2907,N_8833);
or U19264 (N_19264,N_4291,N_5490);
nand U19265 (N_19265,N_1431,N_2713);
and U19266 (N_19266,N_5173,N_4460);
nor U19267 (N_19267,N_4612,N_1814);
nand U19268 (N_19268,N_7282,N_3678);
or U19269 (N_19269,N_1879,N_644);
nand U19270 (N_19270,N_8214,N_3860);
nand U19271 (N_19271,N_7359,N_8353);
xor U19272 (N_19272,N_4186,N_5034);
or U19273 (N_19273,N_5982,N_3386);
nand U19274 (N_19274,N_3683,N_9240);
and U19275 (N_19275,N_3755,N_1211);
xor U19276 (N_19276,N_8950,N_3793);
or U19277 (N_19277,N_2098,N_4438);
nor U19278 (N_19278,N_5520,N_2150);
or U19279 (N_19279,N_8825,N_6745);
and U19280 (N_19280,N_1589,N_1095);
and U19281 (N_19281,N_1851,N_7128);
or U19282 (N_19282,N_7399,N_8516);
and U19283 (N_19283,N_4660,N_9662);
nand U19284 (N_19284,N_6010,N_5892);
nand U19285 (N_19285,N_7815,N_8425);
nor U19286 (N_19286,N_1018,N_7540);
or U19287 (N_19287,N_5131,N_4751);
and U19288 (N_19288,N_3657,N_772);
and U19289 (N_19289,N_7743,N_4742);
nand U19290 (N_19290,N_4802,N_808);
xor U19291 (N_19291,N_4369,N_2290);
nand U19292 (N_19292,N_9629,N_9637);
and U19293 (N_19293,N_589,N_988);
and U19294 (N_19294,N_1811,N_2324);
or U19295 (N_19295,N_2093,N_3539);
nor U19296 (N_19296,N_1404,N_8625);
nor U19297 (N_19297,N_4608,N_6087);
or U19298 (N_19298,N_4515,N_4948);
nand U19299 (N_19299,N_8123,N_2132);
nor U19300 (N_19300,N_1199,N_1535);
nand U19301 (N_19301,N_1731,N_892);
nand U19302 (N_19302,N_5632,N_844);
xnor U19303 (N_19303,N_4643,N_9693);
nand U19304 (N_19304,N_2009,N_6302);
nor U19305 (N_19305,N_1670,N_3141);
and U19306 (N_19306,N_117,N_2417);
and U19307 (N_19307,N_2304,N_9856);
and U19308 (N_19308,N_259,N_9051);
nand U19309 (N_19309,N_4009,N_3459);
nor U19310 (N_19310,N_8164,N_7000);
nand U19311 (N_19311,N_8110,N_5299);
nand U19312 (N_19312,N_900,N_8931);
nand U19313 (N_19313,N_8198,N_7150);
nor U19314 (N_19314,N_4157,N_8011);
and U19315 (N_19315,N_7850,N_3331);
nand U19316 (N_19316,N_2777,N_3750);
nand U19317 (N_19317,N_4903,N_7917);
nand U19318 (N_19318,N_2986,N_5463);
and U19319 (N_19319,N_7704,N_1896);
nor U19320 (N_19320,N_9995,N_9884);
and U19321 (N_19321,N_7065,N_8219);
nand U19322 (N_19322,N_2437,N_1839);
nor U19323 (N_19323,N_6758,N_9545);
nor U19324 (N_19324,N_9269,N_7514);
nor U19325 (N_19325,N_8488,N_1564);
nor U19326 (N_19326,N_6001,N_4429);
and U19327 (N_19327,N_5708,N_6408);
and U19328 (N_19328,N_3907,N_6267);
nand U19329 (N_19329,N_4522,N_7698);
or U19330 (N_19330,N_8695,N_4663);
and U19331 (N_19331,N_767,N_5473);
nand U19332 (N_19332,N_5531,N_4402);
nor U19333 (N_19333,N_2870,N_5674);
nand U19334 (N_19334,N_8020,N_9659);
and U19335 (N_19335,N_1953,N_7444);
nand U19336 (N_19336,N_5515,N_9610);
and U19337 (N_19337,N_196,N_5614);
xor U19338 (N_19338,N_9061,N_3442);
and U19339 (N_19339,N_2992,N_1126);
nand U19340 (N_19340,N_6161,N_3233);
or U19341 (N_19341,N_6241,N_6713);
nand U19342 (N_19342,N_4535,N_4339);
nor U19343 (N_19343,N_5981,N_9393);
nor U19344 (N_19344,N_6965,N_1172);
nor U19345 (N_19345,N_8983,N_2260);
nor U19346 (N_19346,N_8620,N_407);
and U19347 (N_19347,N_7076,N_7038);
and U19348 (N_19348,N_2037,N_9194);
nand U19349 (N_19349,N_6382,N_2459);
and U19350 (N_19350,N_6592,N_7915);
nor U19351 (N_19351,N_7958,N_6635);
or U19352 (N_19352,N_489,N_5999);
or U19353 (N_19353,N_6701,N_3438);
or U19354 (N_19354,N_6273,N_857);
nand U19355 (N_19355,N_8528,N_1702);
nor U19356 (N_19356,N_6826,N_7283);
or U19357 (N_19357,N_4494,N_3905);
or U19358 (N_19358,N_7527,N_5730);
and U19359 (N_19359,N_9774,N_3562);
nor U19360 (N_19360,N_6125,N_1557);
and U19361 (N_19361,N_2770,N_8864);
and U19362 (N_19362,N_3195,N_2847);
nor U19363 (N_19363,N_5418,N_8017);
xor U19364 (N_19364,N_9681,N_4588);
nor U19365 (N_19365,N_961,N_1716);
and U19366 (N_19366,N_3049,N_2849);
nand U19367 (N_19367,N_9483,N_9705);
and U19368 (N_19368,N_7840,N_1651);
or U19369 (N_19369,N_8987,N_6404);
or U19370 (N_19370,N_1726,N_4198);
nor U19371 (N_19371,N_1370,N_5085);
nand U19372 (N_19372,N_5338,N_5419);
or U19373 (N_19373,N_7907,N_8544);
xor U19374 (N_19374,N_6232,N_8758);
xor U19375 (N_19375,N_3211,N_44);
or U19376 (N_19376,N_3428,N_2959);
and U19377 (N_19377,N_7677,N_8670);
and U19378 (N_19378,N_4545,N_2393);
nand U19379 (N_19379,N_2826,N_1697);
nor U19380 (N_19380,N_2846,N_4736);
or U19381 (N_19381,N_6416,N_9778);
xnor U19382 (N_19382,N_9566,N_985);
nor U19383 (N_19383,N_3834,N_5829);
and U19384 (N_19384,N_6604,N_9844);
and U19385 (N_19385,N_6011,N_757);
xnor U19386 (N_19386,N_574,N_187);
and U19387 (N_19387,N_3597,N_2120);
and U19388 (N_19388,N_6733,N_8629);
and U19389 (N_19389,N_4471,N_5187);
or U19390 (N_19390,N_7711,N_9256);
nor U19391 (N_19391,N_7786,N_136);
nor U19392 (N_19392,N_3457,N_2128);
nor U19393 (N_19393,N_9912,N_1385);
or U19394 (N_19394,N_1798,N_3411);
and U19395 (N_19395,N_7763,N_675);
or U19396 (N_19396,N_3010,N_1220);
nand U19397 (N_19397,N_4182,N_3013);
nand U19398 (N_19398,N_3683,N_1691);
nor U19399 (N_19399,N_6899,N_7111);
or U19400 (N_19400,N_4520,N_5073);
nand U19401 (N_19401,N_8519,N_8097);
and U19402 (N_19402,N_8900,N_9982);
nand U19403 (N_19403,N_3345,N_1011);
xor U19404 (N_19404,N_2072,N_8782);
nand U19405 (N_19405,N_1031,N_432);
xnor U19406 (N_19406,N_2042,N_7554);
nand U19407 (N_19407,N_1920,N_3846);
xnor U19408 (N_19408,N_9378,N_551);
nand U19409 (N_19409,N_1770,N_5095);
nand U19410 (N_19410,N_6318,N_8196);
xnor U19411 (N_19411,N_3257,N_7802);
xnor U19412 (N_19412,N_2891,N_6540);
nand U19413 (N_19413,N_3725,N_564);
nor U19414 (N_19414,N_1040,N_1202);
nand U19415 (N_19415,N_9858,N_5438);
or U19416 (N_19416,N_6578,N_5679);
nand U19417 (N_19417,N_4717,N_806);
or U19418 (N_19418,N_1996,N_4133);
nor U19419 (N_19419,N_9613,N_9586);
nand U19420 (N_19420,N_4454,N_9455);
nor U19421 (N_19421,N_906,N_6103);
nand U19422 (N_19422,N_892,N_3399);
nor U19423 (N_19423,N_4881,N_6744);
nand U19424 (N_19424,N_7265,N_697);
or U19425 (N_19425,N_5298,N_7524);
nor U19426 (N_19426,N_4017,N_6804);
nand U19427 (N_19427,N_8812,N_4430);
nand U19428 (N_19428,N_1055,N_2934);
nor U19429 (N_19429,N_5074,N_605);
nand U19430 (N_19430,N_5781,N_7783);
nor U19431 (N_19431,N_5502,N_3619);
nor U19432 (N_19432,N_4456,N_4156);
xor U19433 (N_19433,N_3310,N_8988);
or U19434 (N_19434,N_8112,N_1213);
or U19435 (N_19435,N_1490,N_7870);
xor U19436 (N_19436,N_9551,N_9108);
or U19437 (N_19437,N_6778,N_3688);
nor U19438 (N_19438,N_2706,N_3540);
and U19439 (N_19439,N_1868,N_8508);
and U19440 (N_19440,N_7264,N_7682);
or U19441 (N_19441,N_3029,N_7776);
nor U19442 (N_19442,N_7752,N_8142);
nand U19443 (N_19443,N_98,N_1821);
nand U19444 (N_19444,N_1976,N_4768);
nor U19445 (N_19445,N_4467,N_9773);
nand U19446 (N_19446,N_8157,N_8124);
nand U19447 (N_19447,N_1803,N_5319);
nor U19448 (N_19448,N_3884,N_21);
and U19449 (N_19449,N_2876,N_6057);
or U19450 (N_19450,N_3446,N_3160);
nor U19451 (N_19451,N_5446,N_9215);
or U19452 (N_19452,N_7976,N_9843);
or U19453 (N_19453,N_3070,N_4038);
nor U19454 (N_19454,N_9423,N_7151);
and U19455 (N_19455,N_712,N_5813);
xnor U19456 (N_19456,N_5003,N_7914);
nand U19457 (N_19457,N_5573,N_4907);
or U19458 (N_19458,N_6866,N_2436);
or U19459 (N_19459,N_2228,N_8808);
nand U19460 (N_19460,N_5736,N_6826);
and U19461 (N_19461,N_1547,N_1413);
and U19462 (N_19462,N_5759,N_2317);
nor U19463 (N_19463,N_2124,N_5658);
nand U19464 (N_19464,N_7116,N_3046);
nor U19465 (N_19465,N_4538,N_6511);
and U19466 (N_19466,N_3092,N_1760);
and U19467 (N_19467,N_5892,N_6347);
nand U19468 (N_19468,N_6646,N_7925);
nand U19469 (N_19469,N_5907,N_9711);
nand U19470 (N_19470,N_9600,N_1604);
or U19471 (N_19471,N_6892,N_8864);
or U19472 (N_19472,N_8448,N_2494);
or U19473 (N_19473,N_4974,N_9948);
nor U19474 (N_19474,N_1243,N_4134);
nor U19475 (N_19475,N_4183,N_1785);
and U19476 (N_19476,N_8811,N_4623);
and U19477 (N_19477,N_1439,N_8912);
nor U19478 (N_19478,N_4728,N_7076);
and U19479 (N_19479,N_3772,N_4197);
nand U19480 (N_19480,N_2688,N_5861);
nand U19481 (N_19481,N_7698,N_9031);
or U19482 (N_19482,N_8671,N_2911);
nand U19483 (N_19483,N_2602,N_4684);
nand U19484 (N_19484,N_6826,N_2234);
nand U19485 (N_19485,N_4491,N_4158);
and U19486 (N_19486,N_3831,N_2229);
nor U19487 (N_19487,N_3197,N_914);
and U19488 (N_19488,N_6417,N_6279);
nor U19489 (N_19489,N_2588,N_4960);
or U19490 (N_19490,N_9731,N_9071);
nand U19491 (N_19491,N_1208,N_555);
nor U19492 (N_19492,N_2752,N_9504);
nor U19493 (N_19493,N_2206,N_2321);
and U19494 (N_19494,N_1628,N_8854);
or U19495 (N_19495,N_1648,N_487);
or U19496 (N_19496,N_1931,N_4684);
or U19497 (N_19497,N_1812,N_731);
nand U19498 (N_19498,N_409,N_6583);
and U19499 (N_19499,N_9652,N_6473);
or U19500 (N_19500,N_2680,N_4265);
and U19501 (N_19501,N_378,N_5309);
nand U19502 (N_19502,N_8117,N_2436);
and U19503 (N_19503,N_747,N_3219);
nor U19504 (N_19504,N_8710,N_5996);
nor U19505 (N_19505,N_4647,N_9182);
and U19506 (N_19506,N_4049,N_4226);
xor U19507 (N_19507,N_5184,N_759);
or U19508 (N_19508,N_1431,N_9427);
nor U19509 (N_19509,N_1728,N_6741);
xnor U19510 (N_19510,N_1015,N_4639);
or U19511 (N_19511,N_5126,N_5763);
nand U19512 (N_19512,N_3469,N_247);
and U19513 (N_19513,N_4265,N_5873);
nor U19514 (N_19514,N_6963,N_7390);
nand U19515 (N_19515,N_4975,N_820);
nor U19516 (N_19516,N_5204,N_4784);
and U19517 (N_19517,N_7406,N_5656);
nor U19518 (N_19518,N_5986,N_727);
nor U19519 (N_19519,N_713,N_3287);
nand U19520 (N_19520,N_4892,N_5448);
nor U19521 (N_19521,N_534,N_3585);
nand U19522 (N_19522,N_2886,N_4840);
nand U19523 (N_19523,N_3462,N_5029);
and U19524 (N_19524,N_6647,N_441);
and U19525 (N_19525,N_5101,N_5901);
and U19526 (N_19526,N_2522,N_6460);
nand U19527 (N_19527,N_760,N_8387);
nand U19528 (N_19528,N_69,N_878);
and U19529 (N_19529,N_2097,N_2646);
nand U19530 (N_19530,N_2883,N_262);
and U19531 (N_19531,N_6911,N_7544);
nand U19532 (N_19532,N_3774,N_3082);
or U19533 (N_19533,N_4471,N_3719);
nor U19534 (N_19534,N_4523,N_6834);
and U19535 (N_19535,N_8277,N_4376);
nor U19536 (N_19536,N_6145,N_243);
xnor U19537 (N_19537,N_1686,N_312);
or U19538 (N_19538,N_8705,N_6569);
nor U19539 (N_19539,N_8040,N_6301);
xnor U19540 (N_19540,N_1843,N_8933);
nor U19541 (N_19541,N_4340,N_6310);
nand U19542 (N_19542,N_5430,N_7729);
nand U19543 (N_19543,N_3704,N_253);
and U19544 (N_19544,N_3626,N_6039);
nand U19545 (N_19545,N_2657,N_1053);
or U19546 (N_19546,N_1979,N_7295);
nand U19547 (N_19547,N_7773,N_9595);
and U19548 (N_19548,N_7358,N_3150);
nor U19549 (N_19549,N_5308,N_851);
or U19550 (N_19550,N_9613,N_3791);
nor U19551 (N_19551,N_8162,N_1072);
nand U19552 (N_19552,N_6347,N_66);
or U19553 (N_19553,N_6063,N_1012);
nor U19554 (N_19554,N_8876,N_4543);
nor U19555 (N_19555,N_8042,N_362);
nand U19556 (N_19556,N_7886,N_3750);
nand U19557 (N_19557,N_8315,N_8529);
or U19558 (N_19558,N_4034,N_5652);
nor U19559 (N_19559,N_5068,N_3714);
and U19560 (N_19560,N_7812,N_2123);
xor U19561 (N_19561,N_7366,N_7754);
nor U19562 (N_19562,N_4997,N_3672);
nand U19563 (N_19563,N_287,N_354);
nand U19564 (N_19564,N_9072,N_6256);
nor U19565 (N_19565,N_1721,N_9479);
nor U19566 (N_19566,N_8547,N_957);
nand U19567 (N_19567,N_1136,N_8421);
nand U19568 (N_19568,N_7158,N_8565);
nand U19569 (N_19569,N_6202,N_9378);
nand U19570 (N_19570,N_6421,N_7305);
or U19571 (N_19571,N_518,N_3262);
and U19572 (N_19572,N_9783,N_1255);
nand U19573 (N_19573,N_8445,N_2463);
and U19574 (N_19574,N_9192,N_7891);
or U19575 (N_19575,N_4572,N_2610);
and U19576 (N_19576,N_4189,N_6329);
and U19577 (N_19577,N_8332,N_7936);
xnor U19578 (N_19578,N_5575,N_1654);
or U19579 (N_19579,N_6251,N_5478);
nor U19580 (N_19580,N_9948,N_2151);
and U19581 (N_19581,N_2977,N_7478);
nor U19582 (N_19582,N_3796,N_1892);
nor U19583 (N_19583,N_2511,N_1174);
xor U19584 (N_19584,N_4314,N_2551);
or U19585 (N_19585,N_5238,N_430);
or U19586 (N_19586,N_2666,N_9873);
nand U19587 (N_19587,N_3879,N_2905);
nand U19588 (N_19588,N_8672,N_3162);
nor U19589 (N_19589,N_6761,N_9904);
nor U19590 (N_19590,N_358,N_6810);
xnor U19591 (N_19591,N_303,N_1820);
xor U19592 (N_19592,N_6748,N_4089);
or U19593 (N_19593,N_7273,N_3908);
xor U19594 (N_19594,N_4968,N_7018);
and U19595 (N_19595,N_6517,N_4773);
or U19596 (N_19596,N_5783,N_8113);
xnor U19597 (N_19597,N_4120,N_1713);
nand U19598 (N_19598,N_5740,N_6695);
nor U19599 (N_19599,N_6043,N_2441);
and U19600 (N_19600,N_4697,N_3477);
or U19601 (N_19601,N_6371,N_9709);
or U19602 (N_19602,N_4904,N_5985);
and U19603 (N_19603,N_8774,N_9560);
nor U19604 (N_19604,N_2183,N_631);
and U19605 (N_19605,N_65,N_8236);
nor U19606 (N_19606,N_5104,N_1247);
nor U19607 (N_19607,N_7370,N_9171);
nor U19608 (N_19608,N_9969,N_1395);
and U19609 (N_19609,N_740,N_7630);
and U19610 (N_19610,N_7851,N_3699);
and U19611 (N_19611,N_9328,N_923);
nor U19612 (N_19612,N_4239,N_8163);
or U19613 (N_19613,N_6971,N_8292);
or U19614 (N_19614,N_750,N_3877);
or U19615 (N_19615,N_9957,N_401);
xor U19616 (N_19616,N_1935,N_9114);
xor U19617 (N_19617,N_6605,N_5500);
xnor U19618 (N_19618,N_9116,N_9517);
nand U19619 (N_19619,N_9556,N_6625);
nor U19620 (N_19620,N_602,N_3471);
nand U19621 (N_19621,N_2695,N_9980);
nand U19622 (N_19622,N_7366,N_7159);
or U19623 (N_19623,N_3063,N_3527);
nor U19624 (N_19624,N_4943,N_8378);
nor U19625 (N_19625,N_6572,N_365);
nand U19626 (N_19626,N_247,N_9000);
nor U19627 (N_19627,N_1941,N_481);
nand U19628 (N_19628,N_1049,N_9977);
or U19629 (N_19629,N_4606,N_2875);
nor U19630 (N_19630,N_413,N_3364);
nor U19631 (N_19631,N_8765,N_7728);
nor U19632 (N_19632,N_1886,N_9818);
nor U19633 (N_19633,N_2109,N_9460);
nand U19634 (N_19634,N_722,N_684);
nor U19635 (N_19635,N_4234,N_8472);
and U19636 (N_19636,N_5451,N_4254);
and U19637 (N_19637,N_3055,N_4191);
nor U19638 (N_19638,N_7415,N_8734);
xnor U19639 (N_19639,N_2048,N_4601);
and U19640 (N_19640,N_9426,N_5569);
nor U19641 (N_19641,N_4334,N_870);
nor U19642 (N_19642,N_6918,N_2330);
nand U19643 (N_19643,N_6047,N_3744);
or U19644 (N_19644,N_1954,N_8482);
xnor U19645 (N_19645,N_6048,N_2549);
xnor U19646 (N_19646,N_5542,N_146);
and U19647 (N_19647,N_1291,N_6984);
nand U19648 (N_19648,N_5444,N_4068);
nand U19649 (N_19649,N_7555,N_4285);
nand U19650 (N_19650,N_715,N_2192);
or U19651 (N_19651,N_2291,N_7633);
nand U19652 (N_19652,N_8410,N_3978);
xor U19653 (N_19653,N_9262,N_1628);
and U19654 (N_19654,N_2236,N_1345);
nor U19655 (N_19655,N_5908,N_2943);
nor U19656 (N_19656,N_6254,N_4704);
and U19657 (N_19657,N_9994,N_2620);
and U19658 (N_19658,N_7519,N_4623);
nor U19659 (N_19659,N_6540,N_5968);
or U19660 (N_19660,N_8194,N_6080);
xor U19661 (N_19661,N_4822,N_2595);
xor U19662 (N_19662,N_2482,N_4669);
and U19663 (N_19663,N_7140,N_2624);
or U19664 (N_19664,N_2273,N_7939);
nand U19665 (N_19665,N_5492,N_6273);
or U19666 (N_19666,N_4095,N_9432);
nor U19667 (N_19667,N_3868,N_3379);
and U19668 (N_19668,N_6940,N_7383);
or U19669 (N_19669,N_9063,N_4659);
or U19670 (N_19670,N_8509,N_8207);
nand U19671 (N_19671,N_2423,N_1146);
xnor U19672 (N_19672,N_9153,N_9056);
nand U19673 (N_19673,N_7357,N_7641);
nand U19674 (N_19674,N_1492,N_4172);
or U19675 (N_19675,N_3614,N_4314);
nor U19676 (N_19676,N_2609,N_7990);
or U19677 (N_19677,N_6125,N_8166);
and U19678 (N_19678,N_2364,N_581);
nor U19679 (N_19679,N_567,N_974);
or U19680 (N_19680,N_7744,N_902);
xnor U19681 (N_19681,N_3469,N_2137);
nand U19682 (N_19682,N_862,N_7218);
and U19683 (N_19683,N_3486,N_8592);
or U19684 (N_19684,N_4722,N_2663);
or U19685 (N_19685,N_9084,N_2303);
nand U19686 (N_19686,N_1314,N_5637);
xnor U19687 (N_19687,N_27,N_7550);
xor U19688 (N_19688,N_6729,N_6739);
nor U19689 (N_19689,N_3579,N_3827);
or U19690 (N_19690,N_5667,N_927);
nor U19691 (N_19691,N_9551,N_7418);
and U19692 (N_19692,N_1458,N_4263);
and U19693 (N_19693,N_9630,N_269);
nor U19694 (N_19694,N_8432,N_2068);
and U19695 (N_19695,N_6856,N_8060);
nor U19696 (N_19696,N_6134,N_4043);
or U19697 (N_19697,N_4878,N_5981);
nand U19698 (N_19698,N_1809,N_4424);
nor U19699 (N_19699,N_4834,N_4384);
nor U19700 (N_19700,N_2359,N_886);
and U19701 (N_19701,N_3617,N_3793);
nor U19702 (N_19702,N_8062,N_7206);
and U19703 (N_19703,N_6101,N_9089);
nand U19704 (N_19704,N_9432,N_4016);
or U19705 (N_19705,N_9668,N_3736);
nor U19706 (N_19706,N_7888,N_3581);
nand U19707 (N_19707,N_146,N_5361);
or U19708 (N_19708,N_8715,N_8652);
or U19709 (N_19709,N_2786,N_9031);
nand U19710 (N_19710,N_2408,N_8157);
xor U19711 (N_19711,N_2058,N_5922);
or U19712 (N_19712,N_8944,N_9486);
and U19713 (N_19713,N_5788,N_7547);
nand U19714 (N_19714,N_8753,N_1992);
or U19715 (N_19715,N_3519,N_6390);
or U19716 (N_19716,N_6997,N_6329);
and U19717 (N_19717,N_8634,N_1273);
nor U19718 (N_19718,N_3333,N_9865);
nand U19719 (N_19719,N_5814,N_8023);
xnor U19720 (N_19720,N_7508,N_7302);
or U19721 (N_19721,N_9367,N_8366);
xor U19722 (N_19722,N_8112,N_5925);
nand U19723 (N_19723,N_8302,N_16);
nand U19724 (N_19724,N_5060,N_336);
nor U19725 (N_19725,N_7105,N_8395);
or U19726 (N_19726,N_7151,N_4404);
nand U19727 (N_19727,N_8375,N_5976);
or U19728 (N_19728,N_1402,N_5822);
nor U19729 (N_19729,N_4775,N_2819);
xnor U19730 (N_19730,N_164,N_5009);
nor U19731 (N_19731,N_1069,N_7078);
nand U19732 (N_19732,N_3021,N_8461);
and U19733 (N_19733,N_495,N_856);
nand U19734 (N_19734,N_6537,N_8387);
nand U19735 (N_19735,N_3836,N_3380);
nand U19736 (N_19736,N_207,N_4271);
nand U19737 (N_19737,N_1794,N_9115);
xnor U19738 (N_19738,N_4416,N_793);
or U19739 (N_19739,N_8616,N_8230);
and U19740 (N_19740,N_4610,N_4180);
and U19741 (N_19741,N_8756,N_7696);
nor U19742 (N_19742,N_3551,N_5451);
and U19743 (N_19743,N_8846,N_6520);
nor U19744 (N_19744,N_7900,N_9620);
nor U19745 (N_19745,N_346,N_9362);
xor U19746 (N_19746,N_192,N_1286);
nand U19747 (N_19747,N_5988,N_798);
or U19748 (N_19748,N_5772,N_3023);
nor U19749 (N_19749,N_6957,N_3016);
and U19750 (N_19750,N_4392,N_8397);
nand U19751 (N_19751,N_3899,N_6944);
or U19752 (N_19752,N_4189,N_3391);
or U19753 (N_19753,N_7419,N_4240);
or U19754 (N_19754,N_6079,N_7881);
or U19755 (N_19755,N_7771,N_3011);
nor U19756 (N_19756,N_7455,N_4399);
nand U19757 (N_19757,N_806,N_2009);
xor U19758 (N_19758,N_1071,N_6346);
and U19759 (N_19759,N_2574,N_8847);
and U19760 (N_19760,N_473,N_6912);
nand U19761 (N_19761,N_1107,N_8563);
nand U19762 (N_19762,N_20,N_3932);
or U19763 (N_19763,N_9603,N_2001);
nand U19764 (N_19764,N_6388,N_3271);
or U19765 (N_19765,N_7414,N_7705);
nand U19766 (N_19766,N_9996,N_2499);
and U19767 (N_19767,N_7944,N_9011);
or U19768 (N_19768,N_8325,N_2718);
or U19769 (N_19769,N_3052,N_6077);
nand U19770 (N_19770,N_1699,N_270);
nand U19771 (N_19771,N_1014,N_5148);
or U19772 (N_19772,N_8099,N_9171);
or U19773 (N_19773,N_8016,N_8329);
nand U19774 (N_19774,N_731,N_4432);
and U19775 (N_19775,N_2722,N_8292);
nor U19776 (N_19776,N_7265,N_4163);
nor U19777 (N_19777,N_6173,N_2614);
nand U19778 (N_19778,N_9061,N_8993);
nor U19779 (N_19779,N_6577,N_7956);
nand U19780 (N_19780,N_2125,N_4958);
and U19781 (N_19781,N_5622,N_8288);
nor U19782 (N_19782,N_7052,N_2941);
nor U19783 (N_19783,N_8458,N_1516);
nand U19784 (N_19784,N_6708,N_8948);
xnor U19785 (N_19785,N_5421,N_4785);
or U19786 (N_19786,N_6765,N_149);
xnor U19787 (N_19787,N_7190,N_2972);
xor U19788 (N_19788,N_2307,N_3902);
nand U19789 (N_19789,N_1522,N_9263);
nor U19790 (N_19790,N_5999,N_7229);
or U19791 (N_19791,N_2027,N_872);
nor U19792 (N_19792,N_8685,N_6380);
nor U19793 (N_19793,N_1849,N_9856);
xnor U19794 (N_19794,N_1557,N_8792);
and U19795 (N_19795,N_6553,N_6296);
and U19796 (N_19796,N_8320,N_8684);
or U19797 (N_19797,N_5052,N_9648);
or U19798 (N_19798,N_4033,N_8960);
and U19799 (N_19799,N_358,N_6397);
nand U19800 (N_19800,N_7610,N_3351);
nor U19801 (N_19801,N_4264,N_6719);
or U19802 (N_19802,N_1168,N_9589);
nor U19803 (N_19803,N_3863,N_5536);
nor U19804 (N_19804,N_4343,N_832);
nor U19805 (N_19805,N_9172,N_5395);
nor U19806 (N_19806,N_9909,N_2722);
or U19807 (N_19807,N_8133,N_6982);
nor U19808 (N_19808,N_4214,N_4037);
and U19809 (N_19809,N_5740,N_8608);
or U19810 (N_19810,N_9490,N_2823);
nand U19811 (N_19811,N_8406,N_3393);
and U19812 (N_19812,N_6780,N_4942);
nor U19813 (N_19813,N_1557,N_9535);
nor U19814 (N_19814,N_9961,N_6731);
or U19815 (N_19815,N_6232,N_9256);
nor U19816 (N_19816,N_1258,N_4576);
or U19817 (N_19817,N_991,N_7001);
nand U19818 (N_19818,N_6602,N_470);
or U19819 (N_19819,N_1259,N_3004);
or U19820 (N_19820,N_9574,N_2899);
nor U19821 (N_19821,N_2239,N_4228);
and U19822 (N_19822,N_6908,N_9897);
nand U19823 (N_19823,N_489,N_279);
or U19824 (N_19824,N_6321,N_5112);
and U19825 (N_19825,N_782,N_4871);
xnor U19826 (N_19826,N_8836,N_6010);
xnor U19827 (N_19827,N_69,N_6964);
nor U19828 (N_19828,N_6048,N_4866);
or U19829 (N_19829,N_6197,N_4669);
and U19830 (N_19830,N_4866,N_6305);
nand U19831 (N_19831,N_9873,N_3806);
and U19832 (N_19832,N_4061,N_2630);
and U19833 (N_19833,N_7734,N_8654);
or U19834 (N_19834,N_5667,N_4838);
nand U19835 (N_19835,N_5293,N_7617);
and U19836 (N_19836,N_2654,N_3496);
nand U19837 (N_19837,N_6502,N_8776);
nand U19838 (N_19838,N_5360,N_7052);
nor U19839 (N_19839,N_4523,N_1387);
nor U19840 (N_19840,N_9454,N_6988);
or U19841 (N_19841,N_7746,N_1545);
and U19842 (N_19842,N_7304,N_4500);
or U19843 (N_19843,N_3924,N_777);
and U19844 (N_19844,N_5986,N_3607);
nand U19845 (N_19845,N_3315,N_1034);
nand U19846 (N_19846,N_3405,N_4327);
nor U19847 (N_19847,N_4697,N_6316);
nand U19848 (N_19848,N_3757,N_8098);
and U19849 (N_19849,N_3451,N_1565);
and U19850 (N_19850,N_6676,N_5143);
or U19851 (N_19851,N_931,N_1306);
and U19852 (N_19852,N_5554,N_5371);
or U19853 (N_19853,N_2927,N_2883);
nand U19854 (N_19854,N_6283,N_7739);
nor U19855 (N_19855,N_2395,N_6738);
and U19856 (N_19856,N_6001,N_6337);
xor U19857 (N_19857,N_6092,N_3208);
and U19858 (N_19858,N_4123,N_9471);
or U19859 (N_19859,N_7516,N_5691);
and U19860 (N_19860,N_9562,N_9927);
or U19861 (N_19861,N_7708,N_5311);
and U19862 (N_19862,N_835,N_2954);
or U19863 (N_19863,N_9211,N_3636);
and U19864 (N_19864,N_789,N_8948);
nand U19865 (N_19865,N_8454,N_7575);
and U19866 (N_19866,N_1988,N_2298);
nor U19867 (N_19867,N_9985,N_5883);
xor U19868 (N_19868,N_303,N_6522);
nor U19869 (N_19869,N_3134,N_4897);
and U19870 (N_19870,N_4321,N_5608);
nor U19871 (N_19871,N_218,N_843);
and U19872 (N_19872,N_9431,N_9248);
nand U19873 (N_19873,N_5620,N_9194);
or U19874 (N_19874,N_7476,N_9763);
nor U19875 (N_19875,N_2531,N_435);
nand U19876 (N_19876,N_8614,N_5176);
and U19877 (N_19877,N_747,N_8862);
xnor U19878 (N_19878,N_928,N_4170);
nand U19879 (N_19879,N_2051,N_4813);
nor U19880 (N_19880,N_8224,N_5720);
nor U19881 (N_19881,N_6541,N_9234);
xor U19882 (N_19882,N_9983,N_4631);
nor U19883 (N_19883,N_8112,N_530);
xnor U19884 (N_19884,N_4171,N_1044);
and U19885 (N_19885,N_7162,N_1227);
nor U19886 (N_19886,N_9194,N_7137);
or U19887 (N_19887,N_8472,N_8390);
and U19888 (N_19888,N_8752,N_9496);
and U19889 (N_19889,N_8346,N_3869);
nand U19890 (N_19890,N_2761,N_1136);
and U19891 (N_19891,N_2919,N_6929);
or U19892 (N_19892,N_6944,N_480);
or U19893 (N_19893,N_7886,N_7805);
and U19894 (N_19894,N_3423,N_4875);
or U19895 (N_19895,N_6936,N_7536);
and U19896 (N_19896,N_678,N_2296);
nand U19897 (N_19897,N_9372,N_3001);
nor U19898 (N_19898,N_6683,N_8596);
nor U19899 (N_19899,N_2619,N_7239);
and U19900 (N_19900,N_5002,N_1744);
nand U19901 (N_19901,N_7384,N_4541);
or U19902 (N_19902,N_2702,N_7776);
and U19903 (N_19903,N_2783,N_6878);
nor U19904 (N_19904,N_9238,N_8678);
or U19905 (N_19905,N_3960,N_4743);
and U19906 (N_19906,N_811,N_339);
and U19907 (N_19907,N_6040,N_6732);
nor U19908 (N_19908,N_1759,N_7689);
and U19909 (N_19909,N_8003,N_3155);
xnor U19910 (N_19910,N_691,N_897);
or U19911 (N_19911,N_7115,N_2206);
and U19912 (N_19912,N_4664,N_2100);
or U19913 (N_19913,N_2586,N_7264);
nor U19914 (N_19914,N_8834,N_1713);
and U19915 (N_19915,N_2841,N_4994);
nand U19916 (N_19916,N_8326,N_7865);
or U19917 (N_19917,N_5016,N_8484);
or U19918 (N_19918,N_1952,N_5678);
or U19919 (N_19919,N_6720,N_8258);
xor U19920 (N_19920,N_108,N_7064);
xor U19921 (N_19921,N_6585,N_5311);
nand U19922 (N_19922,N_3972,N_1083);
nand U19923 (N_19923,N_8700,N_6796);
and U19924 (N_19924,N_3993,N_1388);
nand U19925 (N_19925,N_7017,N_841);
or U19926 (N_19926,N_5905,N_1536);
xor U19927 (N_19927,N_3391,N_5472);
or U19928 (N_19928,N_8412,N_8263);
and U19929 (N_19929,N_7307,N_2061);
and U19930 (N_19930,N_7453,N_8839);
or U19931 (N_19931,N_6819,N_8111);
nand U19932 (N_19932,N_6487,N_4508);
nor U19933 (N_19933,N_1858,N_5919);
or U19934 (N_19934,N_6986,N_1644);
and U19935 (N_19935,N_2425,N_2570);
or U19936 (N_19936,N_7020,N_6934);
or U19937 (N_19937,N_418,N_4702);
or U19938 (N_19938,N_9791,N_5542);
and U19939 (N_19939,N_4998,N_7547);
or U19940 (N_19940,N_6503,N_1627);
nand U19941 (N_19941,N_2139,N_7797);
nor U19942 (N_19942,N_8315,N_7302);
nand U19943 (N_19943,N_4740,N_3692);
nand U19944 (N_19944,N_3953,N_3991);
nor U19945 (N_19945,N_7835,N_513);
and U19946 (N_19946,N_233,N_7039);
or U19947 (N_19947,N_8378,N_1734);
and U19948 (N_19948,N_5425,N_7997);
nor U19949 (N_19949,N_2618,N_7265);
nand U19950 (N_19950,N_7036,N_3685);
or U19951 (N_19951,N_7964,N_4894);
nor U19952 (N_19952,N_1804,N_6453);
nor U19953 (N_19953,N_3059,N_638);
nand U19954 (N_19954,N_2350,N_2119);
and U19955 (N_19955,N_4160,N_7099);
nor U19956 (N_19956,N_9854,N_499);
or U19957 (N_19957,N_3136,N_7970);
and U19958 (N_19958,N_2774,N_6090);
or U19959 (N_19959,N_499,N_3792);
or U19960 (N_19960,N_9797,N_3905);
nor U19961 (N_19961,N_5284,N_6459);
nand U19962 (N_19962,N_6946,N_465);
nor U19963 (N_19963,N_6994,N_3483);
nor U19964 (N_19964,N_9664,N_6787);
nand U19965 (N_19965,N_249,N_2841);
or U19966 (N_19966,N_5512,N_6885);
and U19967 (N_19967,N_48,N_8367);
nor U19968 (N_19968,N_9156,N_244);
nand U19969 (N_19969,N_8616,N_3841);
xnor U19970 (N_19970,N_5375,N_7247);
or U19971 (N_19971,N_5237,N_1568);
and U19972 (N_19972,N_1218,N_622);
nor U19973 (N_19973,N_7575,N_6756);
and U19974 (N_19974,N_1715,N_9722);
xnor U19975 (N_19975,N_3767,N_4862);
and U19976 (N_19976,N_8067,N_6266);
nand U19977 (N_19977,N_5030,N_6400);
nor U19978 (N_19978,N_1632,N_3672);
or U19979 (N_19979,N_440,N_7392);
nand U19980 (N_19980,N_9290,N_8646);
or U19981 (N_19981,N_6990,N_8372);
and U19982 (N_19982,N_5668,N_7709);
or U19983 (N_19983,N_7552,N_221);
or U19984 (N_19984,N_8338,N_4238);
or U19985 (N_19985,N_8607,N_4814);
nand U19986 (N_19986,N_4979,N_7360);
nand U19987 (N_19987,N_1916,N_5186);
nand U19988 (N_19988,N_837,N_6305);
nor U19989 (N_19989,N_4358,N_5744);
nand U19990 (N_19990,N_7691,N_4043);
nor U19991 (N_19991,N_28,N_7170);
nand U19992 (N_19992,N_1892,N_3705);
nor U19993 (N_19993,N_6559,N_9399);
and U19994 (N_19994,N_6763,N_1152);
nor U19995 (N_19995,N_8880,N_116);
or U19996 (N_19996,N_3468,N_3234);
nor U19997 (N_19997,N_9911,N_5272);
nand U19998 (N_19998,N_2237,N_1343);
or U19999 (N_19999,N_1386,N_6822);
nor U20000 (N_20000,N_10622,N_16132);
nor U20001 (N_20001,N_14151,N_18746);
nand U20002 (N_20002,N_17789,N_14241);
and U20003 (N_20003,N_10553,N_19040);
and U20004 (N_20004,N_18493,N_16290);
nand U20005 (N_20005,N_19821,N_11470);
nand U20006 (N_20006,N_16162,N_11220);
nand U20007 (N_20007,N_11729,N_11508);
nor U20008 (N_20008,N_15231,N_12488);
and U20009 (N_20009,N_15956,N_12200);
and U20010 (N_20010,N_12221,N_17062);
nor U20011 (N_20011,N_14650,N_14556);
or U20012 (N_20012,N_10000,N_14861);
xor U20013 (N_20013,N_13517,N_10783);
and U20014 (N_20014,N_16967,N_19938);
xnor U20015 (N_20015,N_19733,N_13593);
and U20016 (N_20016,N_18310,N_11693);
nor U20017 (N_20017,N_18611,N_11192);
nor U20018 (N_20018,N_18191,N_15138);
or U20019 (N_20019,N_16651,N_16098);
nor U20020 (N_20020,N_15950,N_16396);
and U20021 (N_20021,N_10775,N_12465);
nand U20022 (N_20022,N_10781,N_17361);
and U20023 (N_20023,N_18801,N_13451);
xnor U20024 (N_20024,N_13157,N_15073);
nand U20025 (N_20025,N_18932,N_18050);
or U20026 (N_20026,N_11668,N_16536);
xor U20027 (N_20027,N_12461,N_13395);
and U20028 (N_20028,N_13265,N_15514);
nand U20029 (N_20029,N_15429,N_19914);
and U20030 (N_20030,N_14212,N_16552);
nand U20031 (N_20031,N_16569,N_14865);
nand U20032 (N_20032,N_16657,N_12786);
nor U20033 (N_20033,N_14983,N_14124);
nor U20034 (N_20034,N_17324,N_17380);
and U20035 (N_20035,N_18277,N_17948);
nor U20036 (N_20036,N_10458,N_14411);
xor U20037 (N_20037,N_12083,N_10580);
or U20038 (N_20038,N_19120,N_14703);
nor U20039 (N_20039,N_17756,N_18497);
or U20040 (N_20040,N_17744,N_18342);
and U20041 (N_20041,N_12249,N_11580);
and U20042 (N_20042,N_19915,N_10241);
or U20043 (N_20043,N_18551,N_15377);
or U20044 (N_20044,N_13894,N_17214);
nor U20045 (N_20045,N_10739,N_16825);
or U20046 (N_20046,N_17343,N_12150);
or U20047 (N_20047,N_12838,N_16118);
xor U20048 (N_20048,N_10873,N_16330);
and U20049 (N_20049,N_13763,N_17894);
nand U20050 (N_20050,N_16860,N_16479);
nor U20051 (N_20051,N_12394,N_10743);
or U20052 (N_20052,N_16170,N_18414);
nand U20053 (N_20053,N_14791,N_12898);
nand U20054 (N_20054,N_16938,N_14200);
or U20055 (N_20055,N_12926,N_17913);
nand U20056 (N_20056,N_10403,N_16856);
xor U20057 (N_20057,N_10490,N_18311);
nand U20058 (N_20058,N_14425,N_12065);
or U20059 (N_20059,N_19358,N_10409);
or U20060 (N_20060,N_15407,N_15776);
nand U20061 (N_20061,N_11873,N_16289);
nand U20062 (N_20062,N_19691,N_18766);
nor U20063 (N_20063,N_10112,N_10258);
nand U20064 (N_20064,N_10015,N_11970);
xnor U20065 (N_20065,N_12025,N_13022);
xor U20066 (N_20066,N_17386,N_14955);
nand U20067 (N_20067,N_18737,N_10143);
nor U20068 (N_20068,N_10378,N_18641);
nor U20069 (N_20069,N_12193,N_10265);
and U20070 (N_20070,N_12358,N_13514);
or U20071 (N_20071,N_14548,N_14726);
nor U20072 (N_20072,N_10876,N_17503);
nor U20073 (N_20073,N_14447,N_18030);
or U20074 (N_20074,N_19085,N_19012);
nand U20075 (N_20075,N_10726,N_19848);
nor U20076 (N_20076,N_19396,N_16766);
nand U20077 (N_20077,N_16265,N_14175);
nor U20078 (N_20078,N_15541,N_19906);
nand U20079 (N_20079,N_14826,N_14603);
nand U20080 (N_20080,N_15698,N_17546);
nand U20081 (N_20081,N_13787,N_16990);
and U20082 (N_20082,N_10151,N_16325);
or U20083 (N_20083,N_14709,N_13735);
or U20084 (N_20084,N_19555,N_18224);
nand U20085 (N_20085,N_19703,N_13708);
nand U20086 (N_20086,N_15567,N_16919);
or U20087 (N_20087,N_17618,N_15819);
or U20088 (N_20088,N_15097,N_11242);
and U20089 (N_20089,N_15146,N_11350);
xnor U20090 (N_20090,N_10413,N_10847);
nor U20091 (N_20091,N_17346,N_14539);
and U20092 (N_20092,N_15584,N_16636);
xor U20093 (N_20093,N_13709,N_14812);
or U20094 (N_20094,N_17730,N_16204);
nand U20095 (N_20095,N_15659,N_14261);
or U20096 (N_20096,N_19628,N_16586);
or U20097 (N_20097,N_15553,N_18321);
or U20098 (N_20098,N_14992,N_15756);
xnor U20099 (N_20099,N_12149,N_12087);
and U20100 (N_20100,N_13486,N_15374);
nor U20101 (N_20101,N_13634,N_12923);
nand U20102 (N_20102,N_18459,N_16449);
nand U20103 (N_20103,N_12758,N_10688);
and U20104 (N_20104,N_12951,N_11285);
and U20105 (N_20105,N_11473,N_19176);
xor U20106 (N_20106,N_11030,N_17301);
nor U20107 (N_20107,N_13710,N_10609);
or U20108 (N_20108,N_16297,N_15070);
nor U20109 (N_20109,N_10655,N_18851);
nand U20110 (N_20110,N_17281,N_17275);
and U20111 (N_20111,N_13196,N_16571);
nand U20112 (N_20112,N_19936,N_18124);
nand U20113 (N_20113,N_13094,N_14941);
nand U20114 (N_20114,N_17711,N_18078);
nor U20115 (N_20115,N_17824,N_12508);
nor U20116 (N_20116,N_13799,N_18235);
nand U20117 (N_20117,N_16435,N_17011);
or U20118 (N_20118,N_10034,N_12708);
xor U20119 (N_20119,N_14572,N_10001);
or U20120 (N_20120,N_10874,N_11063);
nor U20121 (N_20121,N_13428,N_12403);
or U20122 (N_20122,N_11563,N_16150);
nand U20123 (N_20123,N_15479,N_10954);
nand U20124 (N_20124,N_17757,N_14794);
or U20125 (N_20125,N_14077,N_16584);
and U20126 (N_20126,N_11091,N_13680);
and U20127 (N_20127,N_13838,N_16273);
nor U20128 (N_20128,N_17577,N_17524);
or U20129 (N_20129,N_11309,N_14310);
nand U20130 (N_20130,N_16634,N_12267);
or U20131 (N_20131,N_13847,N_14421);
or U20132 (N_20132,N_17178,N_13633);
and U20133 (N_20133,N_13216,N_17074);
nand U20134 (N_20134,N_18290,N_15169);
nand U20135 (N_20135,N_15155,N_15878);
and U20136 (N_20136,N_10278,N_14185);
nand U20137 (N_20137,N_13726,N_19662);
and U20138 (N_20138,N_14670,N_16528);
nor U20139 (N_20139,N_12459,N_14293);
nand U20140 (N_20140,N_10399,N_13957);
or U20141 (N_20141,N_16519,N_10515);
and U20142 (N_20142,N_13504,N_19722);
or U20143 (N_20143,N_11812,N_15452);
nor U20144 (N_20144,N_12489,N_19226);
or U20145 (N_20145,N_18580,N_12326);
nand U20146 (N_20146,N_10219,N_12308);
and U20147 (N_20147,N_14712,N_14196);
or U20148 (N_20148,N_10928,N_15772);
nor U20149 (N_20149,N_14481,N_14181);
or U20150 (N_20150,N_13746,N_15646);
xnor U20151 (N_20151,N_18096,N_15545);
and U20152 (N_20152,N_14322,N_19910);
or U20153 (N_20153,N_19288,N_18619);
nor U20154 (N_20154,N_18798,N_19311);
nand U20155 (N_20155,N_12294,N_19468);
or U20156 (N_20156,N_10487,N_13788);
nor U20157 (N_20157,N_13817,N_19050);
and U20158 (N_20158,N_12866,N_12142);
nand U20159 (N_20159,N_12530,N_15111);
xor U20160 (N_20160,N_19565,N_10372);
or U20161 (N_20161,N_12713,N_13106);
and U20162 (N_20162,N_10090,N_14725);
nor U20163 (N_20163,N_16037,N_15874);
xor U20164 (N_20164,N_16935,N_15614);
and U20165 (N_20165,N_14041,N_11664);
xor U20166 (N_20166,N_12943,N_16521);
nor U20167 (N_20167,N_15876,N_11833);
xor U20168 (N_20168,N_16844,N_16728);
nand U20169 (N_20169,N_18148,N_17309);
or U20170 (N_20170,N_14119,N_16420);
nor U20171 (N_20171,N_17794,N_10193);
and U20172 (N_20172,N_10664,N_14407);
nor U20173 (N_20173,N_10358,N_15570);
nor U20174 (N_20174,N_15573,N_17403);
xor U20175 (N_20175,N_11561,N_14897);
nand U20176 (N_20176,N_10284,N_12770);
xor U20177 (N_20177,N_18442,N_14155);
nand U20178 (N_20178,N_19297,N_17328);
and U20179 (N_20179,N_13139,N_19184);
or U20180 (N_20180,N_16015,N_15781);
or U20181 (N_20181,N_14283,N_18477);
xnor U20182 (N_20182,N_13720,N_10139);
xor U20183 (N_20183,N_14027,N_10999);
or U20184 (N_20184,N_13542,N_15396);
and U20185 (N_20185,N_18372,N_11409);
nor U20186 (N_20186,N_18444,N_17293);
and U20187 (N_20187,N_16467,N_11355);
nor U20188 (N_20188,N_19015,N_10656);
and U20189 (N_20189,N_12422,N_17976);
nor U20190 (N_20190,N_16862,N_13445);
nor U20191 (N_20191,N_13148,N_16384);
xor U20192 (N_20192,N_16045,N_18591);
nand U20193 (N_20193,N_15746,N_18908);
and U20194 (N_20194,N_14692,N_12409);
xor U20195 (N_20195,N_10018,N_11912);
nor U20196 (N_20196,N_11587,N_17308);
or U20197 (N_20197,N_12888,N_12214);
xor U20198 (N_20198,N_17517,N_13315);
and U20199 (N_20199,N_12098,N_13945);
or U20200 (N_20200,N_19701,N_11365);
xnor U20201 (N_20201,N_18537,N_15962);
and U20202 (N_20202,N_16792,N_18940);
and U20203 (N_20203,N_16134,N_15778);
nand U20204 (N_20204,N_10505,N_15520);
nand U20205 (N_20205,N_16794,N_16007);
xnor U20206 (N_20206,N_18297,N_12338);
xnor U20207 (N_20207,N_14087,N_14017);
or U20208 (N_20208,N_10306,N_15859);
and U20209 (N_20209,N_18804,N_11070);
nand U20210 (N_20210,N_12840,N_14773);
xor U20211 (N_20211,N_13562,N_10389);
nand U20212 (N_20212,N_13862,N_19908);
xnor U20213 (N_20213,N_13205,N_16588);
or U20214 (N_20214,N_18540,N_12885);
nand U20215 (N_20215,N_12890,N_15044);
or U20216 (N_20216,N_15168,N_13575);
nor U20217 (N_20217,N_18958,N_14977);
nand U20218 (N_20218,N_12886,N_12134);
and U20219 (N_20219,N_13429,N_15122);
and U20220 (N_20220,N_16955,N_16771);
and U20221 (N_20221,N_19675,N_15852);
or U20222 (N_20222,N_19907,N_18455);
and U20223 (N_20223,N_18383,N_16211);
nand U20224 (N_20224,N_14048,N_10354);
nor U20225 (N_20225,N_13028,N_18351);
nand U20226 (N_20226,N_13072,N_16915);
or U20227 (N_20227,N_13034,N_13639);
nor U20228 (N_20228,N_12755,N_16814);
nand U20229 (N_20229,N_19725,N_19363);
and U20230 (N_20230,N_17411,N_19882);
nand U20231 (N_20231,N_18892,N_12113);
nor U20232 (N_20232,N_14076,N_19976);
nand U20233 (N_20233,N_17803,N_13398);
nor U20234 (N_20234,N_15658,N_16531);
and U20235 (N_20235,N_11572,N_19290);
xnor U20236 (N_20236,N_12157,N_11374);
and U20237 (N_20237,N_18332,N_18167);
and U20238 (N_20238,N_16994,N_15223);
and U20239 (N_20239,N_15544,N_17205);
or U20240 (N_20240,N_18474,N_16929);
and U20241 (N_20241,N_16733,N_16838);
nand U20242 (N_20242,N_19281,N_14642);
or U20243 (N_20243,N_15324,N_14713);
and U20244 (N_20244,N_10121,N_10115);
nand U20245 (N_20245,N_15613,N_17684);
and U20246 (N_20246,N_15526,N_16700);
or U20247 (N_20247,N_14520,N_16058);
xor U20248 (N_20248,N_13381,N_12628);
and U20249 (N_20249,N_17039,N_11139);
nand U20250 (N_20250,N_15999,N_17088);
nor U20251 (N_20251,N_17065,N_19605);
nor U20252 (N_20252,N_10849,N_10048);
nand U20253 (N_20253,N_14232,N_17516);
nor U20254 (N_20254,N_16933,N_12311);
nor U20255 (N_20255,N_14045,N_13037);
nor U20256 (N_20256,N_15257,N_17480);
nor U20257 (N_20257,N_19153,N_15854);
or U20258 (N_20258,N_15036,N_10508);
nor U20259 (N_20259,N_11719,N_19052);
and U20260 (N_20260,N_16503,N_15931);
nor U20261 (N_20261,N_17042,N_10579);
xnor U20262 (N_20262,N_11277,N_16209);
nand U20263 (N_20263,N_16119,N_16335);
nor U20264 (N_20264,N_19212,N_14590);
nor U20265 (N_20265,N_12588,N_10971);
nand U20266 (N_20266,N_15237,N_11874);
xnor U20267 (N_20267,N_16904,N_16765);
and U20268 (N_20268,N_15065,N_11921);
or U20269 (N_20269,N_13640,N_18969);
or U20270 (N_20270,N_11433,N_19874);
xnor U20271 (N_20271,N_19584,N_13457);
and U20272 (N_20272,N_16830,N_18073);
nor U20273 (N_20273,N_13738,N_19231);
nor U20274 (N_20274,N_15509,N_14253);
nor U20275 (N_20275,N_19702,N_14416);
and U20276 (N_20276,N_15908,N_13365);
or U20277 (N_20277,N_16422,N_17492);
and U20278 (N_20278,N_17831,N_16436);
and U20279 (N_20279,N_16495,N_15376);
xnor U20280 (N_20280,N_13431,N_14609);
nor U20281 (N_20281,N_15592,N_15060);
xnor U20282 (N_20282,N_12675,N_11659);
nand U20283 (N_20283,N_17957,N_11398);
or U20284 (N_20284,N_13682,N_16735);
nor U20285 (N_20285,N_18914,N_19026);
or U20286 (N_20286,N_18971,N_17865);
nand U20287 (N_20287,N_17444,N_18395);
xnor U20288 (N_20288,N_10691,N_11509);
nor U20289 (N_20289,N_10484,N_16544);
nand U20290 (N_20290,N_12378,N_11016);
nor U20291 (N_20291,N_10593,N_17144);
nor U20292 (N_20292,N_18471,N_14627);
or U20293 (N_20293,N_18210,N_18667);
nor U20294 (N_20294,N_12612,N_18231);
nor U20295 (N_20295,N_12121,N_11932);
nand U20296 (N_20296,N_15821,N_11569);
or U20297 (N_20297,N_17268,N_11715);
or U20298 (N_20298,N_10832,N_14504);
and U20299 (N_20299,N_19905,N_17098);
nor U20300 (N_20300,N_16761,N_14435);
nor U20301 (N_20301,N_19615,N_11529);
nand U20302 (N_20302,N_10905,N_16390);
or U20303 (N_20303,N_16646,N_12694);
nor U20304 (N_20304,N_11346,N_13730);
nand U20305 (N_20305,N_11842,N_19021);
nand U20306 (N_20306,N_15163,N_10326);
nand U20307 (N_20307,N_17323,N_17889);
or U20308 (N_20308,N_11266,N_18739);
or U20309 (N_20309,N_10339,N_13992);
nand U20310 (N_20310,N_10247,N_17752);
or U20311 (N_20311,N_17857,N_14203);
or U20312 (N_20312,N_12017,N_11924);
or U20313 (N_20313,N_11655,N_17495);
nor U20314 (N_20314,N_14799,N_19391);
or U20315 (N_20315,N_12303,N_19828);
nor U20316 (N_20316,N_15915,N_14903);
and U20317 (N_20317,N_16487,N_19113);
xor U20318 (N_20318,N_15680,N_10244);
nand U20319 (N_20319,N_15785,N_17839);
and U20320 (N_20320,N_18263,N_17843);
nand U20321 (N_20321,N_16893,N_13474);
nor U20322 (N_20322,N_15714,N_18626);
nand U20323 (N_20323,N_12167,N_14846);
nand U20324 (N_20324,N_11961,N_13659);
or U20325 (N_20325,N_16190,N_10749);
and U20326 (N_20326,N_17798,N_19018);
and U20327 (N_20327,N_14156,N_13439);
and U20328 (N_20328,N_16380,N_17832);
or U20329 (N_20329,N_13740,N_19681);
or U20330 (N_20330,N_18993,N_16721);
or U20331 (N_20331,N_17238,N_11193);
and U20332 (N_20332,N_11009,N_18679);
nand U20333 (N_20333,N_15358,N_18600);
or U20334 (N_20334,N_15443,N_18120);
and U20335 (N_20335,N_17988,N_10322);
or U20336 (N_20336,N_18658,N_13966);
and U20337 (N_20337,N_12274,N_17313);
nor U20338 (N_20338,N_10562,N_15599);
or U20339 (N_20339,N_19028,N_15232);
nor U20340 (N_20340,N_11361,N_15523);
nor U20341 (N_20341,N_13518,N_13473);
nor U20342 (N_20342,N_11238,N_16180);
nor U20343 (N_20343,N_15547,N_19934);
xnor U20344 (N_20344,N_11828,N_18312);
or U20345 (N_20345,N_19951,N_16871);
nor U20346 (N_20346,N_14032,N_19765);
nand U20347 (N_20347,N_15216,N_15483);
xnor U20348 (N_20348,N_12699,N_11612);
xor U20349 (N_20349,N_17555,N_10223);
and U20350 (N_20350,N_11468,N_14282);
xor U20351 (N_20351,N_14433,N_14137);
or U20352 (N_20352,N_12350,N_12278);
nand U20353 (N_20353,N_19233,N_10697);
nand U20354 (N_20354,N_14101,N_15059);
nand U20355 (N_20355,N_11151,N_13753);
and U20356 (N_20356,N_17505,N_15591);
and U20357 (N_20357,N_13806,N_15243);
nand U20358 (N_20358,N_18531,N_17081);
and U20359 (N_20359,N_14570,N_15919);
nor U20360 (N_20360,N_14182,N_19454);
nand U20361 (N_20361,N_14498,N_14299);
nor U20362 (N_20362,N_15035,N_10509);
and U20363 (N_20363,N_17931,N_16579);
nor U20364 (N_20364,N_10871,N_11362);
or U20365 (N_20365,N_18162,N_12990);
xnor U20366 (N_20366,N_12637,N_12922);
nor U20367 (N_20367,N_13328,N_10452);
nor U20368 (N_20368,N_19413,N_14662);
and U20369 (N_20369,N_14904,N_19710);
and U20370 (N_20370,N_10363,N_10541);
and U20371 (N_20371,N_13875,N_15311);
xor U20372 (N_20372,N_19469,N_15089);
nor U20373 (N_20373,N_10410,N_11641);
or U20374 (N_20374,N_13481,N_11185);
nor U20375 (N_20375,N_14956,N_18122);
and U20376 (N_20376,N_15976,N_13396);
nand U20377 (N_20377,N_16873,N_19292);
nand U20378 (N_20378,N_11040,N_15234);
xor U20379 (N_20379,N_18519,N_14177);
or U20380 (N_20380,N_13463,N_10721);
and U20381 (N_20381,N_11753,N_17439);
xnor U20382 (N_20382,N_17086,N_15985);
nor U20383 (N_20383,N_11537,N_17868);
nand U20384 (N_20384,N_15172,N_12145);
and U20385 (N_20385,N_16398,N_15422);
nand U20386 (N_20386,N_13025,N_19794);
and U20387 (N_20387,N_12024,N_19479);
nor U20388 (N_20388,N_19131,N_18408);
or U20389 (N_20389,N_18748,N_17958);
xor U20390 (N_20390,N_12380,N_19495);
nor U20391 (N_20391,N_15389,N_19077);
nor U20392 (N_20392,N_14034,N_16438);
nand U20393 (N_20393,N_12205,N_17816);
and U20394 (N_20394,N_13342,N_10331);
nand U20395 (N_20395,N_15677,N_17502);
and U20396 (N_20396,N_11756,N_10450);
or U20397 (N_20397,N_17992,N_18413);
and U20398 (N_20398,N_13215,N_15409);
nor U20399 (N_20399,N_16527,N_16633);
and U20400 (N_20400,N_15270,N_12797);
nor U20401 (N_20401,N_18238,N_17415);
and U20402 (N_20402,N_13599,N_11697);
or U20403 (N_20403,N_10799,N_13357);
or U20404 (N_20404,N_19369,N_18381);
nor U20405 (N_20405,N_15220,N_11243);
nand U20406 (N_20406,N_14952,N_15966);
nand U20407 (N_20407,N_18956,N_19896);
nor U20408 (N_20408,N_17440,N_19280);
or U20409 (N_20409,N_16514,N_10311);
or U20410 (N_20410,N_10757,N_10826);
and U20411 (N_20411,N_11438,N_18943);
nor U20412 (N_20412,N_17610,N_12561);
and U20413 (N_20413,N_14171,N_14775);
nor U20414 (N_20414,N_10689,N_14136);
or U20415 (N_20415,N_18208,N_15972);
and U20416 (N_20416,N_14499,N_10332);
xnor U20417 (N_20417,N_12442,N_16130);
or U20418 (N_20418,N_18164,N_10011);
and U20419 (N_20419,N_10973,N_10519);
nor U20420 (N_20420,N_11599,N_10910);
and U20421 (N_20421,N_19006,N_16757);
nand U20422 (N_20422,N_15087,N_13796);
and U20423 (N_20423,N_14976,N_19782);
nor U20424 (N_20424,N_15152,N_10118);
or U20425 (N_20425,N_13406,N_16294);
and U20426 (N_20426,N_18712,N_19846);
xor U20427 (N_20427,N_15296,N_14094);
xor U20428 (N_20428,N_11223,N_15536);
nand U20429 (N_20429,N_14902,N_15125);
and U20430 (N_20430,N_15153,N_14660);
xor U20431 (N_20431,N_16206,N_12671);
or U20432 (N_20432,N_17344,N_11547);
or U20433 (N_20433,N_12987,N_10304);
nor U20434 (N_20434,N_11839,N_19692);
and U20435 (N_20435,N_15989,N_11304);
and U20436 (N_20436,N_11399,N_12624);
nor U20437 (N_20437,N_13133,N_11847);
nor U20438 (N_20438,N_13324,N_15625);
nand U20439 (N_20439,N_16522,N_16441);
and U20440 (N_20440,N_11460,N_13573);
nor U20441 (N_20441,N_18639,N_17421);
and U20442 (N_20442,N_16827,N_19024);
or U20443 (N_20443,N_19174,N_17680);
nand U20444 (N_20444,N_19823,N_10945);
xor U20445 (N_20445,N_15388,N_17221);
or U20446 (N_20446,N_18990,N_12367);
or U20447 (N_20447,N_14894,N_19715);
xor U20448 (N_20448,N_17892,N_17878);
nand U20449 (N_20449,N_19988,N_16755);
nand U20450 (N_20450,N_10791,N_19850);
nor U20451 (N_20451,N_19510,N_12366);
nor U20452 (N_20452,N_13921,N_15191);
or U20453 (N_20453,N_18004,N_12035);
xor U20454 (N_20454,N_19554,N_19003);
or U20455 (N_20455,N_18646,N_18254);
and U20456 (N_20456,N_13092,N_12373);
and U20457 (N_20457,N_12985,N_17382);
and U20458 (N_20458,N_12947,N_11130);
nand U20459 (N_20459,N_11786,N_11585);
and U20460 (N_20460,N_15894,N_17647);
and U20461 (N_20461,N_11218,N_14989);
and U20462 (N_20462,N_14138,N_18759);
nor U20463 (N_20463,N_18479,N_11504);
nand U20464 (N_20464,N_16279,N_10785);
or U20465 (N_20465,N_13433,N_18979);
nand U20466 (N_20466,N_19880,N_14934);
nand U20467 (N_20467,N_10242,N_17859);
or U20468 (N_20468,N_13908,N_13302);
and U20469 (N_20469,N_17899,N_18451);
or U20470 (N_20470,N_10211,N_11295);
xor U20471 (N_20471,N_13656,N_19862);
and U20472 (N_20472,N_14718,N_19103);
or U20473 (N_20473,N_16036,N_19116);
or U20474 (N_20474,N_13507,N_17360);
nand U20475 (N_20475,N_13340,N_12438);
nor U20476 (N_20476,N_19055,N_15902);
and U20477 (N_20477,N_16821,N_10426);
nand U20478 (N_20478,N_13166,N_14595);
nand U20479 (N_20479,N_19505,N_12164);
and U20480 (N_20480,N_11213,N_16235);
and U20481 (N_20481,N_16085,N_13974);
and U20482 (N_20482,N_12891,N_18830);
or U20483 (N_20483,N_19169,N_15936);
or U20484 (N_20484,N_17120,N_11094);
and U20485 (N_20485,N_18930,N_15954);
nor U20486 (N_20486,N_19478,N_18834);
nor U20487 (N_20487,N_11256,N_19923);
nand U20488 (N_20488,N_17551,N_13551);
nand U20489 (N_20489,N_11224,N_18685);
nor U20490 (N_20490,N_13516,N_13030);
nor U20491 (N_20491,N_11336,N_15427);
nor U20492 (N_20492,N_15442,N_17575);
nand U20493 (N_20493,N_19795,N_16686);
nor U20494 (N_20494,N_17142,N_16629);
nand U20495 (N_20495,N_19561,N_11886);
and U20496 (N_20496,N_18610,N_19797);
nor U20497 (N_20497,N_18787,N_13690);
nor U20498 (N_20498,N_13745,N_12707);
nand U20499 (N_20499,N_12253,N_10779);
or U20500 (N_20500,N_10843,N_14057);
xor U20501 (N_20501,N_19098,N_11302);
nor U20502 (N_20502,N_18329,N_14303);
and U20503 (N_20503,N_10901,N_15380);
nor U20504 (N_20504,N_18846,N_18326);
nor U20505 (N_20505,N_18575,N_15091);
nor U20506 (N_20506,N_12547,N_18555);
and U20507 (N_20507,N_19225,N_12654);
nand U20508 (N_20508,N_19501,N_18618);
nor U20509 (N_20509,N_11505,N_16979);
or U20510 (N_20510,N_16040,N_11624);
and U20511 (N_20511,N_19684,N_16254);
nand U20512 (N_20512,N_16502,N_17376);
or U20513 (N_20513,N_12578,N_12506);
and U20514 (N_20514,N_15678,N_18154);
nor U20515 (N_20515,N_16428,N_15653);
nand U20516 (N_20516,N_13865,N_12822);
or U20517 (N_20517,N_16537,N_19407);
and U20518 (N_20518,N_14569,N_14251);
and U20519 (N_20519,N_14368,N_13073);
and U20520 (N_20520,N_13203,N_15255);
nand U20521 (N_20521,N_19064,N_12485);
nor U20522 (N_20522,N_17228,N_10627);
and U20523 (N_20523,N_11306,N_13938);
nor U20524 (N_20524,N_14466,N_17371);
xor U20525 (N_20525,N_19583,N_18242);
or U20526 (N_20526,N_16474,N_15532);
nand U20527 (N_20527,N_12571,N_15150);
and U20528 (N_20528,N_10525,N_15779);
nor U20529 (N_20529,N_16252,N_14002);
or U20530 (N_20530,N_14021,N_19654);
nand U20531 (N_20531,N_12469,N_17491);
xor U20532 (N_20532,N_17493,N_11863);
nor U20533 (N_20533,N_17701,N_15394);
nand U20534 (N_20534,N_11826,N_15688);
nor U20535 (N_20535,N_15297,N_18197);
and U20536 (N_20536,N_13240,N_14677);
and U20537 (N_20537,N_12499,N_13425);
and U20538 (N_20538,N_12522,N_17280);
and U20539 (N_20539,N_16851,N_19634);
nor U20540 (N_20540,N_14736,N_11542);
nor U20541 (N_20541,N_19200,N_13822);
nand U20542 (N_20542,N_13951,N_10885);
and U20543 (N_20543,N_14684,N_11783);
xor U20544 (N_20544,N_16102,N_18549);
and U20545 (N_20545,N_16219,N_10310);
or U20546 (N_20546,N_12116,N_18923);
xor U20547 (N_20547,N_13842,N_11972);
nand U20548 (N_20548,N_12878,N_12780);
nand U20549 (N_20549,N_12096,N_11170);
nor U20550 (N_20550,N_16981,N_14316);
nor U20551 (N_20551,N_19740,N_17874);
and U20552 (N_20552,N_13597,N_18654);
nor U20553 (N_20553,N_14095,N_10275);
and U20554 (N_20554,N_13187,N_16641);
nand U20555 (N_20555,N_19484,N_10208);
or U20556 (N_20556,N_12073,N_19697);
nor U20557 (N_20557,N_10154,N_15921);
nand U20558 (N_20558,N_11119,N_14749);
nor U20559 (N_20559,N_14475,N_19417);
and U20560 (N_20560,N_19631,N_17699);
nor U20561 (N_20561,N_12196,N_11609);
or U20562 (N_20562,N_18789,N_14078);
and U20563 (N_20563,N_10878,N_14839);
nor U20564 (N_20564,N_14065,N_12130);
nor U20565 (N_20565,N_17237,N_11291);
or U20566 (N_20566,N_11848,N_18563);
nor U20567 (N_20567,N_12042,N_10674);
nor U20568 (N_20568,N_10730,N_13150);
or U20569 (N_20569,N_19640,N_10391);
and U20570 (N_20570,N_18012,N_17597);
and U20571 (N_20571,N_11669,N_18294);
or U20572 (N_20572,N_16658,N_12106);
or U20573 (N_20573,N_12598,N_19053);
nand U20574 (N_20574,N_12263,N_11206);
or U20575 (N_20575,N_13074,N_18412);
nand U20576 (N_20576,N_17627,N_11423);
nand U20577 (N_20577,N_19258,N_18699);
nor U20578 (N_20578,N_17266,N_17819);
and U20579 (N_20579,N_14510,N_13591);
or U20580 (N_20580,N_17457,N_18637);
and U20581 (N_20581,N_13692,N_18015);
or U20582 (N_20582,N_13627,N_10728);
and U20583 (N_20583,N_12076,N_12958);
nor U20584 (N_20584,N_15612,N_18420);
or U20585 (N_20585,N_19661,N_16468);
nor U20586 (N_20586,N_16430,N_19952);
or U20587 (N_20587,N_10263,N_14217);
xnor U20588 (N_20588,N_19800,N_12348);
or U20589 (N_20589,N_15643,N_11048);
or U20590 (N_20590,N_13561,N_17920);
nand U20591 (N_20591,N_12553,N_17729);
nor U20592 (N_20592,N_16179,N_10070);
xnor U20593 (N_20593,N_18648,N_11946);
or U20594 (N_20594,N_10897,N_13722);
nand U20595 (N_20595,N_18110,N_13050);
and U20596 (N_20596,N_19381,N_17749);
xnor U20597 (N_20597,N_17038,N_13455);
nor U20598 (N_20598,N_15912,N_15828);
nor U20599 (N_20599,N_15048,N_16443);
and U20600 (N_20600,N_18710,N_12784);
or U20601 (N_20601,N_11247,N_17675);
nand U20602 (N_20602,N_19776,N_10844);
nand U20603 (N_20603,N_17141,N_18880);
nor U20604 (N_20604,N_16240,N_16156);
and U20605 (N_20605,N_19214,N_19749);
nand U20606 (N_20606,N_17014,N_14222);
or U20607 (N_20607,N_18153,N_15982);
nand U20608 (N_20608,N_19086,N_10863);
xor U20609 (N_20609,N_17506,N_18386);
and U20610 (N_20610,N_11722,N_10836);
nor U20611 (N_20611,N_11616,N_15626);
or U20612 (N_20612,N_19582,N_17035);
and U20613 (N_20613,N_15400,N_11269);
nand U20614 (N_20614,N_12037,N_12976);
or U20615 (N_20615,N_18344,N_17006);
nand U20616 (N_20616,N_16622,N_10958);
nand U20617 (N_20617,N_16866,N_13693);
and U20618 (N_20618,N_13075,N_15318);
nand U20619 (N_20619,N_12734,N_11014);
or U20620 (N_20620,N_15105,N_11493);
xor U20621 (N_20621,N_17020,N_14859);
xnor U20622 (N_20622,N_13351,N_11914);
and U20623 (N_20623,N_12596,N_18862);
nand U20624 (N_20624,N_16116,N_13643);
nor U20625 (N_20625,N_14104,N_13675);
xor U20626 (N_20626,N_12203,N_13033);
xor U20627 (N_20627,N_19992,N_18349);
xor U20628 (N_20628,N_16212,N_14772);
nand U20629 (N_20629,N_12112,N_14195);
and U20630 (N_20630,N_11766,N_17201);
nor U20631 (N_20631,N_15069,N_19339);
nor U20632 (N_20632,N_16613,N_16748);
nand U20633 (N_20633,N_18097,N_18053);
nor U20634 (N_20634,N_13809,N_18803);
nor U20635 (N_20635,N_16108,N_13715);
xnor U20636 (N_20636,N_14531,N_14071);
xor U20637 (N_20637,N_11353,N_17594);
nand U20638 (N_20638,N_19743,N_15334);
nor U20639 (N_20639,N_16005,N_16504);
or U20640 (N_20640,N_17147,N_17246);
and U20641 (N_20641,N_17656,N_13850);
nand U20642 (N_20642,N_14686,N_10169);
nand U20643 (N_20643,N_19436,N_11076);
nand U20644 (N_20644,N_16855,N_15149);
nor U20645 (N_20645,N_15371,N_11706);
nand U20646 (N_20646,N_16885,N_11096);
nand U20647 (N_20647,N_10134,N_16455);
and U20648 (N_20648,N_14553,N_10328);
and U20649 (N_20649,N_12028,N_14698);
nor U20650 (N_20650,N_10764,N_19277);
nor U20651 (N_20651,N_14981,N_16126);
or U20652 (N_20652,N_19074,N_16216);
or U20653 (N_20653,N_15629,N_17291);
and U20654 (N_20654,N_19842,N_15865);
nand U20655 (N_20655,N_19298,N_19178);
or U20656 (N_20656,N_13636,N_10022);
nand U20657 (N_20657,N_18098,N_12406);
and U20658 (N_20658,N_18027,N_19409);
and U20659 (N_20659,N_11241,N_14511);
or U20660 (N_20660,N_14367,N_19164);
or U20661 (N_20661,N_17530,N_11662);
or U20662 (N_20662,N_11037,N_15205);
nor U20663 (N_20663,N_14876,N_12245);
or U20664 (N_20664,N_18615,N_18130);
or U20665 (N_20665,N_17230,N_10895);
or U20666 (N_20666,N_14765,N_19679);
nor U20667 (N_20667,N_17937,N_11384);
or U20668 (N_20668,N_11250,N_18425);
or U20669 (N_20669,N_16702,N_18520);
or U20670 (N_20670,N_15928,N_12243);
or U20671 (N_20671,N_14849,N_14250);
nand U20672 (N_20672,N_10608,N_11114);
or U20673 (N_20673,N_14116,N_19071);
or U20674 (N_20674,N_11221,N_15602);
xnor U20675 (N_20675,N_15433,N_17375);
nor U20676 (N_20676,N_14109,N_13012);
nand U20677 (N_20677,N_11294,N_13385);
and U20678 (N_20678,N_12315,N_17207);
and U20679 (N_20679,N_17838,N_14349);
xor U20680 (N_20680,N_19361,N_16954);
or U20681 (N_20681,N_18826,N_16573);
xor U20682 (N_20682,N_13929,N_12925);
and U20683 (N_20683,N_12462,N_18019);
and U20684 (N_20684,N_19774,N_19332);
or U20685 (N_20685,N_11118,N_19274);
nand U20686 (N_20686,N_17726,N_13949);
nand U20687 (N_20687,N_16987,N_17092);
xor U20688 (N_20688,N_14172,N_10780);
nand U20689 (N_20689,N_13758,N_17409);
or U20690 (N_20690,N_13782,N_15691);
or U20691 (N_20691,N_17471,N_11582);
nor U20692 (N_20692,N_16192,N_15188);
and U20693 (N_20693,N_12321,N_19751);
nor U20694 (N_20694,N_13155,N_18280);
or U20695 (N_20695,N_17110,N_19004);
nor U20696 (N_20696,N_13789,N_14522);
nand U20697 (N_20697,N_15052,N_14245);
nand U20698 (N_20698,N_13147,N_12431);
and U20699 (N_20699,N_17054,N_11920);
and U20700 (N_20700,N_17807,N_19856);
or U20701 (N_20701,N_10616,N_14080);
xor U20702 (N_20702,N_15115,N_18182);
and U20703 (N_20703,N_15475,N_13568);
nor U20704 (N_20704,N_16724,N_18772);
nor U20705 (N_20705,N_16006,N_10368);
nor U20706 (N_20706,N_18644,N_11112);
and U20707 (N_20707,N_19238,N_18652);
xnor U20708 (N_20708,N_12693,N_12663);
or U20709 (N_20709,N_14830,N_11373);
nor U20710 (N_20710,N_12144,N_10993);
nor U20711 (N_20711,N_18786,N_14715);
and U20712 (N_20712,N_17985,N_13254);
and U20713 (N_20713,N_19353,N_19607);
nor U20714 (N_20714,N_13243,N_17888);
nand U20715 (N_20715,N_13023,N_10944);
xor U20716 (N_20716,N_18999,N_17212);
nand U20717 (N_20717,N_14622,N_17648);
xnor U20718 (N_20718,N_12836,N_19947);
xnor U20719 (N_20719,N_19269,N_11386);
xor U20720 (N_20720,N_18394,N_12910);
and U20721 (N_20721,N_12322,N_15473);
and U20722 (N_20722,N_16203,N_14629);
nor U20723 (N_20723,N_14372,N_16541);
xor U20724 (N_20724,N_19333,N_19008);
nor U20725 (N_20725,N_13664,N_11252);
or U20726 (N_20726,N_16245,N_13922);
nand U20727 (N_20727,N_18915,N_10272);
nor U20728 (N_20728,N_19580,N_10865);
nand U20729 (N_20729,N_12212,N_16841);
or U20730 (N_20730,N_18548,N_12559);
xor U20731 (N_20731,N_10731,N_12446);
xor U20732 (N_20732,N_19895,N_13091);
nand U20733 (N_20733,N_11885,N_10716);
or U20734 (N_20734,N_18823,N_16077);
or U20735 (N_20735,N_13773,N_14755);
nor U20736 (N_20736,N_18360,N_14798);
or U20737 (N_20737,N_18428,N_10146);
nor U20738 (N_20738,N_18779,N_19496);
xnor U20739 (N_20739,N_18002,N_18270);
or U20740 (N_20740,N_14312,N_15618);
or U20741 (N_20741,N_13234,N_11635);
or U20742 (N_20742,N_19165,N_16624);
and U20743 (N_20743,N_11690,N_15851);
nand U20744 (N_20744,N_16229,N_14923);
and U20745 (N_20745,N_10995,N_10039);
or U20746 (N_20746,N_13737,N_18886);
and U20747 (N_20747,N_10641,N_18296);
or U20748 (N_20748,N_11643,N_13958);
nor U20749 (N_20749,N_13081,N_10383);
or U20750 (N_20750,N_18187,N_19875);
nand U20751 (N_20751,N_18233,N_19699);
nor U20752 (N_20752,N_18775,N_13142);
and U20753 (N_20753,N_10053,N_14929);
nand U20754 (N_20754,N_13168,N_14383);
or U20755 (N_20755,N_15506,N_19643);
xnor U20756 (N_20756,N_17902,N_13470);
nor U20757 (N_20757,N_12921,N_19275);
or U20758 (N_20758,N_19698,N_13350);
nor U20759 (N_20759,N_11626,N_19806);
and U20760 (N_20760,N_17342,N_15806);
nor U20761 (N_20761,N_19123,N_17252);
and U20762 (N_20762,N_15666,N_11101);
nor U20763 (N_20763,N_13604,N_18628);
nor U20764 (N_20764,N_16388,N_16358);
nand U20765 (N_20765,N_16661,N_14229);
and U20766 (N_20766,N_14474,N_18267);
and U20767 (N_20767,N_18609,N_17624);
and U20768 (N_20768,N_16022,N_10815);
xor U20769 (N_20769,N_19486,N_13366);
nor U20770 (N_20770,N_16151,N_14262);
nor U20771 (N_20771,N_14932,N_10270);
or U20772 (N_20772,N_19093,N_18978);
nand U20773 (N_20773,N_10231,N_16632);
or U20774 (N_20774,N_10589,N_13873);
and U20775 (N_20775,N_18704,N_10330);
nor U20776 (N_20776,N_12169,N_16307);
and U20777 (N_20777,N_12646,N_15310);
xor U20778 (N_20778,N_12819,N_11772);
nor U20779 (N_20779,N_19490,N_12656);
or U20780 (N_20780,N_19205,N_11610);
or U20781 (N_20781,N_13630,N_14259);
nand U20782 (N_20782,N_18048,N_10927);
nor U20783 (N_20783,N_19642,N_11150);
nor U20784 (N_20784,N_16033,N_16169);
xnor U20785 (N_20785,N_13697,N_13432);
or U20786 (N_20786,N_19343,N_10833);
and U20787 (N_20787,N_13707,N_13274);
and U20788 (N_20788,N_12066,N_18962);
nor U20789 (N_20789,N_15221,N_18215);
nor U20790 (N_20790,N_10667,N_11498);
nor U20791 (N_20791,N_11472,N_12510);
or U20792 (N_20792,N_18334,N_18422);
xnor U20793 (N_20793,N_14051,N_12440);
nand U20794 (N_20794,N_15019,N_18916);
nand U20795 (N_20795,N_12495,N_19248);
nand U20796 (N_20796,N_17599,N_15178);
xor U20797 (N_20797,N_13802,N_17396);
or U20798 (N_20798,N_10031,N_16493);
xor U20799 (N_20799,N_11802,N_14789);
and U20800 (N_20800,N_17223,N_10846);
and U20801 (N_20801,N_18393,N_11069);
nand U20802 (N_20802,N_11377,N_18084);
or U20803 (N_20803,N_14361,N_10737);
and U20804 (N_20804,N_11058,N_19588);
or U20805 (N_20805,N_16349,N_12156);
nor U20806 (N_20806,N_16110,N_12209);
and U20807 (N_20807,N_10422,N_11244);
and U20808 (N_20808,N_10659,N_10578);
or U20809 (N_20809,N_13249,N_11777);
or U20810 (N_20810,N_11807,N_12779);
nor U20811 (N_20811,N_11275,N_13371);
nor U20812 (N_20812,N_13401,N_11771);
and U20813 (N_20813,N_12404,N_16014);
nand U20814 (N_20814,N_11755,N_12614);
or U20815 (N_20815,N_12483,N_19270);
and U20816 (N_20816,N_11054,N_18833);
and U20817 (N_20817,N_16129,N_12515);
or U20818 (N_20818,N_13870,N_16481);
nand U20819 (N_20819,N_16674,N_13962);
nor U20820 (N_20820,N_18401,N_17393);
nand U20821 (N_20821,N_11287,N_12724);
nand U20822 (N_20822,N_16669,N_16182);
nor U20823 (N_20823,N_12874,N_18807);
xnor U20824 (N_20824,N_18668,N_14564);
nor U20825 (N_20825,N_19730,N_15468);
and U20826 (N_20826,N_18336,N_19889);
or U20827 (N_20827,N_17745,N_17335);
nand U20828 (N_20828,N_16863,N_16220);
or U20829 (N_20829,N_15457,N_12132);
nor U20830 (N_20830,N_19175,N_16261);
nand U20831 (N_20831,N_16193,N_17776);
or U20832 (N_20832,N_14842,N_10681);
nor U20833 (N_20833,N_18426,N_14050);
or U20834 (N_20834,N_11323,N_14933);
and U20835 (N_20835,N_17193,N_18031);
nand U20836 (N_20836,N_18176,N_11057);
and U20837 (N_20837,N_18416,N_17580);
nand U20838 (N_20838,N_16907,N_18695);
nor U20839 (N_20839,N_18740,N_10959);
nor U20840 (N_20840,N_16393,N_14461);
nand U20841 (N_20841,N_11432,N_19991);
xnor U20842 (N_20842,N_13876,N_16275);
or U20843 (N_20843,N_13232,N_19954);
nand U20844 (N_20844,N_18883,N_18529);
or U20845 (N_20845,N_10497,N_10511);
xnor U20846 (N_20846,N_11111,N_19393);
nor U20847 (N_20847,N_17463,N_17614);
and U20848 (N_20848,N_17596,N_11031);
nor U20849 (N_20849,N_11829,N_18891);
or U20850 (N_20850,N_18897,N_14272);
and U20851 (N_20851,N_10943,N_16988);
nand U20852 (N_20852,N_19220,N_19463);
nor U20853 (N_20853,N_13192,N_14768);
nand U20854 (N_20854,N_14405,N_13140);
nand U20855 (N_20855,N_17778,N_17204);
nand U20856 (N_20856,N_19927,N_15568);
and U20857 (N_20857,N_11598,N_17671);
nor U20858 (N_20858,N_13887,N_10013);
and U20859 (N_20859,N_13886,N_15968);
nand U20860 (N_20860,N_13637,N_11831);
and U20861 (N_20861,N_16214,N_11564);
and U20862 (N_20862,N_17245,N_10522);
xnor U20863 (N_20863,N_17584,N_15210);
xnor U20864 (N_20864,N_12392,N_16743);
and U20865 (N_20865,N_10707,N_19466);
nor U20866 (N_20866,N_19734,N_14154);
nand U20867 (N_20867,N_10150,N_18169);
or U20868 (N_20868,N_19753,N_11571);
nor U20869 (N_20869,N_18665,N_12828);
or U20870 (N_20870,N_11919,N_19548);
nand U20871 (N_20871,N_10257,N_16845);
and U20872 (N_20872,N_11452,N_19898);
nand U20873 (N_20873,N_19676,N_13087);
nor U20874 (N_20874,N_15049,N_16816);
or U20875 (N_20875,N_13687,N_16131);
nor U20876 (N_20876,N_14126,N_14013);
and U20877 (N_20877,N_12010,N_11698);
nand U20878 (N_20878,N_16259,N_15783);
nor U20879 (N_20879,N_16232,N_19294);
nand U20880 (N_20880,N_19614,N_15351);
nor U20881 (N_20881,N_16857,N_14503);
or U20882 (N_20882,N_17723,N_18278);
or U20883 (N_20883,N_10406,N_10772);
and U20884 (N_20884,N_15883,N_13237);
or U20885 (N_20885,N_11862,N_16891);
and U20886 (N_20886,N_17912,N_19902);
nand U20887 (N_20887,N_10137,N_18678);
and U20888 (N_20888,N_16876,N_12339);
xor U20889 (N_20889,N_19957,N_16730);
nand U20890 (N_20890,N_14139,N_17983);
nand U20891 (N_20891,N_10520,N_12879);
xor U20892 (N_20892,N_16810,N_15440);
or U20893 (N_20893,N_11264,N_10732);
or U20894 (N_20894,N_12812,N_10360);
or U20895 (N_20895,N_10558,N_14997);
nand U20896 (N_20896,N_11464,N_12213);
nor U20897 (N_20897,N_15793,N_15903);
nand U20898 (N_20898,N_19450,N_12397);
nor U20899 (N_20899,N_15926,N_12413);
and U20900 (N_20900,N_15993,N_12091);
nand U20901 (N_20901,N_19935,N_13725);
and U20902 (N_20902,N_12340,N_12621);
nor U20903 (N_20903,N_18017,N_19360);
nor U20904 (N_20904,N_16074,N_13225);
or U20905 (N_20905,N_19335,N_16303);
and U20906 (N_20906,N_19959,N_14541);
nand U20907 (N_20907,N_15379,N_17975);
xor U20908 (N_20908,N_14751,N_19092);
or U20909 (N_20909,N_14679,N_14398);
xor U20910 (N_20910,N_14114,N_16196);
nor U20911 (N_20911,N_16607,N_16070);
nand U20912 (N_20912,N_15197,N_12070);
nand U20913 (N_20913,N_10059,N_19660);
nand U20914 (N_20914,N_10167,N_15539);
and U20915 (N_20915,N_15560,N_16831);
nor U20916 (N_20916,N_13767,N_14888);
or U20917 (N_20917,N_16357,N_14221);
nand U20918 (N_20918,N_16288,N_13419);
and U20919 (N_20919,N_11149,N_15664);
or U20920 (N_20920,N_17626,N_17553);
nand U20921 (N_20921,N_19517,N_19869);
and U20922 (N_20922,N_13984,N_13784);
nand U20923 (N_20923,N_14706,N_12814);
and U20924 (N_20924,N_15730,N_11844);
or U20925 (N_20925,N_10386,N_10194);
and U20926 (N_20926,N_18421,N_16985);
or U20927 (N_20927,N_16939,N_13739);
nand U20928 (N_20928,N_10548,N_14790);
nor U20929 (N_20929,N_19170,N_15474);
or U20930 (N_20930,N_14388,N_14852);
nand U20931 (N_20931,N_19859,N_18062);
or U20932 (N_20932,N_19788,N_18964);
nor U20933 (N_20933,N_12398,N_17666);
nand U20934 (N_20934,N_10030,N_15193);
and U20935 (N_20935,N_10488,N_10228);
and U20936 (N_20936,N_19706,N_18599);
and U20937 (N_20937,N_16731,N_19576);
or U20938 (N_20938,N_12750,N_19313);
nand U20939 (N_20939,N_19097,N_16342);
and U20940 (N_20940,N_19714,N_19054);
nor U20941 (N_20941,N_15805,N_13161);
or U20942 (N_20942,N_15731,N_17478);
nor U20943 (N_20943,N_11935,N_17128);
nand U20944 (N_20944,N_19644,N_11858);
nand U20945 (N_20945,N_17698,N_12018);
nand U20946 (N_20946,N_18323,N_18243);
xor U20947 (N_20947,N_16548,N_14769);
nand U20948 (N_20948,N_14302,N_15766);
nand U20949 (N_20949,N_17564,N_11915);
nor U20950 (N_20950,N_17140,N_19787);
nand U20951 (N_20951,N_11644,N_19439);
or U20952 (N_20952,N_12977,N_14682);
xor U20953 (N_20953,N_18980,N_11300);
nand U20954 (N_20954,N_15495,N_10574);
and U20955 (N_20955,N_10400,N_16711);
nor U20956 (N_20956,N_16773,N_16934);
xor U20957 (N_20957,N_10486,N_14039);
and U20958 (N_20958,N_12558,N_13003);
and U20959 (N_20959,N_19072,N_12030);
nor U20960 (N_20960,N_19506,N_10902);
nand U20961 (N_20961,N_16336,N_19172);
or U20962 (N_20962,N_15361,N_12419);
nand U20963 (N_20963,N_16431,N_11619);
and U20964 (N_20964,N_11317,N_18396);
nor U20965 (N_20965,N_19930,N_10500);
nand U20966 (N_20966,N_17910,N_18490);
nor U20967 (N_20967,N_19737,N_12927);
and U20968 (N_20968,N_10862,N_10572);
nand U20969 (N_20969,N_10784,N_17809);
and U20970 (N_20970,N_15317,N_15747);
or U20971 (N_20971,N_14552,N_12080);
and U20972 (N_20972,N_17678,N_11739);
and U20973 (N_20973,N_11074,N_16578);
or U20974 (N_20974,N_11534,N_15010);
xnor U20975 (N_20975,N_18281,N_19209);
xor U20976 (N_20976,N_14776,N_15716);
nor U20977 (N_20977,N_18076,N_18213);
or U20978 (N_20978,N_15660,N_15470);
nor U20979 (N_20979,N_11923,N_13552);
nand U20980 (N_20980,N_19516,N_18733);
nor U20981 (N_20981,N_17562,N_13384);
nand U20982 (N_20982,N_19574,N_12047);
nand U20983 (N_20983,N_13408,N_12247);
nor U20984 (N_20984,N_17504,N_12391);
and U20985 (N_20985,N_10227,N_15832);
nand U20986 (N_20986,N_10443,N_17996);
nand U20987 (N_20987,N_15444,N_13368);
xor U20988 (N_20988,N_18560,N_12335);
nor U20989 (N_20989,N_10639,N_15762);
xnor U20990 (N_20990,N_15505,N_16249);
nor U20991 (N_20991,N_17196,N_11992);
or U20992 (N_20992,N_15610,N_12870);
and U20993 (N_20993,N_15557,N_15007);
or U20994 (N_20994,N_17785,N_14604);
xor U20995 (N_20995,N_14184,N_10577);
nand U20996 (N_20996,N_14544,N_16318);
or U20997 (N_20997,N_13519,N_11790);
xnor U20998 (N_20998,N_17764,N_15627);
xnor U20999 (N_20999,N_13387,N_12847);
and U21000 (N_21000,N_17262,N_10098);
xor U21001 (N_21001,N_11793,N_18533);
or U21002 (N_21002,N_13567,N_14500);
nor U21003 (N_21003,N_19034,N_17064);
nand U21004 (N_21004,N_16786,N_14583);
or U21005 (N_21005,N_12933,N_19744);
and U21006 (N_21006,N_13099,N_12349);
or U21007 (N_21007,N_13301,N_15303);
or U21008 (N_21008,N_19187,N_14741);
xor U21009 (N_21009,N_19322,N_18601);
nor U21010 (N_21010,N_17467,N_11898);
nor U21011 (N_21011,N_13420,N_19591);
nor U21012 (N_21012,N_15620,N_10900);
or U21013 (N_21013,N_14120,N_15603);
nor U21014 (N_21014,N_11776,N_13210);
nor U21015 (N_21015,N_14473,N_14351);
or U21016 (N_21016,N_13620,N_16032);
nor U21017 (N_21017,N_11846,N_19911);
nor U21018 (N_21018,N_12688,N_16165);
xor U21019 (N_21019,N_10613,N_12930);
and U21020 (N_21020,N_19845,N_18907);
nand U21021 (N_21021,N_11896,N_18663);
nand U21022 (N_21022,N_12181,N_11539);
and U21023 (N_21023,N_13248,N_18850);
nor U21024 (N_21024,N_18295,N_15171);
and U21025 (N_21025,N_12562,N_14097);
nand U21026 (N_21026,N_11471,N_19635);
and U21027 (N_21027,N_19649,N_18237);
and U21028 (N_21028,N_14117,N_11229);
or U21029 (N_21029,N_15922,N_17032);
or U21030 (N_21030,N_11820,N_13322);
or U21031 (N_21031,N_18345,N_14183);
nand U21032 (N_21032,N_11785,N_14493);
nor U21033 (N_21033,N_19423,N_17327);
xor U21034 (N_21034,N_14680,N_14141);
nor U21035 (N_21035,N_12377,N_19603);
and U21036 (N_21036,N_12883,N_17926);
xnor U21037 (N_21037,N_13964,N_14360);
nand U21038 (N_21038,N_18587,N_17486);
or U21039 (N_21039,N_17454,N_18703);
nand U21040 (N_21040,N_16448,N_13791);
or U21041 (N_21041,N_18631,N_17929);
nand U21042 (N_21042,N_13089,N_11116);
nand U21043 (N_21043,N_16188,N_19863);
nand U21044 (N_21044,N_13488,N_10853);
nor U21045 (N_21045,N_16740,N_16992);
nor U21046 (N_21046,N_11435,N_18175);
nand U21047 (N_21047,N_14804,N_13136);
nor U21048 (N_21048,N_10556,N_18155);
and U21049 (N_21049,N_13927,N_15339);
and U21050 (N_21050,N_19514,N_15009);
and U21051 (N_21051,N_12617,N_10481);
and U21052 (N_21052,N_10966,N_13246);
and U21053 (N_21053,N_13471,N_16411);
xnor U21054 (N_21054,N_16997,N_16818);
xnor U21055 (N_21055,N_11871,N_11758);
and U21056 (N_21056,N_18424,N_15590);
nor U21057 (N_21057,N_16292,N_15487);
or U21058 (N_21058,N_12793,N_18315);
nand U21059 (N_21059,N_15588,N_10969);
nor U21060 (N_21060,N_10128,N_19609);
and U21061 (N_21061,N_15622,N_10575);
nor U21062 (N_21062,N_14853,N_13933);
nor U21063 (N_21063,N_14206,N_10366);
xor U21064 (N_21064,N_16713,N_10675);
or U21065 (N_21065,N_15173,N_17867);
and U21066 (N_21066,N_12678,N_10750);
nor U21067 (N_21067,N_11215,N_15476);
nand U21068 (N_21068,N_14938,N_14867);
nor U21069 (N_21069,N_15676,N_12368);
nand U21070 (N_21070,N_10290,N_18945);
or U21071 (N_21071,N_19234,N_18010);
or U21072 (N_21072,N_13913,N_14815);
nand U21073 (N_21073,N_13153,N_15914);
and U21074 (N_21074,N_12841,N_15253);
nor U21075 (N_21075,N_18114,N_18624);
and U21076 (N_21076,N_18013,N_11711);
or U21077 (N_21077,N_14691,N_12717);
or U21078 (N_21078,N_15413,N_19532);
nor U21079 (N_21079,N_17823,N_17652);
nand U21080 (N_21080,N_13005,N_17688);
nor U21081 (N_21081,N_18638,N_16574);
and U21082 (N_21082,N_18066,N_18366);
or U21083 (N_21083,N_16374,N_17307);
xnor U21084 (N_21084,N_17195,N_18664);
xnor U21085 (N_21085,N_19340,N_12632);
nor U21086 (N_21086,N_13179,N_13417);
and U21087 (N_21087,N_17273,N_18261);
and U21088 (N_21088,N_19325,N_10709);
or U21089 (N_21089,N_14502,N_16897);
or U21090 (N_21090,N_13629,N_18106);
xnor U21091 (N_21091,N_17116,N_18133);
xor U21092 (N_21092,N_17274,N_16140);
nor U21093 (N_21093,N_15101,N_17790);
and U21094 (N_21094,N_13045,N_19664);
nand U21095 (N_21095,N_12723,N_16345);
nand U21096 (N_21096,N_18047,N_18071);
or U21097 (N_21097,N_16918,N_10390);
xnor U21098 (N_21098,N_15417,N_12299);
or U21099 (N_21099,N_19161,N_18904);
or U21100 (N_21100,N_11176,N_17623);
nor U21101 (N_21101,N_10698,N_10714);
xnor U21102 (N_21102,N_12086,N_18046);
nand U21103 (N_21103,N_11773,N_19265);
or U21104 (N_21104,N_13495,N_18571);
nand U21105 (N_21105,N_13982,N_10605);
nor U21106 (N_21106,N_19160,N_11175);
nor U21107 (N_21107,N_11271,N_14356);
and U21108 (N_21108,N_18797,N_10083);
nand U21109 (N_21109,N_10158,N_16847);
xnor U21110 (N_21110,N_10984,N_18918);
nor U21111 (N_21111,N_14914,N_15942);
nor U21112 (N_21112,N_13327,N_18279);
nand U21113 (N_21113,N_10057,N_11454);
or U21114 (N_21114,N_15594,N_19403);
and U21115 (N_21115,N_18677,N_12698);
nand U21116 (N_21116,N_18841,N_18785);
and U21117 (N_21117,N_11933,N_16485);
and U21118 (N_21118,N_19946,N_15694);
nand U21119 (N_21119,N_10014,N_18584);
or U21120 (N_21120,N_19901,N_15668);
and U21121 (N_21121,N_17722,N_11943);
nand U21122 (N_21122,N_17956,N_12897);
and U21123 (N_21123,N_14160,N_10705);
nor U21124 (N_21124,N_16332,N_13548);
and U21125 (N_21125,N_15266,N_19262);
nand U21126 (N_21126,N_10524,N_15661);
nor U21127 (N_21127,N_17963,N_19724);
nor U21128 (N_21128,N_10594,N_13496);
nor U21129 (N_21129,N_13297,N_15596);
or U21130 (N_21130,N_10388,N_15924);
and U21131 (N_21131,N_10094,N_18287);
nor U21132 (N_21132,N_14634,N_13522);
nor U21133 (N_21133,N_19962,N_10179);
and U21134 (N_21134,N_18613,N_10961);
or U21135 (N_21135,N_16048,N_13691);
nand U21136 (N_21136,N_17036,N_11387);
xor U21137 (N_21137,N_18864,N_12740);
or U21138 (N_21138,N_13478,N_11005);
or U21139 (N_21139,N_14656,N_16347);
and U21140 (N_21140,N_15856,N_14827);
or U21141 (N_21141,N_12638,N_18588);
and U21142 (N_21142,N_14053,N_11476);
nor U21143 (N_21143,N_15994,N_15228);
and U21144 (N_21144,N_16244,N_19352);
or U21145 (N_21145,N_17287,N_18388);
and U21146 (N_21146,N_14857,N_18756);
and U21147 (N_21147,N_15669,N_13611);
or U21148 (N_21148,N_11897,N_11330);
nand U21149 (N_21149,N_13930,N_18216);
or U21150 (N_21150,N_19143,N_18258);
nand U21151 (N_21151,N_15961,N_13831);
or U21152 (N_21152,N_15356,N_10021);
nor U21153 (N_21153,N_10302,N_10604);
nand U21154 (N_21154,N_17320,N_13154);
nor U21155 (N_21155,N_14515,N_19014);
nor U21156 (N_21156,N_14885,N_18723);
nand U21157 (N_21157,N_18328,N_16057);
and U21158 (N_21158,N_12546,N_13523);
nand U21159 (N_21159,N_18750,N_19933);
xnor U21160 (N_21160,N_19671,N_19694);
or U21161 (N_21161,N_11225,N_12785);
nor U21162 (N_21162,N_17639,N_11449);
nor U21163 (N_21163,N_18693,N_10023);
or U21164 (N_21164,N_10956,N_10027);
nor U21165 (N_21165,N_10886,N_17413);
and U21166 (N_21166,N_16931,N_12955);
or U21167 (N_21167,N_17687,N_14364);
nor U21168 (N_21168,N_18673,N_12593);
and U21169 (N_21169,N_18933,N_11519);
or U21170 (N_21170,N_14640,N_16146);
nor U21171 (N_21171,N_15980,N_15373);
or U21172 (N_21172,N_12043,N_14348);
or U21173 (N_21173,N_15312,N_11157);
nor U21174 (N_21174,N_12719,N_13652);
or U21175 (N_21175,N_16484,N_12468);
or U21176 (N_21176,N_17255,N_11052);
and U21177 (N_21177,N_18573,N_17741);
nor U21178 (N_21178,N_14591,N_16158);
and U21179 (N_21179,N_11674,N_11403);
or U21180 (N_21180,N_10877,N_11678);
nor U21181 (N_21181,N_15390,N_19854);
xor U21182 (N_21182,N_19449,N_13380);
or U21183 (N_21183,N_14948,N_12146);
and U21184 (N_21184,N_18847,N_14075);
xnor U21185 (N_21185,N_14547,N_15813);
xor U21186 (N_21186,N_13555,N_14879);
nor U21187 (N_21187,N_15644,N_12407);
and U21188 (N_21188,N_14480,N_11349);
nand U21189 (N_21189,N_12550,N_12914);
nand U21190 (N_21190,N_18866,N_17629);
nor U21191 (N_21191,N_13018,N_11780);
or U21192 (N_21192,N_13412,N_14384);
nand U21193 (N_21193,N_18170,N_19617);
nor U21194 (N_21194,N_12265,N_11512);
nor U21195 (N_21195,N_13250,N_13097);
nand U21196 (N_21196,N_19593,N_19657);
nand U21197 (N_21197,N_13654,N_10161);
nand U21198 (N_21198,N_15329,N_16350);
nor U21199 (N_21199,N_19110,N_10661);
nor U21200 (N_21200,N_13311,N_18669);
and U21201 (N_21201,N_19186,N_11752);
or U21202 (N_21202,N_12261,N_15037);
nand U21203 (N_21203,N_11692,N_12937);
or U21204 (N_21204,N_19035,N_16690);
nand U21205 (N_21205,N_15032,N_14146);
nor U21206 (N_21206,N_11622,N_19530);
xor U21207 (N_21207,N_15615,N_16490);
nor U21208 (N_21208,N_10557,N_14540);
and U21209 (N_21209,N_18207,N_18570);
nand U21210 (N_21210,N_16655,N_10970);
nand U21211 (N_21211,N_14377,N_14783);
or U21212 (N_21212,N_15764,N_10805);
nor U21213 (N_21213,N_12768,N_19537);
and U21214 (N_21214,N_10889,N_14006);
xnor U21215 (N_21215,N_17841,N_14326);
xnor U21216 (N_21216,N_17153,N_18788);
nand U21217 (N_21217,N_16069,N_19193);
nand U21218 (N_21218,N_10898,N_13214);
and U21219 (N_21219,N_18717,N_13016);
or U21220 (N_21220,N_15798,N_17241);
or U21221 (N_21221,N_12701,N_17971);
nor U21222 (N_21222,N_13851,N_19418);
and U21223 (N_21223,N_15248,N_18760);
nand U21224 (N_21224,N_11126,N_16812);
xnor U21225 (N_21225,N_17990,N_18515);
nor U21226 (N_21226,N_13024,N_18112);
or U21227 (N_21227,N_17645,N_19918);
or U21228 (N_21228,N_15319,N_14805);
nand U21229 (N_21229,N_15462,N_11694);
nor U21230 (N_21230,N_18467,N_18140);
and U21231 (N_21231,N_17934,N_14513);
nand U21232 (N_21232,N_11791,N_13856);
and U21233 (N_21233,N_14201,N_14760);
and U21234 (N_21234,N_11699,N_19904);
and U21235 (N_21235,N_17477,N_11333);
nor U21236 (N_21236,N_18100,N_17395);
xor U21237 (N_21237,N_15278,N_10506);
or U21238 (N_21238,N_14494,N_17423);
or U21239 (N_21239,N_12916,N_15271);
and U21240 (N_21240,N_10751,N_13582);
nand U21241 (N_21241,N_12452,N_14334);
nor U21242 (N_21242,N_15984,N_14129);
and U21243 (N_21243,N_18947,N_12610);
or U21244 (N_21244,N_18214,N_14478);
nand U21245 (N_21245,N_12835,N_14445);
and U21246 (N_21246,N_10657,N_11573);
xnor U21247 (N_21247,N_10067,N_13145);
and U21248 (N_21248,N_12370,N_12776);
nand U21249 (N_21249,N_12272,N_16667);
nor U21250 (N_21250,N_13937,N_17410);
nor U21251 (N_21251,N_16575,N_19658);
and U21252 (N_21252,N_11051,N_17348);
or U21253 (N_21253,N_11289,N_12313);
or U21254 (N_21254,N_13191,N_16775);
nand U21255 (N_21255,N_17125,N_16996);
nor U21256 (N_21256,N_17294,N_16957);
nand U21257 (N_21257,N_18843,N_13329);
and U21258 (N_21258,N_16980,N_11499);
and U21259 (N_21259,N_15110,N_19136);
nor U21260 (N_21260,N_10597,N_19458);
and U21261 (N_21261,N_11478,N_10264);
nor U21262 (N_21262,N_13300,N_17412);
nand U21263 (N_21263,N_12545,N_14455);
nor U21264 (N_21264,N_18681,N_15744);
or U21265 (N_21265,N_12005,N_11865);
or U21266 (N_21266,N_16238,N_16567);
xnor U21267 (N_21267,N_17483,N_13549);
or U21268 (N_21268,N_14007,N_14937);
nand U21269 (N_21269,N_10581,N_17337);
or U21270 (N_21270,N_11044,N_12625);
or U21271 (N_21271,N_13444,N_16018);
nand U21272 (N_21272,N_14683,N_14631);
xor U21273 (N_21273,N_14759,N_15504);
nand U21274 (N_21274,N_18156,N_14453);
or U21275 (N_21275,N_10887,N_13547);
and U21276 (N_21276,N_10825,N_19884);
or U21277 (N_21277,N_19546,N_10696);
nor U21278 (N_21278,N_16696,N_19612);
xnor U21279 (N_21279,N_17351,N_14714);
or U21280 (N_21280,N_15428,N_15964);
nor U21281 (N_21281,N_11994,N_12644);
and U21282 (N_21282,N_15204,N_11135);
or U21283 (N_21283,N_18268,N_19695);
nand U21284 (N_21284,N_16762,N_12861);
and U21285 (N_21285,N_14374,N_18948);
and U21286 (N_21286,N_10387,N_14247);
and U21287 (N_21287,N_13069,N_19199);
and U21288 (N_21288,N_11062,N_13364);
xor U21289 (N_21289,N_13700,N_19133);
and U21290 (N_21290,N_11342,N_11503);
nand U21291 (N_21291,N_13316,N_18869);
or U21292 (N_21292,N_19646,N_15424);
or U21293 (N_21293,N_18714,N_18832);
or U21294 (N_21294,N_13532,N_11875);
xnor U21295 (N_21295,N_16553,N_10502);
nand U21296 (N_21296,N_12238,N_18384);
or U21297 (N_21297,N_13195,N_13330);
and U21298 (N_21298,N_15583,N_14330);
xor U21299 (N_21299,N_15309,N_11584);
nand U21300 (N_21300,N_19420,N_15572);
or U21301 (N_21301,N_15561,N_16928);
or U21302 (N_21302,N_10864,N_15959);
or U21303 (N_21303,N_14966,N_16147);
and U21304 (N_21304,N_16530,N_15269);
or U21305 (N_21305,N_16127,N_16253);
and U21306 (N_21306,N_16263,N_16152);
nand U21307 (N_21307,N_18056,N_16973);
nand U21308 (N_21308,N_14468,N_11267);
nand U21309 (N_21309,N_15991,N_12375);
nand U21310 (N_21310,N_11379,N_18691);
and U21311 (N_21311,N_19633,N_11172);
nor U21312 (N_21312,N_15628,N_15251);
nand U21313 (N_21313,N_15261,N_13298);
nand U21314 (N_21314,N_11535,N_16609);
or U21315 (N_21315,N_17970,N_17469);
or U21316 (N_21316,N_12081,N_15872);
nand U21317 (N_21317,N_19475,N_16889);
nor U21318 (N_21318,N_15151,N_10492);
or U21319 (N_21319,N_17397,N_12851);
or U21320 (N_21320,N_17229,N_16059);
and U21321 (N_21321,N_13258,N_17903);
or U21322 (N_21322,N_16184,N_13171);
or U21323 (N_21323,N_16874,N_16846);
or U21324 (N_21324,N_19149,N_15554);
nor U21325 (N_21325,N_14863,N_13267);
or U21326 (N_21326,N_14309,N_15823);
and U21327 (N_21327,N_16173,N_17775);
nor U21328 (N_21328,N_17067,N_13163);
or U21329 (N_21329,N_10220,N_10364);
or U21330 (N_21330,N_12908,N_16589);
or U21331 (N_21331,N_14122,N_15033);
and U21332 (N_21332,N_12463,N_10153);
nand U21333 (N_21333,N_18251,N_19865);
nand U21334 (N_21334,N_11018,N_18008);
and U21335 (N_21335,N_15997,N_14900);
nor U21336 (N_21336,N_11827,N_18307);
or U21337 (N_21337,N_10029,N_16019);
nor U21338 (N_21338,N_15363,N_18304);
or U21339 (N_21339,N_19446,N_18608);
nor U21340 (N_21340,N_17712,N_12104);
xor U21341 (N_21341,N_11642,N_14314);
or U21342 (N_21342,N_13820,N_17448);
or U21343 (N_21343,N_11144,N_12177);
nor U21344 (N_21344,N_19081,N_16953);
or U21345 (N_21345,N_18219,N_12251);
nor U21346 (N_21346,N_16781,N_15016);
nor U21347 (N_21347,N_15420,N_18016);
or U21348 (N_21348,N_11419,N_14081);
nand U21349 (N_21349,N_15454,N_11666);
or U21350 (N_21350,N_16699,N_10568);
nand U21351 (N_21351,N_13724,N_10840);
nand U21352 (N_21352,N_14793,N_17936);
or U21353 (N_21353,N_14313,N_17946);
or U21354 (N_21354,N_16720,N_17676);
or U21355 (N_21355,N_16148,N_12053);
or U21356 (N_21356,N_13352,N_15886);
nor U21357 (N_21357,N_16602,N_18720);
xnor U21358 (N_21358,N_14459,N_17573);
xnor U21359 (N_21359,N_12002,N_11736);
and U21360 (N_21360,N_12597,N_12842);
nand U21361 (N_21361,N_15723,N_10831);
nor U21362 (N_21362,N_14986,N_15833);
xor U21363 (N_21363,N_16949,N_10882);
or U21364 (N_21364,N_14443,N_12616);
nor U21365 (N_21365,N_12549,N_13897);
and U21366 (N_21366,N_15770,N_11249);
or U21367 (N_21367,N_10790,N_11408);
nand U21368 (N_21368,N_12533,N_12481);
nand U21369 (N_21369,N_16875,N_11475);
or U21370 (N_21370,N_11488,N_18627);
and U21371 (N_21371,N_18135,N_18566);
nor U21372 (N_21372,N_11216,N_10704);
xnor U21373 (N_21373,N_11515,N_18144);
or U21374 (N_21374,N_14516,N_10513);
xnor U21375 (N_21375,N_10745,N_18684);
or U21376 (N_21376,N_11815,N_11429);
or U21377 (N_21377,N_10531,N_14518);
nor U21378 (N_21378,N_13117,N_15601);
and U21379 (N_21379,N_13510,N_13997);
nand U21380 (N_21380,N_13441,N_10672);
nand U21381 (N_21381,N_15670,N_18526);
and U21382 (N_21382,N_17601,N_16716);
nand U21383 (N_21383,N_14121,N_17921);
nor U21384 (N_21384,N_16099,N_19528);
or U21385 (N_21385,N_18086,N_10183);
nand U21386 (N_21386,N_17244,N_18767);
xnor U21387 (N_21387,N_17484,N_12980);
nand U21388 (N_21388,N_11421,N_12721);
and U21389 (N_21389,N_17700,N_11492);
or U21390 (N_21390,N_14822,N_16155);
or U21391 (N_21391,N_17260,N_17768);
nand U21392 (N_21392,N_13527,N_12587);
nand U21393 (N_21393,N_13447,N_17387);
and U21394 (N_21394,N_12902,N_10498);
or U21395 (N_21395,N_14974,N_10964);
and U21396 (N_21396,N_18721,N_12382);
nor U21397 (N_21397,N_16368,N_13890);
nor U21398 (N_21398,N_15795,N_15891);
nor U21399 (N_21399,N_11405,N_11750);
nor U21400 (N_21400,N_18814,N_19365);
nor U21401 (N_21401,N_11631,N_14285);
and U21402 (N_21402,N_11147,N_15799);
nand U21403 (N_21403,N_19404,N_16751);
or U21404 (N_21404,N_18057,N_18543);
nand U21405 (N_21405,N_18651,N_18835);
nand U21406 (N_21406,N_11082,N_16822);
nor U21407 (N_21407,N_18716,N_16518);
nand U21408 (N_21408,N_10637,N_11901);
nand U21409 (N_21409,N_15498,N_18457);
nor U21410 (N_21410,N_10875,N_18565);
nor U21411 (N_21411,N_13946,N_10504);
nor U21412 (N_21412,N_10803,N_14482);
nand U21413 (N_21413,N_14072,N_18432);
xor U21414 (N_21414,N_12722,N_10041);
and U21415 (N_21415,N_17093,N_10702);
or U21416 (N_21416,N_16723,N_10226);
and U21417 (N_21417,N_12494,N_18645);
nor U21418 (N_21418,N_12986,N_13977);
or U21419 (N_21419,N_12069,N_16670);
and U21420 (N_21420,N_11469,N_14716);
or U21421 (N_21421,N_10236,N_17779);
and U21422 (N_21422,N_16582,N_18359);
and U21423 (N_21423,N_10824,N_16222);
xnor U21424 (N_21424,N_19462,N_14179);
nand U21425 (N_21425,N_19929,N_19337);
or U21426 (N_21426,N_17704,N_18407);
or U21427 (N_21427,N_10788,N_16262);
nor U21428 (N_21428,N_17235,N_15820);
nand U21429 (N_21429,N_17638,N_16808);
nor U21430 (N_21430,N_18200,N_10345);
and U21431 (N_21431,N_10793,N_12634);
and U21432 (N_21432,N_11725,N_11661);
and U21433 (N_21433,N_15043,N_19587);
or U21434 (N_21434,N_15952,N_13843);
xnor U21435 (N_21435,N_10249,N_10972);
or U21436 (N_21436,N_11877,N_17303);
or U21437 (N_21437,N_10625,N_18472);
or U21438 (N_21438,N_16452,N_14778);
nor U21439 (N_21439,N_12206,N_17980);
nor U21440 (N_21440,N_13866,N_15325);
xor U21441 (N_21441,N_16446,N_10251);
or U21442 (N_21442,N_18225,N_16642);
nor U21443 (N_21443,N_17508,N_11788);
and U21444 (N_21444,N_13067,N_13132);
nand U21445 (N_21445,N_17333,N_18269);
and U21446 (N_21446,N_14647,N_10062);
or U21447 (N_21447,N_17941,N_14555);
or U21448 (N_21448,N_13595,N_12423);
xor U21449 (N_21449,N_11893,N_10660);
and U21450 (N_21450,N_17111,N_19455);
or U21451 (N_21451,N_17973,N_15604);
or U21452 (N_21452,N_12738,N_15811);
xnor U21453 (N_21453,N_16337,N_13456);
xor U21454 (N_21454,N_13370,N_18453);
xnor U21455 (N_21455,N_11544,N_18927);
xor U21456 (N_21456,N_15222,N_18234);
or U21457 (N_21457,N_16026,N_19105);
or U21458 (N_21458,N_13259,N_11268);
nor U21459 (N_21459,N_16526,N_12974);
nand U21460 (N_21460,N_18928,N_16872);
nor U21461 (N_21461,N_12605,N_16867);
xnor U21462 (N_21462,N_19017,N_10812);
or U21463 (N_21463,N_18518,N_12425);
nor U21464 (N_21464,N_12420,N_15488);
xnor U21465 (N_21465,N_19720,N_19421);
nand U21466 (N_21466,N_10997,N_13469);
and U21467 (N_21467,N_13443,N_16789);
and U21468 (N_21468,N_18825,N_17906);
nor U21469 (N_21469,N_14779,N_12548);
and U21470 (N_21470,N_17476,N_12730);
nand U21471 (N_21471,N_14533,N_18749);
nor U21472 (N_21472,N_11084,N_17076);
or U21473 (N_21473,N_16488,N_10653);
nor U21474 (N_21474,N_12314,N_19945);
nand U21475 (N_21475,N_11905,N_11958);
nand U21476 (N_21476,N_15745,N_15406);
nor U21477 (N_21477,N_14614,N_11751);
nand U21478 (N_21478,N_10133,N_17414);
nor U21479 (N_21479,N_17558,N_14049);
nor U21480 (N_21480,N_17586,N_19197);
or U21481 (N_21481,N_19758,N_16717);
nor U21482 (N_21482,N_17373,N_14178);
nor U21483 (N_21483,N_13247,N_13906);
or U21484 (N_21484,N_14530,N_14209);
or U21485 (N_21485,N_10283,N_13694);
or U21486 (N_21486,N_13541,N_12337);
and U21487 (N_21487,N_18761,N_12327);
nor U21488 (N_21488,N_11594,N_18350);
nor U21489 (N_21489,N_14317,N_10043);
nor U21490 (N_21490,N_14236,N_16044);
or U21491 (N_21491,N_19760,N_17231);
nand U21492 (N_21492,N_10536,N_11310);
xor U21493 (N_21493,N_13765,N_18952);
nand U21494 (N_21494,N_17060,N_14380);
nand U21495 (N_21495,N_14365,N_16543);
nor U21496 (N_21496,N_16512,N_18977);
nand U21497 (N_21497,N_19128,N_16687);
nor U21498 (N_21498,N_17822,N_12754);
nand U21499 (N_21499,N_18858,N_19618);
xor U21500 (N_21500,N_19367,N_18256);
nor U21501 (N_21501,N_10801,N_13503);
and U21502 (N_21502,N_17496,N_11768);
nand U21503 (N_21503,N_17330,N_13621);
or U21504 (N_21504,N_10828,N_14644);
nand U21505 (N_21505,N_16381,N_17148);
and U21506 (N_21506,N_10190,N_12575);
xnor U21507 (N_21507,N_14074,N_10010);
or U21508 (N_21508,N_13999,N_17795);
nand U21509 (N_21509,N_14130,N_14654);
nor U21510 (N_21510,N_18021,N_11681);
and U21511 (N_21511,N_15262,N_17155);
nor U21512 (N_21512,N_12505,N_16008);
or U21513 (N_21513,N_15735,N_16835);
nand U21514 (N_21514,N_14987,N_16937);
xor U21515 (N_21515,N_13121,N_16344);
or U21516 (N_21516,N_10723,N_16406);
and U21517 (N_21517,N_16864,N_18232);
nor U21518 (N_21518,N_14549,N_14260);
and U21519 (N_21519,N_19250,N_18126);
nor U21520 (N_21520,N_15758,N_12802);
nand U21521 (N_21521,N_10229,N_17158);
or U21522 (N_21522,N_19254,N_11700);
nand U21523 (N_21523,N_10892,N_13667);
nand U21524 (N_21524,N_14167,N_19549);
or U21525 (N_21525,N_14255,N_15315);
nand U21526 (N_21526,N_18650,N_11962);
nand U21527 (N_21527,N_10911,N_12586);
or U21528 (N_21528,N_18806,N_16896);
nor U21529 (N_21529,N_12473,N_10412);
nor U21530 (N_21530,N_18799,N_10044);
nand U21531 (N_21531,N_14305,N_18702);
xnor U21532 (N_21532,N_16508,N_12170);
nand U21533 (N_21533,N_18991,N_14427);
nor U21534 (N_21534,N_17446,N_14014);
or U21535 (N_21535,N_12111,N_12480);
nor U21536 (N_21536,N_17103,N_14343);
and U21537 (N_21537,N_17621,N_14550);
nand U21538 (N_21538,N_13209,N_17127);
and U21539 (N_21539,N_14219,N_14291);
or U21540 (N_21540,N_14580,N_16627);
xnor U21541 (N_21541,N_12855,N_14301);
or U21542 (N_21542,N_14452,N_10695);
or U21543 (N_21543,N_14391,N_14190);
nand U21544 (N_21544,N_14315,N_11001);
nand U21545 (N_21545,N_15707,N_17765);
xor U21546 (N_21546,N_11368,N_18132);
nor U21547 (N_21547,N_12953,N_15521);
or U21548 (N_21548,N_17461,N_13525);
nor U21549 (N_21549,N_14344,N_12302);
and U21550 (N_21550,N_15083,N_18116);
and U21551 (N_21551,N_17721,N_17377);
nor U21552 (N_21552,N_11173,N_14589);
and U21553 (N_21553,N_10246,N_11956);
and U21554 (N_21554,N_14000,N_18968);
and U21555 (N_21555,N_13919,N_18781);
nor U21556 (N_21556,N_10114,N_16647);
or U21557 (N_21557,N_11290,N_12965);
xor U21558 (N_21558,N_18876,N_16302);
nand U21559 (N_21559,N_15533,N_10012);
xor U21560 (N_21560,N_14208,N_14917);
or U21561 (N_21561,N_13647,N_16746);
and U21562 (N_21562,N_18330,N_13183);
or U21563 (N_21563,N_17070,N_16476);
nand U21564 (N_21564,N_15355,N_15683);
or U21565 (N_21565,N_12681,N_18910);
xor U21566 (N_21566,N_11904,N_11925);
nand U21567 (N_21567,N_14079,N_19925);
nor U21568 (N_21568,N_16800,N_18489);
or U21569 (N_21569,N_17363,N_16494);
and U21570 (N_21570,N_16532,N_14571);
and U21571 (N_21571,N_13852,N_12424);
nand U21572 (N_21572,N_14699,N_14211);
xnor U21573 (N_21573,N_12197,N_14869);
nand U21574 (N_21574,N_18152,N_13934);
nor U21575 (N_21575,N_17023,N_14829);
or U21576 (N_21576,N_18168,N_16382);
nor U21577 (N_21577,N_12296,N_12554);
and U21578 (N_21578,N_19688,N_14739);
or U21579 (N_21579,N_16387,N_19058);
or U21580 (N_21580,N_13061,N_13612);
and U21581 (N_21581,N_17709,N_15333);
xnor U21582 (N_21582,N_12001,N_15958);
nor U21583 (N_21583,N_17862,N_13397);
nand U21584 (N_21584,N_15353,N_18790);
or U21585 (N_21585,N_18885,N_13011);
and U21586 (N_21586,N_11325,N_11903);
nor U21587 (N_21587,N_15144,N_12796);
nand U21588 (N_21588,N_10669,N_12387);
or U21589 (N_21589,N_15564,N_10414);
nand U21590 (N_21590,N_11187,N_11095);
and U21591 (N_21591,N_16625,N_19894);
nand U21592 (N_21592,N_12818,N_19235);
and U21593 (N_21593,N_17777,N_10977);
or U21594 (N_21594,N_11041,N_18285);
or U21595 (N_21595,N_13383,N_14786);
or U21596 (N_21596,N_17981,N_19956);
nand U21597 (N_21597,N_16951,N_11286);
or U21598 (N_21598,N_17519,N_13043);
or U21599 (N_21599,N_15418,N_16727);
or U21600 (N_21600,N_14971,N_13217);
and U21601 (N_21601,N_13219,N_14281);
and U21602 (N_21602,N_10401,N_11663);
or U21603 (N_21603,N_15119,N_19577);
or U21604 (N_21604,N_18435,N_18800);
and U21605 (N_21605,N_13373,N_12490);
nor U21606 (N_21606,N_15039,N_13236);
and U21607 (N_21607,N_11462,N_10960);
or U21608 (N_21608,N_11027,N_11822);
and U21609 (N_21609,N_12859,N_11516);
and U21610 (N_21610,N_11940,N_17715);
xor U21611 (N_21611,N_11567,N_15685);
nand U21612 (N_21612,N_16486,N_19041);
nor U21613 (N_21613,N_17552,N_17805);
and U21614 (N_21614,N_16360,N_16039);
and U21615 (N_21615,N_13760,N_14690);
or U21616 (N_21616,N_17881,N_19068);
nand U21617 (N_21617,N_11757,N_12702);
and U21618 (N_21618,N_17791,N_11311);
nor U21619 (N_21619,N_14244,N_17732);
nor U21620 (N_21620,N_14664,N_12045);
nor U21621 (N_21621,N_13010,N_16373);
nand U21622 (N_21622,N_19470,N_12837);
or U21623 (N_21623,N_16594,N_18616);
nand U21624 (N_21624,N_12913,N_19648);
nor U21625 (N_21625,N_17170,N_19851);
or U21626 (N_21626,N_19167,N_11651);
or U21627 (N_21627,N_14568,N_16176);
nand U21628 (N_21628,N_13124,N_14257);
and U21629 (N_21629,N_12726,N_11025);
nand U21630 (N_21630,N_11707,N_12630);
or U21631 (N_21631,N_10789,N_18777);
nand U21632 (N_21632,N_13466,N_13007);
nor U21633 (N_21633,N_16736,N_15207);
and U21634 (N_21634,N_13332,N_14845);
nor U21635 (N_21635,N_14785,N_19236);
or U21636 (N_21636,N_14215,N_13811);
nor U21637 (N_21637,N_16054,N_15895);
nand U21638 (N_21638,N_10369,N_14728);
xnor U21639 (N_21639,N_16752,N_15028);
nand U21640 (N_21640,N_13772,N_10478);
and U21641 (N_21641,N_12036,N_19230);
xor U21642 (N_21642,N_17961,N_10217);
xor U21643 (N_21643,N_18791,N_13602);
nand U21644 (N_21644,N_15551,N_12664);
xnor U21645 (N_21645,N_16234,N_19155);
and U21646 (N_21646,N_18075,N_19611);
and U21647 (N_21647,N_18884,N_19552);
nand U21648 (N_21648,N_17693,N_18603);
nor U21649 (N_21649,N_16712,N_19844);
or U21650 (N_21650,N_18996,N_16744);
nand U21651 (N_21651,N_11479,N_10017);
nand U21652 (N_21652,N_15986,N_14575);
or U21653 (N_21653,N_17568,N_13382);
and U21654 (N_21654,N_12810,N_14448);
xor U21655 (N_21655,N_11574,N_19380);
xnor U21656 (N_21656,N_13673,N_18392);
nand U21657 (N_21657,N_13293,N_10771);
and U21658 (N_21658,N_12555,N_11769);
nor U21659 (N_21659,N_15949,N_11701);
nand U21660 (N_21660,N_16600,N_17248);
or U21661 (N_21661,N_14574,N_10076);
and U21662 (N_21662,N_17355,N_18101);
xnor U21663 (N_21663,N_18128,N_15585);
nor U21664 (N_21664,N_16457,N_11337);
nor U21665 (N_21665,N_10407,N_14287);
or U21666 (N_21666,N_16819,N_14653);
nand U21667 (N_21667,N_17426,N_19864);
nor U21668 (N_21668,N_11521,N_18136);
nor U21669 (N_21669,N_10087,N_17072);
and U21670 (N_21670,N_16489,N_17104);
nand U21671 (N_21671,N_17304,N_16533);
and U21672 (N_21672,N_14431,N_18542);
or U21673 (N_21673,N_13879,N_13837);
and U21674 (N_21674,N_18984,N_12252);
nor U21675 (N_21675,N_17422,N_17814);
nor U21676 (N_21676,N_12744,N_14926);
nand U21677 (N_21677,N_15180,N_11105);
or U21678 (N_21678,N_12674,N_13264);
nand U21679 (N_21679,N_15179,N_10694);
nand U21680 (N_21680,N_15414,N_12899);
nor U21681 (N_21681,N_17462,N_16189);
nand U21682 (N_21682,N_18820,N_12729);
or U21683 (N_21683,N_16153,N_13112);
nand U21684 (N_21684,N_13266,N_16538);
and U21685 (N_21685,N_16224,N_11595);
xnor U21686 (N_21686,N_10248,N_17771);
nor U21687 (N_21687,N_14742,N_17435);
or U21688 (N_21688,N_18491,N_15408);
nand U21689 (N_21689,N_12306,N_19567);
nand U21690 (N_21690,N_19402,N_19101);
and U21691 (N_21691,N_15849,N_12565);
nor U21692 (N_21692,N_10106,N_15375);
and U21693 (N_21693,N_15378,N_10442);
nand U21694 (N_21694,N_19152,N_17550);
nand U21695 (N_21695,N_18406,N_16500);
nand U21696 (N_21696,N_11060,N_15814);
or U21697 (N_21697,N_11284,N_18470);
and U21698 (N_21698,N_15938,N_18042);
and U21699 (N_21699,N_19287,N_16585);
nor U21700 (N_21700,N_12983,N_13869);
or U21701 (N_21701,N_13963,N_10417);
nor U21702 (N_21702,N_15904,N_13819);
nor U21703 (N_21703,N_18211,N_12372);
and U21704 (N_21704,N_14858,N_13116);
or U21705 (N_21705,N_18817,N_10501);
nor U21706 (N_21706,N_13701,N_13807);
xor U21707 (N_21707,N_15242,N_19379);
or U21708 (N_21708,N_10189,N_17870);
nor U21709 (N_21709,N_17319,N_15360);
nand U21710 (N_21710,N_18043,N_10205);
or U21711 (N_21711,N_19623,N_10175);
and U21712 (N_21712,N_15977,N_11712);
nor U21713 (N_21713,N_14266,N_16551);
nor U21714 (N_21714,N_17189,N_10746);
nor U21715 (N_21715,N_13189,N_16276);
xnor U21716 (N_21716,N_14707,N_11335);
and U21717 (N_21717,N_13531,N_13538);
xnor U21718 (N_21718,N_11636,N_11672);
or U21719 (N_21719,N_13178,N_12539);
and U21720 (N_21720,N_18633,N_19534);
nand U21721 (N_21721,N_14096,N_16883);
nand U21722 (N_21722,N_14333,N_19812);
nor U21723 (N_21723,N_16217,N_10518);
and U21724 (N_21724,N_16051,N_11667);
or U21725 (N_21725,N_12903,N_19166);
and U21726 (N_21726,N_16082,N_13356);
or U21727 (N_21727,N_18988,N_11259);
or U21728 (N_21728,N_19885,N_14404);
or U21729 (N_21729,N_12830,N_19122);
nand U21730 (N_21730,N_13392,N_19913);
nor U21731 (N_21731,N_17835,N_19056);
xnor U21732 (N_21732,N_15342,N_15693);
and U21733 (N_21733,N_18398,N_11128);
xor U21734 (N_21734,N_17909,N_17739);
or U21735 (N_21735,N_13543,N_10634);
and U21736 (N_21736,N_19831,N_15246);
xor U21737 (N_21737,N_12516,N_11200);
nor U21738 (N_21738,N_14643,N_19099);
nand U21739 (N_21739,N_16404,N_19886);
and U21740 (N_21740,N_15302,N_17703);
xnor U21741 (N_21741,N_10357,N_18011);
nand U21742 (N_21742,N_18362,N_13902);
nor U21743 (N_21743,N_12592,N_16884);
xnor U21744 (N_21744,N_17634,N_11194);
or U21745 (N_21745,N_15260,N_19645);
or U21746 (N_21746,N_19408,N_18859);
nand U21747 (N_21747,N_15074,N_12798);
or U21748 (N_21748,N_11320,N_17993);
and U21749 (N_21749,N_16003,N_11816);
or U21750 (N_21750,N_12180,N_12264);
or U21751 (N_21751,N_14615,N_12609);
nand U21752 (N_21752,N_13500,N_17369);
or U21753 (N_21753,N_19437,N_17161);
nor U21754 (N_21754,N_19810,N_17340);
or U21755 (N_21755,N_16041,N_19993);
xor U21756 (N_21756,N_14187,N_16353);
nor U21757 (N_21757,N_15751,N_17735);
nor U21758 (N_21758,N_19203,N_15344);
nand U21759 (N_21759,N_16492,N_14777);
and U21760 (N_21760,N_18899,N_15861);
nand U21761 (N_21761,N_17710,N_13642);
nor U21762 (N_21762,N_19355,N_19922);
nand U21763 (N_21763,N_16796,N_15863);
xnor U21764 (N_21764,N_16767,N_10567);
or U21765 (N_21765,N_14973,N_18283);
nor U21766 (N_21766,N_15439,N_17539);
xor U21767 (N_21767,N_15979,N_10009);
and U21768 (N_21768,N_14082,N_17206);
and U21769 (N_21769,N_15129,N_15000);
nand U21770 (N_21770,N_11158,N_18199);
nand U21771 (N_21771,N_12441,N_18196);
nand U21772 (N_21772,N_13844,N_12055);
nor U21773 (N_21773,N_17806,N_16688);
xor U21774 (N_21774,N_14161,N_11562);
nor U21775 (N_21775,N_13422,N_18536);
or U21776 (N_21776,N_18987,N_16020);
and U21777 (N_21777,N_10666,N_16278);
nand U21778 (N_21778,N_14460,N_18443);
nand U21779 (N_21779,N_16695,N_13423);
nor U21780 (N_21780,N_18938,N_15648);
or U21781 (N_21781,N_18024,N_12074);
nand U21782 (N_21782,N_13818,N_19536);
and U21783 (N_21783,N_13859,N_13491);
and U21784 (N_21784,N_13771,N_14663);
and U21785 (N_21785,N_19341,N_13128);
xor U21786 (N_21786,N_18762,N_19585);
and U21787 (N_21787,N_18123,N_18774);
or U21788 (N_21788,N_17523,N_13421);
nor U21789 (N_21789,N_10717,N_14202);
nor U21790 (N_21790,N_17570,N_10074);
and U21791 (N_21791,N_11282,N_10468);
nand U21792 (N_21792,N_10782,N_18188);
nand U21793 (N_21793,N_16861,N_17434);
nand U21794 (N_21794,N_10543,N_13704);
and U21795 (N_21795,N_12961,N_17796);
nand U21796 (N_21796,N_11441,N_15522);
nor U21797 (N_21797,N_16961,N_13415);
nor U21798 (N_21798,N_16375,N_12304);
xor U21799 (N_21799,N_12573,N_11440);
nand U21800 (N_21800,N_19626,N_16405);
and U21801 (N_21801,N_12769,N_10174);
or U21802 (N_21802,N_15137,N_16950);
or U21803 (N_21803,N_14543,N_16759);
or U21804 (N_21804,N_17433,N_14696);
or U21805 (N_21805,N_18400,N_15392);
xor U21806 (N_21806,N_17154,N_16425);
or U21807 (N_21807,N_17075,N_11463);
or U21808 (N_21808,N_13998,N_19533);
nor U21809 (N_21809,N_10626,N_14809);
and U21810 (N_21810,N_17534,N_19762);
or U21811 (N_21811,N_19888,N_12915);
or U21812 (N_21812,N_13816,N_12523);
or U21813 (N_21813,N_19158,N_10308);
nor U21814 (N_21814,N_13173,N_14969);
and U21815 (N_21815,N_16715,N_11553);
nor U21816 (N_21816,N_16828,N_16916);
nand U21817 (N_21817,N_15885,N_17855);
nor U21818 (N_21818,N_17400,N_10361);
xnor U21819 (N_21819,N_10777,N_10038);
and U21820 (N_21820,N_13152,N_14844);
or U21821 (N_21821,N_18903,N_19076);
and U21822 (N_21822,N_18437,N_16031);
or U21823 (N_21823,N_11929,N_17664);
xor U21824 (N_21824,N_19216,N_14735);
and U21825 (N_21825,N_16491,N_10185);
xnor U21826 (N_21826,N_19512,N_17717);
nor U21827 (N_21827,N_10376,N_17891);
nand U21828 (N_21828,N_13256,N_18436);
nor U21829 (N_21829,N_19429,N_15434);
nand U21830 (N_21830,N_12509,N_12312);
nand U21831 (N_21831,N_18065,N_15686);
and U21832 (N_21832,N_11677,N_13980);
nand U21833 (N_21833,N_18358,N_16972);
and U21834 (N_21834,N_10734,N_14667);
nor U21835 (N_21835,N_11003,N_16136);
xor U21836 (N_21836,N_15051,N_15372);
nor U21837 (N_21837,N_12960,N_12049);
or U21838 (N_21838,N_19785,N_15917);
or U21839 (N_21839,N_15981,N_14921);
nand U21840 (N_21840,N_19917,N_15412);
or U21841 (N_21841,N_19538,N_15206);
nor U21842 (N_21842,N_19188,N_12360);
nor U21843 (N_21843,N_16419,N_11695);
or U21844 (N_21844,N_19524,N_13987);
xor U21845 (N_21845,N_18532,N_12400);
nand U21846 (N_21846,N_17672,N_18000);
and U21847 (N_21847,N_14454,N_19394);
or U21848 (N_21848,N_19632,N_13076);
or U21849 (N_21849,N_17405,N_10957);
or U21850 (N_21850,N_13785,N_17251);
and U21851 (N_21851,N_16096,N_11415);
nor U21852 (N_21852,N_16046,N_17849);
nor U21853 (N_21853,N_11494,N_14586);
nor U21854 (N_21854,N_15702,N_10842);
xor U21855 (N_21855,N_11742,N_19700);
xor U21856 (N_21856,N_17134,N_18189);
nor U21857 (N_21857,N_13198,N_16346);
and U21858 (N_21858,N_18783,N_12604);
and U21859 (N_21859,N_11359,N_18670);
nor U21860 (N_21860,N_19255,N_10429);
nor U21861 (N_21861,N_11741,N_19433);
nand U21862 (N_21862,N_18246,N_12667);
or U21863 (N_21863,N_19273,N_12344);
or U21864 (N_21864,N_18819,N_13909);
nand U21865 (N_21865,N_10398,N_18244);
or U21866 (N_21866,N_10920,N_10007);
nand U21867 (N_21867,N_15759,N_14621);
and U21868 (N_21868,N_19414,N_10297);
or U21869 (N_21869,N_12449,N_11613);
or U21870 (N_21870,N_16560,N_13235);
nand U21871 (N_21871,N_16859,N_13751);
xor U21872 (N_21872,N_18605,N_13925);
and U21873 (N_21873,N_19824,N_19529);
nor U21874 (N_21874,N_17512,N_13339);
and U21875 (N_21875,N_13437,N_19222);
nor U21876 (N_21876,N_11183,N_19111);
or U21877 (N_21877,N_17171,N_16392);
nor U21878 (N_21878,N_10526,N_13402);
nor U21879 (N_21879,N_15846,N_15527);
nand U21880 (N_21880,N_15458,N_19037);
or U21881 (N_21881,N_13990,N_12829);
and U21882 (N_21882,N_14018,N_13928);
and U21883 (N_21883,N_13468,N_10768);
nor U21884 (N_21884,N_13393,N_11276);
xor U21885 (N_21885,N_16086,N_14611);
nor U21886 (N_21886,N_10077,N_12230);
or U21887 (N_21887,N_10807,N_11202);
nand U21888 (N_21888,N_14567,N_10690);
nand U21889 (N_21889,N_19996,N_19948);
and U21890 (N_21890,N_12991,N_19622);
and U21891 (N_21891,N_19336,N_18081);
nand U21892 (N_21892,N_10816,N_17288);
nor U21893 (N_21893,N_10191,N_18217);
nor U21894 (N_21894,N_15492,N_18410);
nand U21895 (N_21895,N_14205,N_19542);
and U21896 (N_21896,N_16395,N_15562);
and U21897 (N_21897,N_11620,N_19990);
nand U21898 (N_21898,N_10127,N_14457);
or U21899 (N_21899,N_18465,N_18378);
nor U21900 (N_21900,N_17136,N_16753);
and U21901 (N_21901,N_13748,N_14517);
and U21902 (N_21902,N_15456,N_17151);
or U21903 (N_21903,N_16112,N_14213);
nor U21904 (N_21904,N_15647,N_12848);
or U21905 (N_21905,N_12746,N_12984);
and U21906 (N_21906,N_17826,N_17871);
nor U21907 (N_21907,N_19185,N_18994);
nand U21908 (N_21908,N_13585,N_17978);
or U21909 (N_21909,N_12557,N_13699);
nor U21910 (N_21910,N_12525,N_18622);
xnor U21911 (N_21911,N_18815,N_18397);
and U21912 (N_21912,N_19855,N_13427);
nor U21913 (N_21913,N_16025,N_14893);
nor U21914 (N_21914,N_11952,N_19539);
xor U21915 (N_21915,N_14290,N_11974);
and U21916 (N_21916,N_10906,N_12191);
and U21917 (N_21917,N_12456,N_15120);
and U21918 (N_21918,N_15834,N_18331);
or U21919 (N_21919,N_17542,N_11558);
xnor U21920 (N_21920,N_16813,N_17474);
and U21921 (N_21921,N_15581,N_13319);
nor U21922 (N_21922,N_14150,N_18385);
or U21923 (N_21923,N_10362,N_11555);
or U21924 (N_21924,N_15162,N_17876);
nand U21925 (N_21925,N_12470,N_19115);
nand U21926 (N_21926,N_12160,N_13903);
or U21927 (N_21927,N_16043,N_19295);
nor U21928 (N_21928,N_11568,N_14637);
and U21929 (N_21929,N_15737,N_12115);
nor U21930 (N_21930,N_12184,N_18163);
nor U21931 (N_21931,N_15898,N_15467);
or U21932 (N_21932,N_10720,N_15578);
and U21933 (N_21933,N_12163,N_10446);
and U21934 (N_21934,N_15503,N_10974);
and U21935 (N_21935,N_12147,N_15971);
or U21936 (N_21936,N_14265,N_10507);
nand U21937 (N_21937,N_19498,N_15712);
nand U21938 (N_21938,N_13535,N_10904);
and U21939 (N_21939,N_19218,N_10131);
nand U21940 (N_21940,N_12059,N_11817);
nor U21941 (N_21941,N_15186,N_14485);
nor U21942 (N_21942,N_19610,N_16408);
or U21943 (N_21943,N_10156,N_14359);
xor U21944 (N_21944,N_16295,N_14856);
and U21945 (N_21945,N_19253,N_12044);
nand U21946 (N_21946,N_18026,N_10054);
nand U21947 (N_21947,N_11623,N_12725);
nand U21948 (N_21948,N_14465,N_17263);
or U21949 (N_21949,N_17190,N_16998);
nor U21950 (N_21950,N_17219,N_15957);
nor U21951 (N_21951,N_16157,N_11434);
and U21952 (N_21952,N_14490,N_13029);
nor U21953 (N_21953,N_12853,N_19667);
and U21954 (N_21954,N_19048,N_18495);
nor U21955 (N_21955,N_16260,N_10456);
or U21956 (N_21956,N_12346,N_19181);
and U21957 (N_21957,N_13932,N_13200);
nor U21958 (N_21958,N_16123,N_14599);
nand U21959 (N_21959,N_14565,N_10546);
nand U21960 (N_21960,N_16902,N_13096);
nand U21961 (N_21961,N_14685,N_18494);
or U21962 (N_21962,N_15499,N_17265);
and U21963 (N_21963,N_17254,N_15405);
nand U21964 (N_21964,N_19928,N_11231);
nand U21965 (N_21965,N_10135,N_17866);
and U21966 (N_21966,N_16166,N_17637);
nand U21967 (N_21967,N_10268,N_13333);
nand U21968 (N_21968,N_18596,N_13610);
and U21969 (N_21969,N_11055,N_13353);
or U21970 (N_21970,N_15796,N_15254);
nand U21971 (N_21971,N_12650,N_11656);
nand U21972 (N_21972,N_18035,N_12154);
or U21973 (N_21973,N_11908,N_19693);
or U21974 (N_21974,N_18607,N_15023);
nand U21975 (N_21975,N_14598,N_11258);
or U21976 (N_21976,N_10396,N_18319);
or U21977 (N_21977,N_13238,N_13978);
nor U21978 (N_21978,N_15998,N_14936);
and U21979 (N_21979,N_17286,N_11298);
and U21980 (N_21980,N_18538,N_19386);
nor U21981 (N_21981,N_17583,N_17554);
nand U21982 (N_21982,N_11077,N_18186);
xnor U21983 (N_21983,N_13002,N_13181);
nor U21984 (N_21984,N_18812,N_18265);
nor U21985 (N_21985,N_12307,N_16316);
or U21986 (N_21986,N_19431,N_14366);
nand U21987 (N_21987,N_12131,N_17240);
nor U21988 (N_21988,N_14890,N_16513);
nor U21989 (N_21989,N_14557,N_11345);
and U21990 (N_21990,N_10547,N_14059);
or U21991 (N_21991,N_12868,N_13348);
and U21992 (N_21992,N_11066,N_11397);
nand U21993 (N_21993,N_18068,N_17593);
or U21994 (N_21994,N_10046,N_16908);
and U21995 (N_21995,N_11843,N_17689);
xnor U21996 (N_21996,N_19219,N_18018);
and U21997 (N_21997,N_16171,N_14803);
or U21998 (N_21998,N_14419,N_18963);
nor U21999 (N_21999,N_16104,N_13881);
nand U22000 (N_22000,N_19775,N_12816);
nand U22001 (N_22001,N_16960,N_11834);
xnor U22002 (N_22002,N_15655,N_14489);
nor U22003 (N_22003,N_13592,N_10109);
or U22004 (N_22004,N_16080,N_18275);
nand U22005 (N_22005,N_11113,N_19321);
nor U22006 (N_22006,N_13485,N_15132);
nand U22007 (N_22007,N_14689,N_15830);
and U22008 (N_22008,N_15722,N_15556);
nand U22009 (N_22009,N_13484,N_11455);
or U22010 (N_22010,N_10592,N_16145);
and U22011 (N_22011,N_19624,N_15524);
nand U22012 (N_22012,N_16922,N_16038);
nand U22013 (N_22013,N_17365,N_18870);
and U22014 (N_22014,N_11059,N_10555);
or U22015 (N_22015,N_13159,N_10813);
nor U22016 (N_22016,N_18586,N_16540);
or U22017 (N_22017,N_13493,N_10564);
nor U22018 (N_22018,N_13628,N_14409);
and U22019 (N_22019,N_13841,N_14545);
or U22020 (N_22020,N_17808,N_17642);
and U22021 (N_22021,N_13995,N_11024);
nor U22022 (N_22022,N_11299,N_15304);
xnor U22023 (N_22023,N_16445,N_17057);
or U22024 (N_22024,N_14587,N_18742);
or U22025 (N_22025,N_19937,N_16683);
or U22026 (N_22026,N_18036,N_19836);
nand U22027 (N_22027,N_12171,N_16840);
xor U22028 (N_22028,N_11743,N_15657);
and U22029 (N_22029,N_17683,N_10610);
and U22030 (N_22030,N_19244,N_10628);
and U22031 (N_22031,N_18680,N_10529);
or U22032 (N_22032,N_18738,N_15230);
and U22033 (N_22033,N_16120,N_14814);
nand U22034 (N_22034,N_15875,N_14995);
xor U22035 (N_22035,N_17782,N_19485);
nand U22036 (N_22036,N_17641,N_11211);
nand U22037 (N_22037,N_11818,N_16075);
or U22038 (N_22038,N_19500,N_16081);
nor U22039 (N_22039,N_10028,N_16458);
and U22040 (N_22040,N_11197,N_19739);
nand U22041 (N_22041,N_19513,N_17549);
nand U22042 (N_22042,N_13846,N_18831);
nand U22043 (N_22043,N_11207,N_12092);
or U22044 (N_22044,N_13577,N_19967);
and U22045 (N_22045,N_12945,N_19441);
nand U22046 (N_22046,N_17954,N_19284);
and U22047 (N_22047,N_19621,N_12531);
and U22048 (N_22048,N_17336,N_16105);
and U22049 (N_22049,N_13648,N_10585);
nand U22050 (N_22050,N_11540,N_10089);
and U22051 (N_22051,N_18922,N_18291);
or U22052 (N_22052,N_15552,N_12416);
or U22053 (N_22053,N_17300,N_14953);
or U22054 (N_22054,N_14963,N_19213);
or U22055 (N_22055,N_14896,N_16848);
and U22056 (N_22056,N_14488,N_11196);
and U22057 (N_22057,N_19738,N_18936);
or U22058 (N_22058,N_11388,N_14410);
or U22059 (N_22059,N_17499,N_13564);
nor U22060 (N_22060,N_18585,N_13728);
nand U22061 (N_22061,N_10611,N_18260);
and U22062 (N_22062,N_19979,N_17968);
xnor U22063 (N_22063,N_17967,N_18322);
nor U22064 (N_22064,N_17366,N_19655);
nor U22065 (N_22065,N_15548,N_12222);
and U22066 (N_22066,N_10987,N_12085);
nor U22067 (N_22067,N_13578,N_13662);
nand U22068 (N_22068,N_12207,N_16677);
nand U22069 (N_22069,N_16969,N_13144);
nand U22070 (N_22070,N_10199,N_14341);
nor U22071 (N_22071,N_12125,N_18795);
nand U22072 (N_22072,N_14597,N_17404);
and U22073 (N_22073,N_17359,N_16849);
nor U22074 (N_22074,N_10282,N_15139);
nor U22075 (N_22075,N_11107,N_14950);
xnor U22076 (N_22076,N_11006,N_16510);
and U22077 (N_22077,N_11607,N_13825);
nand U22078 (N_22078,N_13968,N_17830);
nand U22079 (N_22079,N_15995,N_18780);
and U22080 (N_22080,N_13127,N_15637);
and U22081 (N_22081,N_12934,N_11042);
or U22082 (N_22082,N_17459,N_14939);
and U22083 (N_22083,N_16315,N_16921);
or U22084 (N_22084,N_10740,N_11588);
xor U22085 (N_22085,N_15298,N_18590);
and U22086 (N_22086,N_10967,N_10218);
nor U22087 (N_22087,N_11963,N_10213);
and U22088 (N_22088,N_13747,N_13262);
and U22089 (N_22089,N_11606,N_15534);
or U22090 (N_22090,N_17399,N_15701);
nand U22091 (N_22091,N_10256,N_11278);
xor U22092 (N_22092,N_16581,N_18955);
nand U22093 (N_22093,N_19707,N_12631);
nor U22094 (N_22094,N_13814,N_15034);
or U22095 (N_22095,N_17660,N_13058);
nor U22096 (N_22096,N_15884,N_18158);
nor U22097 (N_22097,N_11941,N_18901);
nand U22098 (N_22098,N_10591,N_16565);
xor U22099 (N_22099,N_14899,N_16355);
nand U22100 (N_22100,N_18690,N_19389);
or U22101 (N_22101,N_15515,N_12803);
and U22102 (N_22102,N_14105,N_11835);
or U22103 (N_22103,N_14886,N_15227);
or U22104 (N_22104,N_12824,N_11448);
and U22105 (N_22105,N_14083,N_10075);
xnor U22106 (N_22106,N_13971,N_18972);
nor U22107 (N_22107,N_16704,N_12775);
and U22108 (N_22108,N_19735,N_13405);
nand U22109 (N_22109,N_14694,N_16407);
or U22110 (N_22110,N_12287,N_17326);
nand U22111 (N_22111,N_16525,N_15794);
and U22112 (N_22112,N_17692,N_16470);
nand U22113 (N_22113,N_15825,N_14311);
or U22114 (N_22114,N_11966,N_12823);
nor U22115 (N_22115,N_11303,N_15249);
and U22116 (N_22116,N_16788,N_11093);
and U22117 (N_22117,N_11034,N_13681);
nor U22118 (N_22118,N_13394,N_18368);
or U22119 (N_22119,N_14496,N_18487);
nor U22120 (N_22120,N_18476,N_12563);
or U22121 (N_22121,N_10935,N_17261);
xnor U22122 (N_22122,N_16801,N_18865);
xnor U22123 (N_22123,N_13872,N_16568);
nand U22124 (N_22124,N_16339,N_10978);
nor U22125 (N_22125,N_16466,N_11527);
nor U22126 (N_22126,N_12242,N_16168);
nand U22127 (N_22127,N_15463,N_17950);
and U22128 (N_22128,N_14458,N_19377);
nand U22129 (N_22129,N_17123,N_18682);
nand U22130 (N_22130,N_11366,N_11518);
nor U22131 (N_22131,N_14582,N_18625);
and U22132 (N_22132,N_15784,N_15935);
xor U22133 (N_22133,N_16659,N_16920);
xor U22134 (N_22134,N_14618,N_12046);
or U22135 (N_22135,N_15308,N_15061);
nor U22136 (N_22136,N_17585,N_16517);
and U22137 (N_22137,N_17842,N_12182);
or U22138 (N_22138,N_12333,N_12800);
xnor U22139 (N_22139,N_19346,N_10186);
and U22140 (N_22140,N_13477,N_16205);
nor U22141 (N_22141,N_12732,N_18674);
nor U22142 (N_22142,N_12228,N_16806);
nand U22143 (N_22143,N_13060,N_10159);
xor U22144 (N_22144,N_16397,N_16901);
nor U22145 (N_22145,N_17949,N_15703);
and U22146 (N_22146,N_16073,N_19942);
nor U22147 (N_22147,N_17571,N_15871);
and U22148 (N_22148,N_17331,N_15519);
xor U22149 (N_22149,N_13031,N_19748);
or U22150 (N_22150,N_10315,N_11763);
nand U22151 (N_22151,N_12317,N_10384);
nand U22152 (N_22152,N_18998,N_19581);
xor U22153 (N_22153,N_18095,N_19843);
and U22154 (N_22154,N_18441,N_12077);
or U22155 (N_22155,N_19452,N_11856);
nand U22156 (N_22156,N_17548,N_11424);
and U22157 (N_22157,N_17854,N_11390);
nand U22158 (N_22158,N_18692,N_10820);
nor U22159 (N_22159,N_11976,N_12703);
nand U22160 (N_22160,N_14270,N_13390);
nand U22161 (N_22161,N_13169,N_15484);
and U22162 (N_22162,N_10576,N_11143);
xnor U22163 (N_22163,N_14062,N_11008);
xnor U22164 (N_22164,N_17655,N_13713);
or U22165 (N_22165,N_15385,N_11389);
nor U22166 (N_22166,N_11022,N_10427);
nor U22167 (N_22167,N_12009,N_18478);
nor U22168 (N_22168,N_10699,N_12645);
and U22169 (N_22169,N_19668,N_16913);
and U22170 (N_22170,N_18911,N_16331);
nand U22171 (N_22171,N_12256,N_11279);
nand U22172 (N_22172,N_16202,N_11627);
nand U22173 (N_22173,N_19460,N_19638);
nor U22174 (N_22174,N_19550,N_11980);
and U22175 (N_22175,N_16550,N_13959);
nand U22176 (N_22176,N_13509,N_14307);
and U22177 (N_22177,N_14998,N_13436);
and U22178 (N_22178,N_15789,N_17533);
or U22179 (N_22179,N_11996,N_18671);
and U22180 (N_22180,N_11906,N_17644);
nand U22181 (N_22181,N_11385,N_12286);
nor U22182 (N_22182,N_16903,N_10107);
or U22183 (N_22183,N_14563,N_16230);
and U22184 (N_22184,N_16385,N_14542);
nor U22185 (N_22185,N_10754,N_14770);
and U22186 (N_22186,N_10708,N_17283);
nand U22187 (N_22187,N_17940,N_18961);
nor U22188 (N_22188,N_18676,N_17959);
and U22189 (N_22189,N_19560,N_16817);
and U22190 (N_22190,N_14745,N_16313);
and U22191 (N_22191,N_12743,N_11689);
and U22192 (N_22192,N_15200,N_12118);
nand U22193 (N_22193,N_18905,N_15130);
nor U22194 (N_22194,N_15879,N_14028);
or U22195 (N_22195,N_13557,N_10811);
xnor U22196 (N_22196,N_12959,N_12345);
xnor U22197 (N_22197,N_12099,N_17691);
and U22198 (N_22198,N_18594,N_14055);
or U22199 (N_22199,N_18346,N_11483);
nor U22200 (N_22200,N_11357,N_11978);
and U22201 (N_22201,N_10177,N_16737);
or U22202 (N_22202,N_15277,N_19138);
xor U22203 (N_22203,N_18810,N_13270);
or U22204 (N_22204,N_13372,N_13278);
and U22205 (N_22205,N_19717,N_16729);
nand U22206 (N_22206,N_19777,N_17697);
nor U22207 (N_22207,N_15907,N_13877);
nor U22208 (N_22208,N_14638,N_18981);
or U22209 (N_22209,N_17213,N_15290);
xor U22210 (N_22210,N_12411,N_13360);
and U22211 (N_22211,N_18808,N_16877);
nand U22212 (N_22212,N_10439,N_15728);
or U22213 (N_22213,N_14877,N_19997);
nand U22214 (N_22214,N_13409,N_10851);
xnor U22215 (N_22215,N_12421,N_17048);
xor U22216 (N_22216,N_13362,N_15528);
nand U22217 (N_22217,N_13589,N_15866);
nor U22218 (N_22218,N_16372,N_16064);
or U22219 (N_22219,N_13489,N_18063);
xnor U22220 (N_22220,N_11910,N_13867);
nand U22221 (N_22221,N_14970,N_19457);
xnor U22222 (N_22222,N_19659,N_19544);
and U22223 (N_22223,N_18499,N_17746);
and U22224 (N_22224,N_17095,N_17720);
nand U22225 (N_22225,N_12661,N_14787);
and U22226 (N_22226,N_11089,N_11137);
or U22227 (N_22227,N_15718,N_18473);
nor U22228 (N_22228,N_13513,N_13337);
or U22229 (N_22229,N_12640,N_10453);
or U22230 (N_22230,N_12966,N_14526);
and U22231 (N_22231,N_15410,N_18793);
or U22232 (N_22232,N_11436,N_15072);
or U22233 (N_22233,N_18072,N_16270);
nor U22234 (N_22234,N_19931,N_10929);
nand U22235 (N_22235,N_16675,N_11628);
and U22236 (N_22236,N_19868,N_16091);
nand U22237 (N_22237,N_13905,N_14243);
xnor U22238 (N_22238,N_19820,N_11687);
nand U22239 (N_22239,N_10774,N_17592);
or U22240 (N_22240,N_17759,N_11975);
nand U22241 (N_22241,N_16948,N_15226);
or U22242 (N_22242,N_19608,N_13515);
and U22243 (N_22243,N_18935,N_17897);
xnor U22244 (N_22244,N_11778,N_18309);
nor U22245 (N_22245,N_16590,N_19307);
and U22246 (N_22246,N_11957,N_16968);
or U22247 (N_22247,N_12363,N_19718);
and U22248 (N_22248,N_18848,N_18612);
and U22249 (N_22249,N_13644,N_12381);
nand U22250 (N_22250,N_12161,N_18347);
nand U22251 (N_22251,N_16666,N_15681);
nor U22252 (N_22252,N_17907,N_15367);
or U22253 (N_22253,N_13048,N_15748);
nand U22254 (N_22254,N_13137,N_18131);
nor U22255 (N_22255,N_14978,N_17955);
and U22256 (N_22256,N_10996,N_11226);
or U22257 (N_22257,N_16117,N_10116);
nand U22258 (N_22258,N_15195,N_14225);
nand U22259 (N_22259,N_12384,N_11615);
nand U22260 (N_22260,N_18111,N_10295);
nor U22261 (N_22261,N_10718,N_13677);
or U22262 (N_22262,N_12839,N_11162);
nand U22263 (N_22263,N_18647,N_12998);
xor U22264 (N_22264,N_17407,N_17591);
or U22265 (N_22265,N_14284,N_10939);
nor U22266 (N_22266,N_10365,N_12240);
nor U22267 (N_22267,N_12920,N_13853);
or U22268 (N_22268,N_12864,N_12078);
nand U22269 (N_22269,N_14673,N_13649);
nand U22270 (N_22270,N_14884,N_19224);
nor U22271 (N_22271,N_19416,N_11049);
nor U22272 (N_22272,N_11523,N_19665);
nor U22273 (N_22273,N_17758,N_19141);
or U22274 (N_22274,N_11849,N_17106);
or U22275 (N_22275,N_12194,N_18982);
nand U22276 (N_22276,N_11417,N_17220);
nand U22277 (N_22277,N_18228,N_12300);
nor U22278 (N_22278,N_19556,N_11029);
or U22279 (N_22279,N_16970,N_12343);
nand U22280 (N_22280,N_17942,N_15845);
nor U22281 (N_22281,N_11611,N_19596);
nor U22282 (N_22282,N_12767,N_15027);
nor U22283 (N_22283,N_12997,N_10965);
and U22284 (N_22284,N_13407,N_18354);
nand U22285 (N_22285,N_18335,N_12229);
or U22286 (N_22286,N_10060,N_15645);
and U22287 (N_22287,N_14506,N_16228);
nand U22288 (N_22288,N_19594,N_13440);
nand U22289 (N_22289,N_10086,N_13544);
or U22290 (N_22290,N_14731,N_12658);
nor U22291 (N_22291,N_10990,N_10480);
and U22292 (N_22292,N_13263,N_14532);
and U22293 (N_22293,N_11727,N_14906);
nor U22294 (N_22294,N_10976,N_15771);
nor U22295 (N_22295,N_16942,N_19201);
or U22296 (N_22296,N_18706,N_11148);
nand U22297 (N_22297,N_12924,N_14288);
nand U22298 (N_22298,N_16272,N_14792);
nand U22299 (N_22299,N_11165,N_10706);
and U22300 (N_22300,N_11036,N_10953);
or U22301 (N_22301,N_11208,N_17243);
or U22302 (N_22302,N_10395,N_18854);
and U22303 (N_22303,N_18931,N_10320);
and U22304 (N_22304,N_18711,N_12931);
nor U22305 (N_22305,N_15161,N_18764);
nand U22306 (N_22306,N_15387,N_15937);
or U22307 (N_22307,N_11716,N_18997);
and U22308 (N_22308,N_11543,N_10424);
and U22309 (N_22309,N_19602,N_14279);
nand U22310 (N_22310,N_14566,N_19109);
nand U22311 (N_22311,N_15576,N_17612);
xnor U22312 (N_22312,N_16306,N_14227);
nand U22313 (N_22313,N_15053,N_16611);
and U22314 (N_22314,N_11703,N_18165);
or U22315 (N_22315,N_11738,N_15430);
or U22316 (N_22316,N_12954,N_14676);
and U22317 (N_22317,N_12904,N_10334);
nor U22318 (N_22318,N_16386,N_19759);
or U22319 (N_22319,N_14576,N_18088);
and U22320 (N_22320,N_16899,N_12978);
or U22321 (N_22321,N_11770,N_14472);
nor U22322 (N_22322,N_15370,N_16389);
nor U22323 (N_22323,N_19578,N_19043);
nand U22324 (N_22324,N_12210,N_16616);
nand U22325 (N_22325,N_13346,N_15882);
and U22326 (N_22326,N_13188,N_18765);
nor U22327 (N_22327,N_17589,N_11068);
nand U22328 (N_22328,N_13804,N_18773);
nor U22329 (N_22329,N_19271,N_19673);
nor U22330 (N_22330,N_10379,N_15960);
or U22331 (N_22331,N_15322,N_11977);
nor U22332 (N_22332,N_17143,N_15650);
nand U22333 (N_22333,N_16024,N_15268);
or U22334 (N_22334,N_12714,N_11188);
or U22335 (N_22335,N_15674,N_10298);
nor U22336 (N_22336,N_19839,N_10975);
and U22337 (N_22337,N_13965,N_11453);
nand U22338 (N_22338,N_13566,N_11280);
nor U22339 (N_22339,N_10343,N_11261);
and U22340 (N_22340,N_12715,N_10744);
and U22341 (N_22341,N_10477,N_17322);
nand U22342 (N_22342,N_12579,N_17350);
and U22343 (N_22343,N_18758,N_12434);
nor U22344 (N_22344,N_15078,N_14296);
and U22345 (N_22345,N_17356,N_14012);
nor U22346 (N_22346,N_16880,N_11621);
nand U22347 (N_22347,N_13900,N_19625);
nand U22348 (N_22348,N_15925,N_15582);
nand U22349 (N_22349,N_16858,N_19597);
and U22350 (N_22350,N_13487,N_11514);
nand U22351 (N_22351,N_15345,N_13377);
and U22352 (N_22352,N_10632,N_16597);
or U22353 (N_22353,N_11857,N_16426);
xnor U22354 (N_22354,N_19260,N_15135);
or U22355 (N_22355,N_17974,N_13400);
xnor U22356 (N_22356,N_14949,N_16197);
nor U22357 (N_22357,N_12771,N_19778);
nand U22358 (N_22358,N_16610,N_18511);
and U22359 (N_22359,N_12739,N_10786);
nand U22360 (N_22360,N_15250,N_14029);
nor U22361 (N_22361,N_17352,N_12215);
nand U22362 (N_22362,N_19790,N_12464);
nor U22363 (N_22363,N_12949,N_17257);
xor U22364 (N_22364,N_18103,N_17695);
or U22365 (N_22365,N_19151,N_11487);
or U22366 (N_22366,N_11032,N_19067);
and U22367 (N_22367,N_11456,N_12061);
nor U22368 (N_22368,N_15743,N_19973);
nand U22369 (N_22369,N_13768,N_16412);
and U22370 (N_22370,N_10350,N_14756);
and U22371 (N_22371,N_13857,N_15742);
nor U22372 (N_22372,N_18272,N_11418);
nor U22373 (N_22373,N_18469,N_10145);
and U22374 (N_22374,N_19650,N_11731);
nor U22375 (N_22375,N_18816,N_17727);
nand U22376 (N_22376,N_11823,N_19696);
and U22377 (N_22377,N_18146,N_19480);
or U22378 (N_22378,N_17102,N_18090);
nor U22379 (N_22379,N_13017,N_11120);
and U22380 (N_22380,N_14935,N_18844);
nor U22381 (N_22381,N_13172,N_19980);
nor U22382 (N_22382,N_19789,N_11560);
nor U22383 (N_22383,N_13308,N_10673);
nand U22384 (N_22384,N_13684,N_13533);
or U22385 (N_22385,N_15525,N_19816);
nand U22386 (N_22386,N_14127,N_15235);
or U22387 (N_22387,N_12491,N_11926);
and U22388 (N_22388,N_14577,N_13868);
or U22389 (N_22389,N_13295,N_17738);
or U22390 (N_22390,N_15905,N_12014);
and U22391 (N_22391,N_11263,N_16707);
nor U22392 (N_22392,N_11230,N_14535);
nor U22393 (N_22393,N_15899,N_19780);
nand U22394 (N_22394,N_15847,N_13646);
nand U22395 (N_22395,N_12088,N_17918);
nand U22396 (N_22396,N_18861,N_17590);
nor U22397 (N_22397,N_18059,N_15933);
nor U22398 (N_22398,N_19348,N_12606);
nor U22399 (N_22399,N_13160,N_10037);
nor U22400 (N_22400,N_12396,N_12486);
nand U22401 (N_22401,N_16779,N_15397);
nand U22402 (N_22402,N_12220,N_18805);
nor U22403 (N_22403,N_17080,N_10003);
nand U22404 (N_22404,N_18303,N_13190);
or U22405 (N_22405,N_11740,N_14331);
nand U22406 (N_22406,N_14358,N_15725);
and U22407 (N_22407,N_10983,N_13688);
nand U22408 (N_22408,N_18160,N_14635);
and U22409 (N_22409,N_17663,N_19442);
nor U22410 (N_22410,N_16679,N_13617);
xnor U22411 (N_22411,N_10333,N_11439);
and U22412 (N_22412,N_13434,N_15704);
or U22413 (N_22413,N_19970,N_16608);
xnor U22414 (N_22414,N_14389,N_14807);
or U22415 (N_22415,N_19061,N_11081);
or U22416 (N_22416,N_13135,N_10020);
or U22417 (N_22417,N_17846,N_11466);
nor U22418 (N_22418,N_10045,N_16201);
nand U22419 (N_22419,N_18082,N_12862);
or U22420 (N_22420,N_11883,N_19425);
or U22421 (N_22421,N_12865,N_19709);
nor U22422 (N_22422,N_12831,N_15107);
or U22423 (N_22423,N_11979,N_16021);
nor U22424 (N_22424,N_16682,N_16914);
nor U22425 (N_22425,N_17760,N_10476);
or U22426 (N_22426,N_17135,N_17595);
or U22427 (N_22427,N_12745,N_19121);
or U22428 (N_22428,N_15215,N_17315);
or U22429 (N_22429,N_10238,N_15740);
nor U22430 (N_22430,N_11444,N_19073);
or U22431 (N_22431,N_12834,N_12122);
nor U22432 (N_22432,N_19830,N_13975);
or U22433 (N_22433,N_16678,N_16995);
nor U22434 (N_22434,N_15750,N_16061);
nand U22435 (N_22435,N_10773,N_17017);
xor U22436 (N_22436,N_18504,N_14320);
or U22437 (N_22437,N_11121,N_14319);
nor U22438 (N_22438,N_13204,N_10499);
and U22439 (N_22439,N_18672,N_13901);
nor U22440 (N_22440,N_17965,N_16887);
or U22441 (N_22441,N_18325,N_19240);
and U22442 (N_22442,N_17900,N_16317);
or U22443 (N_22443,N_14753,N_15455);
or U22444 (N_22444,N_12023,N_11154);
or U22445 (N_22445,N_14771,N_18223);
or U22446 (N_22446,N_19826,N_18602);
or U22447 (N_22447,N_12969,N_10810);
and U22448 (N_22448,N_15671,N_12166);
xor U22449 (N_22449,N_10096,N_19215);
nor U22450 (N_22450,N_12700,N_17441);
nor U22451 (N_22451,N_14501,N_15642);
and U22452 (N_22452,N_12975,N_14064);
nand U22453 (N_22453,N_17357,N_12940);
nand U22454 (N_22454,N_16456,N_18688);
or U22455 (N_22455,N_17740,N_17162);
nand U22456 (N_22456,N_10040,N_10936);
nor U22457 (N_22457,N_16286,N_13052);
xor U22458 (N_22458,N_18890,N_19142);
or U22459 (N_22459,N_16078,N_14207);
and U22460 (N_22460,N_13310,N_19419);
xnor U22461 (N_22461,N_12994,N_19832);
or U22462 (N_22462,N_18508,N_16266);
and U22463 (N_22463,N_11718,N_14340);
and U22464 (N_22464,N_16615,N_15362);
and U22465 (N_22465,N_13776,N_19887);
nand U22466 (N_22466,N_10259,N_19807);
and U22467 (N_22467,N_11733,N_17112);
and U22468 (N_22468,N_13601,N_18198);
and U22469 (N_22469,N_11228,N_17049);
xor U22470 (N_22470,N_12517,N_12972);
nor U22471 (N_22471,N_16940,N_17559);
and U22472 (N_22472,N_15275,N_10276);
or U22473 (N_22473,N_16250,N_10899);
nand U22474 (N_22474,N_19316,N_16870);
nand U22475 (N_22475,N_13078,N_13220);
or U22476 (N_22476,N_11991,N_17679);
and U22477 (N_22477,N_16076,N_18583);
nand U22478 (N_22478,N_13292,N_13343);
nand U22479 (N_22479,N_14538,N_18324);
or U22480 (N_22480,N_12513,N_15348);
nor U22481 (N_22481,N_14766,N_16507);
nand U22482 (N_22482,N_13521,N_15700);
and U22483 (N_22483,N_13598,N_10856);
and U22484 (N_22484,N_11640,N_14774);
nand U22485 (N_22485,N_18104,N_14033);
nor U22486 (N_22486,N_18614,N_10200);
and U22487 (N_22487,N_13961,N_18439);
or U22488 (N_22488,N_17368,N_18222);
nor U22489 (N_22489,N_15543,N_18771);
and U22490 (N_22490,N_16563,N_18502);
xor U22491 (N_22491,N_17793,N_16592);
nand U22492 (N_22492,N_11334,N_10686);
nor U22493 (N_22493,N_13685,N_15022);
nand U22494 (N_22494,N_17719,N_12105);
and U22495 (N_22495,N_13943,N_14655);
or U22496 (N_22496,N_10989,N_11913);
nor U22497 (N_22497,N_19630,N_10891);
and U22498 (N_22498,N_12514,N_16072);
xnor U22499 (N_22499,N_10538,N_11092);
or U22500 (N_22500,N_16403,N_16542);
nand U22501 (N_22501,N_17233,N_11854);
or U22502 (N_22502,N_19891,N_10544);
or U22503 (N_22503,N_15031,N_16213);
xnor U22504 (N_22504,N_11023,N_18660);
xor U22505 (N_22505,N_19595,N_17270);
xnor U22506 (N_22506,N_13666,N_13174);
and U22507 (N_22507,N_13194,N_13506);
nand U22508 (N_22508,N_18125,N_13134);
and U22509 (N_22509,N_17311,N_13085);
nor U22510 (N_22510,N_14602,N_11363);
nand U22511 (N_22511,N_15131,N_16516);
nor U22512 (N_22512,N_13098,N_14350);
xnor U22513 (N_22513,N_18875,N_19488);
or U22514 (N_22514,N_11382,N_14395);
and U22515 (N_22515,N_15024,N_19745);
nor U22516 (N_22516,N_11760,N_11533);
nand U22517 (N_22517,N_17267,N_13120);
nor U22518 (N_22518,N_10795,N_13065);
and U22519 (N_22519,N_10646,N_15328);
nor U22520 (N_22520,N_14159,N_11138);
nand U22521 (N_22521,N_14242,N_13754);
nor U22522 (N_22522,N_18390,N_19492);
and U22523 (N_22523,N_10948,N_15313);
nor U22524 (N_22524,N_11146,N_19011);
xnor U22525 (N_22525,N_12185,N_19453);
nand U22526 (N_22526,N_13954,N_11485);
xor U22527 (N_22527,N_18190,N_18568);
nand U22528 (N_22528,N_11907,N_17511);
xnor U22529 (N_22529,N_13211,N_10346);
nand U22530 (N_22530,N_19553,N_11872);
nor U22531 (N_22531,N_12765,N_10136);
or U22532 (N_22532,N_12788,N_12447);
and U22533 (N_22533,N_18151,N_11939);
and U22534 (N_22534,N_18107,N_19838);
nand U22535 (N_22535,N_15395,N_18399);
nor U22536 (N_22536,N_14733,N_12692);
nor U22537 (N_22537,N_18446,N_12117);
nand U22538 (N_22538,N_16328,N_11227);
or U22539 (N_22539,N_11045,N_11132);
and U22540 (N_22540,N_12457,N_13013);
nor U22541 (N_22541,N_16888,N_14438);
and U22542 (N_22542,N_15969,N_12520);
nand U22543 (N_22543,N_13059,N_19057);
nor U22544 (N_22544,N_11590,N_19100);
nor U22545 (N_22545,N_18636,N_15076);
nor U22546 (N_22546,N_15421,N_13540);
nor U22547 (N_22547,N_10234,N_19521);
and U22548 (N_22548,N_16580,N_14984);
xor U22549 (N_22549,N_14641,N_15077);
nand U22550 (N_22550,N_14321,N_16515);
nand U22551 (N_22551,N_15788,N_11824);
or U22552 (N_22552,N_13520,N_12620);
xnor U22553 (N_22553,N_10110,N_13742);
nand U22554 (N_22554,N_12727,N_12071);
or U22555 (N_22555,N_11017,N_19666);
nor U22556 (N_22556,N_16673,N_14394);
xor U22557 (N_22557,N_15705,N_16185);
or U22558 (N_22558,N_10299,N_15489);
and U22559 (N_22559,N_10496,N_10047);
nor U22560 (N_22560,N_10926,N_15855);
nor U22561 (N_22561,N_13182,N_18029);
xor U22562 (N_22562,N_17880,N_16769);
nor U22563 (N_22563,N_19757,N_15041);
nor U22564 (N_22564,N_19264,N_13358);
and U22565 (N_22565,N_19985,N_18194);
nand U22566 (N_22566,N_18253,N_11395);
or U22567 (N_22567,N_17633,N_15901);
and U22568 (N_22568,N_14681,N_19809);
and U22569 (N_22569,N_12056,N_14975);
nor U22570 (N_22570,N_18404,N_11670);
nand U22571 (N_22571,N_10273,N_18643);
and U22572 (N_22572,N_16595,N_18149);
xor U22573 (N_22573,N_19999,N_13184);
or U22574 (N_22574,N_17105,N_11710);
and U22575 (N_22575,N_18732,N_14415);
and U22576 (N_22576,N_18642,N_13221);
or U22577 (N_22577,N_15352,N_11426);
or U22578 (N_22578,N_17010,N_14132);
nand U22579 (N_22579,N_10147,N_11495);
nand U22580 (N_22580,N_16945,N_13291);
nand U22581 (N_22581,N_14294,N_10459);
and U22582 (N_22582,N_10394,N_13848);
or U22583 (N_22583,N_18080,N_17133);
nand U22584 (N_22584,N_15067,N_10444);
and U22585 (N_22585,N_12988,N_18415);
nor U22586 (N_22586,N_10870,N_11705);
xor U22587 (N_22587,N_13088,N_10261);
and U22588 (N_22588,N_15555,N_16274);
nand U22589 (N_22589,N_18621,N_19331);
nand U22590 (N_22590,N_19306,N_18118);
nand U22591 (N_22591,N_13528,N_13222);
nor U22592 (N_22592,N_16524,N_18250);
and U22593 (N_22593,N_12689,N_13063);
nand U22594 (N_22594,N_12537,N_19476);
or U22595 (N_22595,N_17218,N_19045);
or U22596 (N_22596,N_10890,N_11026);
or U22597 (N_22597,N_13631,N_14982);
and U22598 (N_22598,N_11546,N_11020);
and U22599 (N_22599,N_10130,N_10818);
and U22600 (N_22600,N_15081,N_10097);
xnor U22601 (N_22601,N_12437,N_19849);
or U22602 (N_22602,N_13245,N_18941);
and U22603 (N_22603,N_12410,N_15767);
nand U22604 (N_22604,N_17498,N_11782);
or U22605 (N_22605,N_10068,N_18960);
nand U22606 (N_22606,N_18306,N_15690);
or U22607 (N_22607,N_17905,N_16351);
or U22608 (N_22608,N_16878,N_12849);
and U22609 (N_22609,N_15075,N_15493);
xnor U22610 (N_22610,N_18460,N_18726);
nor U22611 (N_22611,N_14464,N_19994);
xnor U22612 (N_22612,N_12843,N_17901);
nor U22613 (N_22613,N_11708,N_14197);
xor U22614 (N_22614,N_19756,N_12809);
and U22615 (N_22615,N_11891,N_11490);
and U22616 (N_22616,N_17724,N_18037);
nand U22617 (N_22617,N_11186,N_11380);
xor U22618 (N_22618,N_11928,N_13861);
and U22619 (N_22619,N_14537,N_10724);
and U22620 (N_22620,N_11106,N_12227);
or U22621 (N_22621,N_14624,N_16042);
and U22622 (N_22622,N_16163,N_19944);
or U22623 (N_22623,N_16635,N_10195);
nor U22624 (N_22624,N_16932,N_12679);
xnor U22625 (N_22625,N_12218,N_13918);
nor U22626 (N_22626,N_16777,N_13109);
or U22627 (N_22627,N_10668,N_15291);
or U22628 (N_22628,N_10759,N_13233);
or U22629 (N_22629,N_14073,N_11376);
or U22630 (N_22630,N_14128,N_16837);
and U22631 (N_22631,N_12067,N_15213);
nor U22632 (N_22632,N_12995,N_17186);
or U22633 (N_22633,N_18367,N_10883);
nand U22634 (N_22634,N_13378,N_14999);
nor U22635 (N_22635,N_11431,N_19351);
nand U22636 (N_22636,N_18102,N_14286);
or U22637 (N_22637,N_19191,N_17935);
or U22638 (N_22638,N_13734,N_17482);
nor U22639 (N_22639,N_11646,N_12496);
nand U22640 (N_22640,N_18293,N_17381);
or U22641 (N_22641,N_10896,N_16394);
and U22642 (N_22642,N_19036,N_10586);
nand U22643 (N_22643,N_19210,N_17256);
nand U22644 (N_22644,N_18516,N_17090);
or U22645 (N_22645,N_14091,N_11104);
and U22646 (N_22646,N_12894,N_18300);
or U22647 (N_22647,N_13749,N_18069);
nand U22648 (N_22648,N_16978,N_12477);
nor U22649 (N_22649,N_18119,N_12946);
or U22650 (N_22650,N_10755,N_14636);
nand U22651 (N_22651,N_16944,N_19764);
or U22652 (N_22652,N_19817,N_13674);
nor U22653 (N_22653,N_13056,N_17792);
nand U22654 (N_22654,N_10036,N_15118);
or U22655 (N_22655,N_12618,N_11720);
or U22656 (N_22656,N_15708,N_17507);
nor U22657 (N_22657,N_10839,N_13750);
nand U22658 (N_22658,N_12399,N_14166);
nor U22659 (N_22659,N_19434,N_15128);
nand U22660 (N_22660,N_19246,N_14192);
nor U22661 (N_22661,N_19721,N_15634);
or U22662 (N_22662,N_15240,N_14386);
or U22663 (N_22663,N_15202,N_11749);
or U22664 (N_22664,N_17200,N_12622);
and U22665 (N_22665,N_13545,N_13563);
xnor U22666 (N_22666,N_11559,N_19781);
nand U22667 (N_22667,N_17418,N_10342);
nor U22668 (N_22668,N_14376,N_18147);
nand U22669 (N_22669,N_16471,N_17179);
or U22670 (N_22670,N_13572,N_10559);
or U22671 (N_22671,N_10909,N_11364);
and U22672 (N_22672,N_16477,N_15877);
or U22673 (N_22673,N_15459,N_11730);
nor U22674 (N_22674,N_10537,N_19535);
nand U22675 (N_22675,N_16664,N_12361);
and U22676 (N_22676,N_10209,N_13623);
and U22677 (N_22677,N_18348,N_10539);
or U22678 (N_22678,N_15252,N_19916);
nor U22679 (N_22679,N_16917,N_16284);
nor U22680 (N_22680,N_11630,N_19124);
nand U22681 (N_22681,N_16483,N_19144);
or U22682 (N_22682,N_11236,N_13711);
xnor U22683 (N_22683,N_12690,N_15803);
nand U22684 (N_22684,N_11986,N_16231);
and U22685 (N_22685,N_15732,N_12471);
and U22686 (N_22686,N_14440,N_16440);
nand U22687 (N_22687,N_15403,N_14040);
nor U22688 (N_22688,N_17914,N_17026);
and U22689 (N_22689,N_18483,N_11354);
or U22690 (N_22690,N_14462,N_15008);
nor U22691 (N_22691,N_16199,N_10647);
and U22692 (N_22692,N_13686,N_18896);
nor U22693 (N_22693,N_13446,N_15720);
nor U22694 (N_22694,N_13663,N_11714);
and U22695 (N_22695,N_15662,N_12039);
xor U22696 (N_22696,N_14909,N_14625);
nand U22697 (N_22697,N_18649,N_14841);
nor U22698 (N_22698,N_18546,N_15565);
or U22699 (N_22699,N_16143,N_11608);
and U22700 (N_22700,N_16475,N_15184);
nand U22701 (N_22701,N_11331,N_16366);
xnor U22702 (N_22702,N_13051,N_18089);
nand U22703 (N_22703,N_16631,N_16898);
and U22704 (N_22704,N_15480,N_14724);
xor U22705 (N_22705,N_13588,N_10992);
and U22706 (N_22706,N_10171,N_17079);
or U22707 (N_22707,N_11033,N_14924);
nor U22708 (N_22708,N_15285,N_19276);
nor U22709 (N_22709,N_17658,N_10475);
or U22710 (N_22710,N_12535,N_12427);
xor U22711 (N_22711,N_10122,N_11007);
nand U22712 (N_22712,N_13981,N_16718);
or U22713 (N_22713,N_16125,N_17122);
and U22714 (N_22714,N_10019,N_12458);
nor U22715 (N_22715,N_16034,N_16559);
or U22716 (N_22716,N_14125,N_18909);
or U22717 (N_22717,N_17887,N_18040);
nand U22718 (N_22718,N_15332,N_18995);
nor U22719 (N_22719,N_16472,N_17947);
nand U22720 (N_22720,N_13036,N_16734);
nor U22721 (N_22721,N_16612,N_13670);
and U22722 (N_22722,N_13780,N_16177);
or U22723 (N_22723,N_13090,N_19330);
or U22724 (N_22724,N_17535,N_15992);
nand U22725 (N_22725,N_16304,N_17181);
or U22726 (N_22726,N_11746,N_10535);
nor U22727 (N_22727,N_14672,N_15932);
nand U22728 (N_22728,N_19926,N_15983);
xor U22729 (N_22729,N_17465,N_17389);
nand U22730 (N_22730,N_10719,N_17908);
and U22731 (N_22731,N_18708,N_14905);
or U22732 (N_22732,N_12364,N_17582);
nand U22733 (N_22733,N_16308,N_19140);
nand U22734 (N_22734,N_13464,N_18975);
nand U22735 (N_22735,N_13156,N_11401);
nor U22736 (N_22736,N_13057,N_15265);
nor U22737 (N_22737,N_15955,N_18734);
nand U22738 (N_22738,N_12503,N_17833);
and U22739 (N_22739,N_11813,N_10915);
and U22740 (N_22740,N_15112,N_15589);
or U22741 (N_22741,N_16463,N_14252);
nor U22742 (N_22742,N_15218,N_12289);
and U22743 (N_22743,N_12353,N_16562);
and U22744 (N_22744,N_18697,N_12126);
xor U22745 (N_22745,N_11809,N_18481);
nor U22746 (N_22746,N_13450,N_14651);
xnor U22747 (N_22747,N_11931,N_18273);
and U22748 (N_22748,N_15316,N_16001);
xnor U22749 (N_22749,N_19456,N_19783);
nand U22750 (N_22750,N_12748,N_12807);
xor U22751 (N_22751,N_14916,N_14424);
nor U22752 (N_22752,N_11115,N_11316);
nor U22753 (N_22753,N_14346,N_15880);
xor U22754 (N_22754,N_11866,N_17113);
nand U22755 (N_22755,N_18550,N_15665);
nand U22756 (N_22756,N_16924,N_17879);
nor U22757 (N_22757,N_13878,N_10408);
nor U22758 (N_22758,N_17091,N_13201);
nand U22759 (N_22759,N_14968,N_11204);
xnor U22760 (N_22760,N_16691,N_17117);
nor U22761 (N_22761,N_11064,N_19383);
nand U22762 (N_22762,N_18683,N_17069);
xor U22763 (N_22763,N_10512,N_19349);
or U22764 (N_22764,N_16053,N_15366);
or U22765 (N_22765,N_10940,N_17334);
nor U22766 (N_22766,N_17848,N_19060);
or U22767 (N_22767,N_16501,N_10601);
nor U22768 (N_22768,N_16160,N_15211);
nand U22769 (N_22769,N_19791,N_12259);
nor U22770 (N_22770,N_18006,N_11676);
or U22771 (N_22771,N_12068,N_16890);
nand U22772 (N_22772,N_15689,N_10563);
nand U22773 (N_22773,N_14871,N_19206);
and U22774 (N_22774,N_14613,N_13413);
nand U22775 (N_22775,N_10423,N_15247);
xnor U22776 (N_22776,N_12938,N_18266);
nor U22777 (N_22777,N_12290,N_12498);
xor U22778 (N_22778,N_17781,N_17509);
nand U22779 (N_22779,N_11999,N_10741);
and U22780 (N_22780,N_15437,N_12611);
nand U22781 (N_22781,N_14521,N_11735);
nand U22782 (N_22782,N_13268,N_10684);
xor U22783 (N_22783,N_15276,N_11169);
nor U22784 (N_22784,N_13576,N_16618);
nand U22785 (N_22785,N_11551,N_17827);
xor U22786 (N_22786,N_17617,N_19239);
nor U22787 (N_22787,N_10352,N_16063);
nor U22788 (N_22788,N_14801,N_15699);
nor U22789 (N_22789,N_10113,N_16268);
nand U22790 (N_22790,N_13122,N_14414);
or U22791 (N_22791,N_12223,N_13208);
nand U22792 (N_22792,N_15326,N_12389);
nand U22793 (N_22793,N_16598,N_11071);
xor U22794 (N_22794,N_17289,N_14951);
nor U22795 (N_22795,N_17425,N_15575);
or U22796 (N_22796,N_16154,N_10281);
and U22797 (N_22797,N_15617,N_10126);
nor U22798 (N_22798,N_10998,N_11556);
nor U22799 (N_22799,N_14873,N_18094);
nand U22800 (N_22800,N_18085,N_10101);
nor U22801 (N_22801,N_14834,N_12564);
nor U22802 (N_22802,N_13571,N_19114);
or U22803 (N_22803,N_16709,N_19879);
nand U22804 (N_22804,N_10587,N_13494);
or U22805 (N_22805,N_12341,N_12102);
nand U22806 (N_22806,N_19308,N_12319);
and U22807 (N_22807,N_16111,N_12393);
nand U22808 (N_22808,N_13565,N_18239);
nand U22809 (N_22809,N_10215,N_16097);
nand U22810 (N_22810,N_10985,N_18926);
or U22811 (N_22811,N_12850,N_17885);
and U22812 (N_22812,N_18736,N_15123);
and U22813 (N_22813,N_12357,N_19566);
nor U22814 (N_22814,N_19267,N_10004);
nand U22815 (N_22815,N_11960,N_15280);
nand U22816 (N_22816,N_17953,N_18920);
nor U22817 (N_22817,N_17528,N_12342);
nand U22818 (N_22818,N_11085,N_17284);
nor U22819 (N_22819,N_14931,N_11679);
nand U22820 (N_22820,N_17008,N_13583);
and U22821 (N_22821,N_18313,N_16749);
nand U22822 (N_22822,N_18539,N_16982);
nor U22823 (N_22823,N_19451,N_15518);
nor U22824 (N_22824,N_15873,N_13100);
xnor U22825 (N_22825,N_12301,N_16299);
xnor U22826 (N_22826,N_14850,N_18557);
nor U22827 (N_22827,N_13305,N_11673);
and U22828 (N_22828,N_15279,N_12761);
nand U22829 (N_22829,N_14666,N_14088);
or U22830 (N_22830,N_11067,N_17598);
and U22831 (N_22831,N_16605,N_10618);
and U22832 (N_22832,N_12224,N_14275);
nand U22833 (N_22833,N_19148,N_19601);
and U22834 (N_22834,N_16280,N_11632);
and U22835 (N_22835,N_10916,N_19686);
or U22836 (N_22836,N_17302,N_15710);
or U22837 (N_22837,N_15605,N_11155);
nand U22838 (N_22838,N_14060,N_12652);
nor U22839 (N_22839,N_10071,N_11050);
or U22840 (N_22840,N_19162,N_14750);
nor U22841 (N_22841,N_14606,N_13001);
nor U22842 (N_22842,N_19950,N_15001);
nor U22843 (N_22843,N_10380,N_18496);
or U22844 (N_22844,N_15079,N_19183);
xor U22845 (N_22845,N_17012,N_19860);
and U22846 (N_22846,N_11629,N_13416);
and U22847 (N_22847,N_18289,N_10837);
or U22848 (N_22848,N_11593,N_10002);
nor U22849 (N_22849,N_12412,N_12041);
nor U22850 (N_22850,N_19266,N_10123);
or U22851 (N_22851,N_12011,N_10222);
and U22852 (N_22852,N_14234,N_18976);
nor U22853 (N_22853,N_11880,N_13635);
nand U22854 (N_22854,N_14831,N_19319);
nor U22855 (N_22855,N_18617,N_17681);
nand U22856 (N_22856,N_13338,N_17047);
or U22857 (N_22857,N_17208,N_17640);
and U22858 (N_22858,N_16644,N_10319);
nand U22859 (N_22859,N_16807,N_12089);
or U22860 (N_22860,N_12297,N_13896);
and U22861 (N_22861,N_10652,N_15267);
and U22862 (N_22862,N_15109,N_16141);
xor U22863 (N_22863,N_15448,N_13223);
and U22864 (N_22864,N_16341,N_14559);
and U22865 (N_22865,N_12325,N_16776);
or U22866 (N_22866,N_19955,N_19392);
or U22867 (N_22867,N_18606,N_16895);
nor U22868 (N_22868,N_16084,N_14705);
nand U22869 (N_22869,N_12906,N_14847);
and U22870 (N_22870,N_13296,N_10614);
and U22871 (N_22871,N_12871,N_13889);
nor U22872 (N_22872,N_10324,N_10703);
or U22873 (N_22873,N_17538,N_19619);
and U22874 (N_22874,N_17077,N_19541);
nand U22875 (N_22875,N_12619,N_16138);
nor U22876 (N_22876,N_14810,N_11281);
or U22877 (N_22877,N_12443,N_13186);
nand U22878 (N_22878,N_17447,N_18023);
or U22879 (N_22879,N_14534,N_14484);
nor U22880 (N_22880,N_16421,N_10980);
nor U22881 (N_22881,N_11794,N_16496);
or U22882 (N_22882,N_11938,N_14090);
and U22883 (N_22883,N_18722,N_14169);
or U22884 (N_22884,N_14883,N_16986);
and U22885 (N_22885,N_18877,N_11019);
and U22886 (N_22886,N_19324,N_11717);
nand U22887 (N_22887,N_14702,N_17646);
nor U22888 (N_22888,N_11810,N_15093);
nand U22889 (N_22889,N_13252,N_10462);
or U22890 (N_22890,N_10132,N_15203);
xor U22891 (N_22891,N_11501,N_16401);
and U22892 (N_22892,N_16764,N_14836);
nand U22893 (N_22893,N_19426,N_14882);
or U22894 (N_22894,N_14901,N_16660);
nand U22895 (N_22895,N_19387,N_15092);
or U22896 (N_22896,N_15157,N_12426);
and U22897 (N_22897,N_18387,N_13661);
and U22898 (N_22898,N_15944,N_19527);
nand U22899 (N_22899,N_13797,N_16927);
or U22900 (N_22900,N_13027,N_18440);
nand U22901 (N_22901,N_10415,N_13948);
or U22902 (N_22902,N_10460,N_19808);
nand U22903 (N_22903,N_14743,N_17234);
nand U22904 (N_22904,N_11338,N_17821);
and U22905 (N_22905,N_15636,N_12352);
and U22906 (N_22906,N_18248,N_11507);
nor U22907 (N_22907,N_14761,N_15133);
nor U22908 (N_22908,N_18276,N_13084);
nand U22909 (N_22909,N_11307,N_12020);
nor U22910 (N_22910,N_17613,N_14061);
and U22911 (N_22911,N_17456,N_15975);
nor U22912 (N_22912,N_13462,N_16183);
and U22913 (N_22913,N_10540,N_14369);
nor U22914 (N_22914,N_14263,N_19815);
or U22915 (N_22915,N_14487,N_12082);
xnor U22916 (N_22916,N_16656,N_11445);
and U22917 (N_22917,N_17728,N_16793);
nor U22918 (N_22918,N_11709,N_10602);
or U22919 (N_22919,N_19443,N_17747);
or U22920 (N_22920,N_17999,N_12856);
nand U22921 (N_22921,N_12852,N_13892);
nor U22922 (N_22922,N_10224,N_16684);
xor U22923 (N_22923,N_11779,N_18337);
and U22924 (N_22924,N_16093,N_15616);
nand U22925 (N_22925,N_16094,N_10599);
and U22926 (N_22926,N_12736,N_14044);
nor U22927 (N_22927,N_11951,N_11944);
and U22928 (N_22928,N_19763,N_14727);
nand U22929 (N_22929,N_16013,N_19406);
nand U22930 (N_22930,N_17787,N_16909);
nand U22931 (N_22931,N_14959,N_19066);
nand U22932 (N_22932,N_14165,N_15934);
nand U22933 (N_22933,N_12929,N_14133);
or U22934 (N_22934,N_16566,N_16797);
nand U22935 (N_22935,N_12928,N_10766);
xor U22936 (N_22936,N_11392,N_13537);
nand U22937 (N_22937,N_17630,N_14928);
or U22938 (N_22938,N_11579,N_16643);
and U22939 (N_22939,N_10701,N_19375);
and U22940 (N_22940,N_11177,N_14304);
xnor U22941 (N_22941,N_10293,N_12219);
nand U22942 (N_22942,N_14189,N_13458);
nand U22943 (N_22943,N_14820,N_18950);
and U22944 (N_22944,N_10566,N_13774);
nor U22945 (N_22945,N_16555,N_19669);
and U22946 (N_22946,N_15734,N_11732);
nor U22947 (N_22947,N_14180,N_15320);
nor U22948 (N_22948,N_10532,N_19547);
or U22949 (N_22949,N_16882,N_12418);
nor U22950 (N_22950,N_18959,N_18117);
nand U22951 (N_22951,N_15143,N_18837);
nor U22952 (N_22952,N_15471,N_19586);
nor U22953 (N_22953,N_19299,N_19784);
nor U22954 (N_22954,N_10908,N_15500);
nand U22955 (N_22955,N_19473,N_10794);
nor U22956 (N_22956,N_15641,N_10933);
nand U22957 (N_22957,N_16103,N_19616);
and U22958 (N_22958,N_15464,N_12677);
or U22959 (N_22959,N_11867,N_15768);
nor U22960 (N_22960,N_18525,N_18418);
nand U22961 (N_22961,N_12487,N_11997);
and U22962 (N_22962,N_13041,N_16115);
or U22963 (N_22963,N_19459,N_12670);
and U22964 (N_22964,N_13702,N_17003);
and U22965 (N_22965,N_15323,N_15965);
nor U22966 (N_22966,N_12246,N_10402);
and U22967 (N_22967,N_15860,N_18623);
nor U22968 (N_22968,N_15913,N_15709);
or U22969 (N_22969,N_17168,N_16599);
nor U22970 (N_22970,N_18205,N_18456);
or U22971 (N_22971,N_11010,N_16557);
nand U22972 (N_22972,N_18134,N_16732);
and U22973 (N_22973,N_17518,N_12808);
nor U22974 (N_22974,N_13082,N_14558);
and U22975 (N_22975,N_15124,N_16010);
xnor U22976 (N_22976,N_16083,N_13047);
and U22977 (N_22977,N_12241,N_18109);
nor U22978 (N_22978,N_15727,N_10470);
nand U22979 (N_22979,N_12320,N_11131);
and U22980 (N_22980,N_17847,N_15045);
and U22981 (N_22981,N_14355,N_11465);
and U22982 (N_22982,N_19767,N_17919);
nand U22983 (N_22983,N_14423,N_18373);
nor U22984 (N_22984,N_14646,N_11671);
and U22985 (N_22985,N_17016,N_14720);
or U22986 (N_22986,N_12095,N_19636);
nor U22987 (N_22987,N_11830,N_12720);
nand U22988 (N_22988,N_15117,N_17451);
nor U22989 (N_22989,N_11245,N_12268);
xor U22990 (N_22990,N_16556,N_15340);
nor U22991 (N_22991,N_18871,N_17812);
nand U22992 (N_22992,N_15098,N_16869);
nand U22993 (N_22993,N_14297,N_13320);
nor U22994 (N_22994,N_14375,N_14868);
nand U22995 (N_22995,N_18091,N_14708);
or U22996 (N_22996,N_10336,N_13326);
nor U22997 (N_22997,N_12844,N_13341);
or U22998 (N_22998,N_16322,N_15085);
nand U22999 (N_22999,N_11945,N_13812);
or U23000 (N_23000,N_11950,N_14274);
or U23001 (N_23001,N_13823,N_19963);
and U23002 (N_23002,N_15274,N_13009);
nor U23003 (N_23003,N_11765,N_19091);
and U23004 (N_23004,N_16639,N_10294);
nand U23005 (N_23005,N_14758,N_17579);
and U23006 (N_23006,N_13836,N_13375);
nand U23007 (N_23007,N_14237,N_19027);
and U23008 (N_23008,N_10058,N_18753);
nand U23009 (N_23009,N_19771,N_15099);
or U23010 (N_23010,N_17813,N_15569);
nor U23011 (N_23011,N_14273,N_15923);
nor U23012 (N_23012,N_14162,N_18828);
nand U23013 (N_23013,N_19296,N_15887);
nand U23014 (N_23014,N_13657,N_12012);
nand U23015 (N_23015,N_15916,N_17121);
and U23016 (N_23016,N_16062,N_14554);
xor U23017 (N_23017,N_16701,N_16640);
or U23018 (N_23018,N_19390,N_12918);
or U23019 (N_23019,N_18178,N_15425);
nand U23020 (N_23020,N_10968,N_12414);
nor U23021 (N_23021,N_18361,N_16714);
nand U23022 (N_23022,N_16242,N_19179);
or U23023 (N_23023,N_19372,N_16868);
and U23024 (N_23024,N_18292,N_14385);
or U23025 (N_23025,N_19159,N_18919);
and U23026 (N_23026,N_19489,N_19570);
and U23027 (N_23027,N_15782,N_14143);
nor U23028 (N_23028,N_13923,N_10061);
nor U23029 (N_23029,N_11949,N_18989);
xnor U23030 (N_23030,N_12460,N_12355);
xor U23031 (N_23031,N_18402,N_14442);
nor U23032 (N_23032,N_17430,N_14988);
or U23033 (N_23033,N_13410,N_16243);
xor U23034 (N_23034,N_17725,N_17250);
nor U23035 (N_23035,N_18954,N_10683);
nand U23036 (N_23036,N_14194,N_13526);
or U23037 (N_23037,N_12208,N_16416);
nand U23038 (N_23038,N_16296,N_12884);
nor U23039 (N_23039,N_17964,N_14528);
nand U23040 (N_23040,N_10375,N_18967);
and U23041 (N_23041,N_10035,N_10670);
nand U23042 (N_23042,N_12660,N_13813);
nand U23043 (N_23043,N_16965,N_15606);
xnor U23044 (N_23044,N_10638,N_14170);
nor U23045 (N_23045,N_12668,N_17199);
nor U23046 (N_23046,N_17895,N_17292);
nand U23047 (N_23047,N_14967,N_15815);
nor U23048 (N_23048,N_18264,N_12731);
and U23049 (N_23049,N_14131,N_11240);
or U23050 (N_23050,N_17438,N_17470);
nor U23051 (N_23051,N_16087,N_12237);
nand U23052 (N_23052,N_14601,N_19030);
nor U23053 (N_23053,N_11747,N_11639);
nand U23054 (N_23054,N_19089,N_15948);
or U23055 (N_23055,N_13280,N_16291);
xnor U23056 (N_23056,N_11174,N_19966);
nand U23057 (N_23057,N_12567,N_14610);
and U23058 (N_23058,N_12192,N_13947);
nor U23059 (N_23059,N_14216,N_10274);
nand U23060 (N_23060,N_15281,N_14479);
and U23061 (N_23061,N_11764,N_15481);
nand U23062 (N_23062,N_12952,N_14230);
xor U23063 (N_23063,N_15321,N_14620);
and U23064 (N_23064,N_13255,N_12753);
and U23065 (N_23065,N_15046,N_13706);
or U23066 (N_23066,N_14872,N_12476);
xnor U23067 (N_23067,N_17247,N_19145);
or U23068 (N_23068,N_18259,N_14446);
nor U23069 (N_23069,N_17085,N_12623);
xnor U23070 (N_23070,N_11341,N_14617);
nor U23071 (N_23071,N_15817,N_18236);
nor U23072 (N_23072,N_17904,N_12544);
or U23073 (N_23073,N_13424,N_12022);
nor U23074 (N_23074,N_12532,N_13197);
nand U23075 (N_23075,N_14278,N_13821);
nor U23076 (N_23076,N_12666,N_19689);
nand U23077 (N_23077,N_12334,N_19972);
nand U23078 (N_23078,N_17314,N_18545);
and U23079 (N_23079,N_15364,N_13917);
nand U23080 (N_23080,N_12165,N_19317);
nand U23081 (N_23081,N_18582,N_16826);
nand U23082 (N_23082,N_12013,N_17783);
and U23083 (N_23083,N_10571,N_19329);
xnor U23084 (N_23084,N_19531,N_12003);
nor U23085 (N_23085,N_18305,N_12395);
or U23086 (N_23086,N_16535,N_12691);
and U23087 (N_23087,N_13824,N_19719);
nand U23088 (N_23088,N_17514,N_17475);
or U23089 (N_23089,N_19685,N_12234);
or U23090 (N_23090,N_16549,N_10309);
and U23091 (N_23091,N_19029,N_16287);
or U23092 (N_23092,N_12581,N_16089);
xnor U23093 (N_23093,N_13777,N_10063);
nor U23094 (N_23094,N_17991,N_19919);
nor U23095 (N_23095,N_13231,N_10913);
nand U23096 (N_23096,N_15108,N_11391);
nor U23097 (N_23097,N_14492,N_12004);
nor U23098 (N_23098,N_16009,N_14763);
or U23099 (N_23099,N_12016,N_19670);
and U23100 (N_23100,N_18127,N_19001);
and U23101 (N_23101,N_12919,N_17603);
nand U23102 (N_23102,N_14352,N_13283);
nor U23103 (N_23103,N_17834,N_18906);
xnor U23104 (N_23104,N_15164,N_11308);
nor U23105 (N_23105,N_13827,N_10196);
and U23106 (N_23106,N_11787,N_15198);
nand U23107 (N_23107,N_17431,N_19499);
nand U23108 (N_23108,N_14813,N_13206);
or U23109 (N_23109,N_12258,N_11653);
nor U23110 (N_23110,N_16617,N_13391);
or U23111 (N_23111,N_11990,N_11832);
xnor U23112 (N_23112,N_17188,N_12964);
nand U23113 (N_23113,N_11804,N_17853);
or U23114 (N_23114,N_11167,N_18556);
nor U23115 (N_23115,N_19921,N_17766);
or U23116 (N_23116,N_16482,N_15399);
nand U23117 (N_23117,N_12651,N_15611);
nand U23118 (N_23118,N_17690,N_17232);
nor U23119 (N_23119,N_10232,N_11602);
and U23120 (N_23120,N_19182,N_16545);
nand U23121 (N_23121,N_12792,N_15451);
nand U23122 (N_23122,N_16719,N_10834);
or U23123 (N_23123,N_15289,N_11166);
and U23124 (N_23124,N_14486,N_12139);
nor U23125 (N_23125,N_10648,N_11209);
xnor U23126 (N_23126,N_10640,N_14818);
and U23127 (N_23127,N_18868,N_19750);
and U23128 (N_23128,N_12402,N_10099);
nand U23129 (N_23129,N_14401,N_11683);
nor U23130 (N_23130,N_19376,N_14005);
or U23131 (N_23131,N_12000,N_10160);
and U23132 (N_23132,N_18713,N_10860);
or U23133 (N_23133,N_15005,N_15176);
or U23134 (N_23134,N_19059,N_18221);
nand U23135 (N_23135,N_13261,N_10643);
or U23136 (N_23136,N_10348,N_11660);
and U23137 (N_23137,N_14298,N_10300);
and U23138 (N_23138,N_12439,N_14248);
xor U23139 (N_23139,N_14198,N_14851);
and U23140 (N_23140,N_11437,N_17118);
and U23141 (N_23141,N_12881,N_17635);
xnor U23142 (N_23142,N_16400,N_18438);
and U23143 (N_23143,N_19126,N_16576);
and U23144 (N_23144,N_18985,N_14797);
nand U23145 (N_23145,N_11484,N_10327);
nor U23146 (N_23146,N_12709,N_15906);
nand U23147 (N_23147,N_13389,N_16068);
and U23148 (N_23148,N_17031,N_13632);
and U23149 (N_23149,N_18009,N_13275);
xnor U23150 (N_23150,N_14392,N_10761);
nor U23151 (N_23151,N_19520,N_16172);
nor U23152 (N_23152,N_16418,N_16133);
or U23153 (N_23153,N_17718,N_13616);
and U23154 (N_23154,N_10523,N_11073);
or U23155 (N_23155,N_17619,N_17002);
and U23156 (N_23156,N_10866,N_14512);
nor U23157 (N_23157,N_19065,N_15166);
or U23158 (N_23158,N_12225,N_19042);
nor U23159 (N_23159,N_19190,N_15840);
or U23160 (N_23160,N_10033,N_17922);
or U23161 (N_23161,N_19471,N_14420);
nand U23162 (N_23162,N_14817,N_18856);
and U23163 (N_23163,N_16017,N_14835);
or U23164 (N_23164,N_13766,N_15126);
and U23165 (N_23165,N_18514,N_11110);
nand U23166 (N_23166,N_19196,N_12704);
nand U23167 (N_23167,N_15580,N_15030);
nand U23168 (N_23168,N_10198,N_14306);
and U23169 (N_23169,N_19447,N_11125);
or U23170 (N_23170,N_18701,N_17367);
nor U23171 (N_23171,N_19232,N_14957);
nor U23172 (N_23172,N_16241,N_11184);
xor U23173 (N_23173,N_11680,N_19870);
and U23174 (N_23174,N_10850,N_11410);
nor U23175 (N_23175,N_12108,N_15014);
and U23176 (N_23176,N_19020,N_10852);
or U23177 (N_23177,N_17513,N_13717);
nand U23178 (N_23178,N_17046,N_16113);
or U23179 (N_23179,N_18630,N_10619);
nor U23180 (N_23180,N_19829,N_11814);
nor U23181 (N_23181,N_12324,N_12168);
or U23182 (N_23182,N_18171,N_17082);
nor U23183 (N_23183,N_18115,N_12895);
xnor U23184 (N_23184,N_14362,N_11805);
nor U23185 (N_23185,N_13004,N_10250);
or U23186 (N_23186,N_16577,N_10359);
nand U23187 (N_23187,N_18033,N_16799);
nor U23188 (N_23188,N_16593,N_12572);
and U23189 (N_23189,N_15416,N_12187);
nor U23190 (N_23190,N_11293,N_19736);
nor U23191 (N_23191,N_14669,N_10084);
or U23192 (N_23192,N_16159,N_15256);
nor U23193 (N_23193,N_18488,N_19242);
nand U23194 (N_23194,N_14157,N_11047);
nor U23195 (N_23195,N_18973,N_16186);
nand U23196 (N_23196,N_12451,N_11850);
xnor U23197 (N_23197,N_16809,N_19354);
nand U23198 (N_23198,N_19562,N_10202);
and U23199 (N_23199,N_10243,N_12385);
nor U23200 (N_23200,N_19047,N_19677);
nor U23201 (N_23201,N_16464,N_10947);
and U23202 (N_23202,N_17024,N_16055);
nor U23203 (N_23203,N_14687,N_14370);
and U23204 (N_23204,N_18567,N_17977);
nand U23205 (N_23205,N_11142,N_14573);
or U23206 (N_23206,N_18099,N_11004);
nor U23207 (N_23207,N_14562,N_13260);
or U23208 (N_23208,N_15640,N_15106);
nor U23209 (N_23209,N_18363,N_11136);
nor U23210 (N_23210,N_19345,N_10756);
and U23211 (N_23211,N_18893,N_14289);
or U23212 (N_23212,N_18025,N_10830);
or U23213 (N_23213,N_16546,N_14233);
nand U23214 (N_23214,N_17581,N_13202);
and U23215 (N_23215,N_10433,N_12686);
or U23216 (N_23216,N_11821,N_18992);
nand U23217 (N_23217,N_17588,N_13936);
xnor U23218 (N_23218,N_12029,N_11890);
nor U23219 (N_23219,N_16239,N_12962);
nor U23220 (N_23220,N_12900,N_19857);
or U23221 (N_23221,N_15354,N_18715);
xor U23222 (N_23222,N_17531,N_12051);
xnor U23223 (N_23223,N_18430,N_10081);
nand U23224 (N_23224,N_13833,N_19279);
nand U23225 (N_23225,N_17282,N_13461);
or U23226 (N_23226,N_11086,N_19941);
and U23227 (N_23227,N_12936,N_14701);
and U23228 (N_23228,N_14860,N_14342);
xor U23229 (N_23229,N_13180,N_15801);
nor U23230 (N_23230,N_15692,N_13044);
nand U23231 (N_23231,N_17966,N_19049);
nor U23232 (N_23232,N_13834,N_13884);
nor U23233 (N_23233,N_16983,N_14507);
nand U23234 (N_23234,N_15857,N_19293);
xor U23235 (N_23235,N_14264,N_15017);
and U23236 (N_23236,N_11589,N_13695);
and U23237 (N_23237,N_13729,N_13855);
and U23238 (N_23238,N_18498,N_15988);
and U23239 (N_23239,N_13920,N_18986);
or U23240 (N_23240,N_17385,N_10303);
nor U23241 (N_23241,N_12680,N_14338);
or U23242 (N_23242,N_10125,N_10758);
and U23243 (N_23243,N_12027,N_19754);
nor U23244 (N_23244,N_11190,N_16703);
or U23245 (N_23245,N_14038,N_12504);
nand U23246 (N_23246,N_15208,N_12973);
nor U23247 (N_23247,N_13554,N_10893);
or U23248 (N_23248,N_11035,N_19428);
nand U23249 (N_23249,N_11577,N_11383);
nor U23250 (N_23250,N_17616,N_11969);
or U23251 (N_23251,N_12379,N_16379);
and U23252 (N_23252,N_11927,N_15890);
nand U23253 (N_23253,N_12127,N_12867);
nand U23254 (N_23254,N_12255,N_10329);
or U23255 (N_23255,N_19359,N_10102);
or U23256 (N_23256,N_12466,N_15301);
nand U23257 (N_23257,N_14828,N_17037);
and U23258 (N_23258,N_15829,N_10371);
and U23259 (N_23259,N_12963,N_10204);
nand U23260 (N_23260,N_10292,N_17670);
nand U23261 (N_23261,N_10260,N_14990);
xnor U23262 (N_23262,N_10682,N_11430);
nand U23263 (N_23263,N_15802,N_19461);
or U23264 (N_23264,N_16956,N_10663);
and U23265 (N_23265,N_14168,N_16363);
or U23266 (N_23266,N_12762,N_10451);
and U23267 (N_23267,N_19613,N_13960);
nand U23268 (N_23268,N_16912,N_10888);
nand U23269 (N_23269,N_19094,N_16676);
nand U23270 (N_23270,N_18895,N_12031);
or U23271 (N_23271,N_18894,N_15749);
or U23272 (N_23272,N_11348,N_13587);
and U23273 (N_23273,N_16910,N_12021);
nor U23274 (N_23274,N_17150,N_12133);
nor U23275 (N_23275,N_14035,N_19641);
nand U23276 (N_23276,N_11324,N_11134);
and U23277 (N_23277,N_15752,N_11597);
and U23278 (N_23278,N_17473,N_12655);
or U23279 (N_23279,N_12063,N_14056);
xor U23280 (N_23280,N_17056,N_17089);
or U23281 (N_23281,N_16802,N_19395);
nor U23282 (N_23282,N_13314,N_17737);
or U23283 (N_23283,N_11565,N_17159);
nor U23284 (N_23284,N_10008,N_13678);
nand U23285 (N_23285,N_16738,N_18874);
nor U23286 (N_23286,N_13793,N_13650);
nor U23287 (N_23287,N_13786,N_19600);
and U23288 (N_23288,N_16572,N_13618);
or U23289 (N_23289,N_15100,N_14428);
nand U23290 (N_23290,N_17299,N_12008);
nor U23291 (N_23291,N_14862,N_12284);
nand U23292 (N_23292,N_16820,N_13895);
and U23293 (N_23293,N_17041,N_14529);
nand U23294 (N_23294,N_11605,N_19977);
nand U23295 (N_23295,N_13239,N_11845);
xnor U23296 (N_23296,N_10838,N_15104);
nand U23297 (N_23297,N_16865,N_10073);
or U23298 (N_23298,N_13228,N_11239);
and U23299 (N_23299,N_17743,N_14107);
and U23300 (N_23300,N_10420,N_10455);
nor U23301 (N_23301,N_12635,N_11427);
nor U23302 (N_23302,N_12728,N_15438);
nand U23303 (N_23303,N_10514,N_11649);
nand U23304 (N_23304,N_10650,N_10635);
nand U23305 (N_23305,N_11413,N_15453);
nand U23306 (N_23306,N_14004,N_12183);
nor U23307 (N_23307,N_17146,N_10374);
or U23308 (N_23308,N_18173,N_10612);
nor U23309 (N_23309,N_16391,N_13288);
nand U23310 (N_23310,N_13511,N_13609);
xnor U23311 (N_23311,N_19629,N_19953);
or U23312 (N_23312,N_10466,N_13185);
and U23313 (N_23313,N_16114,N_19818);
or U23314 (N_23314,N_15839,N_17182);
nand U23315 (N_23315,N_10296,N_18983);
nand U23316 (N_23316,N_18974,N_16852);
xor U23317 (N_23317,N_14408,N_10025);
nand U23318 (N_23318,N_16558,N_14824);
nor U23319 (N_23319,N_11171,N_16028);
and U23320 (N_23320,N_13307,N_11879);
nor U23321 (N_23321,N_16282,N_13829);
nand U23322 (N_23322,N_11645,N_13800);
or U23323 (N_23323,N_10347,N_14979);
and U23324 (N_23324,N_19497,N_13608);
nand U23325 (N_23325,N_16760,N_13826);
xnor U23326 (N_23326,N_14163,N_12536);
nor U23327 (N_23327,N_18592,N_12199);
or U23328 (N_23328,N_16030,N_18298);
or U23329 (N_23329,N_12151,N_13363);
or U23330 (N_23330,N_11360,N_12101);
and U23331 (N_23331,N_15147,N_11532);
xor U23332 (N_23332,N_13482,N_13055);
nand U23333 (N_23333,N_17442,N_16784);
or U23334 (N_23334,N_11203,N_12876);
and U23335 (N_23335,N_13062,N_14449);
or U23336 (N_23336,N_15631,N_10344);
or U23337 (N_23337,N_11301,N_15263);
nand U23338 (N_23338,N_11633,N_16803);
nor U23339 (N_23339,N_15741,N_18513);
and U23340 (N_23340,N_12497,N_18505);
and U23341 (N_23341,N_15638,N_16377);
or U23342 (N_23342,N_17087,N_13068);
nand U23343 (N_23343,N_18898,N_18751);
or U23344 (N_23344,N_13775,N_17276);
or U23345 (N_23345,N_14719,N_12332);
or U23346 (N_23346,N_16354,N_13603);
and U23347 (N_23347,N_15047,N_12190);
or U23348 (N_23348,N_14147,N_15293);
nand U23349 (N_23349,N_11129,N_12493);
nor U23350 (N_23350,N_11881,N_12292);
and U23351 (N_23351,N_14318,N_15141);
nor U23352 (N_23352,N_12143,N_19400);
and U23353 (N_23353,N_13459,N_14191);
and U23354 (N_23354,N_18553,N_18507);
or U23355 (N_23355,N_19592,N_15738);
nor U23356 (N_23356,N_12615,N_11988);
and U23357 (N_23357,N_16362,N_18597);
nand U23358 (N_23358,N_12642,N_16023);
nand U23359 (N_23359,N_11367,N_17873);
and U23360 (N_23360,N_16842,N_11902);
and U23361 (N_23361,N_15978,N_10016);
nand U23362 (N_23362,N_14895,N_10353);
or U23363 (N_23363,N_16637,N_19177);
nor U23364 (N_23364,N_17427,N_15088);
nor U23365 (N_23365,N_18887,N_11985);
nand U23366 (N_23366,N_13277,N_13594);
nand U23367 (N_23367,N_11474,N_15844);
and U23368 (N_23368,N_17815,N_19405);
and U23369 (N_23369,N_19385,N_14144);
nor U23370 (N_23370,N_19802,N_10991);
nor U23371 (N_23371,N_17844,N_19766);
or U23372 (N_23372,N_17310,N_14001);
nor U23373 (N_23373,N_12673,N_15341);
and U23374 (N_23374,N_17800,N_11576);
nor U23375 (N_23375,N_16745,N_10287);
nand U23376 (N_23376,N_18271,N_15258);
xnor U23377 (N_23377,N_14418,N_12075);
xnor U23378 (N_23378,N_18159,N_12529);
and U23379 (N_23379,N_10170,N_10713);
xor U23380 (N_23380,N_17544,N_18113);
nor U23381 (N_23381,N_17339,N_12749);
and U23382 (N_23382,N_16782,N_17318);
nor U23383 (N_23383,N_14220,N_15836);
xor U23384 (N_23384,N_10550,N_11968);
nand U23385 (N_23385,N_10711,N_16409);
nand U23386 (N_23386,N_19982,N_13839);
or U23387 (N_23387,N_12542,N_12390);
and U23388 (N_23388,N_16423,N_11332);
and U23389 (N_23389,N_16671,N_13119);
or U23390 (N_23390,N_16437,N_13049);
or U23391 (N_23391,N_17481,N_17673);
nor U23392 (N_23392,N_16365,N_17191);
and U23393 (N_23393,N_10119,N_18782);
nand U23394 (N_23394,N_19388,N_13176);
or U23395 (N_23395,N_18226,N_18500);
and U23396 (N_23396,N_10277,N_16135);
and U23397 (N_23397,N_10141,N_10848);
or U23398 (N_23398,N_18480,N_17605);
or U23399 (N_23399,N_14134,N_18752);
nand U23400 (N_23400,N_11178,N_10385);
or U23401 (N_23401,N_11909,N_10988);
nand U23402 (N_23402,N_17099,N_13626);
or U23403 (N_23403,N_11657,N_13279);
or U23404 (N_23404,N_19320,N_14964);
nand U23405 (N_23405,N_10765,N_18051);
and U23406 (N_23406,N_15835,N_15529);
or U23407 (N_23407,N_19440,N_18282);
xor U23408 (N_23408,N_16067,N_18145);
nand U23409 (N_23409,N_17772,N_17027);
and U23410 (N_23410,N_16977,N_17316);
and U23411 (N_23411,N_17194,N_13976);
nand U23412 (N_23412,N_16251,N_12845);
nand U23413 (N_23413,N_10922,N_10528);
or U23414 (N_23414,N_10405,N_11039);
nand U23415 (N_23415,N_19984,N_10355);
and U23416 (N_23416,N_14240,N_10464);
and U23417 (N_23417,N_19805,N_12153);
or U23418 (N_23418,N_12201,N_10325);
nand U23419 (N_23419,N_18754,N_18572);
nand U23420 (N_23420,N_10495,N_13282);
and U23421 (N_23421,N_15472,N_13733);
nand U23422 (N_23422,N_18569,N_12957);
or U23423 (N_23423,N_13175,N_12282);
nand U23424 (N_23424,N_10981,N_13736);
nor U23425 (N_23425,N_19069,N_15357);
or U23426 (N_23426,N_18179,N_17754);
and U23427 (N_23427,N_17607,N_10677);
nand U23428 (N_23428,N_10463,N_17932);
xnor U23429 (N_23429,N_14878,N_17668);
xnor U23430 (N_23430,N_15064,N_12310);
and U23431 (N_23431,N_19704,N_11869);
or U23432 (N_23432,N_12760,N_19620);
nor U23433 (N_23433,N_18547,N_14659);
and U23434 (N_23434,N_14186,N_14422);
nand U23435 (N_23435,N_10085,N_12331);
and U23436 (N_23436,N_19106,N_16649);
xnor U23437 (N_23437,N_15025,N_15696);
and U23438 (N_23438,N_17383,N_14397);
or U23439 (N_23439,N_15970,N_14523);
nor U23440 (N_23440,N_11983,N_10069);
and U23441 (N_23441,N_13460,N_15945);
or U23442 (N_23442,N_15633,N_19147);
nor U23443 (N_23443,N_13950,N_10600);
or U23444 (N_23444,N_17788,N_10280);
or U23445 (N_23445,N_18925,N_15697);
and U23446 (N_23446,N_15156,N_19223);
and U23447 (N_23447,N_17372,N_18755);
nand U23448 (N_23448,N_15951,N_17101);
nand U23449 (N_23449,N_14140,N_17851);
nand U23450 (N_23450,N_16706,N_13323);
nand U23451 (N_23451,N_14347,N_12318);
xnor U23452 (N_23452,N_18353,N_19168);
nor U23453 (N_23453,N_15264,N_14671);
and U23454 (N_23454,N_10621,N_17296);
and U23455 (N_23455,N_13064,N_15624);
xor U23456 (N_23456,N_16016,N_11407);
and U23457 (N_23457,N_15535,N_12649);
nor U23458 (N_23458,N_18045,N_18365);
xnor U23459 (N_23459,N_18022,N_15990);
and U23460 (N_23460,N_13581,N_11201);
and U23461 (N_23461,N_12186,N_17216);
and U23462 (N_23462,N_16352,N_19813);
xor U23463 (N_23463,N_18632,N_12216);
or U23464 (N_23464,N_10894,N_16653);
nand U23465 (N_23465,N_15485,N_10606);
nand U23466 (N_23466,N_18433,N_15003);
nand U23467 (N_23467,N_19000,N_17215);
nor U23468 (N_23468,N_11806,N_17604);
and U23469 (N_23469,N_10207,N_17084);
nand U23470 (N_23470,N_10569,N_16763);
and U23471 (N_23471,N_11686,N_16791);
nor U23472 (N_23472,N_14046,N_10418);
and U23473 (N_23473,N_19070,N_19798);
and U23474 (N_23474,N_12825,N_15066);
and U23475 (N_23475,N_13046,N_11255);
or U23476 (N_23476,N_11811,N_18375);
nor U23477 (N_23477,N_15096,N_19741);
nand U23478 (N_23478,N_16109,N_15987);
and U23479 (N_23479,N_19023,N_13114);
or U23480 (N_23480,N_16324,N_13083);
or U23481 (N_23481,N_18429,N_12175);
nand U23482 (N_23482,N_14594,N_16726);
or U23483 (N_23483,N_19082,N_17840);
and U23484 (N_23484,N_15827,N_10925);
nor U23485 (N_23485,N_10533,N_16834);
nor U23486 (N_23486,N_14164,N_10962);
nand U23487 (N_23487,N_12188,N_15170);
nor U23488 (N_23488,N_12093,N_11840);
or U23489 (N_23489,N_11995,N_16587);
and U23490 (N_23490,N_16993,N_10181);
nor U23491 (N_23491,N_15755,N_11497);
and U23492 (N_23492,N_14239,N_12901);
nand U23493 (N_23493,N_13110,N_18464);
xor U23494 (N_23494,N_15194,N_16256);
nor U23495 (N_23495,N_18770,N_12472);
nor U23496 (N_23496,N_10335,N_19247);
and U23497 (N_23497,N_10482,N_13590);
nand U23498 (N_23498,N_11372,N_15284);
xor U23499 (N_23499,N_19300,N_11181);
nand U23500 (N_23500,N_16815,N_10262);
and U23501 (N_23501,N_15086,N_19773);
and U23502 (N_23502,N_14102,N_17401);
nor U23503 (N_23503,N_12309,N_11002);
or U23504 (N_23504,N_16399,N_18379);
nor U23505 (N_23505,N_13586,N_17860);
nor U23506 (N_23506,N_19647,N_11586);
or U23507 (N_23507,N_15797,N_15598);
nor U23508 (N_23508,N_16012,N_10367);
or U23509 (N_23509,N_11182,N_11859);
nor U23510 (N_23510,N_13665,N_14940);
or U23511 (N_23511,N_10821,N_17460);
nor U23512 (N_23512,N_13113,N_11305);
nor U23513 (N_23513,N_18574,N_19682);
nor U23514 (N_23514,N_13676,N_11246);
and U23515 (N_23515,N_12453,N_12270);
or U23516 (N_23516,N_15870,N_19799);
nor U23517 (N_23517,N_16236,N_16029);
or U23518 (N_23518,N_13743,N_15769);
or U23519 (N_23519,N_17751,N_19899);
nand U23520 (N_23520,N_14616,N_11922);
xor U23521 (N_23521,N_15054,N_16741);
or U23522 (N_23522,N_13810,N_16886);
nand U23523 (N_23523,N_11043,N_12540);
nor U23524 (N_23524,N_13230,N_19207);
nor U23525 (N_23525,N_18689,N_14441);
xor U23526 (N_23526,N_14470,N_19971);
or U23527 (N_23527,N_12684,N_12235);
and U23528 (N_23528,N_14268,N_19867);
and U23529 (N_23529,N_18635,N_14946);
nand U23530 (N_23530,N_14436,N_15927);
nor U23531 (N_23531,N_19502,N_11461);
nand U23532 (N_23532,N_17609,N_17222);
nor U23533 (N_23533,N_10607,N_19569);
or U23534 (N_23534,N_18192,N_17370);
nand U23535 (N_23535,N_17836,N_14497);
nor U23536 (N_23536,N_13904,N_18338);
nand U23537 (N_23537,N_17452,N_18202);
or U23538 (N_23538,N_10642,N_10994);
or U23539 (N_23539,N_14353,N_10164);
or U23540 (N_23540,N_12329,N_18657);
and U23541 (N_23541,N_16144,N_13534);
nand U23542 (N_23542,N_17384,N_17520);
nand U23543 (N_23543,N_15337,N_13613);
nor U23544 (N_23544,N_17464,N_12759);
nand U23545 (N_23545,N_15103,N_15369);
or U23546 (N_23546,N_12432,N_17557);
xor U23547 (N_23547,N_12875,N_10431);
nand U23548 (N_23548,N_18558,N_12417);
or U23549 (N_23549,N_15336,N_12647);
xor U23550 (N_23550,N_10093,N_14927);
nor U23551 (N_23551,N_17258,N_12109);
nand U23552 (N_23552,N_11369,N_19305);
xnor U23553 (N_23553,N_12687,N_17278);
or U23554 (N_23554,N_19229,N_16795);
or U23555 (N_23555,N_17488,N_15192);
nor U23556 (N_23556,N_13660,N_16654);
nand U23557 (N_23557,N_18946,N_19761);
and U23558 (N_23558,N_15853,N_10448);
nand U23559 (N_23559,N_16620,N_10792);
and U23560 (N_23560,N_10440,N_14403);
nor U23561 (N_23561,N_15401,N_11422);
nor U23562 (N_23562,N_19237,N_11124);
nand U23563 (N_23563,N_17130,N_11825);
or U23564 (N_23564,N_15350,N_16348);
or U23565 (N_23565,N_14732,N_15236);
nor U23566 (N_23566,N_15812,N_16539);
nor U23567 (N_23567,N_15229,N_15160);
or U23568 (N_23568,N_19847,N_19063);
and U23569 (N_23569,N_17468,N_18937);
or U23570 (N_23570,N_19683,N_12685);
nor U23571 (N_23571,N_13942,N_11984);
nor U23572 (N_23572,N_17416,N_19779);
xnor U23573 (N_23573,N_18731,N_14665);
nor U23574 (N_23574,N_15706,N_10404);
and U23575 (N_23575,N_19852,N_12583);
nand U23576 (N_23576,N_14246,N_15761);
or U23577 (N_23577,N_17600,N_14235);
nor U23578 (N_23578,N_15491,N_15187);
nor U23579 (N_23579,N_13569,N_13849);
nand U23580 (N_23580,N_19861,N_12893);
and U23581 (N_23581,N_10163,N_12305);
and U23582 (N_23582,N_16498,N_18320);
xnor U23583 (N_23583,N_16694,N_18666);
nor U23584 (N_23584,N_13757,N_12507);
or U23585 (N_23585,N_16233,N_13579);
nand U23586 (N_23586,N_14607,N_19890);
nor U23587 (N_23587,N_11416,N_12782);
nor U23588 (N_23588,N_18912,N_13386);
or U23589 (N_23589,N_11344,N_13769);
and U23590 (N_23590,N_14148,N_16124);
nand U23591 (N_23591,N_13167,N_12594);
nor U23592 (N_23592,N_13718,N_16210);
nor U23593 (N_23593,N_19005,N_12662);
nand U23594 (N_23594,N_10091,N_19310);
and U23595 (N_23595,N_15510,N_19084);
nand U23596 (N_23596,N_16778,N_16941);
or U23597 (N_23597,N_14069,N_18180);
and U23598 (N_23598,N_16414,N_10752);
or U23599 (N_23599,N_11156,N_19156);
xnor U23600 (N_23600,N_11917,N_14608);
nand U23601 (N_23601,N_15717,N_15295);
or U23602 (N_23602,N_13808,N_13141);
nand U23603 (N_23603,N_17733,N_19564);
xor U23604 (N_23604,N_18340,N_11087);
and U23605 (N_23605,N_10881,N_16628);
nand U23606 (N_23606,N_10049,N_16376);
nor U23607 (N_23607,N_17952,N_15858);
or U23608 (N_23608,N_18902,N_13778);
nand U23609 (N_23609,N_19134,N_14271);
nand U23610 (N_23610,N_12110,N_14668);
xnor U23611 (N_23611,N_13624,N_11420);
nor U23612 (N_23612,N_11964,N_10914);
and U23613 (N_23613,N_16178,N_10644);
nor U23614 (N_23614,N_12600,N_15465);
and U23615 (N_23615,N_10736,N_11691);
or U23616 (N_23616,N_11762,N_15469);
nor U23617 (N_23617,N_10800,N_18662);
nor U23618 (N_23618,N_12371,N_12429);
and U23619 (N_23619,N_15461,N_15753);
and U23620 (N_23620,N_15042,N_17374);
and U23621 (N_23621,N_11251,N_15537);
and U23622 (N_23622,N_19981,N_19464);
and U23623 (N_23623,N_17750,N_13803);
and U23624 (N_23624,N_11406,N_15201);
nor U23625 (N_23625,N_19723,N_14509);
and U23626 (N_23626,N_12362,N_13448);
nand U23627 (N_23627,N_17100,N_10493);
nor U23628 (N_23628,N_18083,N_10254);
and U23629 (N_23629,N_18872,N_15869);
and U23630 (N_23630,N_11545,N_17657);
nor U23631 (N_23631,N_15550,N_12580);
nor U23632 (N_23632,N_13376,N_14328);
nor U23633 (N_23633,N_13994,N_10921);
or U23634 (N_23634,N_14193,N_10445);
or U23635 (N_23635,N_15511,N_11198);
xor U23636 (N_23636,N_14947,N_11728);
and U23637 (N_23637,N_14945,N_17716);
nand U23638 (N_23638,N_18686,N_11270);
and U23639 (N_23639,N_14417,N_13019);
nor U23640 (N_23640,N_10255,N_19154);
nand U23641 (N_23641,N_19241,N_17659);
nor U23642 (N_23642,N_18743,N_11015);
nand U23643 (N_23643,N_12806,N_12295);
nand U23644 (N_23644,N_10155,N_14047);
and U23645 (N_23645,N_17636,N_17515);
and U23646 (N_23646,N_19652,N_16149);
nor U23647 (N_23647,N_11993,N_10340);
nor U23648 (N_23648,N_11370,N_14996);
or U23649 (N_23649,N_19415,N_18620);
nor U23650 (N_23650,N_12827,N_11145);
and U23651 (N_23651,N_16623,N_15189);
and U23652 (N_23652,N_13530,N_14630);
or U23653 (N_23653,N_16225,N_10841);
nor U23654 (N_23654,N_18485,N_13779);
or U23655 (N_23655,N_19893,N_11550);
and U23656 (N_23656,N_13744,N_15780);
nand U23657 (N_23657,N_13227,N_18184);
nor U23658 (N_23658,N_19467,N_10316);
xor U23659 (N_23659,N_10129,N_10931);
nor U23660 (N_23660,N_14267,N_13138);
nor U23661 (N_23661,N_15190,N_10279);
nand U23662 (N_23662,N_17137,N_19543);
xnor U23663 (N_23663,N_15095,N_18052);
nand U23664 (N_23664,N_17643,N_19117);
or U23665 (N_23665,N_10712,N_10187);
xor U23666 (N_23666,N_18450,N_12657);
and U23667 (N_23667,N_10338,N_18707);
xnor U23668 (N_23668,N_13107,N_14324);
xnor U23669 (N_23669,N_15209,N_11570);
xnor U23670 (N_23670,N_15619,N_10787);
nand U23671 (N_23671,N_19249,N_15530);
nor U23672 (N_23672,N_15183,N_18534);
nor U23673 (N_23673,N_17030,N_12909);
and U23674 (N_23674,N_19573,N_17175);
and U23675 (N_23675,N_17398,N_16454);
nand U23676 (N_23676,N_17073,N_14657);
or U23677 (N_23677,N_16301,N_19025);
or U23678 (N_23678,N_18468,N_12244);
nor U23679 (N_23679,N_18458,N_14757);
xor U23680 (N_23680,N_11179,N_17911);
and U23681 (N_23681,N_18461,N_14426);
and U23682 (N_23682,N_15002,N_17608);
and U23683 (N_23683,N_12152,N_16311);
nor U23684 (N_23684,N_13940,N_12595);
nand U23685 (N_23685,N_13118,N_16285);
nand U23686 (N_23686,N_11133,N_16739);
nand U23687 (N_23687,N_10955,N_10676);
nor U23688 (N_23688,N_15006,N_14855);
and U23689 (N_23689,N_16509,N_10469);
and U23690 (N_23690,N_15679,N_13741);
or U23691 (N_23691,N_13367,N_18174);
xnor U23692 (N_23692,N_17432,N_13430);
nor U23693 (N_23693,N_15512,N_13761);
and U23694 (N_23694,N_11538,N_18879);
and U23695 (N_23695,N_19598,N_18506);
nand U23696 (N_23696,N_11967,N_17762);
nor U23697 (N_23697,N_15939,N_14226);
nor U23698 (N_23698,N_17930,N_15953);
and U23699 (N_23699,N_16832,N_16989);
or U23700 (N_23700,N_16469,N_17525);
nand U23701 (N_23701,N_14037,N_16434);
or U23702 (N_23702,N_14649,N_10942);
or U23703 (N_23703,N_18939,N_13955);
and U23704 (N_23704,N_14519,N_16004);
or U23705 (N_23705,N_15721,N_11536);
nand U23706 (N_23706,N_18252,N_16499);
nand U23707 (N_23707,N_12501,N_14919);
nand U23708 (N_23708,N_12648,N_16327);
nand U23709 (N_23709,N_17197,N_15726);
or U23710 (N_23710,N_17429,N_12757);
or U23711 (N_23711,N_16370,N_11046);
or U23712 (N_23712,N_10530,N_18339);
nor U23713 (N_23713,N_18087,N_12783);
or U23714 (N_23714,N_13625,N_16783);
nand U23715 (N_23715,N_15974,N_14729);
nor U23716 (N_23716,N_13858,N_18634);
nand U23717 (N_23717,N_14054,N_18559);
and U23718 (N_23718,N_16429,N_19357);
or U23719 (N_23719,N_11195,N_15654);
xnor U23720 (N_23720,N_19163,N_16246);
nor U23721 (N_23721,N_18593,N_19146);
and U23722 (N_23722,N_16853,N_17479);
and U23723 (N_23723,N_12524,N_10722);
nand U23724 (N_23724,N_14123,N_11900);
nand U23725 (N_23725,N_12993,N_13669);
nand U23726 (N_23726,N_14142,N_16198);
xnor U23727 (N_23727,N_17667,N_11648);
xnor U23728 (N_23728,N_11638,N_16974);
nand U23729 (N_23729,N_18921,N_12050);
or U23730 (N_23730,N_12735,N_14224);
xnor U23731 (N_23731,N_15587,N_17264);
nand U23732 (N_23732,N_11272,N_12821);
xor U23733 (N_23733,N_18802,N_15233);
or U23734 (N_23734,N_11601,N_16208);
or U23735 (N_23735,N_19903,N_11358);
nand U23736 (N_23736,N_13103,N_19663);
or U23737 (N_23737,N_16333,N_11486);
and U23738 (N_23738,N_14300,N_14277);
xnor U23739 (N_23739,N_12863,N_19627);
or U23740 (N_23740,N_12137,N_16708);
nand U23741 (N_23741,N_12064,N_10461);
nand U23742 (N_23742,N_10671,N_19448);
or U23743 (N_23743,N_11411,N_17290);
or U23744 (N_23744,N_11989,N_15900);
nand U23745 (N_23745,N_17107,N_11851);
and U23746 (N_23746,N_16451,N_17677);
nand U23747 (N_23747,N_10868,N_10867);
or U23748 (N_23748,N_18209,N_17157);
and U23749 (N_23749,N_10859,N_18727);
nor U23750 (N_23750,N_13794,N_19412);
nor U23751 (N_23751,N_18524,N_11072);
or U23752 (N_23752,N_17443,N_10032);
nand U23753 (N_23753,N_12388,N_19344);
or U23754 (N_23754,N_19090,N_16892);
nand U23755 (N_23755,N_12248,N_13312);
xor U23756 (N_23756,N_13361,N_18137);
nor U23757 (N_23757,N_15918,N_19559);
or U23758 (N_23758,N_15121,N_12857);
or U23759 (N_23759,N_14781,N_17167);
or U23760 (N_23760,N_13347,N_17347);
or U23761 (N_23761,N_12141,N_12706);
nor U23762 (N_23762,N_19995,N_18745);
nor U23763 (N_23763,N_15843,N_13272);
nor U23764 (N_23764,N_17109,N_11852);
and U23765 (N_23765,N_17872,N_18454);
nor U23766 (N_23766,N_18889,N_16417);
nor U23767 (N_23767,N_10416,N_19198);
and U23768 (N_23768,N_15910,N_13815);
nand U23769 (N_23769,N_14717,N_15185);
nand U23770 (N_23770,N_10798,N_10623);
nor U23771 (N_23771,N_16200,N_17173);
nand U23772 (N_23772,N_12336,N_18729);
or U23773 (N_23773,N_13622,N_11684);
nand U23774 (N_23774,N_11853,N_15212);
nand U23775 (N_23775,N_11088,N_15080);
nand U23776 (N_23776,N_16839,N_13689);
nand U23777 (N_23777,N_19384,N_14149);
or U23778 (N_23778,N_16947,N_11552);
and U23779 (N_23779,N_16626,N_19137);
nand U23780 (N_23780,N_19653,N_15134);
or U23781 (N_23781,N_10809,N_15549);
nor U23782 (N_23782,N_12383,N_12832);
nand U23783 (N_23783,N_17203,N_17145);
nor U23784 (N_23784,N_12365,N_17420);
or U23785 (N_23785,N_10823,N_13290);
nand U23786 (N_23786,N_11688,N_19368);
nor U23787 (N_23787,N_18093,N_15305);
or U23788 (N_23788,N_13334,N_16971);
nor U23789 (N_23789,N_19371,N_16619);
nand U23790 (N_23790,N_18201,N_14382);
or U23791 (N_23791,N_17696,N_14011);
and U23792 (N_23792,N_15621,N_18377);
or U23793 (N_23793,N_14960,N_19033);
xor U23794 (N_23794,N_11517,N_16453);
and U23795 (N_23795,N_14612,N_11053);
or U23796 (N_23796,N_19445,N_15635);
and U23797 (N_23797,N_17066,N_18195);
xnor U23798 (N_23798,N_12316,N_14808);
xnor U23799 (N_23799,N_10103,N_15672);
or U23800 (N_23800,N_11878,N_19157);
nand U23801 (N_23801,N_10951,N_17192);
nand U23802 (N_23802,N_18661,N_15497);
or U23803 (N_23803,N_11603,N_15711);
and U23804 (N_23804,N_18001,N_11375);
nor U23805 (N_23805,N_19713,N_18143);
nor U23806 (N_23806,N_14249,N_19104);
or U23807 (N_23807,N_17321,N_17529);
nand U23808 (N_23808,N_12710,N_11971);
nor U23809 (N_23809,N_17298,N_10373);
and U23810 (N_23810,N_10108,N_18247);
or U23811 (N_23811,N_11315,N_10510);
and U23812 (N_23812,N_18484,N_14469);
and U23813 (N_23813,N_11214,N_18503);
nand U23814 (N_23814,N_17541,N_10918);
nand U23815 (N_23815,N_13032,N_14870);
nor U23816 (N_23816,N_19708,N_18419);
nand U23817 (N_23817,N_19637,N_16410);
or U23818 (N_23818,N_14764,N_17997);
nor U23819 (N_23819,N_19399,N_18449);
or U23820 (N_23820,N_18157,N_10884);
and U23821 (N_23821,N_16175,N_15148);
or U23822 (N_23822,N_19579,N_13008);
or U23823 (N_23823,N_12627,N_14363);
and U23824 (N_23824,N_14645,N_10937);
or U23825 (N_23825,N_10066,N_10024);
or U23826 (N_23826,N_12120,N_15967);
nand U23827 (N_23827,N_10377,N_13671);
xnor U23828 (N_23828,N_18966,N_19075);
nor U23829 (N_23829,N_11959,N_12804);
and U23830 (N_23830,N_16462,N_18067);
or U23831 (N_23831,N_10665,N_18944);
nand U23832 (N_23832,N_14477,N_14023);
and U23833 (N_23833,N_19483,N_16329);
and U23834 (N_23834,N_19841,N_11767);
and U23835 (N_23835,N_19604,N_12090);
nor U23836 (N_23836,N_13828,N_14444);
or U23837 (N_23837,N_17015,N_13556);
xnor U23838 (N_23838,N_19370,N_15540);
nor U23839 (N_23839,N_18492,N_16936);
nor U23840 (N_23840,N_14695,N_15327);
and U23841 (N_23841,N_11936,N_11652);
xor U23842 (N_23842,N_19366,N_11153);
nor U23843 (N_23843,N_17572,N_16758);
or U23844 (N_23844,N_18034,N_16300);
nand U23845 (N_23845,N_18725,N_16281);
nand U23846 (N_23846,N_12826,N_12880);
xnor U23847 (N_23847,N_12576,N_15239);
and U23848 (N_23848,N_18181,N_11090);
nand U23849 (N_23849,N_11222,N_19968);
nand U23850 (N_23850,N_18427,N_17561);
nor U23851 (N_23851,N_17180,N_19304);
or U23852 (N_23852,N_18604,N_16079);
or U23853 (N_23853,N_15335,N_17537);
nand U23854 (N_23854,N_14505,N_14276);
and U23855 (N_23855,N_16964,N_11097);
nor U23856 (N_23856,N_16833,N_16850);
or U23857 (N_23857,N_11496,N_14825);
nor U23858 (N_23858,N_11530,N_16824);
nor U23859 (N_23859,N_13079,N_12138);
nand U23860 (N_23860,N_14578,N_13798);
nand U23861 (N_23861,N_10733,N_19742);
or U23862 (N_23862,N_19211,N_14811);
nand U23863 (N_23863,N_10545,N_13529);
or U23864 (N_23864,N_19481,N_15402);
and U23865 (N_23865,N_12275,N_11520);
nor U23866 (N_23866,N_14734,N_19769);
nand U23867 (N_23867,N_16323,N_17277);
or U23868 (N_23868,N_12944,N_10203);
nand U23869 (N_23869,N_12178,N_10636);
xnor U23870 (N_23870,N_15307,N_18778);
and U23871 (N_23871,N_14112,N_16071);
nand U23872 (N_23872,N_12330,N_15736);
nand U23873 (N_23873,N_17917,N_15713);
nand U23874 (N_23874,N_11861,N_14238);
xnor U23875 (N_23875,N_15600,N_13969);
nor U23876 (N_23876,N_15816,N_19986);
and U23877 (N_23877,N_12172,N_11318);
or U23878 (N_23878,N_16959,N_12374);
nor U23879 (N_23879,N_19866,N_14254);
nand U23880 (N_23880,N_12062,N_15140);
or U23881 (N_23881,N_17325,N_17163);
and U23882 (N_23882,N_15792,N_18768);
and U23883 (N_23883,N_13993,N_12094);
nand U23884 (N_23884,N_19038,N_13066);
nand U23885 (N_23885,N_13218,N_10117);
nand U23886 (N_23886,N_19127,N_18341);
nor U23887 (N_23887,N_16060,N_17166);
xnor U23888 (N_23888,N_11326,N_11262);
xor U23889 (N_23889,N_12872,N_11618);
nand U23890 (N_23890,N_11734,N_18318);
and U23891 (N_23891,N_11123,N_15314);
nor U23892 (N_23892,N_11122,N_19687);
nor U23893 (N_23893,N_13379,N_15502);
nand U23894 (N_23894,N_19726,N_16604);
nor U23895 (N_23895,N_18005,N_16343);
or U23896 (N_23896,N_17249,N_18541);
and U23897 (N_23897,N_10797,N_11482);
nand U23898 (N_23898,N_14258,N_11522);
or U23899 (N_23899,N_17305,N_10903);
nor U23900 (N_23900,N_14335,N_15652);
nand U23901 (N_23901,N_14118,N_16722);
and U23902 (N_23902,N_12124,N_13241);
and U23903 (N_23903,N_13299,N_12799);
nor U23904 (N_23904,N_18728,N_13655);
nor U23905 (N_23905,N_12233,N_10858);
and U23906 (N_23906,N_19705,N_12794);
nand U23907 (N_23907,N_15018,N_19822);
or U23908 (N_23908,N_17115,N_18257);
nand U23909 (N_23909,N_13759,N_18032);
nand U23910 (N_23910,N_11759,N_12907);
or U23911 (N_23911,N_13539,N_15241);
and U23912 (N_23912,N_18629,N_18108);
xor U23913 (N_23913,N_14467,N_19171);
nor U23914 (N_23914,N_10288,N_19900);
and U23915 (N_23915,N_18873,N_11801);
nand U23916 (N_23916,N_17861,N_10382);
nor U23917 (N_23917,N_13912,N_19998);
nand U23918 (N_23918,N_13015,N_13321);
xnor U23919 (N_23919,N_13574,N_13910);
nand U23920 (N_23920,N_10080,N_17388);
nand U23921 (N_23921,N_13213,N_17767);
or U23922 (N_23922,N_14357,N_10201);
or U23923 (N_23923,N_17560,N_16047);
nor U23924 (N_23924,N_13224,N_19118);
and U23925 (N_23925,N_18376,N_17033);
and U23926 (N_23926,N_18371,N_18314);
nand U23927 (N_23927,N_18417,N_19180);
nand U23928 (N_23928,N_11549,N_17034);
or U23929 (N_23929,N_17875,N_15773);
and U23930 (N_23930,N_18462,N_18818);
xnor U23931 (N_23931,N_14833,N_10596);
nand U23932 (N_23932,N_14788,N_11654);
and U23933 (N_23933,N_19939,N_14024);
nor U23934 (N_23934,N_15881,N_17989);
nand U23935 (N_23935,N_11233,N_15182);
nor U23936 (N_23936,N_13020,N_14832);
nand U23937 (N_23937,N_19837,N_10180);
nand U23938 (N_23938,N_13731,N_15608);
or U23939 (N_23939,N_13498,N_13130);
and U23940 (N_23940,N_19312,N_13162);
and U23941 (N_23941,N_14025,N_16564);
xnor U23942 (N_23942,N_19835,N_13313);
and U23943 (N_23943,N_19909,N_17987);
nand U23944 (N_23944,N_11930,N_13465);
nand U23945 (N_23945,N_12084,N_18028);
and U23946 (N_23946,N_12742,N_12386);
xnor U23947 (N_23947,N_18763,N_14450);
nor U23948 (N_23948,N_19430,N_15159);
or U23949 (N_23949,N_19526,N_18074);
and U23950 (N_23950,N_11506,N_10770);
or U23951 (N_23951,N_10551,N_11892);
nor U23952 (N_23952,N_10056,N_13638);
or U23953 (N_23953,N_13944,N_17969);
or U23954 (N_23954,N_11451,N_19130);
nor U23955 (N_23955,N_18724,N_14115);
or U23956 (N_23956,N_17129,N_12643);
xnor U23957 (N_23957,N_13536,N_14437);
xnor U23958 (N_23958,N_16478,N_17995);
nand U23959 (N_23959,N_15384,N_11887);
nand U23960 (N_23960,N_14546,N_16754);
and U23961 (N_23961,N_16320,N_18951);
or U23962 (N_23962,N_11726,N_18836);
nand U23963 (N_23963,N_14944,N_16002);
nor U23964 (N_23964,N_18581,N_15181);
nor U23965 (N_23965,N_13472,N_16267);
or U23966 (N_23966,N_16900,N_12543);
nand U23967 (N_23967,N_17176,N_18411);
nand U23968 (N_23968,N_15649,N_18423);
nand U23969 (N_23969,N_12582,N_12179);
and U23970 (N_23970,N_13164,N_19286);
nand U23971 (N_23971,N_11481,N_10176);
or U23972 (N_23972,N_11260,N_15477);
or U23973 (N_23973,N_14043,N_17271);
nor U23974 (N_23974,N_11784,N_13403);
and U23975 (N_23975,N_12636,N_15841);
and U23976 (N_23976,N_12528,N_17124);
nor U23977 (N_23977,N_15423,N_12811);
or U23978 (N_23978,N_16461,N_17253);
nor U23979 (N_23979,N_11675,N_19732);
and U23980 (N_23980,N_19364,N_18014);
and U23981 (N_23981,N_14942,N_11737);
or U23982 (N_23982,N_19044,N_12787);
and U23983 (N_23983,N_10762,N_12376);
and U23984 (N_23984,N_18929,N_13129);
and U23985 (N_23985,N_17982,N_10912);
and U23986 (N_23986,N_18249,N_11257);
or U23987 (N_23987,N_19568,N_18653);
or U23988 (N_23988,N_13727,N_17172);
nor U23989 (N_23989,N_16340,N_19873);
nor U23990 (N_23990,N_14711,N_17083);
or U23991 (N_23991,N_18949,N_17925);
or U23992 (N_23992,N_17536,N_19883);
nand U23993 (N_23993,N_14030,N_18757);
nand U23994 (N_23994,N_14463,N_18463);
or U23995 (N_23995,N_10776,N_15343);
or U23996 (N_23996,N_10725,N_12527);
nand U23997 (N_23997,N_16926,N_11425);
nor U23998 (N_23998,N_13452,N_16770);
nand U23999 (N_23999,N_17071,N_18881);
nand U24000 (N_24000,N_15450,N_17774);
and U24001 (N_24001,N_15478,N_15196);
nor U24002 (N_24002,N_12639,N_18598);
nor U24003 (N_24003,N_15862,N_10485);
and U24004 (N_24004,N_17052,N_14915);
xnor U24005 (N_24005,N_12589,N_12521);
or U24006 (N_24006,N_11477,N_14837);
and U24007 (N_24007,N_13000,N_18061);
xnor U24008 (N_24008,N_10197,N_12351);
and U24009 (N_24009,N_17497,N_11443);
xor U24010 (N_24010,N_11781,N_17864);
nor U24011 (N_24011,N_17108,N_18527);
or U24012 (N_24012,N_18431,N_17239);
nor U24013 (N_24013,N_11467,N_18299);
nand U24014 (N_24014,N_17202,N_11205);
nand U24015 (N_24015,N_10072,N_18953);
or U24016 (N_24016,N_11312,N_17898);
and U24017 (N_24017,N_12569,N_13893);
or U24018 (N_24018,N_14336,N_10924);
or U24019 (N_24019,N_10100,N_18357);
or U24020 (N_24020,N_13915,N_16663);
and U24021 (N_24021,N_11954,N_11987);
or U24022 (N_24022,N_10435,N_10729);
nor U24023 (N_24023,N_17650,N_13926);
nor U24024 (N_24024,N_11340,N_17490);
nand U24025 (N_24025,N_12633,N_19256);
or U24026 (N_24026,N_13080,N_18719);
and U24027 (N_24027,N_10679,N_14009);
nor U24028 (N_24028,N_17226,N_11982);
nand U24029 (N_24029,N_10952,N_15868);
nand U24030 (N_24030,N_11457,N_10817);
nand U24031 (N_24031,N_13285,N_15842);
or U24032 (N_24032,N_15167,N_10808);
nand U24033 (N_24033,N_11721,N_13874);
nand U24034 (N_24034,N_10321,N_10854);
or U24035 (N_24035,N_14721,N_10603);
or U24036 (N_24036,N_12896,N_12204);
nand U24037 (N_24037,N_18121,N_15675);
nand U24038 (N_24038,N_17453,N_10658);
nand U24039 (N_24039,N_14429,N_14588);
or U24040 (N_24040,N_19016,N_12591);
nand U24041 (N_24041,N_19983,N_11541);
xor U24042 (N_24042,N_15623,N_13331);
xor U24043 (N_24043,N_19494,N_10005);
nor U24044 (N_24044,N_18403,N_19482);
nor U24045 (N_24045,N_10286,N_14912);
nor U24046 (N_24046,N_15300,N_14323);
xor U24047 (N_24047,N_15347,N_18020);
nand U24048 (N_24048,N_17685,N_15531);
or U24049 (N_24049,N_14084,N_18445);
and U24050 (N_24050,N_14379,N_18409);
or U24051 (N_24051,N_12195,N_12231);
and U24052 (N_24052,N_14188,N_16356);
nand U24053 (N_24053,N_11347,N_15445);
nand U24054 (N_24054,N_11548,N_12752);
and U24055 (N_24055,N_10042,N_17556);
nand U24056 (N_24056,N_10521,N_18809);
and U24057 (N_24057,N_11841,N_17748);
or U24058 (N_24058,N_16591,N_18659);
nor U24059 (N_24059,N_14796,N_10397);
or U24060 (N_24060,N_19819,N_12052);
xor U24061 (N_24061,N_11021,N_10266);
nor U24062 (N_24062,N_11489,N_11948);
nor U24063 (N_24063,N_12613,N_18274);
nand U24064 (N_24064,N_11319,N_19135);
nor U24065 (N_24065,N_10588,N_12328);
xnor U24066 (N_24066,N_10649,N_17114);
nor U24067 (N_24067,N_19793,N_12941);
nor U24068 (N_24068,N_19969,N_10857);
or U24069 (N_24069,N_11450,N_12672);
or U24070 (N_24070,N_13502,N_13449);
nor U24071 (N_24071,N_19768,N_10474);
and U24072 (N_24072,N_11314,N_19651);
and U24073 (N_24073,N_17804,N_16271);
and U24074 (N_24074,N_12763,N_19518);
or U24075 (N_24075,N_19303,N_10370);
and U24076 (N_24076,N_19227,N_11394);
nor U24077 (N_24077,N_18142,N_13860);
nor U24078 (N_24078,N_14961,N_13335);
nor U24079 (N_24079,N_10467,N_11775);
or U24080 (N_24080,N_19397,N_17487);
xnor U24081 (N_24081,N_11947,N_13418);
nor U24082 (N_24082,N_17526,N_12607);
or U24083 (N_24083,N_19007,N_10760);
nand U24084 (N_24084,N_10105,N_12560);
xor U24085 (N_24085,N_18792,N_19672);
nor U24086 (N_24086,N_15739,N_15724);
and U24087 (N_24087,N_10465,N_17119);
or U24088 (N_24088,N_17653,N_17702);
xor U24089 (N_24089,N_16361,N_13721);
nor U24090 (N_24090,N_12653,N_11253);
xnor U24091 (N_24091,N_14802,N_15687);
or U24092 (N_24092,N_15368,N_19678);
xnor U24093 (N_24093,N_18829,N_13505);
nor U24094 (N_24094,N_18092,N_11894);
or U24095 (N_24095,N_16191,N_18512);
nand U24096 (N_24096,N_12435,N_18744);
xnor U24097 (N_24097,N_16603,N_12484);
nand U24098 (N_24098,N_18475,N_15331);
nand U24099 (N_24099,N_13070,N_17714);
nand U24100 (N_24100,N_14943,N_17126);
or U24101 (N_24101,N_15867,N_16529);
and U24102 (N_24102,N_13832,N_13835);
and U24103 (N_24103,N_16128,N_12982);
nand U24104 (N_24104,N_15888,N_16223);
xnor U24105 (N_24105,N_16621,N_15760);
and U24106 (N_24106,N_16906,N_14524);
nand U24107 (N_24107,N_15398,N_18317);
and U24108 (N_24108,N_17686,N_19716);
nand U24109 (N_24109,N_14561,N_13756);
nor U24110 (N_24110,N_19949,N_18849);
and U24111 (N_24111,N_19796,N_17708);
or U24112 (N_24112,N_14780,N_10225);
xnor U24113 (N_24113,N_10651,N_11774);
xnor U24114 (N_24114,N_14980,N_16685);
nand U24115 (N_24115,N_10026,N_19563);
nor U24116 (N_24116,N_17797,N_13863);
nor U24117 (N_24117,N_10188,N_12323);
nand U24118 (N_24118,N_10630,N_14256);
nor U24119 (N_24119,N_13991,N_13123);
nand U24120 (N_24120,N_13126,N_13269);
or U24121 (N_24121,N_17979,N_15349);
or U24122 (N_24122,N_16174,N_16823);
and U24123 (N_24123,N_19509,N_18913);
xor U24124 (N_24124,N_16413,N_12526);
or U24125 (N_24125,N_10313,N_15338);
nor U24126 (N_24126,N_19032,N_11459);
and U24127 (N_24127,N_18286,N_11212);
nor U24128 (N_24128,N_16984,N_14387);
or U24129 (N_24129,N_17628,N_12534);
and U24130 (N_24130,N_16662,N_15294);
xnor U24131 (N_24131,N_16088,N_16139);
nand U24132 (N_24132,N_18776,N_18316);
and U24133 (N_24133,N_17763,N_19792);
or U24134 (N_24134,N_13143,N_15940);
nand U24135 (N_24135,N_14015,N_11168);
and U24136 (N_24136,N_16181,N_17540);
nand U24137 (N_24137,N_18521,N_13014);
xnor U24138 (N_24138,N_17198,N_16107);
nor U24139 (N_24139,N_17184,N_19432);
and U24140 (N_24140,N_18389,N_17362);
and U24141 (N_24141,N_14723,N_12445);
or U24142 (N_24142,N_16319,N_19087);
or U24143 (N_24143,N_17354,N_15597);
xor U24144 (N_24144,N_18262,N_18448);
or U24145 (N_24145,N_11510,N_14093);
nor U24146 (N_24146,N_18838,N_15177);
and U24147 (N_24147,N_10006,N_12718);
xor U24148 (N_24148,N_15102,N_13093);
or U24149 (N_24149,N_12159,N_12119);
nor U24150 (N_24150,N_16402,N_15695);
nor U24151 (N_24151,N_15114,N_13560);
nor U24152 (N_24152,N_15386,N_12479);
and U24153 (N_24153,N_17661,N_12584);
nor U24154 (N_24154,N_17007,N_11273);
or U24155 (N_24155,N_17984,N_12669);
nor U24156 (N_24156,N_12570,N_11237);
or U24157 (N_24157,N_18900,N_18917);
nor U24158 (N_24158,N_17877,N_12257);
and U24159 (N_24159,N_19272,N_12629);
or U24160 (N_24160,N_18355,N_10645);
nor U24161 (N_24161,N_11400,N_13467);
or U24162 (N_24162,N_11152,N_17419);
nor U24163 (N_24163,N_19599,N_12283);
nor U24164 (N_24164,N_11011,N_14036);
nor U24165 (N_24165,N_10678,N_11491);
or U24166 (N_24166,N_16277,N_17001);
nand U24167 (N_24167,N_11876,N_12135);
nand U24168 (N_24168,N_11837,N_15259);
xnor U24169 (N_24169,N_14471,N_17004);
nor U24170 (N_24170,N_16672,N_13165);
or U24171 (N_24171,N_19960,N_15538);
nand U24172 (N_24172,N_10434,N_15774);
or U24173 (N_24173,N_15566,N_11744);
nand U24174 (N_24174,N_12989,N_19002);
nor U24175 (N_24175,N_18535,N_17428);
nand U24176 (N_24176,N_12756,N_14639);
nand U24177 (N_24177,N_10317,N_16371);
nand U24178 (N_24178,N_11581,N_13286);
nor U24179 (N_24179,N_16161,N_17131);
nand U24180 (N_24180,N_13888,N_13935);
and U24181 (N_24181,N_13973,N_19964);
or U24182 (N_24182,N_16606,N_12696);
or U24183 (N_24183,N_12291,N_13988);
or U24184 (N_24184,N_14907,N_14560);
nor U24185 (N_24185,N_12815,N_18218);
nand U24186 (N_24186,N_17051,N_15056);
and U24187 (N_24187,N_10381,N_11428);
nand U24188 (N_24188,N_16298,N_13369);
nor U24189 (N_24189,N_14746,N_18055);
and U24190 (N_24190,N_14821,N_13705);
and U24191 (N_24191,N_13151,N_12999);
nor U24192 (N_24192,N_10192,N_14704);
and U24193 (N_24193,N_14145,N_15787);
or U24194 (N_24194,N_17165,N_12015);
nand U24195 (N_24195,N_15419,N_14581);
and U24196 (N_24196,N_11109,N_10861);
nor U24197 (N_24197,N_17028,N_17939);
or U24198 (N_24198,N_17259,N_11614);
nor U24199 (N_24199,N_17882,N_14648);
or U24200 (N_24200,N_19411,N_10419);
and U24201 (N_24201,N_10050,N_18730);
nand U24202 (N_24202,N_11140,N_12846);
or U24203 (N_24203,N_10285,N_13102);
or U24204 (N_24204,N_12751,N_11159);
nand U24205 (N_24205,N_19590,N_19302);
nor U24206 (N_24206,N_10963,N_10184);
nand U24207 (N_24207,N_11180,N_15850);
nand U24208 (N_24208,N_15154,N_14153);
and U24209 (N_24209,N_10941,N_17631);
nor U24210 (N_24210,N_17587,N_16958);
or U24211 (N_24211,N_16742,N_19515);
nor U24212 (N_24212,N_16167,N_19975);
nand U24213 (N_24213,N_11981,N_18509);
nand U24214 (N_24214,N_16991,N_14223);
nand U24215 (N_24215,N_11658,N_14228);
or U24216 (N_24216,N_15809,N_17063);
and U24217 (N_24217,N_18544,N_16645);
nor U24218 (N_24218,N_15663,N_12148);
nand U24219 (N_24219,N_15501,N_12058);
nand U24220 (N_24220,N_17632,N_16092);
and U24221 (N_24221,N_17829,N_14633);
nor U24222 (N_24222,N_11916,N_17364);
nand U24223 (N_24223,N_19080,N_10237);
or U24224 (N_24224,N_14327,N_16293);
or U24225 (N_24225,N_17510,N_19374);
nor U24226 (N_24226,N_15040,N_16221);
nand U24227 (N_24227,N_18356,N_15393);
and U24228 (N_24228,N_18857,N_13619);
and U24229 (N_24229,N_17810,N_13442);
nor U24230 (N_24230,N_16447,N_11704);
and U24231 (N_24231,N_11918,N_19503);
xor U24232 (N_24232,N_14354,N_12601);
or U24233 (N_24233,N_12285,N_17332);
nand U24234 (N_24234,N_11864,N_12603);
nand U24235 (N_24235,N_12741,N_11789);
or U24236 (N_24236,N_14887,N_10165);
nand U24237 (N_24237,N_17501,N_19342);
nor U24238 (N_24238,N_15563,N_13931);
nand U24239 (N_24239,N_16100,N_17753);
xor U24240 (N_24240,N_17392,N_18204);
or U24241 (N_24241,N_18434,N_12541);
nor U24242 (N_24242,N_13501,N_12369);
and U24243 (N_24243,N_19872,N_19912);
or U24244 (N_24244,N_15436,N_10271);
nor U24245 (N_24245,N_10982,N_12979);
nor U24246 (N_24246,N_19558,N_19871);
or U24247 (N_24247,N_10454,N_18064);
nand U24248 (N_24248,N_12789,N_10425);
or U24249 (N_24249,N_12764,N_17545);
xor U24250 (N_24250,N_18675,N_12040);
nor U24251 (N_24251,N_15943,N_15225);
or U24252 (N_24252,N_13226,N_14854);
and U24253 (N_24253,N_17615,N_11098);
or U24254 (N_24254,N_11000,N_10323);
and U24255 (N_24255,N_18888,N_16367);
or U24256 (N_24256,N_19731,N_14693);
or U24257 (N_24257,N_18517,N_16596);
or U24258 (N_24258,N_18079,N_18193);
and U24259 (N_24259,N_18058,N_18038);
nor U24260 (N_24260,N_10516,N_19251);
nand U24261 (N_24261,N_18240,N_17402);
nand U24262 (N_24262,N_19263,N_11524);
nand U24263 (N_24263,N_15490,N_10230);
or U24264 (N_24264,N_11103,N_19924);
nor U24265 (N_24265,N_10934,N_14875);
nand U24266 (N_24266,N_19318,N_11292);
or U24267 (N_24267,N_14722,N_19195);
nand U24268 (N_24268,N_17924,N_16050);
or U24269 (N_24269,N_15214,N_17927);
or U24270 (N_24270,N_17096,N_11265);
and U24271 (N_24271,N_12128,N_17329);
nand U24272 (N_24272,N_11566,N_15217);
nor U24273 (N_24273,N_17850,N_16415);
nand U24274 (N_24274,N_13038,N_15777);
and U24275 (N_24275,N_11798,N_12813);
nand U24276 (N_24276,N_13244,N_17858);
or U24277 (N_24277,N_11557,N_10441);
and U24278 (N_24278,N_14439,N_13880);
nor U24279 (N_24279,N_17602,N_10166);
nand U24280 (N_24280,N_13253,N_11102);
and U24281 (N_24281,N_18561,N_17799);
nor U24282 (N_24282,N_15715,N_11160);
nand U24283 (N_24283,N_15021,N_15029);
and U24284 (N_24284,N_14579,N_11446);
or U24285 (N_24285,N_16378,N_19192);
and U24286 (N_24286,N_19747,N_18369);
nand U24287 (N_24287,N_15245,N_17998);
and U24288 (N_24288,N_14016,N_13158);
nand U24289 (N_24289,N_12454,N_19876);
xnor U24290 (N_24290,N_19259,N_19283);
xor U24291 (N_24291,N_11870,N_19301);
nor U24292 (N_24292,N_15946,N_12939);
and U24293 (N_24293,N_19268,N_19892);
and U24294 (N_24294,N_17013,N_14108);
nand U24295 (N_24295,N_10491,N_12359);
and U24296 (N_24296,N_19540,N_10534);
and U24297 (N_24297,N_15810,N_16570);
or U24298 (N_24298,N_10938,N_11895);
or U24299 (N_24299,N_17022,N_17574);
and U24300 (N_24300,N_15288,N_18522);
or U24301 (N_24301,N_16963,N_13149);
xnor U24302 (N_24302,N_15090,N_11108);
nand U24303 (N_24303,N_18769,N_16772);
nand U24304 (N_24304,N_14737,N_12436);
xnor U24305 (N_24305,N_10560,N_14972);
and U24306 (N_24306,N_17224,N_17761);
or U24307 (N_24307,N_10124,N_18229);
nand U24308 (N_24308,N_15431,N_18333);
and U24309 (N_24309,N_12347,N_17097);
nor U24310 (N_24310,N_17185,N_16432);
nor U24311 (N_24311,N_15055,N_16480);
and U24312 (N_24312,N_17450,N_13399);
nand U24313 (N_24313,N_14700,N_14111);
xnor U24314 (N_24314,N_15359,N_17472);
nand U24315 (N_24315,N_14678,N_12189);
and U24316 (N_24316,N_15116,N_19523);
and U24317 (N_24317,N_14838,N_16312);
or U24318 (N_24318,N_10307,N_11797);
nand U24319 (N_24319,N_17297,N_14063);
nor U24320 (N_24320,N_14400,N_15632);
nand U24321 (N_24321,N_13039,N_16444);
or U24322 (N_24322,N_14052,N_11882);
nand U24323 (N_24323,N_16255,N_12791);
nand U24324 (N_24324,N_12034,N_16052);
xor U24325 (N_24325,N_10301,N_11528);
nor U24326 (N_24326,N_11511,N_12048);
or U24327 (N_24327,N_12097,N_12288);
or U24328 (N_24328,N_14067,N_16787);
nor U24329 (N_24329,N_12103,N_16035);
and U24330 (N_24330,N_10923,N_13956);
xor U24331 (N_24331,N_12585,N_19257);
and U24332 (N_24332,N_15775,N_19940);
xor U24333 (N_24333,N_19326,N_19958);
nor U24334 (N_24334,N_18049,N_12774);
or U24335 (N_24335,N_17801,N_17358);
and U24336 (N_24336,N_11724,N_12552);
nand U24337 (N_24337,N_16790,N_17994);
or U24338 (N_24338,N_17068,N_11321);
or U24339 (N_24339,N_19228,N_11761);
or U24340 (N_24340,N_10629,N_18705);
and U24341 (N_24341,N_11080,N_11889);
and U24342 (N_24342,N_19129,N_10356);
or U24343 (N_24343,N_16911,N_17928);
and U24344 (N_24344,N_13426,N_10738);
and U24345 (N_24345,N_15763,N_19507);
nand U24346 (N_24346,N_15848,N_10436);
nand U24347 (N_24347,N_12518,N_10778);
or U24348 (N_24348,N_17494,N_17606);
or U24349 (N_24349,N_10269,N_12500);
nor U24350 (N_24350,N_15733,N_15175);
and U24351 (N_24351,N_14451,N_15404);
nor U24352 (N_24352,N_19046,N_10796);
nor U24353 (N_24353,N_19125,N_19051);
or U24354 (N_24354,N_14430,N_17424);
nand U24355 (N_24355,N_18405,N_12778);
nor U24356 (N_24356,N_11803,N_17915);
nand U24357 (N_24357,N_10430,N_10584);
and U24358 (N_24358,N_11796,N_19350);
nor U24359 (N_24359,N_13411,N_18595);
and U24360 (N_24360,N_13916,N_19853);
nand U24361 (N_24361,N_11356,N_16905);
nand U24362 (N_24362,N_15896,N_17734);
nor U24363 (N_24363,N_11836,N_13672);
or U24364 (N_24364,N_10095,N_15460);
nand U24365 (N_24365,N_12905,N_11378);
nor U24366 (N_24366,N_12475,N_19491);
or U24367 (N_24367,N_11682,N_19278);
or U24368 (N_24368,N_14173,N_18655);
xnor U24369 (N_24369,N_19139,N_12556);
or U24370 (N_24370,N_17890,N_11412);
or U24371 (N_24371,N_17817,N_11942);
nor U24372 (N_24372,N_14864,N_16090);
and U24373 (N_24373,N_13580,N_17565);
or U24374 (N_24374,N_13170,N_14345);
nand U24375 (N_24375,N_16442,N_18523);
or U24376 (N_24376,N_17078,N_19095);
nor U24377 (N_24377,N_19291,N_17138);
and U24378 (N_24378,N_12173,N_14762);
nand U24379 (N_24379,N_12202,N_10549);
or U24380 (N_24380,N_15038,N_10245);
or U24381 (N_24381,N_10142,N_14806);
xnor U24382 (N_24382,N_15929,N_18784);
nand U24383 (N_24383,N_13454,N_19572);
nor U24384 (N_24384,N_11065,N_15273);
or U24385 (N_24385,N_19674,N_12293);
nand U24386 (N_24386,N_17050,N_11127);
nand U24387 (N_24387,N_14042,N_17651);
nor U24388 (N_24388,N_13374,N_10178);
nor U24389 (N_24389,N_11888,N_19897);
xnor U24390 (N_24390,N_17755,N_16195);
and U24391 (N_24391,N_17547,N_10582);
or U24392 (N_24392,N_10318,N_15822);
and U24393 (N_24393,N_10421,N_19557);
xor U24394 (N_24394,N_12538,N_17863);
nand U24395 (N_24395,N_15684,N_12455);
or U24396 (N_24396,N_10092,N_14866);
and U24397 (N_24397,N_12659,N_14697);
nor U24398 (N_24398,N_10819,N_14086);
nor U24399 (N_24399,N_16520,N_11637);
or U24400 (N_24400,N_16805,N_14022);
nor U24401 (N_24401,N_19401,N_12889);
or U24402 (N_24402,N_15559,N_16095);
and U24403 (N_24403,N_10240,N_17489);
nor U24404 (N_24404,N_14092,N_13986);
nor U24405 (N_24405,N_15577,N_14922);
nand U24406 (N_24406,N_12682,N_10267);
nor U24407 (N_24407,N_13898,N_17458);
nand U24408 (N_24408,N_16652,N_13414);
and U24409 (N_24409,N_17654,N_10727);
nand U24410 (N_24410,N_12833,N_15441);
nand U24411 (N_24411,N_10216,N_14740);
xor U24412 (N_24412,N_19221,N_12626);
and U24413 (N_24413,N_16383,N_14269);
nand U24414 (N_24414,N_19712,N_12566);
and U24415 (N_24415,N_18245,N_12478);
nand U24416 (N_24416,N_11799,N_12405);
nor U24417 (N_24417,N_17869,N_19194);
xnor U24418 (N_24418,N_16065,N_13790);
and U24419 (N_24419,N_12992,N_15546);
or U24420 (N_24420,N_17784,N_15831);
nor U24421 (N_24421,N_10561,N_18794);
nor U24422 (N_24422,N_18370,N_12006);
nor U24423 (N_24423,N_17285,N_16681);
nand U24424 (N_24424,N_18177,N_14231);
and U24425 (N_24425,N_15165,N_13294);
nand U24426 (N_24426,N_11800,N_10210);
nor U24427 (N_24427,N_19202,N_16648);
xnor U24428 (N_24428,N_11013,N_18863);
or U24429 (N_24429,N_10517,N_16705);
nand U24430 (N_24430,N_13480,N_17543);
xnor U24431 (N_24431,N_12026,N_10565);
and U24432 (N_24432,N_18172,N_10489);
and U24433 (N_24433,N_15286,N_12401);
nand U24434 (N_24434,N_16638,N_19243);
nor U24435 (N_24435,N_14623,N_14730);
nor U24436 (N_24436,N_18302,N_17943);
nor U24437 (N_24437,N_19108,N_14010);
and U24438 (N_24438,N_17349,N_18579);
xnor U24439 (N_24439,N_14898,N_11328);
nand U24440 (N_24440,N_12273,N_16523);
or U24441 (N_24441,N_15050,N_11329);
or U24442 (N_24442,N_10341,N_12568);
nor U24443 (N_24443,N_12415,N_17649);
nor U24444 (N_24444,N_19435,N_19504);
or U24445 (N_24445,N_16798,N_13668);
nand U24446 (N_24446,N_17893,N_14600);
nand U24447 (N_24447,N_18212,N_19690);
xor U24448 (N_24448,N_16194,N_16000);
nor U24449 (N_24449,N_12932,N_18640);
or U24450 (N_24450,N_19551,N_15920);
and U24451 (N_24451,N_18343,N_10088);
nand U24452 (N_24452,N_17802,N_10835);
nand U24453 (N_24453,N_11754,N_13125);
nor U24454 (N_24454,N_14483,N_16747);
nand U24455 (N_24455,N_12236,N_15082);
xnor U24456 (N_24456,N_11232,N_17183);
nand U24457 (N_24457,N_10687,N_17705);
nor U24458 (N_24458,N_17883,N_15719);
xnor U24459 (N_24459,N_19323,N_12917);
and U24460 (N_24460,N_15071,N_17236);
or U24461 (N_24461,N_19804,N_11745);
nand U24462 (N_24462,N_15593,N_13712);
xor U24463 (N_24463,N_18577,N_14218);
or U24464 (N_24464,N_13199,N_17567);
nor U24465 (N_24465,N_19356,N_19119);
xnor U24466 (N_24466,N_11339,N_19920);
and U24467 (N_24467,N_10869,N_13042);
or U24468 (N_24468,N_13284,N_16264);
or U24469 (N_24469,N_15057,N_13941);
and U24470 (N_24470,N_16668,N_10693);
nor U24471 (N_24471,N_14619,N_17040);
nor U24472 (N_24472,N_18054,N_12198);
nor U24473 (N_24473,N_12887,N_13703);
nand U24474 (N_24474,N_14396,N_17164);
or U24475 (N_24475,N_12950,N_13679);
or U24476 (N_24476,N_19289,N_14652);
nor U24477 (N_24477,N_12176,N_17972);
or U24478 (N_24478,N_11199,N_16804);
or U24479 (N_24479,N_17408,N_18220);
nor U24480 (N_24480,N_13193,N_15272);
and U24481 (N_24481,N_12114,N_18230);
or U24482 (N_24482,N_19013,N_14747);
nor U24483 (N_24483,N_13483,N_13304);
nor U24484 (N_24484,N_12948,N_16338);
nand U24485 (N_24485,N_12100,N_15068);
and U24486 (N_24486,N_17174,N_18552);
or U24487 (N_24487,N_14068,N_17770);
nand U24488 (N_24488,N_12854,N_17279);
nand U24489 (N_24489,N_14784,N_16056);
and U24490 (N_24490,N_14632,N_17611);
or U24491 (N_24491,N_16943,N_19858);
nor U24492 (N_24492,N_12129,N_16680);
nor U24493 (N_24493,N_15607,N_12716);
or U24494 (N_24494,N_19727,N_13570);
and U24495 (N_24495,N_11038,N_14688);
or U24496 (N_24496,N_17061,N_10917);
nor U24497 (N_24497,N_18822,N_17059);
xor U24498 (N_24498,N_14920,N_12162);
xor U24499 (N_24499,N_15558,N_10064);
and U24500 (N_24500,N_18530,N_11075);
and U24501 (N_24501,N_11274,N_17152);
and U24502 (N_24502,N_16314,N_18241);
nor U24503 (N_24503,N_15084,N_12817);
xnor U24504 (N_24504,N_19261,N_13864);
and U24505 (N_24505,N_11248,N_14058);
nor U24506 (N_24506,N_11625,N_15595);
or U24507 (N_24507,N_12971,N_13104);
nand U24508 (N_24508,N_13698,N_18138);
xnor U24509 (N_24509,N_14754,N_11592);
or U24510 (N_24510,N_10949,N_11458);
or U24511 (N_24511,N_17828,N_14962);
nand U24512 (N_24512,N_17394,N_13276);
nand U24513 (N_24513,N_18934,N_12773);
and U24514 (N_24514,N_10172,N_19328);
nand U24515 (N_24515,N_10104,N_18105);
nand U24516 (N_24516,N_14994,N_11327);
and U24517 (N_24517,N_17662,N_17169);
or U24518 (N_24518,N_12641,N_13546);
and U24519 (N_24519,N_16066,N_13354);
nor U24520 (N_24520,N_15435,N_17045);
or U24521 (N_24521,N_12032,N_10845);
xor U24522 (N_24522,N_19444,N_11234);
xnor U24523 (N_24523,N_11393,N_11191);
and U24524 (N_24524,N_15244,N_11028);
nand U24525 (N_24525,N_17029,N_11696);
and U24526 (N_24526,N_18139,N_18860);
and U24527 (N_24527,N_12279,N_11525);
and U24528 (N_24528,N_19062,N_15094);
nor U24529 (N_24529,N_15238,N_18129);
or U24530 (N_24530,N_11163,N_16364);
nor U24531 (N_24531,N_14514,N_14110);
nor U24532 (N_24532,N_11288,N_12892);
xnor U24533 (N_24533,N_13289,N_11161);
nand U24534 (N_24534,N_16756,N_13996);
nor U24535 (N_24535,N_16237,N_13871);
nand U24536 (N_24536,N_14308,N_11396);
and U24537 (N_24537,N_15113,N_14908);
nand U24538 (N_24538,N_17951,N_11371);
nand U24539 (N_24539,N_10291,N_14089);
or U24540 (N_24540,N_14399,N_17295);
and U24541 (N_24541,N_12665,N_14782);
xor U24542 (N_24542,N_11665,N_16424);
nand U24543 (N_24543,N_10880,N_19961);
and U24544 (N_24544,N_13732,N_10349);
and U24545 (N_24545,N_15791,N_19519);
and U24546 (N_24546,N_15011,N_18039);
or U24547 (N_24547,N_13651,N_11078);
and U24548 (N_24548,N_11189,N_13967);
or U24549 (N_24549,N_16164,N_13077);
or U24550 (N_24550,N_14889,N_10814);
or U24551 (N_24551,N_12123,N_12858);
and U24552 (N_24552,N_18301,N_16359);
nor U24553 (N_24553,N_16027,N_10437);
and U24554 (N_24554,N_19022,N_17820);
nor U24555 (N_24555,N_12695,N_10438);
and U24556 (N_24556,N_16326,N_14280);
and U24557 (N_24557,N_11647,N_13021);
nand U24558 (N_24558,N_11219,N_12805);
nand U24559 (N_24559,N_19078,N_13146);
and U24560 (N_24560,N_14113,N_10827);
and U24561 (N_24561,N_14675,N_10449);
and U24562 (N_24562,N_16750,N_15026);
or U24563 (N_24563,N_11442,N_10685);
nor U24564 (N_24564,N_13989,N_19009);
or U24565 (N_24565,N_10221,N_14325);
or U24566 (N_24566,N_13801,N_13325);
nor U24567 (N_24567,N_13553,N_13605);
or U24568 (N_24568,N_12226,N_18824);
and U24569 (N_24569,N_19204,N_12482);
nand U24570 (N_24570,N_12217,N_19606);
nor U24571 (N_24571,N_15381,N_15486);
and U24572 (N_24572,N_15199,N_16465);
xnor U24573 (N_24573,N_10393,N_11578);
nand U24574 (N_24574,N_17786,N_13108);
nor U24575 (N_24575,N_14339,N_17005);
nor U24576 (N_24576,N_17532,N_13524);
or U24577 (N_24577,N_19711,N_17682);
or U24578 (N_24578,N_11596,N_17674);
or U24579 (N_24579,N_11965,N_10950);
and U24580 (N_24580,N_11297,N_18735);
nor U24581 (N_24581,N_17707,N_12474);
xnor U24582 (N_24582,N_18694,N_13891);
nor U24583 (N_24583,N_18827,N_15897);
nand U24584 (N_24584,N_17417,N_16248);
nand U24585 (N_24585,N_13006,N_14434);
or U24586 (N_24586,N_10598,N_19508);
nand U24587 (N_24587,N_17852,N_15838);
nand U24588 (N_24588,N_16305,N_14954);
nand U24589 (N_24589,N_17500,N_12408);
and U24590 (N_24590,N_18374,N_18811);
nand U24591 (N_24591,N_16227,N_10662);
nor U24592 (N_24592,N_14098,N_11117);
nor U24593 (N_24593,N_14373,N_18382);
or U24594 (N_24594,N_14204,N_15012);
or U24595 (N_24595,N_14019,N_15346);
nor U24596 (N_24596,N_12911,N_10314);
or U24597 (N_24597,N_12266,N_10483);
and U24598 (N_24598,N_18576,N_15432);
and U24599 (N_24599,N_13830,N_16725);
nand U24600 (N_24600,N_18882,N_17938);
nor U24601 (N_24601,N_16511,N_17217);
or U24602 (N_24602,N_12107,N_13550);
nand U24603 (N_24603,N_15382,N_19987);
nor U24604 (N_24604,N_13497,N_15893);
and U24605 (N_24605,N_13271,N_18452);
or U24606 (N_24606,N_16310,N_16106);
or U24607 (N_24607,N_16999,N_11617);
nand U24608 (N_24608,N_15754,N_18183);
or U24609 (N_24609,N_12912,N_11352);
nor U24610 (N_24610,N_15656,N_12820);
nor U24611 (N_24611,N_16952,N_10351);
or U24612 (N_24612,N_10212,N_15447);
xnor U24613 (N_24613,N_10289,N_13359);
nand U24614 (N_24614,N_14874,N_15818);
nor U24615 (N_24615,N_18077,N_11061);
nand U24616 (N_24616,N_14158,N_18206);
nor U24617 (N_24617,N_17466,N_19398);
nand U24618 (N_24618,N_19477,N_13479);
or U24619 (N_24619,N_18942,N_15287);
nor U24620 (N_24620,N_17449,N_13105);
or U24621 (N_24621,N_17811,N_11343);
nor U24622 (N_24622,N_15219,N_15449);
xnor U24623 (N_24623,N_13762,N_12935);
or U24624 (N_24624,N_14661,N_17706);
nand U24625 (N_24625,N_15020,N_12433);
nand U24626 (N_24626,N_12250,N_11934);
and U24627 (N_24627,N_18965,N_15804);
nor U24628 (N_24628,N_19285,N_13899);
and U24629 (N_24629,N_13696,N_10747);
nand U24630 (N_24630,N_14892,N_16257);
and U24631 (N_24631,N_10879,N_18698);
and U24632 (N_24632,N_14748,N_17021);
nand U24633 (N_24633,N_18852,N_10305);
nor U24634 (N_24634,N_17578,N_11973);
nand U24635 (N_24635,N_18447,N_10233);
or U24636 (N_24636,N_15889,N_14031);
and U24637 (N_24637,N_14085,N_17187);
nor U24638 (N_24638,N_12519,N_13719);
nor U24639 (N_24639,N_10055,N_10692);
nor U24640 (N_24640,N_15507,N_12781);
or U24641 (N_24641,N_17742,N_14508);
and U24642 (N_24642,N_18166,N_16697);
nor U24643 (N_24643,N_11998,N_12232);
and U24644 (N_24644,N_16218,N_10473);
or U24645 (N_24645,N_12712,N_11141);
nor U24646 (N_24646,N_15639,N_19132);
or U24647 (N_24647,N_18486,N_17886);
and U24648 (N_24648,N_12450,N_19096);
or U24649 (N_24649,N_15996,N_11381);
and U24650 (N_24650,N_10590,N_16698);
nor U24651 (N_24651,N_13438,N_15330);
nor U24652 (N_24652,N_10471,N_15158);
nand U24653 (N_24653,N_19575,N_12356);
nand U24654 (N_24654,N_15517,N_18391);
and U24655 (N_24655,N_17132,N_17437);
nand U24656 (N_24656,N_19752,N_16843);
or U24657 (N_24657,N_16547,N_19803);
nor U24658 (N_24658,N_11911,N_10872);
or U24659 (N_24659,N_17527,N_19974);
xor U24660 (N_24660,N_19728,N_16321);
or U24661 (N_24661,N_10253,N_10148);
nor U24662 (N_24662,N_18853,N_15786);
nand U24663 (N_24663,N_17160,N_12280);
nand U24664 (N_24664,N_18696,N_13645);
and U24665 (N_24665,N_13559,N_17177);
nand U24666 (N_24666,N_14605,N_14456);
nor U24667 (N_24667,N_15482,N_15930);
and U24668 (N_24668,N_11254,N_13251);
nand U24669 (N_24669,N_17521,N_19217);
or U24670 (N_24670,N_12140,N_10082);
nand U24671 (N_24671,N_16923,N_18327);
nor U24672 (N_24672,N_17884,N_13939);
and U24673 (N_24673,N_18842,N_13229);
nand U24674 (N_24674,N_17960,N_14491);
nand U24675 (N_24675,N_19989,N_11351);
nand U24676 (N_24676,N_12057,N_13345);
or U24677 (N_24677,N_15542,N_13318);
and U24678 (N_24678,N_13054,N_19039);
or U24679 (N_24679,N_14106,N_18003);
and U24680 (N_24680,N_10767,N_10570);
nand U24681 (N_24681,N_13071,N_13596);
or U24682 (N_24682,N_11713,N_10907);
and U24683 (N_24683,N_11526,N_17896);
nor U24684 (N_24684,N_17055,N_17945);
and U24685 (N_24685,N_18185,N_13476);
nor U24686 (N_24686,N_10583,N_14985);
nor U24687 (N_24687,N_15224,N_17149);
nand U24688 (N_24688,N_18878,N_11685);
xor U24689 (N_24689,N_13755,N_19770);
nor U24690 (N_24690,N_17345,N_17916);
nor U24691 (N_24691,N_19729,N_19571);
nand U24692 (N_24692,N_18855,N_17043);
nor U24693 (N_24693,N_11531,N_17210);
or U24694 (N_24694,N_12877,N_15630);
xnor U24695 (N_24695,N_14843,N_18845);
or U24696 (N_24696,N_18141,N_12996);
nand U24697 (N_24697,N_12492,N_12511);
nor U24698 (N_24698,N_19680,N_17211);
and U24699 (N_24699,N_19112,N_16561);
and U24700 (N_24700,N_11322,N_10140);
or U24701 (N_24701,N_18501,N_12737);
and U24702 (N_24702,N_13512,N_13883);
nor U24703 (N_24703,N_14406,N_11480);
or U24704 (N_24704,N_12981,N_14628);
and U24705 (N_24705,N_12072,N_12599);
or U24706 (N_24706,N_14993,N_14100);
nor U24707 (N_24707,N_13854,N_16975);
nor U24708 (N_24708,N_18709,N_14958);
xor U24709 (N_24709,N_15911,N_14292);
or U24710 (N_24710,N_17338,N_12574);
and U24711 (N_24711,N_15306,N_18840);
or U24712 (N_24712,N_17341,N_17019);
or U24713 (N_24713,N_17731,N_17665);
nor U24714 (N_24714,N_19282,N_10979);
xor U24715 (N_24715,N_18796,N_17933);
xor U24716 (N_24716,N_18466,N_17009);
nand U24717 (N_24717,N_14848,N_10620);
nand U24718 (N_24718,N_14795,N_15145);
and U24719 (N_24719,N_19746,N_17845);
and U24720 (N_24720,N_15963,N_12276);
nor U24721 (N_24721,N_15973,N_16692);
nor U24722 (N_24722,N_18352,N_16121);
and U24723 (N_24723,N_19102,N_12967);
nand U24724 (N_24724,N_11575,N_12136);
or U24725 (N_24725,N_10633,N_18718);
nor U24726 (N_24726,N_13924,N_18813);
and U24727 (N_24727,N_12801,N_12772);
nand U24728 (N_24728,N_19801,N_14913);
or U24729 (N_24729,N_19208,N_16473);
or U24730 (N_24730,N_16207,N_18041);
xor U24731 (N_24731,N_16630,N_14658);
nor U24732 (N_24732,N_12054,N_11600);
or U24733 (N_24733,N_14584,N_15837);
nor U24734 (N_24734,N_19382,N_13101);
and U24735 (N_24735,N_18150,N_15892);
xor U24736 (N_24736,N_19881,N_10162);
and U24737 (N_24737,N_15574,N_19472);
nand U24738 (N_24738,N_15299,N_13453);
nor U24739 (N_24739,N_10595,N_13716);
and U24740 (N_24740,N_11604,N_11079);
or U24741 (N_24741,N_15516,N_14910);
nand U24742 (N_24742,N_12239,N_10542);
or U24743 (N_24743,N_14881,N_15142);
xnor U24744 (N_24744,N_16583,N_17353);
nand U24745 (N_24745,N_14329,N_16101);
xor U24746 (N_24746,N_10157,N_11868);
nand U24747 (N_24747,N_14880,N_16976);
or U24748 (N_24748,N_17837,N_17669);
nor U24749 (N_24749,N_11554,N_10152);
or U24750 (N_24750,N_10631,N_12942);
and U24751 (N_24751,N_15673,N_19465);
and U24752 (N_24752,N_11899,N_13355);
nor U24753 (N_24753,N_11953,N_18044);
and U24754 (N_24754,N_12683,N_11748);
or U24755 (N_24755,N_16433,N_10919);
nor U24756 (N_24756,N_15808,N_17094);
or U24757 (N_24757,N_13606,N_11283);
or U24758 (N_24758,N_10239,N_14413);
nand U24759 (N_24759,N_13683,N_15682);
and U24760 (N_24760,N_19827,N_16811);
nand U24761 (N_24761,N_13344,N_12747);
xor U24762 (N_24762,N_13273,N_12430);
nand U24763 (N_24763,N_12007,N_10206);
or U24764 (N_24764,N_17856,N_18308);
nand U24765 (N_24765,N_19362,N_12211);
and U24766 (N_24766,N_13435,N_14592);
nor U24767 (N_24767,N_16460,N_18687);
and U24768 (N_24768,N_17620,N_14930);
or U24769 (N_24769,N_13972,N_16710);
nor U24770 (N_24770,N_10337,N_10715);
and U24771 (N_24771,N_11591,N_18227);
and U24772 (N_24772,N_14337,N_17139);
or U24773 (N_24773,N_19811,N_13979);
or U24774 (N_24774,N_19833,N_18288);
nor U24775 (N_24775,N_10432,N_15062);
and U24776 (N_24776,N_16049,N_15466);
or U24777 (N_24777,N_13641,N_16450);
nand U24778 (N_24778,N_16283,N_13475);
nor U24779 (N_24779,N_15790,N_11099);
nand U24780 (N_24780,N_19189,N_15383);
or U24781 (N_24781,N_14390,N_13281);
and U24782 (N_24782,N_13840,N_16427);
or U24783 (N_24783,N_19834,N_13026);
and U24784 (N_24784,N_18060,N_14402);
nor U24785 (N_24785,N_19786,N_10182);
or U24786 (N_24786,N_13040,N_17317);
nor U24787 (N_24787,N_15513,N_19755);
and U24788 (N_24788,N_16269,N_10855);
or U24789 (N_24789,N_19487,N_19315);
nand U24790 (N_24790,N_13752,N_15864);
and U24791 (N_24791,N_14135,N_17312);
nor U24792 (N_24792,N_11955,N_14925);
or U24793 (N_24793,N_13723,N_19010);
and U24794 (N_24794,N_14710,N_12254);
nor U24795 (N_24795,N_16854,N_12882);
nand U24796 (N_24796,N_19173,N_15729);
or U24797 (N_24797,N_10802,N_17156);
nor U24798 (N_24798,N_17436,N_14536);
nand U24799 (N_24799,N_13953,N_18482);
nor U24800 (N_24800,N_17569,N_19347);
xor U24801 (N_24801,N_12033,N_10986);
or U24802 (N_24802,N_10700,N_13257);
and U24803 (N_24803,N_15586,N_17818);
nor U24804 (N_24804,N_10494,N_17306);
nor U24805 (N_24805,N_13242,N_12590);
xnor U24806 (N_24806,N_14551,N_16534);
nor U24807 (N_24807,N_13985,N_17825);
nor U24808 (N_24808,N_13770,N_11056);
nand U24809 (N_24809,N_13499,N_10149);
xnor U24810 (N_24810,N_15365,N_14816);
or U24811 (N_24811,N_14432,N_14738);
or U24812 (N_24812,N_17576,N_12444);
and U24813 (N_24813,N_16122,N_13035);
nor U24814 (N_24814,N_15426,N_18528);
and U24815 (N_24815,N_19814,N_19079);
xor U24816 (N_24816,N_12158,N_18747);
nand U24817 (N_24817,N_14020,N_14214);
or U24818 (N_24818,N_15579,N_15282);
and U24819 (N_24819,N_14891,N_11855);
or U24820 (N_24820,N_15807,N_15757);
nand U24821 (N_24821,N_19511,N_16780);
and U24822 (N_24822,N_15174,N_10680);
nor U24823 (N_24823,N_14527,N_16142);
and U24824 (N_24824,N_13952,N_16925);
nand U24825 (N_24825,N_13914,N_18741);
nand U24826 (N_24826,N_10654,N_13600);
xnor U24827 (N_24827,N_10554,N_13783);
or U24828 (N_24828,N_15015,N_12019);
nor U24829 (N_24829,N_14412,N_16309);
nor U24830 (N_24830,N_18284,N_18821);
or U24831 (N_24831,N_10735,N_13303);
and U24832 (N_24832,N_12060,N_13795);
nand U24833 (N_24833,N_14026,N_12174);
or U24834 (N_24834,N_16439,N_18255);
or U24835 (N_24835,N_17000,N_11860);
nor U24836 (N_24836,N_10710,N_10144);
nand U24837 (N_24837,N_16459,N_14393);
nand U24838 (N_24838,N_14823,N_14991);
or U24839 (N_24839,N_17769,N_19932);
nor U24840 (N_24840,N_19965,N_17025);
and U24841 (N_24841,N_13558,N_11447);
or U24842 (N_24842,N_14008,N_19422);
nand U24843 (N_24843,N_12676,N_14744);
nand U24844 (N_24844,N_19545,N_12262);
and U24845 (N_24845,N_10573,N_18589);
and U24846 (N_24846,N_19150,N_10173);
and U24847 (N_24847,N_19877,N_10111);
or U24848 (N_24848,N_14174,N_17391);
xnor U24849 (N_24849,N_10065,N_14819);
or U24850 (N_24850,N_14070,N_14495);
nor U24851 (N_24851,N_15058,N_14525);
and U24852 (N_24852,N_10617,N_12790);
xor U24853 (N_24853,N_11884,N_17694);
or U24854 (N_24854,N_12873,N_13349);
or U24855 (N_24855,N_16601,N_17390);
and U24856 (N_24856,N_15136,N_16829);
or U24857 (N_24857,N_16774,N_11634);
nand U24858 (N_24858,N_19309,N_13615);
nor U24859 (N_24859,N_11792,N_12705);
nand U24860 (N_24860,N_15941,N_19424);
nor U24861 (N_24861,N_11217,N_11502);
nand U24862 (N_24862,N_15800,N_10748);
nand U24863 (N_24863,N_16946,N_11819);
nand U24864 (N_24864,N_13885,N_19252);
nor U24865 (N_24865,N_18957,N_13714);
nor U24866 (N_24866,N_19825,N_12733);
and U24867 (N_24867,N_16966,N_15063);
and U24868 (N_24868,N_17227,N_17053);
xnor U24869 (N_24869,N_14210,N_17566);
or U24870 (N_24870,N_12298,N_18578);
nor U24871 (N_24871,N_18564,N_13653);
nor U24872 (N_24872,N_12860,N_17378);
or U24873 (N_24873,N_10235,N_13306);
and U24874 (N_24874,N_19525,N_12602);
nor U24875 (N_24875,N_19943,N_13131);
xnor U24876 (N_24876,N_10932,N_11313);
nor U24877 (N_24877,N_15496,N_19314);
or U24878 (N_24878,N_12869,N_12777);
or U24879 (N_24879,N_13882,N_14378);
nor U24880 (N_24880,N_17622,N_15667);
and U24881 (N_24881,N_11795,N_11164);
or U24882 (N_24882,N_11937,N_10552);
or U24883 (N_24883,N_18203,N_12697);
nand U24884 (N_24884,N_12038,N_18656);
or U24885 (N_24885,N_11404,N_10822);
nand U24886 (N_24886,N_12608,N_11235);
xnor U24887 (N_24887,N_10763,N_19522);
or U24888 (N_24888,N_18700,N_19772);
and U24889 (N_24889,N_11402,N_13086);
xnor U24890 (N_24890,N_10742,N_10138);
nor U24891 (N_24891,N_14800,N_12448);
or U24892 (N_24892,N_17058,N_13508);
nor U24893 (N_24893,N_16962,N_12970);
nand U24894 (N_24894,N_16226,N_10472);
nand U24895 (N_24895,N_12956,N_13095);
or U24896 (N_24896,N_17272,N_13492);
nand U24897 (N_24897,N_17269,N_19378);
or U24898 (N_24898,N_17379,N_13404);
nor U24899 (N_24899,N_15415,N_15283);
nand U24900 (N_24900,N_14965,N_16137);
xor U24901 (N_24901,N_16011,N_13212);
or U24902 (N_24902,N_19840,N_13388);
xnor U24903 (N_24903,N_13336,N_16894);
and U24904 (N_24904,N_15127,N_13658);
nor U24905 (N_24905,N_14596,N_16689);
or U24906 (N_24906,N_10829,N_13845);
and U24907 (N_24907,N_10479,N_11296);
nor U24908 (N_24908,N_15765,N_14840);
nor U24909 (N_24909,N_17986,N_12577);
nand U24910 (N_24910,N_13115,N_17485);
nor U24911 (N_24911,N_15651,N_14626);
and U24912 (N_24912,N_15508,N_19474);
and U24913 (N_24913,N_15411,N_19338);
nor U24914 (N_24914,N_14152,N_19031);
or U24915 (N_24915,N_10078,N_12968);
or U24916 (N_24916,N_19427,N_18161);
xnor U24917 (N_24917,N_14476,N_10428);
and U24918 (N_24918,N_18562,N_10447);
nand U24919 (N_24919,N_16505,N_16497);
or U24920 (N_24920,N_19245,N_14911);
or U24921 (N_24921,N_11500,N_14003);
or U24922 (N_24922,N_19334,N_13584);
nor U24923 (N_24923,N_11838,N_13287);
nand U24924 (N_24924,N_11808,N_16768);
or U24925 (N_24925,N_14176,N_12551);
nand U24926 (N_24926,N_10503,N_10804);
and U24927 (N_24927,N_18924,N_15826);
or U24928 (N_24928,N_15013,N_13805);
nand U24929 (N_24929,N_17522,N_10753);
and U24930 (N_24930,N_16930,N_17225);
nor U24931 (N_24931,N_10312,N_18554);
nand U24932 (N_24932,N_14585,N_12795);
and U24933 (N_24933,N_14066,N_16650);
nor U24934 (N_24934,N_19493,N_15909);
nand U24935 (N_24935,N_17713,N_16785);
and U24936 (N_24936,N_19978,N_12269);
or U24937 (N_24937,N_14381,N_15004);
nor U24938 (N_24938,N_17625,N_11583);
nand U24939 (N_24939,N_10411,N_12502);
xnor U24940 (N_24940,N_11650,N_16693);
or U24941 (N_24941,N_14918,N_19438);
and U24942 (N_24942,N_14674,N_10930);
or U24943 (N_24943,N_18867,N_16881);
nor U24944 (N_24944,N_17923,N_18364);
and U24945 (N_24945,N_15391,N_17773);
or U24946 (N_24946,N_12766,N_19373);
and U24947 (N_24947,N_17044,N_10769);
nor U24948 (N_24948,N_17563,N_14295);
nand U24949 (N_24949,N_14767,N_13792);
nand U24950 (N_24950,N_12467,N_12428);
and U24951 (N_24951,N_19878,N_19589);
nor U24952 (N_24952,N_10527,N_11012);
or U24953 (N_24953,N_12512,N_17780);
and U24954 (N_24954,N_17736,N_15292);
nor U24955 (N_24955,N_10168,N_10214);
nor U24956 (N_24956,N_13970,N_11702);
or U24957 (N_24957,N_13764,N_12711);
nand U24958 (N_24958,N_18007,N_12079);
and U24959 (N_24959,N_11083,N_10946);
nor U24960 (N_24960,N_14371,N_13177);
or U24961 (N_24961,N_18970,N_13907);
and U24962 (N_24962,N_10051,N_10052);
xor U24963 (N_24963,N_11100,N_10252);
or U24964 (N_24964,N_10457,N_16614);
xor U24965 (N_24965,N_11414,N_10079);
nor U24966 (N_24966,N_13490,N_16554);
or U24967 (N_24967,N_15571,N_18839);
nand U24968 (N_24968,N_12277,N_10392);
nand U24969 (N_24969,N_10615,N_17406);
or U24970 (N_24970,N_11513,N_19107);
and U24971 (N_24971,N_17018,N_16879);
xor U24972 (N_24972,N_15609,N_14103);
nand U24973 (N_24973,N_13911,N_15824);
nand U24974 (N_24974,N_15446,N_14199);
nor U24975 (N_24975,N_13614,N_14752);
or U24976 (N_24976,N_16506,N_16247);
or U24977 (N_24977,N_14099,N_19088);
nand U24978 (N_24978,N_13607,N_14332);
nand U24979 (N_24979,N_13207,N_12271);
nor U24980 (N_24980,N_17944,N_12354);
xor U24981 (N_24981,N_15494,N_13053);
and U24982 (N_24982,N_19639,N_19656);
and U24983 (N_24983,N_13317,N_19019);
xor U24984 (N_24984,N_16187,N_13309);
nand U24985 (N_24985,N_16258,N_17209);
and U24986 (N_24986,N_18070,N_19410);
nor U24987 (N_24987,N_14593,N_12155);
or U24988 (N_24988,N_17455,N_16215);
nand U24989 (N_24989,N_13983,N_17962);
and U24990 (N_24990,N_16665,N_10624);
and U24991 (N_24991,N_19327,N_11210);
or U24992 (N_24992,N_18380,N_19083);
or U24993 (N_24993,N_12260,N_11723);
nor U24994 (N_24994,N_13781,N_17445);
and U24995 (N_24995,N_17242,N_13111);
and U24996 (N_24996,N_16334,N_10120);
xor U24997 (N_24997,N_10806,N_18510);
and U24998 (N_24998,N_16836,N_16369);
or U24999 (N_24999,N_12281,N_15947);
and U25000 (N_25000,N_11720,N_14231);
and U25001 (N_25001,N_13229,N_17683);
nand U25002 (N_25002,N_14050,N_13059);
nor U25003 (N_25003,N_19613,N_16525);
nand U25004 (N_25004,N_11829,N_10984);
or U25005 (N_25005,N_17338,N_10526);
nor U25006 (N_25006,N_15087,N_12436);
nor U25007 (N_25007,N_19432,N_11102);
xor U25008 (N_25008,N_11918,N_11040);
nor U25009 (N_25009,N_12927,N_17190);
nand U25010 (N_25010,N_12688,N_10131);
and U25011 (N_25011,N_18609,N_16898);
nand U25012 (N_25012,N_19595,N_16579);
nand U25013 (N_25013,N_18209,N_17541);
or U25014 (N_25014,N_13413,N_10725);
or U25015 (N_25015,N_19830,N_11194);
and U25016 (N_25016,N_10272,N_10921);
xor U25017 (N_25017,N_15023,N_17814);
or U25018 (N_25018,N_18832,N_16473);
nand U25019 (N_25019,N_19443,N_13439);
nor U25020 (N_25020,N_12274,N_18234);
or U25021 (N_25021,N_19481,N_13393);
nor U25022 (N_25022,N_10894,N_16193);
nand U25023 (N_25023,N_16273,N_16801);
and U25024 (N_25024,N_10852,N_11958);
nor U25025 (N_25025,N_17057,N_10668);
or U25026 (N_25026,N_11854,N_12526);
nor U25027 (N_25027,N_10756,N_19018);
nand U25028 (N_25028,N_15906,N_19866);
xor U25029 (N_25029,N_11543,N_13499);
xnor U25030 (N_25030,N_19056,N_10799);
and U25031 (N_25031,N_10123,N_14601);
and U25032 (N_25032,N_12923,N_19925);
nor U25033 (N_25033,N_18433,N_18974);
nor U25034 (N_25034,N_10402,N_19374);
nor U25035 (N_25035,N_10355,N_19865);
nand U25036 (N_25036,N_13294,N_18782);
and U25037 (N_25037,N_12696,N_17020);
nor U25038 (N_25038,N_14094,N_15735);
or U25039 (N_25039,N_19683,N_12712);
or U25040 (N_25040,N_19928,N_15785);
or U25041 (N_25041,N_16057,N_18312);
xor U25042 (N_25042,N_14166,N_10432);
and U25043 (N_25043,N_19067,N_10020);
xor U25044 (N_25044,N_10820,N_10053);
nand U25045 (N_25045,N_15793,N_13174);
and U25046 (N_25046,N_16194,N_18170);
or U25047 (N_25047,N_11687,N_16150);
nor U25048 (N_25048,N_14432,N_12834);
xor U25049 (N_25049,N_11948,N_10725);
nor U25050 (N_25050,N_19512,N_11135);
nor U25051 (N_25051,N_18087,N_18124);
nand U25052 (N_25052,N_15197,N_15998);
or U25053 (N_25053,N_13644,N_19926);
and U25054 (N_25054,N_15946,N_14978);
nand U25055 (N_25055,N_15205,N_10306);
and U25056 (N_25056,N_15064,N_17020);
or U25057 (N_25057,N_15771,N_14669);
xnor U25058 (N_25058,N_17786,N_14767);
nor U25059 (N_25059,N_16046,N_18296);
or U25060 (N_25060,N_15880,N_16161);
nand U25061 (N_25061,N_13262,N_18667);
or U25062 (N_25062,N_18970,N_12050);
xnor U25063 (N_25063,N_16597,N_12302);
and U25064 (N_25064,N_16581,N_18615);
and U25065 (N_25065,N_19392,N_11645);
or U25066 (N_25066,N_11752,N_10700);
nand U25067 (N_25067,N_18668,N_14292);
and U25068 (N_25068,N_13697,N_14690);
nand U25069 (N_25069,N_13138,N_12765);
and U25070 (N_25070,N_19374,N_11463);
nand U25071 (N_25071,N_12997,N_13641);
xor U25072 (N_25072,N_10165,N_17048);
and U25073 (N_25073,N_11721,N_15040);
or U25074 (N_25074,N_10182,N_18577);
nor U25075 (N_25075,N_10364,N_17692);
or U25076 (N_25076,N_12493,N_18560);
nand U25077 (N_25077,N_13916,N_15613);
nor U25078 (N_25078,N_13916,N_18119);
nor U25079 (N_25079,N_10872,N_19268);
xnor U25080 (N_25080,N_17638,N_13461);
xor U25081 (N_25081,N_16243,N_13670);
nand U25082 (N_25082,N_10833,N_15488);
xnor U25083 (N_25083,N_18622,N_19436);
nand U25084 (N_25084,N_12116,N_16029);
and U25085 (N_25085,N_12702,N_11503);
nor U25086 (N_25086,N_10400,N_10481);
nand U25087 (N_25087,N_14900,N_13906);
or U25088 (N_25088,N_15942,N_19379);
nand U25089 (N_25089,N_15197,N_12109);
and U25090 (N_25090,N_17613,N_15285);
nor U25091 (N_25091,N_10216,N_15060);
nor U25092 (N_25092,N_18721,N_18690);
nand U25093 (N_25093,N_14277,N_15074);
and U25094 (N_25094,N_15202,N_15971);
nand U25095 (N_25095,N_12993,N_15159);
nand U25096 (N_25096,N_11392,N_16017);
nor U25097 (N_25097,N_13544,N_17281);
xnor U25098 (N_25098,N_19314,N_17866);
or U25099 (N_25099,N_10646,N_15491);
and U25100 (N_25100,N_14188,N_14833);
nand U25101 (N_25101,N_18835,N_13772);
and U25102 (N_25102,N_11541,N_14052);
or U25103 (N_25103,N_13320,N_11506);
nand U25104 (N_25104,N_14925,N_13773);
nor U25105 (N_25105,N_14367,N_18439);
nand U25106 (N_25106,N_13065,N_12458);
nor U25107 (N_25107,N_15999,N_14895);
and U25108 (N_25108,N_19274,N_14463);
xnor U25109 (N_25109,N_11051,N_14545);
nor U25110 (N_25110,N_16919,N_17333);
nor U25111 (N_25111,N_19198,N_17996);
nand U25112 (N_25112,N_17413,N_14755);
or U25113 (N_25113,N_17829,N_11881);
and U25114 (N_25114,N_14789,N_17886);
nor U25115 (N_25115,N_19737,N_15670);
nor U25116 (N_25116,N_16947,N_19803);
or U25117 (N_25117,N_13877,N_13810);
or U25118 (N_25118,N_14216,N_14247);
xnor U25119 (N_25119,N_15179,N_11360);
nor U25120 (N_25120,N_13881,N_14936);
and U25121 (N_25121,N_16898,N_16311);
and U25122 (N_25122,N_15374,N_13845);
or U25123 (N_25123,N_15052,N_18974);
nor U25124 (N_25124,N_11390,N_17249);
and U25125 (N_25125,N_14399,N_10257);
nand U25126 (N_25126,N_13244,N_17687);
nand U25127 (N_25127,N_11334,N_11780);
nor U25128 (N_25128,N_17849,N_14013);
or U25129 (N_25129,N_15200,N_11959);
nor U25130 (N_25130,N_11127,N_19755);
nand U25131 (N_25131,N_11504,N_12300);
nand U25132 (N_25132,N_16011,N_16632);
or U25133 (N_25133,N_11674,N_13343);
nor U25134 (N_25134,N_14581,N_15663);
and U25135 (N_25135,N_15572,N_15063);
nand U25136 (N_25136,N_17658,N_16862);
or U25137 (N_25137,N_12478,N_18747);
and U25138 (N_25138,N_19455,N_18406);
nor U25139 (N_25139,N_17218,N_10342);
or U25140 (N_25140,N_15087,N_18942);
and U25141 (N_25141,N_13353,N_17920);
and U25142 (N_25142,N_13371,N_18561);
nand U25143 (N_25143,N_16683,N_13099);
and U25144 (N_25144,N_18657,N_13249);
or U25145 (N_25145,N_13697,N_15049);
or U25146 (N_25146,N_18080,N_13292);
nor U25147 (N_25147,N_13205,N_18175);
nor U25148 (N_25148,N_19799,N_17674);
nand U25149 (N_25149,N_16682,N_19039);
or U25150 (N_25150,N_18492,N_16666);
nand U25151 (N_25151,N_19247,N_13246);
or U25152 (N_25152,N_17162,N_12326);
and U25153 (N_25153,N_14335,N_16016);
nor U25154 (N_25154,N_14750,N_19918);
and U25155 (N_25155,N_17876,N_18619);
nor U25156 (N_25156,N_19223,N_13157);
nand U25157 (N_25157,N_10153,N_10495);
nand U25158 (N_25158,N_17361,N_16014);
and U25159 (N_25159,N_11344,N_19697);
or U25160 (N_25160,N_15772,N_14246);
nand U25161 (N_25161,N_19734,N_11101);
or U25162 (N_25162,N_13399,N_18770);
or U25163 (N_25163,N_16803,N_17263);
nand U25164 (N_25164,N_10356,N_10134);
nand U25165 (N_25165,N_14899,N_18224);
nor U25166 (N_25166,N_16155,N_18268);
nand U25167 (N_25167,N_12648,N_16225);
or U25168 (N_25168,N_12176,N_15348);
or U25169 (N_25169,N_17614,N_19199);
or U25170 (N_25170,N_16195,N_16284);
or U25171 (N_25171,N_18575,N_11261);
xor U25172 (N_25172,N_15786,N_15620);
and U25173 (N_25173,N_15011,N_18652);
and U25174 (N_25174,N_12337,N_15331);
and U25175 (N_25175,N_13395,N_10608);
nor U25176 (N_25176,N_18008,N_19345);
or U25177 (N_25177,N_19764,N_17203);
or U25178 (N_25178,N_11935,N_17024);
nor U25179 (N_25179,N_10345,N_18801);
or U25180 (N_25180,N_19565,N_19038);
nand U25181 (N_25181,N_13466,N_18040);
and U25182 (N_25182,N_13949,N_16814);
xor U25183 (N_25183,N_14557,N_16373);
or U25184 (N_25184,N_10030,N_13561);
xnor U25185 (N_25185,N_14432,N_17421);
and U25186 (N_25186,N_12797,N_15290);
nor U25187 (N_25187,N_16989,N_11664);
nor U25188 (N_25188,N_14812,N_16408);
and U25189 (N_25189,N_15008,N_17648);
or U25190 (N_25190,N_19747,N_19656);
xor U25191 (N_25191,N_14506,N_13278);
nor U25192 (N_25192,N_15050,N_12485);
nor U25193 (N_25193,N_17680,N_16863);
and U25194 (N_25194,N_15592,N_18786);
nand U25195 (N_25195,N_14757,N_13895);
nor U25196 (N_25196,N_17953,N_14241);
nor U25197 (N_25197,N_15568,N_12210);
xor U25198 (N_25198,N_17090,N_10805);
nor U25199 (N_25199,N_10887,N_13626);
and U25200 (N_25200,N_10301,N_14751);
and U25201 (N_25201,N_11524,N_12978);
or U25202 (N_25202,N_12519,N_17487);
or U25203 (N_25203,N_17624,N_10099);
xor U25204 (N_25204,N_10159,N_11452);
nand U25205 (N_25205,N_19291,N_14310);
and U25206 (N_25206,N_10174,N_18867);
xor U25207 (N_25207,N_14331,N_18896);
nand U25208 (N_25208,N_16522,N_13337);
and U25209 (N_25209,N_16332,N_17496);
nor U25210 (N_25210,N_13899,N_19145);
nor U25211 (N_25211,N_18089,N_17673);
xnor U25212 (N_25212,N_18280,N_18763);
and U25213 (N_25213,N_14271,N_17525);
xor U25214 (N_25214,N_12068,N_17206);
nand U25215 (N_25215,N_11552,N_13886);
nor U25216 (N_25216,N_16465,N_16715);
and U25217 (N_25217,N_10351,N_18633);
and U25218 (N_25218,N_13028,N_18973);
nand U25219 (N_25219,N_18350,N_11497);
xor U25220 (N_25220,N_17640,N_15952);
and U25221 (N_25221,N_15562,N_13198);
nor U25222 (N_25222,N_15366,N_12879);
nor U25223 (N_25223,N_16325,N_18856);
nor U25224 (N_25224,N_19245,N_19021);
and U25225 (N_25225,N_19904,N_17703);
xnor U25226 (N_25226,N_17271,N_15184);
nand U25227 (N_25227,N_11474,N_19521);
or U25228 (N_25228,N_14709,N_13432);
and U25229 (N_25229,N_16670,N_16401);
or U25230 (N_25230,N_10069,N_15757);
nand U25231 (N_25231,N_10434,N_16185);
xor U25232 (N_25232,N_10424,N_10792);
nor U25233 (N_25233,N_14105,N_12535);
and U25234 (N_25234,N_18401,N_19540);
nor U25235 (N_25235,N_12187,N_10031);
or U25236 (N_25236,N_18531,N_13203);
or U25237 (N_25237,N_19484,N_12027);
and U25238 (N_25238,N_10503,N_10261);
and U25239 (N_25239,N_11358,N_16015);
nand U25240 (N_25240,N_10637,N_11021);
nand U25241 (N_25241,N_10880,N_10744);
nor U25242 (N_25242,N_14013,N_10682);
or U25243 (N_25243,N_18234,N_12760);
nand U25244 (N_25244,N_15652,N_11512);
nand U25245 (N_25245,N_19027,N_15920);
nand U25246 (N_25246,N_13838,N_14644);
or U25247 (N_25247,N_18488,N_17306);
and U25248 (N_25248,N_19502,N_18675);
or U25249 (N_25249,N_11565,N_14971);
xor U25250 (N_25250,N_15052,N_16867);
or U25251 (N_25251,N_13604,N_17079);
or U25252 (N_25252,N_18892,N_17921);
xor U25253 (N_25253,N_13006,N_19356);
and U25254 (N_25254,N_11708,N_17208);
nor U25255 (N_25255,N_17989,N_11465);
and U25256 (N_25256,N_15024,N_13716);
or U25257 (N_25257,N_17418,N_17237);
or U25258 (N_25258,N_11396,N_11182);
nor U25259 (N_25259,N_12518,N_15591);
nand U25260 (N_25260,N_19926,N_11234);
nor U25261 (N_25261,N_15491,N_10000);
and U25262 (N_25262,N_17661,N_11433);
and U25263 (N_25263,N_10601,N_13763);
and U25264 (N_25264,N_13026,N_11020);
or U25265 (N_25265,N_13174,N_12080);
or U25266 (N_25266,N_18882,N_15063);
and U25267 (N_25267,N_13160,N_13362);
nor U25268 (N_25268,N_15012,N_10121);
and U25269 (N_25269,N_18671,N_10272);
and U25270 (N_25270,N_11561,N_19449);
and U25271 (N_25271,N_15986,N_16620);
xnor U25272 (N_25272,N_13984,N_18760);
nor U25273 (N_25273,N_12966,N_10833);
and U25274 (N_25274,N_16978,N_17605);
nand U25275 (N_25275,N_17451,N_17961);
xor U25276 (N_25276,N_17879,N_13087);
or U25277 (N_25277,N_12456,N_15738);
nand U25278 (N_25278,N_12179,N_14983);
or U25279 (N_25279,N_11884,N_17233);
and U25280 (N_25280,N_15390,N_10180);
and U25281 (N_25281,N_13231,N_10388);
and U25282 (N_25282,N_19444,N_11583);
nand U25283 (N_25283,N_17769,N_14641);
or U25284 (N_25284,N_14197,N_14084);
xnor U25285 (N_25285,N_15889,N_18828);
nor U25286 (N_25286,N_11896,N_13585);
nor U25287 (N_25287,N_15712,N_11716);
or U25288 (N_25288,N_16025,N_19082);
nor U25289 (N_25289,N_13670,N_16887);
xor U25290 (N_25290,N_14863,N_18385);
and U25291 (N_25291,N_18743,N_14339);
xnor U25292 (N_25292,N_17240,N_11329);
or U25293 (N_25293,N_16629,N_17336);
nor U25294 (N_25294,N_16363,N_14357);
xor U25295 (N_25295,N_12297,N_15217);
nor U25296 (N_25296,N_18700,N_11961);
or U25297 (N_25297,N_11637,N_12024);
and U25298 (N_25298,N_13179,N_16133);
nor U25299 (N_25299,N_17378,N_16152);
and U25300 (N_25300,N_15935,N_17892);
nor U25301 (N_25301,N_17897,N_10181);
or U25302 (N_25302,N_17980,N_13092);
or U25303 (N_25303,N_18744,N_14549);
or U25304 (N_25304,N_11767,N_18075);
or U25305 (N_25305,N_14036,N_14343);
xnor U25306 (N_25306,N_16724,N_17519);
nor U25307 (N_25307,N_11355,N_10539);
or U25308 (N_25308,N_10953,N_14233);
nor U25309 (N_25309,N_19060,N_16854);
and U25310 (N_25310,N_13944,N_12701);
nand U25311 (N_25311,N_12995,N_16995);
or U25312 (N_25312,N_15310,N_10715);
nand U25313 (N_25313,N_10703,N_11460);
and U25314 (N_25314,N_18762,N_19771);
nand U25315 (N_25315,N_10362,N_14751);
xnor U25316 (N_25316,N_13188,N_10397);
xnor U25317 (N_25317,N_15700,N_17045);
nor U25318 (N_25318,N_10964,N_17833);
or U25319 (N_25319,N_13568,N_18218);
nor U25320 (N_25320,N_19552,N_12768);
nand U25321 (N_25321,N_12049,N_15391);
nor U25322 (N_25322,N_18907,N_17487);
or U25323 (N_25323,N_12956,N_17570);
nor U25324 (N_25324,N_13712,N_19430);
and U25325 (N_25325,N_18085,N_19351);
or U25326 (N_25326,N_10582,N_12326);
nor U25327 (N_25327,N_16828,N_17426);
or U25328 (N_25328,N_18824,N_12564);
nand U25329 (N_25329,N_18006,N_15916);
or U25330 (N_25330,N_13879,N_14285);
nor U25331 (N_25331,N_17428,N_14586);
nor U25332 (N_25332,N_12482,N_18924);
or U25333 (N_25333,N_10628,N_14031);
and U25334 (N_25334,N_19500,N_13405);
or U25335 (N_25335,N_17010,N_10494);
nand U25336 (N_25336,N_19647,N_16293);
xor U25337 (N_25337,N_13856,N_10427);
or U25338 (N_25338,N_12374,N_16947);
or U25339 (N_25339,N_16806,N_10363);
nand U25340 (N_25340,N_19797,N_12653);
nor U25341 (N_25341,N_13373,N_10881);
nor U25342 (N_25342,N_18282,N_13954);
or U25343 (N_25343,N_13932,N_11344);
nor U25344 (N_25344,N_14313,N_12740);
or U25345 (N_25345,N_11842,N_13283);
and U25346 (N_25346,N_11369,N_12700);
nor U25347 (N_25347,N_11980,N_10677);
and U25348 (N_25348,N_13986,N_18239);
nand U25349 (N_25349,N_13964,N_14246);
or U25350 (N_25350,N_17449,N_14573);
and U25351 (N_25351,N_17376,N_19706);
nand U25352 (N_25352,N_14991,N_11067);
xnor U25353 (N_25353,N_14903,N_14507);
xor U25354 (N_25354,N_15357,N_19418);
nand U25355 (N_25355,N_15964,N_11795);
and U25356 (N_25356,N_17306,N_12798);
and U25357 (N_25357,N_17366,N_16467);
or U25358 (N_25358,N_11561,N_19120);
or U25359 (N_25359,N_17808,N_13426);
or U25360 (N_25360,N_17436,N_14725);
nor U25361 (N_25361,N_16375,N_15686);
xor U25362 (N_25362,N_17744,N_17798);
nand U25363 (N_25363,N_16415,N_17181);
nand U25364 (N_25364,N_11714,N_18162);
xnor U25365 (N_25365,N_13413,N_10166);
nor U25366 (N_25366,N_11411,N_16688);
nor U25367 (N_25367,N_11578,N_15161);
nand U25368 (N_25368,N_15756,N_10702);
nor U25369 (N_25369,N_11027,N_16784);
or U25370 (N_25370,N_19410,N_13712);
and U25371 (N_25371,N_17998,N_10326);
nor U25372 (N_25372,N_14418,N_10620);
nand U25373 (N_25373,N_12463,N_12636);
or U25374 (N_25374,N_15500,N_15189);
nor U25375 (N_25375,N_15392,N_19042);
or U25376 (N_25376,N_16317,N_11088);
and U25377 (N_25377,N_13999,N_16870);
nor U25378 (N_25378,N_13828,N_15316);
nor U25379 (N_25379,N_12754,N_11528);
xor U25380 (N_25380,N_14308,N_16010);
and U25381 (N_25381,N_10149,N_12761);
nor U25382 (N_25382,N_16580,N_10335);
or U25383 (N_25383,N_16346,N_18633);
nor U25384 (N_25384,N_17635,N_10811);
xnor U25385 (N_25385,N_11117,N_12784);
nor U25386 (N_25386,N_16130,N_12321);
or U25387 (N_25387,N_14651,N_18711);
and U25388 (N_25388,N_17863,N_19909);
or U25389 (N_25389,N_19050,N_17304);
nor U25390 (N_25390,N_18091,N_11100);
nand U25391 (N_25391,N_14013,N_14896);
and U25392 (N_25392,N_16998,N_14255);
and U25393 (N_25393,N_18686,N_13454);
xnor U25394 (N_25394,N_15800,N_14253);
xor U25395 (N_25395,N_14156,N_18594);
nand U25396 (N_25396,N_12467,N_17677);
nand U25397 (N_25397,N_11199,N_19404);
xnor U25398 (N_25398,N_14306,N_16174);
nor U25399 (N_25399,N_12106,N_11379);
nor U25400 (N_25400,N_11229,N_11958);
and U25401 (N_25401,N_18620,N_15421);
nand U25402 (N_25402,N_14761,N_13114);
nor U25403 (N_25403,N_19352,N_14146);
or U25404 (N_25404,N_15617,N_10061);
nor U25405 (N_25405,N_10379,N_19763);
nor U25406 (N_25406,N_13268,N_17255);
nand U25407 (N_25407,N_11928,N_19165);
and U25408 (N_25408,N_18293,N_15457);
or U25409 (N_25409,N_10570,N_13420);
nor U25410 (N_25410,N_19836,N_11149);
nor U25411 (N_25411,N_18615,N_11922);
or U25412 (N_25412,N_17529,N_16447);
nand U25413 (N_25413,N_13420,N_16543);
and U25414 (N_25414,N_12036,N_11617);
nand U25415 (N_25415,N_16003,N_10321);
nor U25416 (N_25416,N_19338,N_12399);
nor U25417 (N_25417,N_12925,N_12869);
and U25418 (N_25418,N_19303,N_11700);
or U25419 (N_25419,N_12577,N_15846);
and U25420 (N_25420,N_12953,N_10602);
nor U25421 (N_25421,N_17314,N_19430);
xnor U25422 (N_25422,N_15402,N_16333);
nor U25423 (N_25423,N_11584,N_12381);
or U25424 (N_25424,N_13116,N_16056);
nand U25425 (N_25425,N_19827,N_17671);
nor U25426 (N_25426,N_15862,N_12533);
or U25427 (N_25427,N_10128,N_16906);
nand U25428 (N_25428,N_15442,N_15064);
or U25429 (N_25429,N_19489,N_14004);
xor U25430 (N_25430,N_10549,N_12783);
or U25431 (N_25431,N_10754,N_16185);
nand U25432 (N_25432,N_11009,N_13207);
nor U25433 (N_25433,N_14558,N_19487);
nor U25434 (N_25434,N_11944,N_18226);
nand U25435 (N_25435,N_13165,N_11656);
nand U25436 (N_25436,N_18945,N_19122);
nand U25437 (N_25437,N_11028,N_10328);
or U25438 (N_25438,N_17449,N_12266);
nand U25439 (N_25439,N_18704,N_13787);
or U25440 (N_25440,N_14784,N_16368);
nand U25441 (N_25441,N_12918,N_11343);
and U25442 (N_25442,N_19047,N_14274);
and U25443 (N_25443,N_16529,N_19896);
and U25444 (N_25444,N_13328,N_12913);
or U25445 (N_25445,N_18022,N_18709);
or U25446 (N_25446,N_18663,N_19450);
nor U25447 (N_25447,N_18003,N_17114);
and U25448 (N_25448,N_16379,N_11324);
or U25449 (N_25449,N_19384,N_16964);
nand U25450 (N_25450,N_12246,N_15340);
nor U25451 (N_25451,N_15651,N_12532);
nor U25452 (N_25452,N_17303,N_17578);
or U25453 (N_25453,N_13151,N_11422);
nor U25454 (N_25454,N_11136,N_14426);
nor U25455 (N_25455,N_19378,N_15403);
xnor U25456 (N_25456,N_13604,N_13179);
nand U25457 (N_25457,N_17174,N_13344);
xnor U25458 (N_25458,N_12135,N_18246);
nor U25459 (N_25459,N_13070,N_19090);
xor U25460 (N_25460,N_13660,N_12173);
xnor U25461 (N_25461,N_13931,N_19420);
and U25462 (N_25462,N_14725,N_10350);
nor U25463 (N_25463,N_18384,N_14653);
xor U25464 (N_25464,N_18065,N_15062);
and U25465 (N_25465,N_17750,N_16023);
and U25466 (N_25466,N_19150,N_11754);
or U25467 (N_25467,N_12284,N_15704);
or U25468 (N_25468,N_19589,N_18805);
nor U25469 (N_25469,N_10781,N_18094);
or U25470 (N_25470,N_12642,N_18068);
and U25471 (N_25471,N_14216,N_12373);
and U25472 (N_25472,N_12822,N_14840);
or U25473 (N_25473,N_10085,N_12774);
nand U25474 (N_25474,N_19402,N_17047);
xnor U25475 (N_25475,N_16820,N_16248);
nor U25476 (N_25476,N_17332,N_13179);
xor U25477 (N_25477,N_17087,N_15786);
nand U25478 (N_25478,N_12670,N_16256);
or U25479 (N_25479,N_11348,N_19860);
and U25480 (N_25480,N_19706,N_13158);
nand U25481 (N_25481,N_11110,N_10995);
xnor U25482 (N_25482,N_10433,N_18271);
nand U25483 (N_25483,N_10096,N_18867);
and U25484 (N_25484,N_16272,N_13392);
and U25485 (N_25485,N_12948,N_11348);
or U25486 (N_25486,N_10461,N_19703);
and U25487 (N_25487,N_19522,N_17994);
nor U25488 (N_25488,N_19750,N_17445);
nor U25489 (N_25489,N_14071,N_12135);
or U25490 (N_25490,N_14652,N_11858);
and U25491 (N_25491,N_10365,N_17519);
or U25492 (N_25492,N_14751,N_16264);
or U25493 (N_25493,N_13670,N_15327);
and U25494 (N_25494,N_16120,N_11693);
nand U25495 (N_25495,N_10490,N_10177);
nand U25496 (N_25496,N_18409,N_10609);
xor U25497 (N_25497,N_11619,N_17553);
or U25498 (N_25498,N_10630,N_13915);
or U25499 (N_25499,N_14786,N_10291);
or U25500 (N_25500,N_16715,N_17078);
nor U25501 (N_25501,N_11768,N_10336);
nor U25502 (N_25502,N_12700,N_14541);
or U25503 (N_25503,N_15119,N_18183);
nand U25504 (N_25504,N_14222,N_18472);
or U25505 (N_25505,N_15795,N_10748);
nor U25506 (N_25506,N_17330,N_15703);
nand U25507 (N_25507,N_17882,N_18430);
nand U25508 (N_25508,N_13626,N_12806);
nor U25509 (N_25509,N_16447,N_19710);
and U25510 (N_25510,N_11876,N_14502);
nand U25511 (N_25511,N_15913,N_18887);
or U25512 (N_25512,N_11830,N_15725);
or U25513 (N_25513,N_10631,N_19033);
nor U25514 (N_25514,N_19986,N_18249);
and U25515 (N_25515,N_14795,N_18462);
nor U25516 (N_25516,N_18530,N_16386);
or U25517 (N_25517,N_17386,N_14699);
nor U25518 (N_25518,N_13739,N_15739);
and U25519 (N_25519,N_11177,N_10932);
nand U25520 (N_25520,N_16606,N_12280);
and U25521 (N_25521,N_18136,N_15339);
nand U25522 (N_25522,N_17290,N_16775);
nand U25523 (N_25523,N_18663,N_11980);
nor U25524 (N_25524,N_12008,N_18209);
and U25525 (N_25525,N_17446,N_12970);
and U25526 (N_25526,N_17571,N_18742);
or U25527 (N_25527,N_15513,N_10396);
nor U25528 (N_25528,N_13596,N_11797);
nor U25529 (N_25529,N_16599,N_11576);
nand U25530 (N_25530,N_10796,N_15456);
nor U25531 (N_25531,N_19243,N_19170);
nand U25532 (N_25532,N_17413,N_17384);
nor U25533 (N_25533,N_11260,N_14358);
nor U25534 (N_25534,N_18032,N_10050);
or U25535 (N_25535,N_16192,N_10291);
or U25536 (N_25536,N_10051,N_12138);
nand U25537 (N_25537,N_12899,N_19984);
nand U25538 (N_25538,N_14568,N_14394);
and U25539 (N_25539,N_14704,N_19053);
or U25540 (N_25540,N_19936,N_14200);
nor U25541 (N_25541,N_14151,N_13587);
nor U25542 (N_25542,N_14315,N_12475);
xor U25543 (N_25543,N_17809,N_14910);
and U25544 (N_25544,N_10404,N_14092);
and U25545 (N_25545,N_17948,N_19634);
nor U25546 (N_25546,N_11387,N_12560);
or U25547 (N_25547,N_11213,N_11152);
nand U25548 (N_25548,N_15168,N_12113);
nand U25549 (N_25549,N_12638,N_10890);
nor U25550 (N_25550,N_14317,N_16985);
and U25551 (N_25551,N_19947,N_10088);
and U25552 (N_25552,N_15913,N_11416);
and U25553 (N_25553,N_10253,N_15544);
and U25554 (N_25554,N_14084,N_18000);
nor U25555 (N_25555,N_11378,N_18904);
xnor U25556 (N_25556,N_18276,N_16821);
and U25557 (N_25557,N_10675,N_15521);
or U25558 (N_25558,N_11699,N_19237);
nand U25559 (N_25559,N_14170,N_12676);
nor U25560 (N_25560,N_10779,N_11791);
or U25561 (N_25561,N_11195,N_12291);
nand U25562 (N_25562,N_12064,N_10111);
or U25563 (N_25563,N_14102,N_16223);
or U25564 (N_25564,N_12499,N_12178);
nor U25565 (N_25565,N_10433,N_14792);
and U25566 (N_25566,N_18964,N_17000);
xor U25567 (N_25567,N_15693,N_11185);
and U25568 (N_25568,N_12754,N_10699);
nor U25569 (N_25569,N_10907,N_14443);
nor U25570 (N_25570,N_15497,N_19798);
and U25571 (N_25571,N_11696,N_10746);
nor U25572 (N_25572,N_15755,N_10486);
nor U25573 (N_25573,N_16723,N_15452);
or U25574 (N_25574,N_17432,N_11087);
nand U25575 (N_25575,N_15932,N_14959);
and U25576 (N_25576,N_11465,N_18006);
or U25577 (N_25577,N_17874,N_14850);
or U25578 (N_25578,N_13721,N_18616);
nor U25579 (N_25579,N_17027,N_13605);
nand U25580 (N_25580,N_14233,N_12820);
or U25581 (N_25581,N_13384,N_16565);
and U25582 (N_25582,N_10866,N_17478);
nor U25583 (N_25583,N_17388,N_18881);
or U25584 (N_25584,N_14813,N_18681);
nand U25585 (N_25585,N_14371,N_19846);
and U25586 (N_25586,N_12787,N_18603);
nor U25587 (N_25587,N_17144,N_10805);
nor U25588 (N_25588,N_15610,N_13009);
nor U25589 (N_25589,N_15777,N_13707);
or U25590 (N_25590,N_10829,N_14081);
nor U25591 (N_25591,N_18833,N_13983);
or U25592 (N_25592,N_18513,N_14376);
or U25593 (N_25593,N_14408,N_12823);
nand U25594 (N_25594,N_17666,N_15514);
and U25595 (N_25595,N_10232,N_12170);
nand U25596 (N_25596,N_12715,N_10682);
and U25597 (N_25597,N_18860,N_12013);
xnor U25598 (N_25598,N_16311,N_14935);
or U25599 (N_25599,N_18308,N_14220);
or U25600 (N_25600,N_13088,N_18141);
nor U25601 (N_25601,N_17469,N_16852);
nand U25602 (N_25602,N_13424,N_12323);
nor U25603 (N_25603,N_10572,N_14517);
nor U25604 (N_25604,N_14549,N_12556);
nand U25605 (N_25605,N_14725,N_14759);
nand U25606 (N_25606,N_13402,N_15324);
nand U25607 (N_25607,N_10075,N_11268);
and U25608 (N_25608,N_14592,N_16721);
nor U25609 (N_25609,N_17590,N_15185);
xnor U25610 (N_25610,N_10255,N_16808);
nor U25611 (N_25611,N_15578,N_19984);
or U25612 (N_25612,N_10886,N_15852);
or U25613 (N_25613,N_16007,N_16591);
nor U25614 (N_25614,N_15080,N_16893);
and U25615 (N_25615,N_11423,N_14597);
and U25616 (N_25616,N_16874,N_16190);
nand U25617 (N_25617,N_11136,N_11133);
and U25618 (N_25618,N_16129,N_12086);
xnor U25619 (N_25619,N_10501,N_16443);
nor U25620 (N_25620,N_18846,N_11063);
and U25621 (N_25621,N_18268,N_11706);
nor U25622 (N_25622,N_15439,N_18785);
nand U25623 (N_25623,N_10213,N_15123);
or U25624 (N_25624,N_12082,N_13434);
and U25625 (N_25625,N_17994,N_16563);
nor U25626 (N_25626,N_12730,N_13242);
nand U25627 (N_25627,N_12363,N_16661);
nor U25628 (N_25628,N_13356,N_15155);
and U25629 (N_25629,N_18119,N_15780);
nand U25630 (N_25630,N_15384,N_14580);
nor U25631 (N_25631,N_19010,N_14254);
nand U25632 (N_25632,N_12887,N_15910);
or U25633 (N_25633,N_18332,N_10567);
or U25634 (N_25634,N_11843,N_14522);
nor U25635 (N_25635,N_13750,N_16787);
xnor U25636 (N_25636,N_19485,N_11065);
and U25637 (N_25637,N_10112,N_16756);
xor U25638 (N_25638,N_13764,N_18055);
or U25639 (N_25639,N_13016,N_14875);
nor U25640 (N_25640,N_18412,N_13295);
xor U25641 (N_25641,N_13412,N_16371);
nor U25642 (N_25642,N_17293,N_14661);
nand U25643 (N_25643,N_15351,N_10479);
nand U25644 (N_25644,N_11939,N_16574);
nand U25645 (N_25645,N_18744,N_11750);
nand U25646 (N_25646,N_12646,N_15931);
and U25647 (N_25647,N_10334,N_17343);
and U25648 (N_25648,N_10892,N_18427);
and U25649 (N_25649,N_18133,N_12981);
xnor U25650 (N_25650,N_19270,N_17989);
xor U25651 (N_25651,N_14233,N_10816);
or U25652 (N_25652,N_18697,N_19460);
nand U25653 (N_25653,N_15919,N_19680);
or U25654 (N_25654,N_19778,N_11122);
or U25655 (N_25655,N_11750,N_14341);
nand U25656 (N_25656,N_13834,N_19238);
and U25657 (N_25657,N_14817,N_13008);
nand U25658 (N_25658,N_11069,N_15357);
and U25659 (N_25659,N_18798,N_13033);
and U25660 (N_25660,N_18423,N_19765);
nor U25661 (N_25661,N_13072,N_18485);
nand U25662 (N_25662,N_14605,N_19007);
nand U25663 (N_25663,N_12833,N_12859);
nor U25664 (N_25664,N_14791,N_19323);
nor U25665 (N_25665,N_13950,N_10702);
and U25666 (N_25666,N_13811,N_11352);
nand U25667 (N_25667,N_18704,N_10352);
and U25668 (N_25668,N_10787,N_13121);
nand U25669 (N_25669,N_19033,N_14587);
and U25670 (N_25670,N_15324,N_10035);
nand U25671 (N_25671,N_18341,N_14265);
or U25672 (N_25672,N_16240,N_19634);
and U25673 (N_25673,N_12414,N_16391);
nor U25674 (N_25674,N_14710,N_16217);
or U25675 (N_25675,N_16382,N_15946);
nand U25676 (N_25676,N_14718,N_18847);
nand U25677 (N_25677,N_11431,N_13722);
or U25678 (N_25678,N_15042,N_11561);
nor U25679 (N_25679,N_19494,N_19621);
or U25680 (N_25680,N_14061,N_14245);
or U25681 (N_25681,N_18264,N_16657);
xnor U25682 (N_25682,N_10994,N_14112);
and U25683 (N_25683,N_10752,N_16411);
or U25684 (N_25684,N_12612,N_17483);
or U25685 (N_25685,N_13120,N_13899);
nor U25686 (N_25686,N_11003,N_18223);
and U25687 (N_25687,N_19346,N_14577);
nor U25688 (N_25688,N_15923,N_13650);
or U25689 (N_25689,N_19156,N_12231);
nor U25690 (N_25690,N_16368,N_10346);
and U25691 (N_25691,N_18818,N_15070);
nand U25692 (N_25692,N_14311,N_12574);
nand U25693 (N_25693,N_17404,N_17564);
nand U25694 (N_25694,N_15361,N_12431);
nand U25695 (N_25695,N_12973,N_16701);
and U25696 (N_25696,N_18751,N_15092);
or U25697 (N_25697,N_11725,N_15192);
and U25698 (N_25698,N_19269,N_12258);
or U25699 (N_25699,N_19115,N_13378);
nand U25700 (N_25700,N_11813,N_13653);
nand U25701 (N_25701,N_16838,N_18789);
and U25702 (N_25702,N_18866,N_10551);
nor U25703 (N_25703,N_11540,N_14605);
or U25704 (N_25704,N_12218,N_11200);
nand U25705 (N_25705,N_13586,N_17501);
or U25706 (N_25706,N_12517,N_18684);
nor U25707 (N_25707,N_14995,N_12277);
nand U25708 (N_25708,N_14408,N_13483);
nor U25709 (N_25709,N_19659,N_11916);
or U25710 (N_25710,N_12758,N_12885);
nand U25711 (N_25711,N_14902,N_11493);
and U25712 (N_25712,N_11602,N_11306);
nor U25713 (N_25713,N_15381,N_15429);
or U25714 (N_25714,N_15975,N_15954);
nand U25715 (N_25715,N_19654,N_11426);
nand U25716 (N_25716,N_14391,N_10232);
and U25717 (N_25717,N_13560,N_11787);
nand U25718 (N_25718,N_11417,N_10155);
nor U25719 (N_25719,N_11042,N_11296);
xnor U25720 (N_25720,N_11400,N_12357);
xor U25721 (N_25721,N_10987,N_19555);
nand U25722 (N_25722,N_11661,N_17084);
nor U25723 (N_25723,N_13086,N_13513);
nand U25724 (N_25724,N_18499,N_14977);
or U25725 (N_25725,N_16675,N_18441);
nand U25726 (N_25726,N_19429,N_12694);
xnor U25727 (N_25727,N_10973,N_11269);
and U25728 (N_25728,N_18990,N_12340);
and U25729 (N_25729,N_16660,N_18178);
and U25730 (N_25730,N_17832,N_17860);
nand U25731 (N_25731,N_10871,N_17255);
nand U25732 (N_25732,N_11053,N_15751);
or U25733 (N_25733,N_19965,N_17601);
nor U25734 (N_25734,N_13462,N_18476);
nand U25735 (N_25735,N_10423,N_11582);
or U25736 (N_25736,N_12908,N_15913);
xor U25737 (N_25737,N_10903,N_17564);
and U25738 (N_25738,N_14828,N_15188);
nand U25739 (N_25739,N_10777,N_11692);
and U25740 (N_25740,N_18450,N_16984);
nand U25741 (N_25741,N_16382,N_16866);
or U25742 (N_25742,N_15823,N_11824);
or U25743 (N_25743,N_16286,N_18579);
and U25744 (N_25744,N_14984,N_19441);
or U25745 (N_25745,N_15127,N_10051);
and U25746 (N_25746,N_11411,N_17837);
nor U25747 (N_25747,N_10512,N_18433);
and U25748 (N_25748,N_13876,N_10772);
xnor U25749 (N_25749,N_12370,N_12381);
and U25750 (N_25750,N_13144,N_15215);
nor U25751 (N_25751,N_10577,N_17944);
and U25752 (N_25752,N_12713,N_19664);
or U25753 (N_25753,N_18972,N_18538);
or U25754 (N_25754,N_19286,N_16135);
or U25755 (N_25755,N_15574,N_15127);
or U25756 (N_25756,N_12582,N_15992);
nor U25757 (N_25757,N_13692,N_12963);
nor U25758 (N_25758,N_19395,N_12598);
or U25759 (N_25759,N_13623,N_17191);
and U25760 (N_25760,N_16019,N_13962);
nand U25761 (N_25761,N_11986,N_14497);
xor U25762 (N_25762,N_13146,N_18826);
xor U25763 (N_25763,N_19734,N_14608);
or U25764 (N_25764,N_12528,N_15520);
nor U25765 (N_25765,N_18391,N_16050);
and U25766 (N_25766,N_15234,N_10479);
and U25767 (N_25767,N_10943,N_14872);
nor U25768 (N_25768,N_19701,N_12825);
and U25769 (N_25769,N_19267,N_11032);
nor U25770 (N_25770,N_11991,N_10822);
nand U25771 (N_25771,N_19621,N_13305);
or U25772 (N_25772,N_16950,N_12526);
and U25773 (N_25773,N_16504,N_17237);
and U25774 (N_25774,N_10017,N_14544);
nand U25775 (N_25775,N_15988,N_15285);
nor U25776 (N_25776,N_12282,N_11246);
and U25777 (N_25777,N_12730,N_17138);
or U25778 (N_25778,N_10927,N_13781);
xor U25779 (N_25779,N_14406,N_17087);
nor U25780 (N_25780,N_11931,N_15191);
nor U25781 (N_25781,N_16211,N_18951);
or U25782 (N_25782,N_16322,N_13585);
nand U25783 (N_25783,N_16881,N_17568);
nor U25784 (N_25784,N_17964,N_15845);
and U25785 (N_25785,N_10817,N_16820);
and U25786 (N_25786,N_18788,N_10411);
nand U25787 (N_25787,N_17399,N_18397);
or U25788 (N_25788,N_15638,N_18549);
nand U25789 (N_25789,N_16325,N_18275);
nor U25790 (N_25790,N_18708,N_13042);
nor U25791 (N_25791,N_16184,N_10934);
or U25792 (N_25792,N_16612,N_12223);
xnor U25793 (N_25793,N_17767,N_12664);
or U25794 (N_25794,N_10024,N_16857);
and U25795 (N_25795,N_19478,N_13801);
nor U25796 (N_25796,N_12556,N_14711);
nor U25797 (N_25797,N_12779,N_13552);
nor U25798 (N_25798,N_19485,N_12766);
nor U25799 (N_25799,N_10307,N_16699);
nor U25800 (N_25800,N_10957,N_13760);
nand U25801 (N_25801,N_18860,N_12049);
or U25802 (N_25802,N_13717,N_18827);
nand U25803 (N_25803,N_19411,N_10183);
or U25804 (N_25804,N_11274,N_19020);
nor U25805 (N_25805,N_12135,N_14385);
nor U25806 (N_25806,N_14219,N_10882);
nand U25807 (N_25807,N_11018,N_15108);
nor U25808 (N_25808,N_15911,N_13082);
nor U25809 (N_25809,N_15562,N_16348);
xor U25810 (N_25810,N_19920,N_15806);
nand U25811 (N_25811,N_18647,N_11059);
xor U25812 (N_25812,N_13880,N_15111);
nand U25813 (N_25813,N_17954,N_19991);
or U25814 (N_25814,N_12632,N_13149);
nand U25815 (N_25815,N_15683,N_14310);
or U25816 (N_25816,N_17384,N_11261);
xnor U25817 (N_25817,N_17922,N_16073);
and U25818 (N_25818,N_13001,N_14131);
nand U25819 (N_25819,N_14315,N_13373);
nor U25820 (N_25820,N_13188,N_12691);
nand U25821 (N_25821,N_15655,N_12057);
and U25822 (N_25822,N_16786,N_13090);
and U25823 (N_25823,N_13544,N_10753);
and U25824 (N_25824,N_12322,N_18502);
nand U25825 (N_25825,N_18704,N_12105);
and U25826 (N_25826,N_16743,N_14572);
xor U25827 (N_25827,N_17925,N_16543);
and U25828 (N_25828,N_13045,N_15549);
and U25829 (N_25829,N_10842,N_19300);
nor U25830 (N_25830,N_16847,N_17394);
xnor U25831 (N_25831,N_13303,N_14658);
or U25832 (N_25832,N_12386,N_16303);
or U25833 (N_25833,N_13763,N_10718);
or U25834 (N_25834,N_11789,N_11308);
xnor U25835 (N_25835,N_18348,N_12702);
nor U25836 (N_25836,N_12939,N_13461);
and U25837 (N_25837,N_17524,N_11275);
and U25838 (N_25838,N_19225,N_13152);
nor U25839 (N_25839,N_19744,N_13261);
nor U25840 (N_25840,N_13691,N_18743);
and U25841 (N_25841,N_10121,N_15940);
xnor U25842 (N_25842,N_10620,N_17224);
or U25843 (N_25843,N_11844,N_15074);
and U25844 (N_25844,N_14084,N_17710);
nor U25845 (N_25845,N_11270,N_13699);
nor U25846 (N_25846,N_10730,N_19629);
nand U25847 (N_25847,N_13472,N_12547);
and U25848 (N_25848,N_12258,N_18203);
nand U25849 (N_25849,N_13659,N_18541);
and U25850 (N_25850,N_15357,N_17063);
nand U25851 (N_25851,N_17471,N_10731);
and U25852 (N_25852,N_14260,N_12519);
nand U25853 (N_25853,N_15720,N_12266);
xnor U25854 (N_25854,N_16277,N_13913);
and U25855 (N_25855,N_19004,N_12580);
xnor U25856 (N_25856,N_12994,N_11208);
nand U25857 (N_25857,N_18498,N_15533);
and U25858 (N_25858,N_11593,N_16548);
or U25859 (N_25859,N_16170,N_19876);
nand U25860 (N_25860,N_13242,N_14409);
nor U25861 (N_25861,N_16854,N_11635);
or U25862 (N_25862,N_19733,N_19019);
and U25863 (N_25863,N_16495,N_18209);
or U25864 (N_25864,N_19500,N_15577);
nand U25865 (N_25865,N_12661,N_18602);
nand U25866 (N_25866,N_11315,N_17439);
xor U25867 (N_25867,N_19017,N_11777);
xnor U25868 (N_25868,N_17349,N_15541);
nand U25869 (N_25869,N_16214,N_13345);
or U25870 (N_25870,N_16285,N_19368);
nand U25871 (N_25871,N_16097,N_18626);
or U25872 (N_25872,N_13482,N_12468);
nor U25873 (N_25873,N_19627,N_11856);
nand U25874 (N_25874,N_17733,N_19058);
nor U25875 (N_25875,N_16949,N_16862);
or U25876 (N_25876,N_16921,N_18434);
nand U25877 (N_25877,N_17372,N_11049);
nor U25878 (N_25878,N_10061,N_16602);
xor U25879 (N_25879,N_14284,N_11387);
nor U25880 (N_25880,N_10567,N_16258);
xor U25881 (N_25881,N_14703,N_11362);
nor U25882 (N_25882,N_17069,N_11594);
nor U25883 (N_25883,N_10036,N_16177);
nor U25884 (N_25884,N_14492,N_19771);
xor U25885 (N_25885,N_15003,N_14318);
xnor U25886 (N_25886,N_14713,N_10778);
nor U25887 (N_25887,N_15172,N_15131);
xor U25888 (N_25888,N_10272,N_13377);
nor U25889 (N_25889,N_13693,N_16095);
nand U25890 (N_25890,N_13633,N_10652);
or U25891 (N_25891,N_16544,N_14929);
nor U25892 (N_25892,N_19335,N_18944);
nor U25893 (N_25893,N_14825,N_17116);
or U25894 (N_25894,N_18386,N_12210);
and U25895 (N_25895,N_12281,N_11486);
nand U25896 (N_25896,N_15310,N_13782);
nor U25897 (N_25897,N_16428,N_12340);
or U25898 (N_25898,N_14606,N_18687);
nor U25899 (N_25899,N_18794,N_11933);
and U25900 (N_25900,N_12290,N_11807);
xor U25901 (N_25901,N_19371,N_10582);
nand U25902 (N_25902,N_16806,N_12561);
nand U25903 (N_25903,N_16398,N_12544);
and U25904 (N_25904,N_18641,N_19613);
and U25905 (N_25905,N_19621,N_17148);
xnor U25906 (N_25906,N_13536,N_10663);
nor U25907 (N_25907,N_11658,N_18037);
xor U25908 (N_25908,N_19362,N_19772);
or U25909 (N_25909,N_15654,N_12430);
and U25910 (N_25910,N_14904,N_14934);
or U25911 (N_25911,N_13066,N_13736);
and U25912 (N_25912,N_14089,N_10074);
or U25913 (N_25913,N_10365,N_10883);
and U25914 (N_25914,N_19687,N_17717);
nor U25915 (N_25915,N_19595,N_13380);
nor U25916 (N_25916,N_18077,N_10918);
nor U25917 (N_25917,N_13195,N_18068);
nand U25918 (N_25918,N_18703,N_15211);
or U25919 (N_25919,N_17188,N_11407);
or U25920 (N_25920,N_12201,N_19390);
nand U25921 (N_25921,N_19183,N_15358);
nor U25922 (N_25922,N_13715,N_15494);
nand U25923 (N_25923,N_10500,N_12096);
nand U25924 (N_25924,N_18509,N_10802);
or U25925 (N_25925,N_12010,N_18462);
nand U25926 (N_25926,N_16422,N_12430);
and U25927 (N_25927,N_12515,N_16657);
nand U25928 (N_25928,N_13759,N_18317);
and U25929 (N_25929,N_17560,N_11972);
or U25930 (N_25930,N_11777,N_14729);
or U25931 (N_25931,N_13304,N_11562);
nor U25932 (N_25932,N_11061,N_18242);
and U25933 (N_25933,N_12169,N_13022);
or U25934 (N_25934,N_18682,N_14911);
nor U25935 (N_25935,N_19329,N_12946);
nand U25936 (N_25936,N_13766,N_16751);
and U25937 (N_25937,N_17910,N_19311);
and U25938 (N_25938,N_17087,N_18042);
or U25939 (N_25939,N_11851,N_17951);
nand U25940 (N_25940,N_11679,N_18225);
and U25941 (N_25941,N_11639,N_12549);
or U25942 (N_25942,N_19168,N_17695);
and U25943 (N_25943,N_14577,N_10663);
and U25944 (N_25944,N_19860,N_13477);
nand U25945 (N_25945,N_13835,N_19259);
or U25946 (N_25946,N_18994,N_17091);
nor U25947 (N_25947,N_10686,N_10767);
nor U25948 (N_25948,N_14371,N_19771);
and U25949 (N_25949,N_18377,N_12502);
xor U25950 (N_25950,N_12429,N_17760);
and U25951 (N_25951,N_19475,N_10667);
nand U25952 (N_25952,N_19714,N_13597);
nor U25953 (N_25953,N_14200,N_15824);
and U25954 (N_25954,N_11211,N_18134);
xor U25955 (N_25955,N_19038,N_16189);
xor U25956 (N_25956,N_13117,N_10128);
and U25957 (N_25957,N_10601,N_19382);
xnor U25958 (N_25958,N_11343,N_10275);
nand U25959 (N_25959,N_13905,N_12311);
nand U25960 (N_25960,N_17961,N_16303);
and U25961 (N_25961,N_15256,N_13439);
or U25962 (N_25962,N_10064,N_15227);
xnor U25963 (N_25963,N_16291,N_13086);
or U25964 (N_25964,N_12890,N_16764);
xnor U25965 (N_25965,N_12764,N_10514);
nand U25966 (N_25966,N_17127,N_12605);
or U25967 (N_25967,N_10575,N_14386);
or U25968 (N_25968,N_11415,N_14967);
and U25969 (N_25969,N_19177,N_12442);
nor U25970 (N_25970,N_13836,N_10923);
or U25971 (N_25971,N_11273,N_14321);
and U25972 (N_25972,N_19858,N_16195);
or U25973 (N_25973,N_17943,N_16621);
nand U25974 (N_25974,N_15232,N_13844);
nor U25975 (N_25975,N_10545,N_12663);
or U25976 (N_25976,N_19069,N_10356);
or U25977 (N_25977,N_19275,N_12022);
nor U25978 (N_25978,N_17506,N_12327);
nor U25979 (N_25979,N_14266,N_11716);
nand U25980 (N_25980,N_15451,N_16406);
nor U25981 (N_25981,N_15449,N_19938);
or U25982 (N_25982,N_15197,N_16727);
nand U25983 (N_25983,N_13462,N_13699);
or U25984 (N_25984,N_18623,N_17887);
and U25985 (N_25985,N_12624,N_15802);
nor U25986 (N_25986,N_19539,N_19433);
and U25987 (N_25987,N_19092,N_15645);
nor U25988 (N_25988,N_18908,N_19026);
and U25989 (N_25989,N_16252,N_16352);
nor U25990 (N_25990,N_18788,N_10232);
or U25991 (N_25991,N_19127,N_14285);
nand U25992 (N_25992,N_17274,N_11346);
nand U25993 (N_25993,N_12170,N_11016);
and U25994 (N_25994,N_11978,N_16845);
nand U25995 (N_25995,N_10722,N_10334);
nor U25996 (N_25996,N_10562,N_17212);
or U25997 (N_25997,N_12902,N_19212);
or U25998 (N_25998,N_16990,N_12361);
nand U25999 (N_25999,N_18175,N_17707);
or U26000 (N_26000,N_18456,N_18149);
nand U26001 (N_26001,N_14928,N_18199);
nand U26002 (N_26002,N_11700,N_13455);
nor U26003 (N_26003,N_14466,N_19468);
nor U26004 (N_26004,N_14145,N_18644);
nand U26005 (N_26005,N_18234,N_15172);
nand U26006 (N_26006,N_19768,N_16532);
or U26007 (N_26007,N_10480,N_11107);
and U26008 (N_26008,N_17845,N_13179);
and U26009 (N_26009,N_17647,N_19522);
and U26010 (N_26010,N_17646,N_19246);
nor U26011 (N_26011,N_10547,N_17980);
nand U26012 (N_26012,N_19258,N_13225);
nor U26013 (N_26013,N_17511,N_16157);
xnor U26014 (N_26014,N_18230,N_11350);
nand U26015 (N_26015,N_19521,N_19338);
nor U26016 (N_26016,N_16414,N_13583);
or U26017 (N_26017,N_15026,N_15665);
and U26018 (N_26018,N_13274,N_15386);
nand U26019 (N_26019,N_10124,N_10885);
nor U26020 (N_26020,N_15144,N_19068);
or U26021 (N_26021,N_10098,N_11622);
nand U26022 (N_26022,N_14399,N_18629);
and U26023 (N_26023,N_17299,N_16868);
nand U26024 (N_26024,N_19957,N_14904);
nand U26025 (N_26025,N_10179,N_18790);
nor U26026 (N_26026,N_14245,N_17737);
nor U26027 (N_26027,N_12163,N_11403);
or U26028 (N_26028,N_12557,N_18698);
or U26029 (N_26029,N_15151,N_18887);
xnor U26030 (N_26030,N_16189,N_14760);
or U26031 (N_26031,N_16596,N_15997);
xor U26032 (N_26032,N_15922,N_18595);
and U26033 (N_26033,N_13290,N_11027);
xnor U26034 (N_26034,N_12339,N_19275);
nand U26035 (N_26035,N_13251,N_15984);
xor U26036 (N_26036,N_12510,N_15403);
nand U26037 (N_26037,N_18051,N_12631);
and U26038 (N_26038,N_15929,N_10901);
nor U26039 (N_26039,N_12895,N_17983);
and U26040 (N_26040,N_19254,N_19101);
and U26041 (N_26041,N_16932,N_14069);
or U26042 (N_26042,N_12144,N_15511);
nand U26043 (N_26043,N_11953,N_16937);
nand U26044 (N_26044,N_19178,N_10275);
and U26045 (N_26045,N_16783,N_13905);
nand U26046 (N_26046,N_10534,N_14734);
or U26047 (N_26047,N_13983,N_10672);
nor U26048 (N_26048,N_11987,N_14720);
nor U26049 (N_26049,N_13425,N_13741);
or U26050 (N_26050,N_14764,N_17231);
nor U26051 (N_26051,N_15657,N_11617);
or U26052 (N_26052,N_12382,N_10919);
xor U26053 (N_26053,N_12903,N_13464);
xnor U26054 (N_26054,N_19654,N_15911);
nor U26055 (N_26055,N_11638,N_16586);
and U26056 (N_26056,N_19288,N_19869);
nor U26057 (N_26057,N_11267,N_19955);
or U26058 (N_26058,N_14299,N_18940);
nand U26059 (N_26059,N_15344,N_19122);
nor U26060 (N_26060,N_17986,N_15000);
nand U26061 (N_26061,N_12418,N_17732);
or U26062 (N_26062,N_12393,N_14884);
nand U26063 (N_26063,N_16713,N_17515);
or U26064 (N_26064,N_18721,N_15350);
and U26065 (N_26065,N_19682,N_19354);
nand U26066 (N_26066,N_19033,N_19794);
and U26067 (N_26067,N_12650,N_12160);
nor U26068 (N_26068,N_11046,N_13316);
xor U26069 (N_26069,N_18420,N_16451);
nor U26070 (N_26070,N_17179,N_15038);
or U26071 (N_26071,N_13440,N_16525);
nand U26072 (N_26072,N_13618,N_12263);
and U26073 (N_26073,N_15036,N_18597);
or U26074 (N_26074,N_11137,N_11580);
nand U26075 (N_26075,N_18150,N_17715);
and U26076 (N_26076,N_18129,N_16511);
or U26077 (N_26077,N_15431,N_12400);
nand U26078 (N_26078,N_10164,N_15322);
xor U26079 (N_26079,N_12653,N_14139);
and U26080 (N_26080,N_18851,N_11104);
nand U26081 (N_26081,N_14905,N_14877);
nor U26082 (N_26082,N_12451,N_12470);
nor U26083 (N_26083,N_13111,N_17933);
or U26084 (N_26084,N_13155,N_11858);
nand U26085 (N_26085,N_10990,N_17263);
xnor U26086 (N_26086,N_14943,N_16224);
or U26087 (N_26087,N_15944,N_10521);
or U26088 (N_26088,N_10934,N_10772);
nand U26089 (N_26089,N_14451,N_19327);
xnor U26090 (N_26090,N_15970,N_19902);
xor U26091 (N_26091,N_10091,N_10765);
and U26092 (N_26092,N_11388,N_10200);
nand U26093 (N_26093,N_10332,N_18266);
nand U26094 (N_26094,N_13247,N_17957);
and U26095 (N_26095,N_17193,N_18971);
or U26096 (N_26096,N_15319,N_19636);
nor U26097 (N_26097,N_11025,N_10011);
nor U26098 (N_26098,N_16862,N_11748);
nand U26099 (N_26099,N_15472,N_11400);
nor U26100 (N_26100,N_17730,N_12515);
nand U26101 (N_26101,N_19960,N_12354);
nor U26102 (N_26102,N_15873,N_13634);
nor U26103 (N_26103,N_19053,N_13355);
xnor U26104 (N_26104,N_12505,N_12622);
and U26105 (N_26105,N_16648,N_15270);
and U26106 (N_26106,N_14444,N_15955);
xnor U26107 (N_26107,N_17231,N_10650);
or U26108 (N_26108,N_18228,N_14685);
nor U26109 (N_26109,N_18886,N_16495);
xnor U26110 (N_26110,N_19026,N_18820);
or U26111 (N_26111,N_17238,N_11267);
nor U26112 (N_26112,N_10227,N_16749);
or U26113 (N_26113,N_14162,N_14255);
and U26114 (N_26114,N_18873,N_19522);
or U26115 (N_26115,N_11664,N_14396);
nor U26116 (N_26116,N_17128,N_19044);
nor U26117 (N_26117,N_18391,N_16940);
xor U26118 (N_26118,N_11390,N_19680);
or U26119 (N_26119,N_17565,N_15080);
or U26120 (N_26120,N_14031,N_17523);
or U26121 (N_26121,N_10388,N_18630);
and U26122 (N_26122,N_16436,N_18108);
nor U26123 (N_26123,N_15133,N_18177);
xnor U26124 (N_26124,N_12565,N_12834);
xor U26125 (N_26125,N_14139,N_14448);
and U26126 (N_26126,N_16482,N_10752);
and U26127 (N_26127,N_15765,N_16809);
nor U26128 (N_26128,N_18472,N_13849);
xnor U26129 (N_26129,N_10242,N_12375);
nand U26130 (N_26130,N_19618,N_14947);
or U26131 (N_26131,N_15846,N_10100);
nand U26132 (N_26132,N_19637,N_10044);
nor U26133 (N_26133,N_16469,N_10506);
or U26134 (N_26134,N_18362,N_17057);
or U26135 (N_26135,N_15144,N_13878);
or U26136 (N_26136,N_15228,N_12286);
nor U26137 (N_26137,N_14510,N_17346);
and U26138 (N_26138,N_10816,N_15170);
nand U26139 (N_26139,N_15199,N_18340);
and U26140 (N_26140,N_17675,N_19066);
and U26141 (N_26141,N_10029,N_12234);
nor U26142 (N_26142,N_11429,N_15058);
nor U26143 (N_26143,N_13884,N_13402);
xor U26144 (N_26144,N_12412,N_19007);
and U26145 (N_26145,N_19607,N_15093);
nand U26146 (N_26146,N_11904,N_17518);
nand U26147 (N_26147,N_18235,N_19675);
nor U26148 (N_26148,N_18025,N_14898);
or U26149 (N_26149,N_15959,N_19141);
or U26150 (N_26150,N_17253,N_10921);
or U26151 (N_26151,N_16832,N_18674);
or U26152 (N_26152,N_11528,N_12386);
nand U26153 (N_26153,N_15175,N_12946);
and U26154 (N_26154,N_13315,N_19232);
or U26155 (N_26155,N_15536,N_18211);
and U26156 (N_26156,N_18843,N_19147);
nor U26157 (N_26157,N_12762,N_16228);
and U26158 (N_26158,N_10853,N_14258);
nand U26159 (N_26159,N_15853,N_11246);
nor U26160 (N_26160,N_16103,N_11807);
and U26161 (N_26161,N_18973,N_13141);
and U26162 (N_26162,N_17512,N_15724);
nor U26163 (N_26163,N_17141,N_18948);
nand U26164 (N_26164,N_11399,N_17050);
and U26165 (N_26165,N_18303,N_17044);
and U26166 (N_26166,N_11292,N_17527);
nand U26167 (N_26167,N_14059,N_15224);
nor U26168 (N_26168,N_11927,N_10090);
or U26169 (N_26169,N_12659,N_19334);
nor U26170 (N_26170,N_17594,N_11143);
or U26171 (N_26171,N_13205,N_10746);
nor U26172 (N_26172,N_14665,N_19566);
nor U26173 (N_26173,N_11630,N_19133);
xnor U26174 (N_26174,N_18746,N_13729);
nand U26175 (N_26175,N_14524,N_11934);
nand U26176 (N_26176,N_16468,N_17206);
nand U26177 (N_26177,N_11131,N_15815);
xnor U26178 (N_26178,N_11996,N_18440);
and U26179 (N_26179,N_11724,N_13698);
or U26180 (N_26180,N_16690,N_18487);
and U26181 (N_26181,N_15416,N_19640);
nand U26182 (N_26182,N_16231,N_10802);
nand U26183 (N_26183,N_10609,N_12459);
nor U26184 (N_26184,N_16973,N_15706);
xnor U26185 (N_26185,N_18973,N_12812);
and U26186 (N_26186,N_12213,N_11965);
or U26187 (N_26187,N_10691,N_14457);
nand U26188 (N_26188,N_11136,N_16655);
nor U26189 (N_26189,N_13298,N_11352);
nand U26190 (N_26190,N_12395,N_17400);
or U26191 (N_26191,N_16041,N_17030);
and U26192 (N_26192,N_12189,N_16109);
nand U26193 (N_26193,N_16651,N_14247);
xor U26194 (N_26194,N_12459,N_14479);
and U26195 (N_26195,N_14877,N_15915);
or U26196 (N_26196,N_12360,N_13570);
xor U26197 (N_26197,N_18958,N_15449);
and U26198 (N_26198,N_16630,N_19701);
or U26199 (N_26199,N_17665,N_18948);
nor U26200 (N_26200,N_16122,N_14689);
nand U26201 (N_26201,N_13474,N_18195);
xor U26202 (N_26202,N_16477,N_19320);
nor U26203 (N_26203,N_17401,N_19477);
nor U26204 (N_26204,N_11698,N_11510);
and U26205 (N_26205,N_16427,N_18661);
and U26206 (N_26206,N_12834,N_13307);
nand U26207 (N_26207,N_18863,N_18578);
or U26208 (N_26208,N_15009,N_18434);
and U26209 (N_26209,N_15852,N_11574);
or U26210 (N_26210,N_11962,N_16776);
nand U26211 (N_26211,N_10339,N_19381);
and U26212 (N_26212,N_17001,N_14229);
nand U26213 (N_26213,N_18733,N_10135);
or U26214 (N_26214,N_18731,N_10219);
nor U26215 (N_26215,N_18834,N_15008);
nor U26216 (N_26216,N_12461,N_11373);
and U26217 (N_26217,N_12418,N_11420);
or U26218 (N_26218,N_19890,N_18629);
or U26219 (N_26219,N_16021,N_16948);
or U26220 (N_26220,N_18014,N_11232);
and U26221 (N_26221,N_13950,N_15402);
or U26222 (N_26222,N_13839,N_19989);
nor U26223 (N_26223,N_17153,N_14948);
nor U26224 (N_26224,N_15444,N_10172);
or U26225 (N_26225,N_11647,N_13329);
and U26226 (N_26226,N_15680,N_14807);
xnor U26227 (N_26227,N_12282,N_16776);
xnor U26228 (N_26228,N_15831,N_12963);
nand U26229 (N_26229,N_13874,N_17507);
nand U26230 (N_26230,N_14693,N_13500);
or U26231 (N_26231,N_10155,N_13953);
or U26232 (N_26232,N_18761,N_12683);
xor U26233 (N_26233,N_18086,N_18698);
and U26234 (N_26234,N_13499,N_14004);
xnor U26235 (N_26235,N_16987,N_17326);
nand U26236 (N_26236,N_10085,N_12698);
nor U26237 (N_26237,N_15554,N_16845);
xnor U26238 (N_26238,N_14970,N_10341);
or U26239 (N_26239,N_16775,N_16908);
nand U26240 (N_26240,N_11094,N_17963);
or U26241 (N_26241,N_14171,N_15567);
or U26242 (N_26242,N_15758,N_14356);
and U26243 (N_26243,N_15097,N_15891);
nand U26244 (N_26244,N_13129,N_16211);
nor U26245 (N_26245,N_14472,N_13059);
and U26246 (N_26246,N_13011,N_11204);
and U26247 (N_26247,N_10577,N_12935);
and U26248 (N_26248,N_18201,N_12347);
nand U26249 (N_26249,N_19501,N_17455);
or U26250 (N_26250,N_16374,N_17990);
nand U26251 (N_26251,N_14819,N_14989);
nand U26252 (N_26252,N_10704,N_13933);
nand U26253 (N_26253,N_10821,N_15713);
and U26254 (N_26254,N_13474,N_17869);
xor U26255 (N_26255,N_18082,N_14414);
nor U26256 (N_26256,N_13681,N_10694);
nor U26257 (N_26257,N_13434,N_18352);
and U26258 (N_26258,N_11510,N_12895);
nor U26259 (N_26259,N_18572,N_12546);
xor U26260 (N_26260,N_17482,N_12876);
or U26261 (N_26261,N_10150,N_12888);
nor U26262 (N_26262,N_18192,N_14108);
and U26263 (N_26263,N_16086,N_18065);
nor U26264 (N_26264,N_12972,N_13201);
nor U26265 (N_26265,N_16972,N_12124);
and U26266 (N_26266,N_17321,N_10806);
xor U26267 (N_26267,N_13278,N_12545);
or U26268 (N_26268,N_11558,N_16851);
nor U26269 (N_26269,N_12890,N_17355);
nor U26270 (N_26270,N_10706,N_15232);
nor U26271 (N_26271,N_12928,N_18217);
or U26272 (N_26272,N_16173,N_18317);
xnor U26273 (N_26273,N_10677,N_14577);
xor U26274 (N_26274,N_17343,N_11433);
nand U26275 (N_26275,N_12993,N_14200);
nor U26276 (N_26276,N_10519,N_16280);
xor U26277 (N_26277,N_15746,N_12493);
and U26278 (N_26278,N_10729,N_15540);
and U26279 (N_26279,N_18209,N_10760);
or U26280 (N_26280,N_10504,N_17957);
and U26281 (N_26281,N_11687,N_16650);
nand U26282 (N_26282,N_18163,N_16463);
nor U26283 (N_26283,N_19509,N_11052);
and U26284 (N_26284,N_17229,N_16722);
nand U26285 (N_26285,N_10378,N_19493);
nand U26286 (N_26286,N_13905,N_15624);
or U26287 (N_26287,N_19359,N_17488);
nand U26288 (N_26288,N_12369,N_18703);
or U26289 (N_26289,N_14224,N_16197);
xor U26290 (N_26290,N_16369,N_13073);
nand U26291 (N_26291,N_11217,N_12945);
or U26292 (N_26292,N_10443,N_14614);
and U26293 (N_26293,N_15075,N_14893);
nand U26294 (N_26294,N_12878,N_18692);
nor U26295 (N_26295,N_11208,N_10360);
nand U26296 (N_26296,N_17013,N_11847);
and U26297 (N_26297,N_15020,N_14777);
xor U26298 (N_26298,N_10750,N_11028);
and U26299 (N_26299,N_14956,N_12318);
or U26300 (N_26300,N_10176,N_17772);
nand U26301 (N_26301,N_16035,N_19717);
xnor U26302 (N_26302,N_17178,N_12192);
or U26303 (N_26303,N_16176,N_17880);
nand U26304 (N_26304,N_19388,N_13642);
and U26305 (N_26305,N_11829,N_15322);
and U26306 (N_26306,N_19931,N_14561);
nand U26307 (N_26307,N_16216,N_18026);
nor U26308 (N_26308,N_18167,N_15074);
nand U26309 (N_26309,N_15768,N_16714);
and U26310 (N_26310,N_10395,N_15051);
nor U26311 (N_26311,N_18569,N_19659);
or U26312 (N_26312,N_16646,N_15071);
nor U26313 (N_26313,N_13127,N_16999);
and U26314 (N_26314,N_11187,N_14042);
nor U26315 (N_26315,N_18981,N_15564);
and U26316 (N_26316,N_16252,N_15706);
nor U26317 (N_26317,N_19137,N_12144);
nor U26318 (N_26318,N_18791,N_14284);
nor U26319 (N_26319,N_11214,N_17169);
or U26320 (N_26320,N_18987,N_14412);
nor U26321 (N_26321,N_14008,N_15397);
nor U26322 (N_26322,N_10373,N_17622);
nor U26323 (N_26323,N_19513,N_16492);
nand U26324 (N_26324,N_17692,N_16817);
or U26325 (N_26325,N_12685,N_14115);
and U26326 (N_26326,N_14048,N_15853);
xnor U26327 (N_26327,N_15722,N_16361);
or U26328 (N_26328,N_13806,N_10961);
and U26329 (N_26329,N_18654,N_15611);
xnor U26330 (N_26330,N_11479,N_14176);
nand U26331 (N_26331,N_10781,N_17661);
nor U26332 (N_26332,N_18059,N_19925);
and U26333 (N_26333,N_17667,N_18533);
nor U26334 (N_26334,N_11707,N_17398);
nor U26335 (N_26335,N_16460,N_17585);
and U26336 (N_26336,N_17495,N_16201);
xor U26337 (N_26337,N_14097,N_18198);
nand U26338 (N_26338,N_11396,N_18599);
nand U26339 (N_26339,N_10300,N_15913);
xnor U26340 (N_26340,N_14170,N_19468);
or U26341 (N_26341,N_17625,N_18576);
or U26342 (N_26342,N_16458,N_19931);
and U26343 (N_26343,N_13094,N_11046);
and U26344 (N_26344,N_17619,N_18039);
xnor U26345 (N_26345,N_18926,N_16740);
and U26346 (N_26346,N_19902,N_18014);
nor U26347 (N_26347,N_13411,N_12539);
nand U26348 (N_26348,N_14673,N_17707);
and U26349 (N_26349,N_14228,N_13605);
and U26350 (N_26350,N_16287,N_14318);
nand U26351 (N_26351,N_17428,N_14548);
or U26352 (N_26352,N_18968,N_18846);
xor U26353 (N_26353,N_17063,N_15856);
and U26354 (N_26354,N_12029,N_11029);
nand U26355 (N_26355,N_11247,N_15504);
nor U26356 (N_26356,N_13035,N_15150);
and U26357 (N_26357,N_17070,N_18272);
nor U26358 (N_26358,N_17275,N_12700);
or U26359 (N_26359,N_19545,N_15034);
and U26360 (N_26360,N_17907,N_17308);
or U26361 (N_26361,N_17279,N_11608);
nor U26362 (N_26362,N_11424,N_16552);
nand U26363 (N_26363,N_16840,N_13441);
and U26364 (N_26364,N_17514,N_11446);
or U26365 (N_26365,N_15665,N_16528);
nand U26366 (N_26366,N_17491,N_15681);
or U26367 (N_26367,N_14535,N_16245);
nand U26368 (N_26368,N_12039,N_13825);
or U26369 (N_26369,N_13110,N_15521);
and U26370 (N_26370,N_14657,N_12046);
nand U26371 (N_26371,N_14912,N_12156);
or U26372 (N_26372,N_15237,N_16389);
nand U26373 (N_26373,N_11122,N_16543);
and U26374 (N_26374,N_18746,N_12561);
and U26375 (N_26375,N_16909,N_14679);
nor U26376 (N_26376,N_10990,N_15394);
nand U26377 (N_26377,N_14042,N_13523);
nor U26378 (N_26378,N_13631,N_14193);
nor U26379 (N_26379,N_10274,N_10222);
or U26380 (N_26380,N_12212,N_10716);
nand U26381 (N_26381,N_13670,N_13146);
nand U26382 (N_26382,N_12764,N_15179);
nand U26383 (N_26383,N_17026,N_12989);
and U26384 (N_26384,N_17112,N_14827);
and U26385 (N_26385,N_10719,N_14500);
nand U26386 (N_26386,N_17150,N_15542);
or U26387 (N_26387,N_12699,N_10079);
nor U26388 (N_26388,N_10127,N_10605);
nor U26389 (N_26389,N_19331,N_19727);
and U26390 (N_26390,N_13498,N_12352);
and U26391 (N_26391,N_18730,N_19293);
and U26392 (N_26392,N_10145,N_17587);
and U26393 (N_26393,N_18065,N_13216);
or U26394 (N_26394,N_16190,N_14450);
nand U26395 (N_26395,N_11588,N_10518);
or U26396 (N_26396,N_19296,N_10744);
or U26397 (N_26397,N_16782,N_18094);
nand U26398 (N_26398,N_10856,N_16231);
and U26399 (N_26399,N_16914,N_19901);
nor U26400 (N_26400,N_14072,N_14992);
or U26401 (N_26401,N_15656,N_12267);
and U26402 (N_26402,N_12788,N_19572);
or U26403 (N_26403,N_11216,N_10154);
or U26404 (N_26404,N_15062,N_18885);
nor U26405 (N_26405,N_17272,N_10901);
and U26406 (N_26406,N_13660,N_13301);
nor U26407 (N_26407,N_11751,N_11475);
or U26408 (N_26408,N_16818,N_17999);
nor U26409 (N_26409,N_13161,N_11116);
xor U26410 (N_26410,N_16324,N_12115);
nor U26411 (N_26411,N_10019,N_10158);
nand U26412 (N_26412,N_17063,N_18083);
and U26413 (N_26413,N_12243,N_15390);
and U26414 (N_26414,N_16085,N_13491);
nand U26415 (N_26415,N_13949,N_10534);
nand U26416 (N_26416,N_13614,N_14072);
or U26417 (N_26417,N_13689,N_15782);
or U26418 (N_26418,N_10980,N_11819);
xor U26419 (N_26419,N_10825,N_17320);
nand U26420 (N_26420,N_19972,N_17775);
nor U26421 (N_26421,N_14840,N_10757);
xor U26422 (N_26422,N_12659,N_18219);
nand U26423 (N_26423,N_19562,N_14566);
and U26424 (N_26424,N_10017,N_17188);
nand U26425 (N_26425,N_18038,N_17449);
nor U26426 (N_26426,N_19814,N_15604);
nor U26427 (N_26427,N_10320,N_17851);
xnor U26428 (N_26428,N_16324,N_18531);
and U26429 (N_26429,N_19772,N_11541);
nor U26430 (N_26430,N_17702,N_16243);
or U26431 (N_26431,N_17624,N_19425);
nand U26432 (N_26432,N_18571,N_13628);
and U26433 (N_26433,N_19517,N_19670);
nand U26434 (N_26434,N_15214,N_17151);
nor U26435 (N_26435,N_16381,N_17982);
and U26436 (N_26436,N_14579,N_14069);
nor U26437 (N_26437,N_14050,N_18030);
or U26438 (N_26438,N_18597,N_15215);
nor U26439 (N_26439,N_18580,N_15453);
xor U26440 (N_26440,N_18175,N_13035);
and U26441 (N_26441,N_16928,N_18969);
or U26442 (N_26442,N_17363,N_11446);
nand U26443 (N_26443,N_11788,N_12412);
nand U26444 (N_26444,N_18924,N_11775);
xnor U26445 (N_26445,N_17597,N_18848);
xor U26446 (N_26446,N_16928,N_17065);
or U26447 (N_26447,N_14534,N_16656);
nor U26448 (N_26448,N_12942,N_17274);
nand U26449 (N_26449,N_12484,N_12989);
or U26450 (N_26450,N_16268,N_17979);
nand U26451 (N_26451,N_11173,N_18417);
xnor U26452 (N_26452,N_13539,N_11358);
nor U26453 (N_26453,N_17839,N_16275);
and U26454 (N_26454,N_16136,N_17221);
and U26455 (N_26455,N_16887,N_16899);
nand U26456 (N_26456,N_16634,N_12188);
nand U26457 (N_26457,N_11491,N_11629);
nor U26458 (N_26458,N_13871,N_12769);
and U26459 (N_26459,N_15307,N_15459);
or U26460 (N_26460,N_14333,N_10747);
nand U26461 (N_26461,N_13408,N_18033);
and U26462 (N_26462,N_13838,N_19266);
xnor U26463 (N_26463,N_17240,N_15696);
or U26464 (N_26464,N_19116,N_11128);
nor U26465 (N_26465,N_12973,N_12901);
nor U26466 (N_26466,N_17024,N_10516);
and U26467 (N_26467,N_16444,N_16070);
nand U26468 (N_26468,N_13854,N_18087);
or U26469 (N_26469,N_11481,N_17475);
and U26470 (N_26470,N_10523,N_18055);
or U26471 (N_26471,N_11782,N_19931);
nor U26472 (N_26472,N_10206,N_13157);
nand U26473 (N_26473,N_18075,N_19889);
nand U26474 (N_26474,N_19874,N_15013);
or U26475 (N_26475,N_13451,N_14797);
nor U26476 (N_26476,N_12920,N_16144);
nand U26477 (N_26477,N_17785,N_14192);
or U26478 (N_26478,N_18227,N_14757);
nor U26479 (N_26479,N_18835,N_16802);
and U26480 (N_26480,N_12308,N_11967);
or U26481 (N_26481,N_16606,N_15558);
nor U26482 (N_26482,N_18566,N_11944);
nor U26483 (N_26483,N_17068,N_13646);
and U26484 (N_26484,N_16551,N_15435);
nor U26485 (N_26485,N_11767,N_17096);
nand U26486 (N_26486,N_16872,N_16453);
xnor U26487 (N_26487,N_17009,N_11258);
or U26488 (N_26488,N_12946,N_13726);
nor U26489 (N_26489,N_18960,N_17243);
or U26490 (N_26490,N_14472,N_14040);
nand U26491 (N_26491,N_16239,N_12671);
and U26492 (N_26492,N_16493,N_13986);
or U26493 (N_26493,N_15041,N_19693);
and U26494 (N_26494,N_14155,N_15703);
nor U26495 (N_26495,N_14857,N_12281);
or U26496 (N_26496,N_11203,N_10254);
and U26497 (N_26497,N_17360,N_11182);
or U26498 (N_26498,N_12951,N_16189);
and U26499 (N_26499,N_18834,N_19993);
and U26500 (N_26500,N_13131,N_18994);
and U26501 (N_26501,N_14962,N_18454);
or U26502 (N_26502,N_15787,N_18665);
xnor U26503 (N_26503,N_19437,N_13441);
xnor U26504 (N_26504,N_14859,N_12142);
or U26505 (N_26505,N_13656,N_14424);
and U26506 (N_26506,N_19637,N_13318);
nand U26507 (N_26507,N_17394,N_16728);
and U26508 (N_26508,N_12148,N_15171);
nor U26509 (N_26509,N_10080,N_15380);
nor U26510 (N_26510,N_18503,N_16231);
nor U26511 (N_26511,N_12905,N_18641);
nand U26512 (N_26512,N_19869,N_13377);
nand U26513 (N_26513,N_17260,N_17948);
and U26514 (N_26514,N_13187,N_10341);
nor U26515 (N_26515,N_12199,N_13878);
nor U26516 (N_26516,N_17909,N_16621);
or U26517 (N_26517,N_11617,N_18384);
nand U26518 (N_26518,N_17761,N_15405);
xnor U26519 (N_26519,N_16828,N_11775);
nand U26520 (N_26520,N_16207,N_11395);
nand U26521 (N_26521,N_14651,N_11425);
nand U26522 (N_26522,N_10211,N_15966);
nand U26523 (N_26523,N_14167,N_12034);
nor U26524 (N_26524,N_14986,N_17919);
and U26525 (N_26525,N_10191,N_16999);
or U26526 (N_26526,N_13805,N_14670);
or U26527 (N_26527,N_14918,N_13863);
or U26528 (N_26528,N_15990,N_18559);
or U26529 (N_26529,N_14299,N_16179);
nand U26530 (N_26530,N_17430,N_18897);
or U26531 (N_26531,N_11522,N_10418);
nor U26532 (N_26532,N_18180,N_12097);
or U26533 (N_26533,N_11837,N_11875);
or U26534 (N_26534,N_18457,N_12479);
and U26535 (N_26535,N_15286,N_12404);
nand U26536 (N_26536,N_16800,N_16503);
or U26537 (N_26537,N_16499,N_10411);
and U26538 (N_26538,N_16229,N_16959);
nor U26539 (N_26539,N_18328,N_15055);
and U26540 (N_26540,N_14148,N_16857);
nand U26541 (N_26541,N_15891,N_12504);
or U26542 (N_26542,N_12185,N_19506);
and U26543 (N_26543,N_16800,N_15457);
nor U26544 (N_26544,N_14673,N_10341);
or U26545 (N_26545,N_14426,N_13372);
nor U26546 (N_26546,N_16285,N_19879);
or U26547 (N_26547,N_16576,N_12413);
and U26548 (N_26548,N_13101,N_17161);
nand U26549 (N_26549,N_10944,N_18651);
nand U26550 (N_26550,N_11938,N_16019);
nor U26551 (N_26551,N_11065,N_10360);
nand U26552 (N_26552,N_10545,N_13242);
or U26553 (N_26553,N_14635,N_18050);
or U26554 (N_26554,N_17518,N_17865);
and U26555 (N_26555,N_10159,N_14188);
or U26556 (N_26556,N_13690,N_18704);
and U26557 (N_26557,N_17717,N_11463);
nor U26558 (N_26558,N_12353,N_12389);
nor U26559 (N_26559,N_14203,N_15386);
or U26560 (N_26560,N_14638,N_12174);
nor U26561 (N_26561,N_11919,N_18964);
nand U26562 (N_26562,N_18045,N_14278);
xnor U26563 (N_26563,N_18222,N_11627);
nand U26564 (N_26564,N_16567,N_17844);
nand U26565 (N_26565,N_16414,N_12478);
and U26566 (N_26566,N_12816,N_11819);
and U26567 (N_26567,N_16592,N_12514);
nand U26568 (N_26568,N_19285,N_13001);
nor U26569 (N_26569,N_12210,N_14826);
nand U26570 (N_26570,N_11512,N_11139);
nor U26571 (N_26571,N_19482,N_18095);
or U26572 (N_26572,N_14464,N_12286);
xnor U26573 (N_26573,N_16385,N_19086);
nor U26574 (N_26574,N_12911,N_18257);
and U26575 (N_26575,N_15829,N_11210);
and U26576 (N_26576,N_17288,N_14431);
and U26577 (N_26577,N_18239,N_16295);
or U26578 (N_26578,N_17723,N_12001);
xnor U26579 (N_26579,N_14985,N_14679);
and U26580 (N_26580,N_10567,N_12010);
xor U26581 (N_26581,N_10331,N_16934);
nor U26582 (N_26582,N_15508,N_12584);
and U26583 (N_26583,N_10510,N_14238);
and U26584 (N_26584,N_16514,N_13196);
or U26585 (N_26585,N_19082,N_13779);
nor U26586 (N_26586,N_14023,N_15185);
or U26587 (N_26587,N_12396,N_15105);
nand U26588 (N_26588,N_16460,N_17638);
and U26589 (N_26589,N_10584,N_13600);
and U26590 (N_26590,N_18740,N_15600);
and U26591 (N_26591,N_14281,N_16396);
or U26592 (N_26592,N_13364,N_17253);
nand U26593 (N_26593,N_12617,N_14546);
nand U26594 (N_26594,N_18311,N_16198);
and U26595 (N_26595,N_11926,N_13121);
nor U26596 (N_26596,N_13773,N_17166);
or U26597 (N_26597,N_11351,N_13219);
or U26598 (N_26598,N_11065,N_14566);
or U26599 (N_26599,N_14155,N_15337);
and U26600 (N_26600,N_17073,N_12501);
nand U26601 (N_26601,N_19185,N_18538);
nand U26602 (N_26602,N_14382,N_19240);
nand U26603 (N_26603,N_14767,N_11610);
or U26604 (N_26604,N_19723,N_13288);
nand U26605 (N_26605,N_18102,N_12585);
and U26606 (N_26606,N_14558,N_13482);
nand U26607 (N_26607,N_11898,N_17813);
nand U26608 (N_26608,N_19295,N_16353);
nand U26609 (N_26609,N_16127,N_13172);
or U26610 (N_26610,N_16315,N_18435);
nand U26611 (N_26611,N_17243,N_19481);
and U26612 (N_26612,N_15945,N_19228);
or U26613 (N_26613,N_19869,N_10421);
and U26614 (N_26614,N_14723,N_14107);
and U26615 (N_26615,N_12869,N_10063);
nor U26616 (N_26616,N_18513,N_18120);
nor U26617 (N_26617,N_18190,N_11334);
and U26618 (N_26618,N_18369,N_12845);
or U26619 (N_26619,N_10088,N_13436);
nor U26620 (N_26620,N_13037,N_19156);
or U26621 (N_26621,N_18508,N_15580);
or U26622 (N_26622,N_12967,N_16973);
or U26623 (N_26623,N_18900,N_10812);
nand U26624 (N_26624,N_10701,N_11365);
and U26625 (N_26625,N_12787,N_12108);
or U26626 (N_26626,N_10530,N_16238);
and U26627 (N_26627,N_17435,N_12168);
or U26628 (N_26628,N_10058,N_16012);
nand U26629 (N_26629,N_17837,N_14902);
nor U26630 (N_26630,N_11770,N_16788);
xnor U26631 (N_26631,N_12709,N_13917);
and U26632 (N_26632,N_18248,N_11251);
nand U26633 (N_26633,N_12110,N_13117);
xnor U26634 (N_26634,N_13464,N_18161);
xnor U26635 (N_26635,N_10124,N_18176);
xnor U26636 (N_26636,N_11536,N_19052);
nand U26637 (N_26637,N_19690,N_12846);
and U26638 (N_26638,N_16137,N_19906);
or U26639 (N_26639,N_18951,N_19854);
xor U26640 (N_26640,N_19317,N_18235);
nor U26641 (N_26641,N_13649,N_17895);
nand U26642 (N_26642,N_13008,N_10442);
nand U26643 (N_26643,N_10132,N_11092);
nand U26644 (N_26644,N_10416,N_19641);
nand U26645 (N_26645,N_15631,N_13541);
and U26646 (N_26646,N_11088,N_13612);
and U26647 (N_26647,N_15473,N_15575);
and U26648 (N_26648,N_13145,N_14207);
nand U26649 (N_26649,N_15071,N_16099);
or U26650 (N_26650,N_10357,N_16213);
or U26651 (N_26651,N_17690,N_18362);
nor U26652 (N_26652,N_17577,N_11069);
nor U26653 (N_26653,N_13450,N_12684);
and U26654 (N_26654,N_19809,N_10715);
or U26655 (N_26655,N_10873,N_16101);
and U26656 (N_26656,N_16134,N_16852);
nor U26657 (N_26657,N_13368,N_16932);
nand U26658 (N_26658,N_19581,N_19261);
or U26659 (N_26659,N_19296,N_11174);
and U26660 (N_26660,N_19394,N_14074);
nor U26661 (N_26661,N_11074,N_16575);
nor U26662 (N_26662,N_18671,N_12238);
xor U26663 (N_26663,N_11681,N_19226);
xnor U26664 (N_26664,N_13129,N_18424);
or U26665 (N_26665,N_15626,N_10073);
or U26666 (N_26666,N_18892,N_16834);
and U26667 (N_26667,N_17164,N_11907);
or U26668 (N_26668,N_10758,N_12493);
nor U26669 (N_26669,N_10792,N_13387);
nor U26670 (N_26670,N_11654,N_15249);
and U26671 (N_26671,N_16816,N_17770);
nand U26672 (N_26672,N_10995,N_15342);
nand U26673 (N_26673,N_15851,N_17774);
nand U26674 (N_26674,N_11724,N_16661);
and U26675 (N_26675,N_14762,N_12401);
nor U26676 (N_26676,N_19680,N_12908);
nor U26677 (N_26677,N_19334,N_19913);
or U26678 (N_26678,N_12310,N_11315);
xor U26679 (N_26679,N_18180,N_14898);
nand U26680 (N_26680,N_17698,N_17001);
nor U26681 (N_26681,N_12870,N_10352);
or U26682 (N_26682,N_12067,N_13754);
or U26683 (N_26683,N_13031,N_12911);
and U26684 (N_26684,N_16413,N_18602);
nor U26685 (N_26685,N_17841,N_18553);
or U26686 (N_26686,N_13827,N_14221);
or U26687 (N_26687,N_16961,N_10465);
nor U26688 (N_26688,N_15955,N_19329);
or U26689 (N_26689,N_12754,N_13104);
or U26690 (N_26690,N_19827,N_11885);
or U26691 (N_26691,N_10599,N_13335);
or U26692 (N_26692,N_17807,N_11153);
nor U26693 (N_26693,N_16313,N_10844);
and U26694 (N_26694,N_12306,N_17833);
nand U26695 (N_26695,N_19084,N_17499);
and U26696 (N_26696,N_11719,N_16529);
or U26697 (N_26697,N_13710,N_11710);
nand U26698 (N_26698,N_19743,N_18885);
xnor U26699 (N_26699,N_14107,N_10486);
or U26700 (N_26700,N_13552,N_16560);
xnor U26701 (N_26701,N_16436,N_13271);
or U26702 (N_26702,N_13759,N_13103);
and U26703 (N_26703,N_15021,N_15042);
and U26704 (N_26704,N_19365,N_18056);
and U26705 (N_26705,N_17460,N_14191);
or U26706 (N_26706,N_15198,N_17010);
or U26707 (N_26707,N_16963,N_10267);
nor U26708 (N_26708,N_12234,N_17081);
nor U26709 (N_26709,N_14893,N_10973);
and U26710 (N_26710,N_10827,N_16130);
and U26711 (N_26711,N_13270,N_10704);
and U26712 (N_26712,N_12621,N_17369);
and U26713 (N_26713,N_19173,N_10362);
nor U26714 (N_26714,N_10081,N_15179);
and U26715 (N_26715,N_13854,N_18203);
xnor U26716 (N_26716,N_14642,N_14192);
nor U26717 (N_26717,N_13498,N_13076);
and U26718 (N_26718,N_16796,N_19523);
and U26719 (N_26719,N_14809,N_17595);
nor U26720 (N_26720,N_18786,N_16666);
or U26721 (N_26721,N_12281,N_18051);
and U26722 (N_26722,N_19190,N_10724);
nor U26723 (N_26723,N_13037,N_13128);
nand U26724 (N_26724,N_15533,N_14073);
xnor U26725 (N_26725,N_11626,N_16825);
nand U26726 (N_26726,N_18281,N_19523);
and U26727 (N_26727,N_10611,N_10996);
nand U26728 (N_26728,N_16570,N_13103);
nand U26729 (N_26729,N_12044,N_19636);
nor U26730 (N_26730,N_13058,N_17662);
and U26731 (N_26731,N_16497,N_13884);
xnor U26732 (N_26732,N_15913,N_19687);
nand U26733 (N_26733,N_18151,N_11016);
and U26734 (N_26734,N_14201,N_10154);
or U26735 (N_26735,N_19264,N_19040);
and U26736 (N_26736,N_17644,N_15170);
nand U26737 (N_26737,N_18593,N_14502);
or U26738 (N_26738,N_13711,N_16526);
and U26739 (N_26739,N_17796,N_13367);
and U26740 (N_26740,N_15879,N_19810);
nor U26741 (N_26741,N_17432,N_18312);
nand U26742 (N_26742,N_16691,N_12408);
nand U26743 (N_26743,N_10192,N_11589);
or U26744 (N_26744,N_18767,N_14271);
nor U26745 (N_26745,N_17189,N_11920);
nand U26746 (N_26746,N_18091,N_15296);
nor U26747 (N_26747,N_13746,N_17588);
nand U26748 (N_26748,N_14274,N_17359);
or U26749 (N_26749,N_11644,N_14111);
and U26750 (N_26750,N_19878,N_16127);
nand U26751 (N_26751,N_17729,N_10899);
and U26752 (N_26752,N_10885,N_16507);
nand U26753 (N_26753,N_14478,N_11000);
nand U26754 (N_26754,N_11624,N_12360);
and U26755 (N_26755,N_14319,N_18990);
nand U26756 (N_26756,N_12005,N_18974);
nand U26757 (N_26757,N_14407,N_12788);
nor U26758 (N_26758,N_18776,N_15697);
or U26759 (N_26759,N_19494,N_18932);
nand U26760 (N_26760,N_16730,N_17360);
nor U26761 (N_26761,N_10014,N_12757);
and U26762 (N_26762,N_14101,N_17737);
and U26763 (N_26763,N_10725,N_10737);
or U26764 (N_26764,N_17566,N_13862);
and U26765 (N_26765,N_17802,N_13324);
nor U26766 (N_26766,N_19094,N_19656);
and U26767 (N_26767,N_18991,N_14583);
and U26768 (N_26768,N_12455,N_18700);
nor U26769 (N_26769,N_18331,N_18539);
nand U26770 (N_26770,N_12719,N_16172);
and U26771 (N_26771,N_14840,N_13215);
and U26772 (N_26772,N_19765,N_18865);
nand U26773 (N_26773,N_16046,N_17826);
or U26774 (N_26774,N_19479,N_17933);
nand U26775 (N_26775,N_15451,N_16057);
and U26776 (N_26776,N_11344,N_17761);
or U26777 (N_26777,N_17608,N_16776);
or U26778 (N_26778,N_12607,N_18043);
nand U26779 (N_26779,N_15192,N_13493);
or U26780 (N_26780,N_13705,N_18972);
and U26781 (N_26781,N_12405,N_16329);
nor U26782 (N_26782,N_14890,N_17447);
nor U26783 (N_26783,N_13864,N_16820);
xnor U26784 (N_26784,N_13596,N_10754);
nand U26785 (N_26785,N_15936,N_15117);
and U26786 (N_26786,N_12693,N_10016);
or U26787 (N_26787,N_12291,N_12644);
or U26788 (N_26788,N_16888,N_15052);
and U26789 (N_26789,N_19121,N_14284);
or U26790 (N_26790,N_12851,N_11350);
or U26791 (N_26791,N_18380,N_19620);
nor U26792 (N_26792,N_11093,N_14116);
and U26793 (N_26793,N_10037,N_13148);
nor U26794 (N_26794,N_12996,N_16748);
nor U26795 (N_26795,N_12887,N_18630);
and U26796 (N_26796,N_15174,N_15126);
and U26797 (N_26797,N_10404,N_17409);
nor U26798 (N_26798,N_13668,N_15895);
nor U26799 (N_26799,N_10563,N_15125);
or U26800 (N_26800,N_16600,N_18456);
nor U26801 (N_26801,N_13897,N_11263);
nand U26802 (N_26802,N_15667,N_12793);
and U26803 (N_26803,N_10719,N_17522);
nor U26804 (N_26804,N_16075,N_15704);
or U26805 (N_26805,N_18600,N_11884);
and U26806 (N_26806,N_12438,N_19986);
nand U26807 (N_26807,N_18325,N_15931);
or U26808 (N_26808,N_13217,N_11812);
xnor U26809 (N_26809,N_16160,N_19681);
nor U26810 (N_26810,N_15143,N_10913);
or U26811 (N_26811,N_14915,N_10387);
and U26812 (N_26812,N_12444,N_16166);
nor U26813 (N_26813,N_16974,N_13679);
nand U26814 (N_26814,N_10145,N_12418);
and U26815 (N_26815,N_10655,N_10675);
xnor U26816 (N_26816,N_14932,N_16092);
nor U26817 (N_26817,N_10773,N_13053);
or U26818 (N_26818,N_13877,N_18967);
and U26819 (N_26819,N_19726,N_15398);
or U26820 (N_26820,N_18442,N_19773);
or U26821 (N_26821,N_14136,N_15954);
nor U26822 (N_26822,N_18132,N_17295);
xnor U26823 (N_26823,N_12616,N_12018);
nor U26824 (N_26824,N_19482,N_15246);
nor U26825 (N_26825,N_18032,N_18856);
xnor U26826 (N_26826,N_17626,N_16783);
nand U26827 (N_26827,N_10670,N_11563);
nand U26828 (N_26828,N_17124,N_11094);
nand U26829 (N_26829,N_11017,N_18659);
or U26830 (N_26830,N_16427,N_17921);
or U26831 (N_26831,N_15536,N_19401);
nand U26832 (N_26832,N_12378,N_14433);
and U26833 (N_26833,N_15265,N_13023);
nand U26834 (N_26834,N_13540,N_13868);
nand U26835 (N_26835,N_17651,N_12353);
or U26836 (N_26836,N_14702,N_16216);
nor U26837 (N_26837,N_12254,N_10844);
nor U26838 (N_26838,N_11233,N_17536);
and U26839 (N_26839,N_12659,N_12658);
nand U26840 (N_26840,N_11655,N_15112);
and U26841 (N_26841,N_17094,N_15281);
nand U26842 (N_26842,N_11240,N_11489);
nand U26843 (N_26843,N_14453,N_11857);
nor U26844 (N_26844,N_12452,N_19504);
nor U26845 (N_26845,N_14958,N_14493);
nand U26846 (N_26846,N_18399,N_15169);
and U26847 (N_26847,N_13118,N_12500);
nor U26848 (N_26848,N_15315,N_17003);
nand U26849 (N_26849,N_18838,N_17418);
and U26850 (N_26850,N_12395,N_17742);
nor U26851 (N_26851,N_14227,N_11755);
and U26852 (N_26852,N_14049,N_12156);
xor U26853 (N_26853,N_17546,N_15993);
or U26854 (N_26854,N_18789,N_18771);
and U26855 (N_26855,N_10787,N_15942);
nand U26856 (N_26856,N_10464,N_17659);
xnor U26857 (N_26857,N_19674,N_10006);
and U26858 (N_26858,N_13993,N_10360);
nand U26859 (N_26859,N_17663,N_10116);
xnor U26860 (N_26860,N_18612,N_13472);
xnor U26861 (N_26861,N_14257,N_14025);
nor U26862 (N_26862,N_10291,N_15515);
or U26863 (N_26863,N_14136,N_19492);
nor U26864 (N_26864,N_13268,N_17513);
xnor U26865 (N_26865,N_17259,N_17549);
and U26866 (N_26866,N_17988,N_15118);
xnor U26867 (N_26867,N_16313,N_19474);
or U26868 (N_26868,N_16602,N_11166);
xor U26869 (N_26869,N_14661,N_12667);
nand U26870 (N_26870,N_18411,N_17415);
or U26871 (N_26871,N_18154,N_16977);
and U26872 (N_26872,N_13971,N_18266);
and U26873 (N_26873,N_19243,N_15019);
nand U26874 (N_26874,N_12439,N_15171);
or U26875 (N_26875,N_17169,N_10314);
or U26876 (N_26876,N_10830,N_15196);
nor U26877 (N_26877,N_16731,N_11071);
and U26878 (N_26878,N_17139,N_14593);
nor U26879 (N_26879,N_10882,N_15014);
nand U26880 (N_26880,N_11547,N_12117);
or U26881 (N_26881,N_15748,N_11167);
nor U26882 (N_26882,N_19159,N_10810);
and U26883 (N_26883,N_11555,N_17784);
or U26884 (N_26884,N_11717,N_17628);
nor U26885 (N_26885,N_15918,N_12875);
and U26886 (N_26886,N_15032,N_18773);
nor U26887 (N_26887,N_18694,N_11010);
or U26888 (N_26888,N_11828,N_15680);
or U26889 (N_26889,N_12163,N_12637);
or U26890 (N_26890,N_11077,N_10092);
nor U26891 (N_26891,N_13979,N_10984);
or U26892 (N_26892,N_11867,N_14627);
nor U26893 (N_26893,N_16309,N_17410);
nand U26894 (N_26894,N_15436,N_15520);
or U26895 (N_26895,N_11699,N_11946);
and U26896 (N_26896,N_13964,N_10353);
or U26897 (N_26897,N_13134,N_17886);
and U26898 (N_26898,N_15184,N_16864);
nor U26899 (N_26899,N_19869,N_12986);
and U26900 (N_26900,N_10293,N_11700);
nand U26901 (N_26901,N_15329,N_18551);
nand U26902 (N_26902,N_18457,N_13738);
or U26903 (N_26903,N_11336,N_18182);
and U26904 (N_26904,N_19910,N_12234);
nor U26905 (N_26905,N_11587,N_11206);
nand U26906 (N_26906,N_15306,N_11643);
nor U26907 (N_26907,N_14365,N_11555);
or U26908 (N_26908,N_10419,N_18947);
and U26909 (N_26909,N_15259,N_13657);
nand U26910 (N_26910,N_17238,N_19022);
and U26911 (N_26911,N_13436,N_14841);
or U26912 (N_26912,N_14789,N_12124);
and U26913 (N_26913,N_12748,N_17299);
nand U26914 (N_26914,N_14699,N_16415);
and U26915 (N_26915,N_16654,N_19222);
nand U26916 (N_26916,N_13090,N_17642);
or U26917 (N_26917,N_16196,N_18947);
nor U26918 (N_26918,N_11068,N_14654);
and U26919 (N_26919,N_13910,N_17292);
nor U26920 (N_26920,N_17972,N_19226);
or U26921 (N_26921,N_12684,N_11289);
and U26922 (N_26922,N_17708,N_15770);
nand U26923 (N_26923,N_13770,N_15594);
nor U26924 (N_26924,N_14242,N_10114);
and U26925 (N_26925,N_18545,N_16086);
or U26926 (N_26926,N_15378,N_13626);
nand U26927 (N_26927,N_13657,N_18860);
and U26928 (N_26928,N_14559,N_15094);
nor U26929 (N_26929,N_10917,N_19708);
or U26930 (N_26930,N_16141,N_10259);
or U26931 (N_26931,N_10567,N_13495);
nand U26932 (N_26932,N_11717,N_16014);
and U26933 (N_26933,N_18064,N_16046);
or U26934 (N_26934,N_11714,N_16585);
nand U26935 (N_26935,N_10369,N_16855);
xor U26936 (N_26936,N_17758,N_16277);
nor U26937 (N_26937,N_11207,N_13395);
and U26938 (N_26938,N_12076,N_11823);
or U26939 (N_26939,N_11623,N_17172);
nand U26940 (N_26940,N_17975,N_13175);
nand U26941 (N_26941,N_19110,N_10805);
nand U26942 (N_26942,N_11402,N_17838);
nor U26943 (N_26943,N_18390,N_15719);
nor U26944 (N_26944,N_15269,N_10048);
nor U26945 (N_26945,N_16096,N_18215);
or U26946 (N_26946,N_15697,N_19285);
nand U26947 (N_26947,N_16390,N_13327);
xor U26948 (N_26948,N_14878,N_10917);
nor U26949 (N_26949,N_10246,N_16506);
and U26950 (N_26950,N_13089,N_18493);
and U26951 (N_26951,N_10449,N_13393);
nand U26952 (N_26952,N_16083,N_12304);
and U26953 (N_26953,N_19508,N_12085);
or U26954 (N_26954,N_16403,N_17112);
nor U26955 (N_26955,N_13270,N_19583);
nand U26956 (N_26956,N_12360,N_19348);
nor U26957 (N_26957,N_19686,N_13497);
and U26958 (N_26958,N_17080,N_18877);
nor U26959 (N_26959,N_18069,N_17592);
nand U26960 (N_26960,N_10854,N_12449);
nor U26961 (N_26961,N_18041,N_18424);
xnor U26962 (N_26962,N_17386,N_14824);
nand U26963 (N_26963,N_10637,N_11872);
and U26964 (N_26964,N_19243,N_10452);
nand U26965 (N_26965,N_17744,N_15451);
or U26966 (N_26966,N_18148,N_13662);
and U26967 (N_26967,N_19253,N_19740);
or U26968 (N_26968,N_17242,N_12003);
or U26969 (N_26969,N_14563,N_11781);
nor U26970 (N_26970,N_14338,N_16587);
nor U26971 (N_26971,N_16107,N_11712);
or U26972 (N_26972,N_16264,N_11462);
nand U26973 (N_26973,N_16767,N_16543);
or U26974 (N_26974,N_14610,N_12345);
nor U26975 (N_26975,N_18097,N_10323);
nand U26976 (N_26976,N_19792,N_16493);
and U26977 (N_26977,N_19476,N_12547);
nor U26978 (N_26978,N_19470,N_13885);
and U26979 (N_26979,N_18564,N_18530);
and U26980 (N_26980,N_18992,N_10449);
and U26981 (N_26981,N_19764,N_11294);
xnor U26982 (N_26982,N_19386,N_16896);
xor U26983 (N_26983,N_10729,N_15136);
nor U26984 (N_26984,N_16538,N_16543);
or U26985 (N_26985,N_14767,N_15721);
nand U26986 (N_26986,N_11343,N_10905);
nand U26987 (N_26987,N_15625,N_10192);
xor U26988 (N_26988,N_15461,N_15164);
and U26989 (N_26989,N_19926,N_10098);
and U26990 (N_26990,N_15725,N_16795);
or U26991 (N_26991,N_19852,N_17362);
or U26992 (N_26992,N_10516,N_13121);
xnor U26993 (N_26993,N_16936,N_14557);
nor U26994 (N_26994,N_10999,N_18471);
and U26995 (N_26995,N_16168,N_14899);
or U26996 (N_26996,N_10533,N_11171);
and U26997 (N_26997,N_17972,N_16699);
or U26998 (N_26998,N_13328,N_15380);
nor U26999 (N_26999,N_12060,N_14535);
or U27000 (N_27000,N_11549,N_11116);
nand U27001 (N_27001,N_19539,N_12666);
or U27002 (N_27002,N_10101,N_10304);
or U27003 (N_27003,N_18771,N_18801);
xor U27004 (N_27004,N_11454,N_17580);
or U27005 (N_27005,N_18288,N_10809);
or U27006 (N_27006,N_19413,N_11871);
nand U27007 (N_27007,N_11428,N_19638);
and U27008 (N_27008,N_17931,N_16303);
xnor U27009 (N_27009,N_12899,N_12997);
and U27010 (N_27010,N_18099,N_15723);
or U27011 (N_27011,N_15333,N_18594);
nor U27012 (N_27012,N_10853,N_14400);
or U27013 (N_27013,N_14109,N_10071);
xor U27014 (N_27014,N_17031,N_14922);
and U27015 (N_27015,N_15212,N_17168);
nor U27016 (N_27016,N_10158,N_12255);
nand U27017 (N_27017,N_10625,N_10356);
or U27018 (N_27018,N_17202,N_10152);
and U27019 (N_27019,N_14724,N_10448);
nor U27020 (N_27020,N_12004,N_17216);
nor U27021 (N_27021,N_14543,N_18248);
nor U27022 (N_27022,N_12731,N_14261);
xor U27023 (N_27023,N_10470,N_13361);
nand U27024 (N_27024,N_12125,N_17080);
nor U27025 (N_27025,N_17343,N_12164);
xor U27026 (N_27026,N_10773,N_13386);
nor U27027 (N_27027,N_16236,N_15729);
nor U27028 (N_27028,N_18045,N_18346);
xor U27029 (N_27029,N_16252,N_17186);
nand U27030 (N_27030,N_15101,N_11015);
nand U27031 (N_27031,N_16717,N_11946);
nor U27032 (N_27032,N_11346,N_18040);
and U27033 (N_27033,N_16770,N_12088);
nor U27034 (N_27034,N_13026,N_13102);
or U27035 (N_27035,N_14192,N_16488);
xor U27036 (N_27036,N_17987,N_18891);
nor U27037 (N_27037,N_14131,N_15080);
nand U27038 (N_27038,N_15942,N_11724);
nand U27039 (N_27039,N_15730,N_10614);
or U27040 (N_27040,N_12390,N_16903);
nor U27041 (N_27041,N_14354,N_17427);
xnor U27042 (N_27042,N_19074,N_15063);
or U27043 (N_27043,N_14463,N_17294);
and U27044 (N_27044,N_18727,N_11928);
nand U27045 (N_27045,N_17568,N_17951);
nor U27046 (N_27046,N_13491,N_18754);
and U27047 (N_27047,N_13786,N_18152);
or U27048 (N_27048,N_14644,N_11581);
nor U27049 (N_27049,N_14145,N_11925);
or U27050 (N_27050,N_15288,N_10621);
nand U27051 (N_27051,N_13518,N_17331);
nand U27052 (N_27052,N_13843,N_12648);
and U27053 (N_27053,N_17978,N_19853);
or U27054 (N_27054,N_14215,N_14430);
nand U27055 (N_27055,N_19739,N_14131);
nor U27056 (N_27056,N_10626,N_12373);
and U27057 (N_27057,N_11147,N_10511);
nand U27058 (N_27058,N_10449,N_15588);
or U27059 (N_27059,N_15043,N_17192);
nand U27060 (N_27060,N_16878,N_18117);
and U27061 (N_27061,N_16075,N_18679);
and U27062 (N_27062,N_10769,N_15826);
nor U27063 (N_27063,N_17991,N_10355);
or U27064 (N_27064,N_19420,N_17569);
nand U27065 (N_27065,N_13860,N_17491);
or U27066 (N_27066,N_16948,N_11897);
or U27067 (N_27067,N_12272,N_12931);
or U27068 (N_27068,N_12534,N_16596);
and U27069 (N_27069,N_17078,N_18351);
nor U27070 (N_27070,N_15054,N_11420);
or U27071 (N_27071,N_18490,N_15513);
nand U27072 (N_27072,N_19137,N_16251);
nand U27073 (N_27073,N_19750,N_16472);
or U27074 (N_27074,N_11513,N_14848);
nand U27075 (N_27075,N_19969,N_17854);
and U27076 (N_27076,N_17522,N_11030);
nor U27077 (N_27077,N_12841,N_13218);
nand U27078 (N_27078,N_19210,N_18086);
nor U27079 (N_27079,N_11039,N_11406);
or U27080 (N_27080,N_14880,N_12156);
or U27081 (N_27081,N_11265,N_15978);
nand U27082 (N_27082,N_11930,N_15654);
xnor U27083 (N_27083,N_17641,N_15771);
or U27084 (N_27084,N_17985,N_17987);
or U27085 (N_27085,N_15142,N_19813);
nor U27086 (N_27086,N_11936,N_10904);
nor U27087 (N_27087,N_14252,N_10707);
or U27088 (N_27088,N_18132,N_12853);
and U27089 (N_27089,N_17948,N_12391);
nand U27090 (N_27090,N_10558,N_18634);
nor U27091 (N_27091,N_19816,N_18113);
nand U27092 (N_27092,N_11722,N_16267);
nand U27093 (N_27093,N_16742,N_13947);
nor U27094 (N_27094,N_10133,N_14253);
xor U27095 (N_27095,N_15891,N_11523);
and U27096 (N_27096,N_18719,N_16771);
nor U27097 (N_27097,N_10642,N_18553);
xor U27098 (N_27098,N_14541,N_15589);
or U27099 (N_27099,N_15978,N_17497);
nor U27100 (N_27100,N_18049,N_16613);
or U27101 (N_27101,N_12870,N_11595);
and U27102 (N_27102,N_15551,N_15350);
or U27103 (N_27103,N_12108,N_16812);
xnor U27104 (N_27104,N_13842,N_14396);
nand U27105 (N_27105,N_12307,N_15781);
or U27106 (N_27106,N_12759,N_17232);
nor U27107 (N_27107,N_10646,N_17164);
nand U27108 (N_27108,N_19316,N_11637);
or U27109 (N_27109,N_17525,N_14657);
nor U27110 (N_27110,N_19050,N_19222);
and U27111 (N_27111,N_19006,N_11112);
nand U27112 (N_27112,N_14092,N_13443);
or U27113 (N_27113,N_19930,N_16491);
nand U27114 (N_27114,N_11824,N_15464);
or U27115 (N_27115,N_18098,N_10338);
and U27116 (N_27116,N_11790,N_13765);
and U27117 (N_27117,N_10165,N_15787);
nand U27118 (N_27118,N_12630,N_19363);
nor U27119 (N_27119,N_10022,N_10317);
nor U27120 (N_27120,N_18804,N_12113);
or U27121 (N_27121,N_10653,N_14956);
nor U27122 (N_27122,N_14116,N_12689);
nand U27123 (N_27123,N_16398,N_19805);
nand U27124 (N_27124,N_13853,N_17755);
or U27125 (N_27125,N_18935,N_15046);
and U27126 (N_27126,N_19714,N_14425);
and U27127 (N_27127,N_13629,N_18554);
and U27128 (N_27128,N_18911,N_11803);
and U27129 (N_27129,N_16944,N_16332);
nor U27130 (N_27130,N_11492,N_14718);
or U27131 (N_27131,N_15172,N_11572);
or U27132 (N_27132,N_15936,N_18409);
nand U27133 (N_27133,N_19725,N_17049);
nand U27134 (N_27134,N_14278,N_10961);
nand U27135 (N_27135,N_16301,N_11307);
nor U27136 (N_27136,N_10805,N_17591);
nand U27137 (N_27137,N_15276,N_17488);
or U27138 (N_27138,N_14102,N_11062);
or U27139 (N_27139,N_12213,N_17852);
nor U27140 (N_27140,N_18694,N_17557);
nor U27141 (N_27141,N_17080,N_16046);
and U27142 (N_27142,N_15679,N_19291);
nor U27143 (N_27143,N_15805,N_15325);
nor U27144 (N_27144,N_16904,N_17957);
and U27145 (N_27145,N_11594,N_19737);
nand U27146 (N_27146,N_18673,N_10045);
xnor U27147 (N_27147,N_14178,N_16196);
nor U27148 (N_27148,N_15268,N_11966);
nand U27149 (N_27149,N_19858,N_15399);
xnor U27150 (N_27150,N_11532,N_11444);
nand U27151 (N_27151,N_13247,N_16482);
nor U27152 (N_27152,N_12496,N_19019);
and U27153 (N_27153,N_11214,N_14649);
and U27154 (N_27154,N_18549,N_17949);
and U27155 (N_27155,N_12564,N_18732);
nor U27156 (N_27156,N_17897,N_16163);
or U27157 (N_27157,N_16438,N_18678);
nand U27158 (N_27158,N_10199,N_12680);
or U27159 (N_27159,N_13812,N_14690);
xnor U27160 (N_27160,N_18433,N_18111);
nand U27161 (N_27161,N_17202,N_16788);
or U27162 (N_27162,N_10817,N_14189);
or U27163 (N_27163,N_10761,N_12188);
xor U27164 (N_27164,N_13984,N_10078);
or U27165 (N_27165,N_18154,N_14656);
nand U27166 (N_27166,N_19611,N_12128);
or U27167 (N_27167,N_13549,N_12305);
nand U27168 (N_27168,N_16703,N_14313);
or U27169 (N_27169,N_15824,N_12433);
nor U27170 (N_27170,N_15633,N_18120);
nand U27171 (N_27171,N_11795,N_15949);
nand U27172 (N_27172,N_17153,N_17450);
nor U27173 (N_27173,N_19403,N_12509);
nand U27174 (N_27174,N_14740,N_15117);
and U27175 (N_27175,N_17103,N_11438);
or U27176 (N_27176,N_16261,N_11846);
and U27177 (N_27177,N_12671,N_16766);
xor U27178 (N_27178,N_12826,N_19650);
nor U27179 (N_27179,N_13701,N_13288);
nand U27180 (N_27180,N_11100,N_11716);
nor U27181 (N_27181,N_10534,N_13220);
nand U27182 (N_27182,N_19035,N_13667);
nand U27183 (N_27183,N_19985,N_17717);
nand U27184 (N_27184,N_13808,N_14914);
xor U27185 (N_27185,N_17547,N_11116);
and U27186 (N_27186,N_15800,N_15347);
nor U27187 (N_27187,N_10276,N_15210);
or U27188 (N_27188,N_14030,N_11021);
and U27189 (N_27189,N_12929,N_15684);
or U27190 (N_27190,N_19148,N_11082);
nand U27191 (N_27191,N_14763,N_11510);
nand U27192 (N_27192,N_19949,N_10039);
and U27193 (N_27193,N_15875,N_12798);
nand U27194 (N_27194,N_15741,N_14544);
nand U27195 (N_27195,N_17045,N_11536);
and U27196 (N_27196,N_14949,N_12788);
nand U27197 (N_27197,N_15725,N_15593);
nand U27198 (N_27198,N_12064,N_10443);
and U27199 (N_27199,N_11215,N_17555);
nand U27200 (N_27200,N_12774,N_10410);
and U27201 (N_27201,N_10063,N_16178);
nand U27202 (N_27202,N_15794,N_12146);
xnor U27203 (N_27203,N_13839,N_12116);
or U27204 (N_27204,N_14075,N_17736);
or U27205 (N_27205,N_14976,N_11261);
or U27206 (N_27206,N_18681,N_13973);
nand U27207 (N_27207,N_17343,N_14046);
nand U27208 (N_27208,N_19535,N_10973);
nor U27209 (N_27209,N_14730,N_12976);
or U27210 (N_27210,N_16492,N_15544);
nor U27211 (N_27211,N_15394,N_14901);
or U27212 (N_27212,N_11652,N_10605);
or U27213 (N_27213,N_15761,N_17720);
or U27214 (N_27214,N_19026,N_14490);
or U27215 (N_27215,N_14109,N_15988);
or U27216 (N_27216,N_14161,N_18734);
nand U27217 (N_27217,N_16501,N_11902);
or U27218 (N_27218,N_17886,N_18376);
or U27219 (N_27219,N_11516,N_10650);
and U27220 (N_27220,N_14528,N_11072);
or U27221 (N_27221,N_17604,N_18816);
or U27222 (N_27222,N_10487,N_11889);
xor U27223 (N_27223,N_18615,N_19150);
and U27224 (N_27224,N_17025,N_19647);
and U27225 (N_27225,N_14840,N_15841);
nor U27226 (N_27226,N_18791,N_11564);
or U27227 (N_27227,N_10593,N_19497);
nand U27228 (N_27228,N_12388,N_10946);
and U27229 (N_27229,N_13789,N_14125);
and U27230 (N_27230,N_10053,N_19788);
nor U27231 (N_27231,N_11921,N_17448);
nand U27232 (N_27232,N_12581,N_12542);
and U27233 (N_27233,N_12764,N_14653);
nand U27234 (N_27234,N_10861,N_14978);
and U27235 (N_27235,N_10012,N_17722);
and U27236 (N_27236,N_16345,N_14843);
xor U27237 (N_27237,N_19332,N_10356);
nand U27238 (N_27238,N_15816,N_13043);
nand U27239 (N_27239,N_17323,N_17893);
and U27240 (N_27240,N_19565,N_15327);
nor U27241 (N_27241,N_19952,N_14210);
nand U27242 (N_27242,N_16129,N_12226);
nor U27243 (N_27243,N_18585,N_14644);
or U27244 (N_27244,N_12729,N_13433);
nand U27245 (N_27245,N_11719,N_10039);
nor U27246 (N_27246,N_16769,N_14929);
xor U27247 (N_27247,N_15520,N_15358);
or U27248 (N_27248,N_13012,N_18792);
nand U27249 (N_27249,N_10771,N_15783);
and U27250 (N_27250,N_11131,N_15599);
xnor U27251 (N_27251,N_17678,N_13716);
nand U27252 (N_27252,N_12734,N_16594);
nor U27253 (N_27253,N_16162,N_11985);
nor U27254 (N_27254,N_10568,N_16179);
nor U27255 (N_27255,N_12832,N_11785);
xnor U27256 (N_27256,N_15156,N_19994);
nor U27257 (N_27257,N_16465,N_11572);
or U27258 (N_27258,N_11865,N_16329);
and U27259 (N_27259,N_15312,N_13103);
xnor U27260 (N_27260,N_12303,N_11899);
and U27261 (N_27261,N_19488,N_17280);
and U27262 (N_27262,N_14797,N_12442);
xnor U27263 (N_27263,N_11648,N_13812);
nand U27264 (N_27264,N_11271,N_13579);
and U27265 (N_27265,N_11983,N_13572);
nand U27266 (N_27266,N_16396,N_15447);
nand U27267 (N_27267,N_16061,N_15450);
or U27268 (N_27268,N_16339,N_15988);
or U27269 (N_27269,N_13081,N_17018);
xor U27270 (N_27270,N_16528,N_19676);
and U27271 (N_27271,N_18731,N_14987);
xnor U27272 (N_27272,N_12495,N_12907);
and U27273 (N_27273,N_18515,N_11328);
or U27274 (N_27274,N_12899,N_14291);
and U27275 (N_27275,N_12845,N_15658);
and U27276 (N_27276,N_12391,N_13410);
xor U27277 (N_27277,N_17016,N_18666);
xor U27278 (N_27278,N_14463,N_19748);
nand U27279 (N_27279,N_18985,N_16017);
or U27280 (N_27280,N_12705,N_16223);
or U27281 (N_27281,N_16113,N_13610);
and U27282 (N_27282,N_19358,N_14190);
and U27283 (N_27283,N_15625,N_13292);
nor U27284 (N_27284,N_10670,N_12345);
nand U27285 (N_27285,N_13205,N_13177);
or U27286 (N_27286,N_15446,N_19511);
or U27287 (N_27287,N_11787,N_16149);
nand U27288 (N_27288,N_17906,N_12807);
and U27289 (N_27289,N_19722,N_14254);
and U27290 (N_27290,N_16290,N_16530);
or U27291 (N_27291,N_17870,N_19967);
nor U27292 (N_27292,N_11403,N_15164);
xnor U27293 (N_27293,N_13655,N_18125);
and U27294 (N_27294,N_15306,N_14510);
and U27295 (N_27295,N_16008,N_17820);
nor U27296 (N_27296,N_13558,N_10568);
nor U27297 (N_27297,N_11720,N_16773);
nand U27298 (N_27298,N_10503,N_18600);
and U27299 (N_27299,N_10156,N_14468);
or U27300 (N_27300,N_15769,N_14005);
nand U27301 (N_27301,N_12239,N_11796);
nand U27302 (N_27302,N_10011,N_18913);
and U27303 (N_27303,N_18620,N_15995);
nor U27304 (N_27304,N_13543,N_13930);
nor U27305 (N_27305,N_15008,N_14085);
nand U27306 (N_27306,N_16629,N_16703);
nand U27307 (N_27307,N_19416,N_16201);
xor U27308 (N_27308,N_15272,N_13585);
and U27309 (N_27309,N_12682,N_16558);
and U27310 (N_27310,N_18544,N_17004);
nand U27311 (N_27311,N_16276,N_16136);
nor U27312 (N_27312,N_17976,N_17966);
or U27313 (N_27313,N_16252,N_11344);
nor U27314 (N_27314,N_16650,N_12799);
nand U27315 (N_27315,N_18164,N_15777);
nand U27316 (N_27316,N_16332,N_11775);
nor U27317 (N_27317,N_16294,N_15238);
nor U27318 (N_27318,N_17468,N_13893);
and U27319 (N_27319,N_15957,N_11524);
nand U27320 (N_27320,N_16296,N_17969);
or U27321 (N_27321,N_17412,N_18594);
and U27322 (N_27322,N_15815,N_16145);
nor U27323 (N_27323,N_10482,N_16361);
and U27324 (N_27324,N_11433,N_19194);
and U27325 (N_27325,N_18268,N_16840);
nor U27326 (N_27326,N_15143,N_18730);
nor U27327 (N_27327,N_19802,N_12388);
or U27328 (N_27328,N_10934,N_19526);
and U27329 (N_27329,N_13212,N_11816);
or U27330 (N_27330,N_18852,N_17697);
nand U27331 (N_27331,N_10872,N_10447);
or U27332 (N_27332,N_18664,N_10030);
or U27333 (N_27333,N_19601,N_19684);
or U27334 (N_27334,N_13978,N_12169);
nand U27335 (N_27335,N_13777,N_16386);
nor U27336 (N_27336,N_19215,N_18933);
nand U27337 (N_27337,N_16359,N_17270);
nor U27338 (N_27338,N_12467,N_18396);
or U27339 (N_27339,N_16369,N_13818);
or U27340 (N_27340,N_17683,N_12346);
or U27341 (N_27341,N_16892,N_19441);
or U27342 (N_27342,N_13393,N_15972);
nor U27343 (N_27343,N_14244,N_18131);
nor U27344 (N_27344,N_14570,N_14104);
nor U27345 (N_27345,N_13374,N_18988);
nor U27346 (N_27346,N_14362,N_15086);
and U27347 (N_27347,N_11443,N_15647);
nand U27348 (N_27348,N_18319,N_10626);
nand U27349 (N_27349,N_17789,N_14007);
or U27350 (N_27350,N_18188,N_16743);
nand U27351 (N_27351,N_10934,N_13968);
and U27352 (N_27352,N_16610,N_10307);
nor U27353 (N_27353,N_14908,N_17192);
nor U27354 (N_27354,N_10529,N_16276);
nor U27355 (N_27355,N_14438,N_10222);
and U27356 (N_27356,N_13216,N_12698);
nor U27357 (N_27357,N_17539,N_14587);
nand U27358 (N_27358,N_11593,N_17982);
nor U27359 (N_27359,N_15626,N_12850);
nand U27360 (N_27360,N_18152,N_10749);
or U27361 (N_27361,N_18725,N_15826);
or U27362 (N_27362,N_13324,N_14012);
and U27363 (N_27363,N_14054,N_13468);
and U27364 (N_27364,N_13189,N_16302);
or U27365 (N_27365,N_11905,N_10867);
nor U27366 (N_27366,N_14995,N_15522);
xor U27367 (N_27367,N_18592,N_11718);
or U27368 (N_27368,N_19254,N_19046);
nor U27369 (N_27369,N_12375,N_12420);
or U27370 (N_27370,N_14076,N_15020);
nor U27371 (N_27371,N_18906,N_13369);
nor U27372 (N_27372,N_13808,N_15509);
nand U27373 (N_27373,N_17602,N_18583);
nand U27374 (N_27374,N_14319,N_15778);
and U27375 (N_27375,N_17237,N_19750);
nor U27376 (N_27376,N_13653,N_11734);
xnor U27377 (N_27377,N_10482,N_18492);
and U27378 (N_27378,N_12854,N_19883);
and U27379 (N_27379,N_10094,N_18702);
and U27380 (N_27380,N_10474,N_15855);
and U27381 (N_27381,N_15543,N_19709);
nand U27382 (N_27382,N_13613,N_19602);
nor U27383 (N_27383,N_14192,N_17833);
or U27384 (N_27384,N_15698,N_12298);
or U27385 (N_27385,N_15729,N_18017);
and U27386 (N_27386,N_18017,N_16550);
nand U27387 (N_27387,N_14036,N_10487);
nand U27388 (N_27388,N_11575,N_15279);
nor U27389 (N_27389,N_13202,N_12723);
nand U27390 (N_27390,N_19186,N_15644);
and U27391 (N_27391,N_16568,N_15611);
nor U27392 (N_27392,N_12057,N_13255);
and U27393 (N_27393,N_19598,N_10218);
nor U27394 (N_27394,N_19831,N_11653);
nor U27395 (N_27395,N_19543,N_11471);
xor U27396 (N_27396,N_13010,N_12244);
nand U27397 (N_27397,N_16308,N_16516);
nor U27398 (N_27398,N_18653,N_14990);
and U27399 (N_27399,N_19612,N_17025);
nor U27400 (N_27400,N_10214,N_15537);
or U27401 (N_27401,N_18454,N_11894);
and U27402 (N_27402,N_13950,N_15579);
nor U27403 (N_27403,N_17683,N_13686);
nand U27404 (N_27404,N_10256,N_13457);
and U27405 (N_27405,N_10118,N_12835);
and U27406 (N_27406,N_14833,N_12691);
nor U27407 (N_27407,N_14535,N_12188);
nor U27408 (N_27408,N_16403,N_19285);
nor U27409 (N_27409,N_19066,N_15681);
nor U27410 (N_27410,N_12449,N_10327);
or U27411 (N_27411,N_19252,N_11828);
and U27412 (N_27412,N_16200,N_18804);
or U27413 (N_27413,N_10761,N_10048);
nor U27414 (N_27414,N_11510,N_16213);
nor U27415 (N_27415,N_16686,N_13624);
xor U27416 (N_27416,N_15293,N_12319);
nand U27417 (N_27417,N_14763,N_16000);
xor U27418 (N_27418,N_17612,N_18191);
and U27419 (N_27419,N_13251,N_13442);
or U27420 (N_27420,N_16661,N_16493);
and U27421 (N_27421,N_19741,N_12579);
nor U27422 (N_27422,N_11295,N_12291);
nand U27423 (N_27423,N_11480,N_16602);
nor U27424 (N_27424,N_13209,N_10094);
nand U27425 (N_27425,N_18438,N_19938);
nand U27426 (N_27426,N_17641,N_17226);
or U27427 (N_27427,N_17480,N_10433);
xnor U27428 (N_27428,N_13397,N_16179);
xor U27429 (N_27429,N_18060,N_10606);
or U27430 (N_27430,N_13561,N_10304);
nand U27431 (N_27431,N_14026,N_11009);
nor U27432 (N_27432,N_14210,N_19225);
or U27433 (N_27433,N_18899,N_17727);
and U27434 (N_27434,N_14733,N_12056);
nor U27435 (N_27435,N_19735,N_18188);
and U27436 (N_27436,N_15607,N_13436);
and U27437 (N_27437,N_16812,N_15869);
and U27438 (N_27438,N_17982,N_18709);
and U27439 (N_27439,N_19740,N_13769);
nand U27440 (N_27440,N_16015,N_14610);
nand U27441 (N_27441,N_15457,N_17797);
or U27442 (N_27442,N_14897,N_13264);
and U27443 (N_27443,N_17571,N_17125);
and U27444 (N_27444,N_11529,N_11233);
nor U27445 (N_27445,N_13711,N_16464);
and U27446 (N_27446,N_17612,N_18448);
or U27447 (N_27447,N_10681,N_16582);
nand U27448 (N_27448,N_14261,N_14718);
nor U27449 (N_27449,N_17860,N_14395);
nor U27450 (N_27450,N_14834,N_15253);
nor U27451 (N_27451,N_12446,N_10003);
nor U27452 (N_27452,N_18836,N_17832);
or U27453 (N_27453,N_14721,N_13232);
nand U27454 (N_27454,N_14786,N_15775);
nor U27455 (N_27455,N_10741,N_16748);
nor U27456 (N_27456,N_15905,N_15123);
nor U27457 (N_27457,N_14702,N_10700);
nand U27458 (N_27458,N_16553,N_14631);
or U27459 (N_27459,N_12777,N_14607);
nand U27460 (N_27460,N_14380,N_13544);
nand U27461 (N_27461,N_19533,N_15650);
nor U27462 (N_27462,N_16278,N_17830);
nand U27463 (N_27463,N_19990,N_16915);
xnor U27464 (N_27464,N_17933,N_11925);
or U27465 (N_27465,N_13054,N_18578);
nor U27466 (N_27466,N_13032,N_17989);
or U27467 (N_27467,N_12895,N_16362);
nand U27468 (N_27468,N_10875,N_13759);
or U27469 (N_27469,N_15548,N_17517);
nor U27470 (N_27470,N_18579,N_15120);
nand U27471 (N_27471,N_19508,N_17776);
and U27472 (N_27472,N_13159,N_11893);
nor U27473 (N_27473,N_11350,N_19909);
or U27474 (N_27474,N_19695,N_14353);
nand U27475 (N_27475,N_18053,N_14363);
or U27476 (N_27476,N_14225,N_16689);
or U27477 (N_27477,N_17484,N_17379);
nand U27478 (N_27478,N_10176,N_19783);
nor U27479 (N_27479,N_14296,N_12909);
xnor U27480 (N_27480,N_15938,N_10610);
and U27481 (N_27481,N_16496,N_15372);
and U27482 (N_27482,N_11184,N_10596);
xnor U27483 (N_27483,N_17160,N_12791);
or U27484 (N_27484,N_12290,N_11879);
nand U27485 (N_27485,N_10021,N_11976);
or U27486 (N_27486,N_11842,N_16823);
or U27487 (N_27487,N_16303,N_12089);
nor U27488 (N_27488,N_18372,N_10125);
or U27489 (N_27489,N_13444,N_19573);
and U27490 (N_27490,N_19390,N_14905);
nor U27491 (N_27491,N_19883,N_19726);
nand U27492 (N_27492,N_16199,N_13622);
nand U27493 (N_27493,N_15993,N_15925);
nand U27494 (N_27494,N_13292,N_17540);
and U27495 (N_27495,N_17220,N_10568);
nand U27496 (N_27496,N_17101,N_16886);
or U27497 (N_27497,N_11579,N_11248);
nor U27498 (N_27498,N_13428,N_16721);
nor U27499 (N_27499,N_19818,N_17280);
xnor U27500 (N_27500,N_18644,N_16045);
nand U27501 (N_27501,N_14070,N_17547);
and U27502 (N_27502,N_18794,N_11586);
or U27503 (N_27503,N_18007,N_14739);
or U27504 (N_27504,N_10057,N_17281);
xor U27505 (N_27505,N_17897,N_12695);
and U27506 (N_27506,N_19252,N_10278);
and U27507 (N_27507,N_17546,N_12565);
nor U27508 (N_27508,N_13253,N_18284);
nor U27509 (N_27509,N_11087,N_12008);
or U27510 (N_27510,N_16122,N_11036);
and U27511 (N_27511,N_11187,N_13483);
nor U27512 (N_27512,N_10871,N_15500);
and U27513 (N_27513,N_14470,N_19787);
or U27514 (N_27514,N_16485,N_17141);
nor U27515 (N_27515,N_15114,N_17256);
nor U27516 (N_27516,N_12484,N_10700);
and U27517 (N_27517,N_12148,N_15002);
nor U27518 (N_27518,N_10427,N_15227);
or U27519 (N_27519,N_17590,N_10436);
xnor U27520 (N_27520,N_11402,N_10298);
and U27521 (N_27521,N_18163,N_13133);
nand U27522 (N_27522,N_11057,N_16160);
nor U27523 (N_27523,N_11490,N_17606);
and U27524 (N_27524,N_19604,N_11261);
or U27525 (N_27525,N_17438,N_19616);
nor U27526 (N_27526,N_12383,N_17361);
or U27527 (N_27527,N_16676,N_11401);
nand U27528 (N_27528,N_19618,N_15976);
or U27529 (N_27529,N_13854,N_19129);
or U27530 (N_27530,N_15536,N_13032);
and U27531 (N_27531,N_17174,N_11167);
or U27532 (N_27532,N_12171,N_19977);
nand U27533 (N_27533,N_16820,N_12054);
and U27534 (N_27534,N_15618,N_16082);
and U27535 (N_27535,N_16744,N_12375);
nand U27536 (N_27536,N_17224,N_11142);
nor U27537 (N_27537,N_17403,N_15401);
nand U27538 (N_27538,N_13628,N_14607);
nand U27539 (N_27539,N_15241,N_13534);
or U27540 (N_27540,N_17696,N_19747);
xor U27541 (N_27541,N_12292,N_19220);
and U27542 (N_27542,N_18589,N_14771);
nand U27543 (N_27543,N_13336,N_15896);
nand U27544 (N_27544,N_12279,N_10760);
or U27545 (N_27545,N_13826,N_10971);
and U27546 (N_27546,N_15695,N_12292);
or U27547 (N_27547,N_13102,N_13597);
and U27548 (N_27548,N_18037,N_19470);
and U27549 (N_27549,N_10695,N_11495);
and U27550 (N_27550,N_18783,N_13346);
nand U27551 (N_27551,N_11605,N_14477);
nand U27552 (N_27552,N_16727,N_16593);
nor U27553 (N_27553,N_16259,N_15030);
xor U27554 (N_27554,N_19753,N_15230);
nand U27555 (N_27555,N_12139,N_18412);
and U27556 (N_27556,N_14917,N_16761);
or U27557 (N_27557,N_14799,N_16768);
nand U27558 (N_27558,N_10348,N_14907);
nand U27559 (N_27559,N_14908,N_14458);
or U27560 (N_27560,N_10884,N_12355);
and U27561 (N_27561,N_18939,N_10283);
or U27562 (N_27562,N_19612,N_17677);
and U27563 (N_27563,N_12047,N_14703);
and U27564 (N_27564,N_11344,N_18191);
nor U27565 (N_27565,N_16540,N_11779);
nor U27566 (N_27566,N_18009,N_13725);
or U27567 (N_27567,N_10934,N_14017);
or U27568 (N_27568,N_11924,N_12962);
and U27569 (N_27569,N_12937,N_18405);
nor U27570 (N_27570,N_14638,N_19278);
nor U27571 (N_27571,N_14079,N_18250);
nor U27572 (N_27572,N_10273,N_11388);
and U27573 (N_27573,N_19793,N_13181);
or U27574 (N_27574,N_11521,N_15012);
nand U27575 (N_27575,N_19461,N_12870);
nor U27576 (N_27576,N_11876,N_13899);
nor U27577 (N_27577,N_14444,N_18226);
or U27578 (N_27578,N_19404,N_15985);
nor U27579 (N_27579,N_10014,N_11194);
nor U27580 (N_27580,N_19981,N_18373);
and U27581 (N_27581,N_17367,N_11302);
nor U27582 (N_27582,N_14232,N_16031);
xnor U27583 (N_27583,N_17250,N_14348);
xnor U27584 (N_27584,N_19991,N_10635);
nor U27585 (N_27585,N_16310,N_15492);
nand U27586 (N_27586,N_15540,N_16162);
and U27587 (N_27587,N_17689,N_19093);
xnor U27588 (N_27588,N_11554,N_10970);
or U27589 (N_27589,N_18877,N_17177);
nor U27590 (N_27590,N_19997,N_11602);
nor U27591 (N_27591,N_14658,N_17651);
or U27592 (N_27592,N_17411,N_19067);
and U27593 (N_27593,N_15865,N_12619);
and U27594 (N_27594,N_18492,N_10506);
xor U27595 (N_27595,N_11125,N_13827);
or U27596 (N_27596,N_16362,N_10646);
and U27597 (N_27597,N_15139,N_12756);
nor U27598 (N_27598,N_15241,N_16759);
nor U27599 (N_27599,N_16331,N_14554);
nand U27600 (N_27600,N_14006,N_11329);
nor U27601 (N_27601,N_12110,N_12366);
and U27602 (N_27602,N_11354,N_13847);
nor U27603 (N_27603,N_15924,N_13904);
and U27604 (N_27604,N_11150,N_15943);
or U27605 (N_27605,N_14029,N_17134);
nor U27606 (N_27606,N_11847,N_17752);
xnor U27607 (N_27607,N_15608,N_10742);
nor U27608 (N_27608,N_10507,N_15533);
nand U27609 (N_27609,N_14866,N_15195);
nor U27610 (N_27610,N_19106,N_13526);
and U27611 (N_27611,N_15869,N_11925);
or U27612 (N_27612,N_13623,N_11951);
and U27613 (N_27613,N_18625,N_16986);
nor U27614 (N_27614,N_10527,N_18766);
or U27615 (N_27615,N_19697,N_16890);
and U27616 (N_27616,N_15362,N_12430);
and U27617 (N_27617,N_14686,N_11579);
nand U27618 (N_27618,N_16915,N_15604);
and U27619 (N_27619,N_11576,N_16929);
xor U27620 (N_27620,N_13520,N_19984);
and U27621 (N_27621,N_16061,N_14192);
or U27622 (N_27622,N_16096,N_13024);
nand U27623 (N_27623,N_19654,N_15836);
nor U27624 (N_27624,N_12118,N_19852);
or U27625 (N_27625,N_10186,N_18893);
xnor U27626 (N_27626,N_12741,N_17126);
or U27627 (N_27627,N_15958,N_12605);
nand U27628 (N_27628,N_13006,N_10781);
nand U27629 (N_27629,N_10712,N_19603);
nor U27630 (N_27630,N_15863,N_13651);
xnor U27631 (N_27631,N_16997,N_18662);
or U27632 (N_27632,N_12462,N_14462);
nor U27633 (N_27633,N_15052,N_15969);
nor U27634 (N_27634,N_13302,N_12738);
or U27635 (N_27635,N_19856,N_17572);
or U27636 (N_27636,N_10605,N_15197);
or U27637 (N_27637,N_15331,N_13589);
xor U27638 (N_27638,N_13126,N_11804);
or U27639 (N_27639,N_16452,N_11826);
nor U27640 (N_27640,N_18068,N_15898);
or U27641 (N_27641,N_17671,N_16708);
and U27642 (N_27642,N_19240,N_12521);
nor U27643 (N_27643,N_14319,N_16499);
and U27644 (N_27644,N_11602,N_10725);
nand U27645 (N_27645,N_13316,N_17258);
nor U27646 (N_27646,N_11471,N_10392);
nor U27647 (N_27647,N_11789,N_19007);
nor U27648 (N_27648,N_13802,N_19973);
or U27649 (N_27649,N_10618,N_14176);
and U27650 (N_27650,N_13430,N_17158);
and U27651 (N_27651,N_15640,N_12271);
nand U27652 (N_27652,N_14914,N_11065);
or U27653 (N_27653,N_14254,N_16867);
or U27654 (N_27654,N_10576,N_10704);
nor U27655 (N_27655,N_13448,N_11184);
nand U27656 (N_27656,N_19482,N_14276);
nor U27657 (N_27657,N_10899,N_18731);
and U27658 (N_27658,N_11862,N_12937);
or U27659 (N_27659,N_14858,N_12735);
or U27660 (N_27660,N_15553,N_15077);
xnor U27661 (N_27661,N_13220,N_10903);
nor U27662 (N_27662,N_13095,N_10861);
or U27663 (N_27663,N_12418,N_11403);
xor U27664 (N_27664,N_18557,N_19485);
nor U27665 (N_27665,N_10250,N_19822);
xor U27666 (N_27666,N_12225,N_11672);
or U27667 (N_27667,N_19754,N_10075);
and U27668 (N_27668,N_11174,N_19531);
and U27669 (N_27669,N_11035,N_19065);
or U27670 (N_27670,N_16471,N_13493);
xor U27671 (N_27671,N_10538,N_15198);
nand U27672 (N_27672,N_18782,N_11037);
and U27673 (N_27673,N_17836,N_14494);
or U27674 (N_27674,N_16697,N_15275);
nor U27675 (N_27675,N_19419,N_14549);
and U27676 (N_27676,N_13432,N_13625);
and U27677 (N_27677,N_12960,N_17064);
or U27678 (N_27678,N_17344,N_16869);
and U27679 (N_27679,N_17297,N_11402);
nand U27680 (N_27680,N_16263,N_15964);
nor U27681 (N_27681,N_13666,N_18629);
or U27682 (N_27682,N_12825,N_11181);
and U27683 (N_27683,N_16157,N_11571);
nor U27684 (N_27684,N_15925,N_15613);
nand U27685 (N_27685,N_19011,N_18076);
nand U27686 (N_27686,N_13960,N_16598);
nor U27687 (N_27687,N_10525,N_18787);
nor U27688 (N_27688,N_13822,N_14141);
nand U27689 (N_27689,N_17507,N_17529);
nand U27690 (N_27690,N_12387,N_17254);
or U27691 (N_27691,N_17752,N_11078);
or U27692 (N_27692,N_19589,N_12158);
and U27693 (N_27693,N_12863,N_19194);
and U27694 (N_27694,N_17370,N_12103);
and U27695 (N_27695,N_17833,N_14173);
nand U27696 (N_27696,N_10526,N_13209);
nor U27697 (N_27697,N_12599,N_19963);
xor U27698 (N_27698,N_13477,N_11003);
xnor U27699 (N_27699,N_17647,N_10169);
and U27700 (N_27700,N_14132,N_16547);
nor U27701 (N_27701,N_12070,N_17049);
or U27702 (N_27702,N_18878,N_18087);
nor U27703 (N_27703,N_11633,N_13612);
nand U27704 (N_27704,N_10110,N_11905);
or U27705 (N_27705,N_15835,N_16908);
and U27706 (N_27706,N_14790,N_15421);
nand U27707 (N_27707,N_17378,N_14037);
or U27708 (N_27708,N_13430,N_15383);
or U27709 (N_27709,N_16925,N_15231);
nand U27710 (N_27710,N_11912,N_19048);
or U27711 (N_27711,N_16481,N_15364);
nand U27712 (N_27712,N_14646,N_10297);
and U27713 (N_27713,N_11485,N_15732);
nor U27714 (N_27714,N_18509,N_14443);
and U27715 (N_27715,N_19900,N_10152);
nor U27716 (N_27716,N_15100,N_15986);
or U27717 (N_27717,N_11665,N_14462);
or U27718 (N_27718,N_19186,N_13836);
or U27719 (N_27719,N_14372,N_14145);
or U27720 (N_27720,N_17638,N_16197);
nor U27721 (N_27721,N_17789,N_15160);
nand U27722 (N_27722,N_12291,N_17310);
and U27723 (N_27723,N_11273,N_10904);
nand U27724 (N_27724,N_16181,N_16564);
nand U27725 (N_27725,N_13800,N_16844);
and U27726 (N_27726,N_12777,N_17359);
nand U27727 (N_27727,N_12994,N_15830);
nand U27728 (N_27728,N_10170,N_12105);
or U27729 (N_27729,N_11265,N_14378);
and U27730 (N_27730,N_19847,N_15212);
and U27731 (N_27731,N_14406,N_14337);
or U27732 (N_27732,N_19799,N_17663);
and U27733 (N_27733,N_12834,N_19235);
and U27734 (N_27734,N_19190,N_18228);
xor U27735 (N_27735,N_13517,N_16367);
nor U27736 (N_27736,N_10686,N_10588);
or U27737 (N_27737,N_14467,N_10095);
and U27738 (N_27738,N_10537,N_10342);
nand U27739 (N_27739,N_15984,N_15213);
nand U27740 (N_27740,N_17036,N_13096);
nand U27741 (N_27741,N_10720,N_15478);
nor U27742 (N_27742,N_15678,N_10335);
and U27743 (N_27743,N_15504,N_19660);
or U27744 (N_27744,N_10882,N_11950);
nand U27745 (N_27745,N_13831,N_15949);
nand U27746 (N_27746,N_13397,N_18640);
and U27747 (N_27747,N_16579,N_14368);
nand U27748 (N_27748,N_17596,N_12127);
and U27749 (N_27749,N_15377,N_17083);
and U27750 (N_27750,N_15866,N_17412);
and U27751 (N_27751,N_10989,N_11688);
nand U27752 (N_27752,N_15912,N_13360);
xnor U27753 (N_27753,N_17576,N_14542);
or U27754 (N_27754,N_13259,N_18751);
nor U27755 (N_27755,N_18865,N_12911);
and U27756 (N_27756,N_17667,N_10933);
and U27757 (N_27757,N_18226,N_18105);
xnor U27758 (N_27758,N_15620,N_19231);
nand U27759 (N_27759,N_10405,N_10847);
and U27760 (N_27760,N_15899,N_16844);
and U27761 (N_27761,N_13049,N_12692);
or U27762 (N_27762,N_12555,N_11719);
xor U27763 (N_27763,N_15421,N_15205);
and U27764 (N_27764,N_19065,N_12187);
and U27765 (N_27765,N_10297,N_14036);
or U27766 (N_27766,N_10149,N_12573);
and U27767 (N_27767,N_10445,N_10386);
and U27768 (N_27768,N_19648,N_10278);
nand U27769 (N_27769,N_17130,N_14480);
nor U27770 (N_27770,N_12994,N_13849);
nor U27771 (N_27771,N_17588,N_16732);
nor U27772 (N_27772,N_17846,N_10089);
and U27773 (N_27773,N_10627,N_11393);
or U27774 (N_27774,N_12147,N_10565);
xnor U27775 (N_27775,N_19334,N_13045);
nor U27776 (N_27776,N_19524,N_14249);
or U27777 (N_27777,N_18847,N_18519);
nand U27778 (N_27778,N_17204,N_10690);
or U27779 (N_27779,N_11420,N_15331);
nor U27780 (N_27780,N_18325,N_17159);
nand U27781 (N_27781,N_14126,N_18131);
xor U27782 (N_27782,N_18409,N_19515);
or U27783 (N_27783,N_13814,N_19979);
or U27784 (N_27784,N_15282,N_13258);
or U27785 (N_27785,N_10014,N_10762);
or U27786 (N_27786,N_13297,N_13864);
or U27787 (N_27787,N_11031,N_12776);
or U27788 (N_27788,N_13111,N_18866);
and U27789 (N_27789,N_10618,N_19332);
nor U27790 (N_27790,N_16864,N_12846);
nor U27791 (N_27791,N_19394,N_10416);
nor U27792 (N_27792,N_14585,N_10061);
nand U27793 (N_27793,N_11255,N_19731);
nor U27794 (N_27794,N_10776,N_18043);
or U27795 (N_27795,N_10926,N_19172);
and U27796 (N_27796,N_15444,N_16924);
nand U27797 (N_27797,N_16690,N_16944);
or U27798 (N_27798,N_13657,N_19591);
or U27799 (N_27799,N_11101,N_12436);
nor U27800 (N_27800,N_10328,N_17012);
xnor U27801 (N_27801,N_13267,N_16073);
and U27802 (N_27802,N_14526,N_11541);
nor U27803 (N_27803,N_12290,N_17139);
xor U27804 (N_27804,N_16591,N_14495);
nor U27805 (N_27805,N_10173,N_16224);
or U27806 (N_27806,N_13263,N_12494);
xor U27807 (N_27807,N_14804,N_19703);
and U27808 (N_27808,N_14576,N_19483);
nand U27809 (N_27809,N_13739,N_15850);
or U27810 (N_27810,N_19765,N_16851);
xor U27811 (N_27811,N_11000,N_13254);
nand U27812 (N_27812,N_15942,N_19727);
xnor U27813 (N_27813,N_12360,N_14678);
nor U27814 (N_27814,N_19255,N_19538);
and U27815 (N_27815,N_11291,N_19533);
nand U27816 (N_27816,N_14833,N_17440);
nor U27817 (N_27817,N_15161,N_11806);
or U27818 (N_27818,N_15595,N_18336);
and U27819 (N_27819,N_15576,N_13545);
or U27820 (N_27820,N_12580,N_14233);
or U27821 (N_27821,N_18012,N_15027);
and U27822 (N_27822,N_13395,N_19759);
and U27823 (N_27823,N_11619,N_16682);
or U27824 (N_27824,N_13350,N_15938);
xor U27825 (N_27825,N_19418,N_17352);
and U27826 (N_27826,N_15777,N_19468);
and U27827 (N_27827,N_11157,N_12757);
and U27828 (N_27828,N_12598,N_19273);
and U27829 (N_27829,N_13127,N_11420);
and U27830 (N_27830,N_12995,N_17680);
xnor U27831 (N_27831,N_11598,N_13946);
nand U27832 (N_27832,N_16773,N_11778);
or U27833 (N_27833,N_10405,N_13278);
nand U27834 (N_27834,N_11883,N_13251);
nand U27835 (N_27835,N_10224,N_12473);
nor U27836 (N_27836,N_18409,N_12140);
nor U27837 (N_27837,N_11879,N_11902);
and U27838 (N_27838,N_11289,N_12542);
xnor U27839 (N_27839,N_14127,N_10074);
xor U27840 (N_27840,N_10882,N_10375);
or U27841 (N_27841,N_14786,N_10518);
nor U27842 (N_27842,N_11455,N_13663);
nand U27843 (N_27843,N_12204,N_15189);
nand U27844 (N_27844,N_11796,N_16002);
or U27845 (N_27845,N_19654,N_16094);
nand U27846 (N_27846,N_18584,N_12757);
nor U27847 (N_27847,N_19949,N_17992);
or U27848 (N_27848,N_12770,N_15136);
nor U27849 (N_27849,N_15622,N_10194);
nand U27850 (N_27850,N_16521,N_19987);
nor U27851 (N_27851,N_15465,N_12399);
or U27852 (N_27852,N_10014,N_16240);
nor U27853 (N_27853,N_10566,N_14938);
and U27854 (N_27854,N_19921,N_19670);
or U27855 (N_27855,N_12184,N_11146);
and U27856 (N_27856,N_17041,N_12367);
and U27857 (N_27857,N_13960,N_17848);
xor U27858 (N_27858,N_16008,N_17492);
or U27859 (N_27859,N_14169,N_18998);
and U27860 (N_27860,N_18737,N_19053);
or U27861 (N_27861,N_11074,N_16333);
or U27862 (N_27862,N_14495,N_11930);
or U27863 (N_27863,N_16683,N_16631);
nor U27864 (N_27864,N_16456,N_11847);
nand U27865 (N_27865,N_12510,N_11377);
nand U27866 (N_27866,N_19630,N_17416);
nor U27867 (N_27867,N_17106,N_15885);
and U27868 (N_27868,N_12049,N_12284);
or U27869 (N_27869,N_14349,N_17539);
and U27870 (N_27870,N_15474,N_11131);
xor U27871 (N_27871,N_17627,N_11753);
or U27872 (N_27872,N_18411,N_17544);
or U27873 (N_27873,N_13860,N_11546);
nand U27874 (N_27874,N_10083,N_13013);
or U27875 (N_27875,N_19665,N_10957);
nand U27876 (N_27876,N_17453,N_16471);
xor U27877 (N_27877,N_16167,N_19798);
or U27878 (N_27878,N_18982,N_12878);
or U27879 (N_27879,N_16067,N_11416);
or U27880 (N_27880,N_11941,N_16564);
or U27881 (N_27881,N_18443,N_17562);
nand U27882 (N_27882,N_15361,N_10547);
nor U27883 (N_27883,N_11821,N_16394);
and U27884 (N_27884,N_12292,N_13821);
nand U27885 (N_27885,N_11208,N_15510);
and U27886 (N_27886,N_13165,N_19584);
and U27887 (N_27887,N_16107,N_11408);
nand U27888 (N_27888,N_11263,N_18491);
nor U27889 (N_27889,N_19025,N_10270);
nor U27890 (N_27890,N_17123,N_18854);
nor U27891 (N_27891,N_10137,N_17163);
and U27892 (N_27892,N_14596,N_19763);
nor U27893 (N_27893,N_10077,N_17433);
nor U27894 (N_27894,N_13971,N_13898);
nor U27895 (N_27895,N_15832,N_14685);
nand U27896 (N_27896,N_11603,N_14942);
or U27897 (N_27897,N_11645,N_16685);
nand U27898 (N_27898,N_11179,N_10990);
xor U27899 (N_27899,N_18712,N_17577);
or U27900 (N_27900,N_15669,N_17583);
nand U27901 (N_27901,N_11295,N_17623);
xnor U27902 (N_27902,N_13399,N_16346);
nand U27903 (N_27903,N_11168,N_19264);
nand U27904 (N_27904,N_12020,N_12910);
and U27905 (N_27905,N_11541,N_14624);
nor U27906 (N_27906,N_12503,N_12961);
nand U27907 (N_27907,N_11911,N_10339);
xnor U27908 (N_27908,N_19088,N_14797);
nor U27909 (N_27909,N_19175,N_11688);
or U27910 (N_27910,N_13678,N_10933);
nand U27911 (N_27911,N_16418,N_11726);
or U27912 (N_27912,N_14107,N_12432);
or U27913 (N_27913,N_15939,N_11285);
and U27914 (N_27914,N_18993,N_19319);
nor U27915 (N_27915,N_13491,N_15890);
or U27916 (N_27916,N_12276,N_12795);
or U27917 (N_27917,N_14776,N_16191);
xor U27918 (N_27918,N_12029,N_16475);
nor U27919 (N_27919,N_17241,N_15360);
nand U27920 (N_27920,N_13883,N_18780);
nor U27921 (N_27921,N_11464,N_13371);
and U27922 (N_27922,N_13805,N_17957);
nor U27923 (N_27923,N_18875,N_17019);
nor U27924 (N_27924,N_12711,N_15671);
or U27925 (N_27925,N_17766,N_18304);
nor U27926 (N_27926,N_16442,N_17474);
or U27927 (N_27927,N_13958,N_15700);
or U27928 (N_27928,N_13685,N_12508);
or U27929 (N_27929,N_13387,N_10671);
or U27930 (N_27930,N_13400,N_10392);
xnor U27931 (N_27931,N_10930,N_19725);
nor U27932 (N_27932,N_12699,N_17733);
xnor U27933 (N_27933,N_15039,N_16297);
nor U27934 (N_27934,N_14757,N_12451);
or U27935 (N_27935,N_14514,N_17847);
or U27936 (N_27936,N_11011,N_19571);
nand U27937 (N_27937,N_17978,N_11161);
and U27938 (N_27938,N_15776,N_18472);
nor U27939 (N_27939,N_16300,N_12215);
nor U27940 (N_27940,N_14009,N_16099);
and U27941 (N_27941,N_16515,N_18869);
or U27942 (N_27942,N_16907,N_12517);
nand U27943 (N_27943,N_13667,N_11075);
or U27944 (N_27944,N_14773,N_15214);
nor U27945 (N_27945,N_15605,N_17275);
nor U27946 (N_27946,N_18904,N_19288);
and U27947 (N_27947,N_13446,N_11282);
nor U27948 (N_27948,N_16671,N_13330);
nor U27949 (N_27949,N_15265,N_15239);
nand U27950 (N_27950,N_12823,N_12840);
or U27951 (N_27951,N_16718,N_11723);
nor U27952 (N_27952,N_19712,N_13703);
xnor U27953 (N_27953,N_19052,N_14508);
and U27954 (N_27954,N_13559,N_12239);
nor U27955 (N_27955,N_18751,N_10991);
nand U27956 (N_27956,N_19356,N_18246);
nand U27957 (N_27957,N_17618,N_13187);
or U27958 (N_27958,N_17741,N_16851);
nor U27959 (N_27959,N_10693,N_16742);
or U27960 (N_27960,N_10447,N_12440);
nand U27961 (N_27961,N_11425,N_16740);
nand U27962 (N_27962,N_19544,N_13888);
nor U27963 (N_27963,N_17686,N_16728);
or U27964 (N_27964,N_10075,N_16098);
and U27965 (N_27965,N_16580,N_15945);
or U27966 (N_27966,N_18797,N_18840);
xnor U27967 (N_27967,N_12611,N_18323);
nor U27968 (N_27968,N_18061,N_16280);
nand U27969 (N_27969,N_15226,N_18420);
nand U27970 (N_27970,N_13252,N_11583);
xnor U27971 (N_27971,N_14234,N_17530);
and U27972 (N_27972,N_16878,N_19164);
nor U27973 (N_27973,N_16769,N_19417);
xnor U27974 (N_27974,N_11746,N_10559);
or U27975 (N_27975,N_14102,N_13624);
or U27976 (N_27976,N_19496,N_17080);
nor U27977 (N_27977,N_17144,N_16423);
nand U27978 (N_27978,N_16580,N_14612);
or U27979 (N_27979,N_10988,N_10626);
or U27980 (N_27980,N_15524,N_11319);
nand U27981 (N_27981,N_17748,N_16678);
or U27982 (N_27982,N_11233,N_11296);
and U27983 (N_27983,N_19329,N_18661);
xnor U27984 (N_27984,N_10171,N_11678);
and U27985 (N_27985,N_10840,N_10895);
nand U27986 (N_27986,N_16324,N_12022);
nand U27987 (N_27987,N_16442,N_12012);
nand U27988 (N_27988,N_16149,N_16196);
nand U27989 (N_27989,N_19488,N_15374);
nor U27990 (N_27990,N_10302,N_11804);
or U27991 (N_27991,N_14273,N_16854);
xnor U27992 (N_27992,N_14051,N_12392);
nor U27993 (N_27993,N_17598,N_16164);
or U27994 (N_27994,N_17295,N_18192);
nor U27995 (N_27995,N_16352,N_17708);
nor U27996 (N_27996,N_13653,N_12420);
nor U27997 (N_27997,N_12557,N_14119);
nand U27998 (N_27998,N_11998,N_15704);
or U27999 (N_27999,N_18118,N_13364);
nand U28000 (N_28000,N_11397,N_15827);
or U28001 (N_28001,N_13761,N_14409);
nor U28002 (N_28002,N_12416,N_13336);
and U28003 (N_28003,N_14696,N_19015);
nand U28004 (N_28004,N_15712,N_11008);
nand U28005 (N_28005,N_11792,N_14646);
or U28006 (N_28006,N_17053,N_17542);
nor U28007 (N_28007,N_12464,N_12864);
nor U28008 (N_28008,N_17411,N_16872);
nand U28009 (N_28009,N_15369,N_19726);
nor U28010 (N_28010,N_14201,N_12488);
and U28011 (N_28011,N_14766,N_10622);
and U28012 (N_28012,N_10310,N_18474);
xnor U28013 (N_28013,N_14029,N_18143);
nand U28014 (N_28014,N_14358,N_13954);
and U28015 (N_28015,N_10005,N_11835);
nand U28016 (N_28016,N_16403,N_13487);
nor U28017 (N_28017,N_13519,N_18660);
and U28018 (N_28018,N_16026,N_12100);
xor U28019 (N_28019,N_18427,N_16705);
or U28020 (N_28020,N_18819,N_17186);
nor U28021 (N_28021,N_16848,N_18646);
or U28022 (N_28022,N_16325,N_16398);
or U28023 (N_28023,N_15122,N_19450);
xor U28024 (N_28024,N_19818,N_17808);
nand U28025 (N_28025,N_19773,N_15136);
nor U28026 (N_28026,N_19635,N_18257);
or U28027 (N_28027,N_12685,N_14131);
and U28028 (N_28028,N_17734,N_10752);
nand U28029 (N_28029,N_17900,N_10898);
or U28030 (N_28030,N_12373,N_10709);
nor U28031 (N_28031,N_10202,N_10963);
nor U28032 (N_28032,N_11804,N_16620);
nand U28033 (N_28033,N_16693,N_19122);
nor U28034 (N_28034,N_10204,N_12312);
or U28035 (N_28035,N_17423,N_10039);
and U28036 (N_28036,N_11380,N_14129);
nor U28037 (N_28037,N_11824,N_13646);
and U28038 (N_28038,N_13416,N_17560);
and U28039 (N_28039,N_16918,N_10910);
and U28040 (N_28040,N_14792,N_12216);
nand U28041 (N_28041,N_15983,N_14801);
xor U28042 (N_28042,N_19943,N_10360);
or U28043 (N_28043,N_14600,N_12522);
and U28044 (N_28044,N_16272,N_11662);
or U28045 (N_28045,N_15809,N_18039);
nand U28046 (N_28046,N_15567,N_16111);
nand U28047 (N_28047,N_10142,N_19589);
nor U28048 (N_28048,N_11680,N_17326);
and U28049 (N_28049,N_17161,N_16680);
nand U28050 (N_28050,N_19009,N_10502);
nand U28051 (N_28051,N_19281,N_12626);
and U28052 (N_28052,N_16980,N_16245);
nor U28053 (N_28053,N_18070,N_13384);
or U28054 (N_28054,N_15228,N_14587);
nand U28055 (N_28055,N_10290,N_16837);
nor U28056 (N_28056,N_10961,N_10670);
and U28057 (N_28057,N_19545,N_11939);
nand U28058 (N_28058,N_13628,N_19107);
and U28059 (N_28059,N_14120,N_13797);
xor U28060 (N_28060,N_11102,N_11755);
and U28061 (N_28061,N_16145,N_14013);
and U28062 (N_28062,N_13803,N_11470);
and U28063 (N_28063,N_16665,N_12644);
xor U28064 (N_28064,N_16291,N_11426);
nand U28065 (N_28065,N_14269,N_10632);
or U28066 (N_28066,N_11269,N_19567);
or U28067 (N_28067,N_14468,N_16333);
nor U28068 (N_28068,N_15536,N_18505);
or U28069 (N_28069,N_12034,N_16410);
and U28070 (N_28070,N_13425,N_15830);
and U28071 (N_28071,N_19056,N_15737);
nand U28072 (N_28072,N_12282,N_12449);
xnor U28073 (N_28073,N_13602,N_14779);
nor U28074 (N_28074,N_15691,N_16879);
nand U28075 (N_28075,N_15010,N_19983);
xor U28076 (N_28076,N_14761,N_17366);
nor U28077 (N_28077,N_18319,N_12733);
xor U28078 (N_28078,N_18046,N_19167);
nor U28079 (N_28079,N_18882,N_12100);
xnor U28080 (N_28080,N_10928,N_16510);
xnor U28081 (N_28081,N_18427,N_10299);
or U28082 (N_28082,N_10247,N_18606);
or U28083 (N_28083,N_12924,N_13125);
and U28084 (N_28084,N_12639,N_18512);
nand U28085 (N_28085,N_18081,N_11944);
nor U28086 (N_28086,N_17416,N_17500);
and U28087 (N_28087,N_16163,N_10425);
nor U28088 (N_28088,N_11177,N_15580);
and U28089 (N_28089,N_10972,N_15345);
or U28090 (N_28090,N_11901,N_19272);
nor U28091 (N_28091,N_14322,N_17642);
or U28092 (N_28092,N_10060,N_15691);
and U28093 (N_28093,N_19895,N_19613);
nor U28094 (N_28094,N_10717,N_19004);
or U28095 (N_28095,N_16006,N_16785);
or U28096 (N_28096,N_11265,N_19560);
nand U28097 (N_28097,N_14997,N_12868);
nor U28098 (N_28098,N_17591,N_18719);
nor U28099 (N_28099,N_10074,N_17172);
nor U28100 (N_28100,N_11744,N_10975);
nor U28101 (N_28101,N_19898,N_17051);
nor U28102 (N_28102,N_18368,N_15634);
nand U28103 (N_28103,N_15461,N_15050);
and U28104 (N_28104,N_16558,N_13228);
nand U28105 (N_28105,N_18692,N_14211);
or U28106 (N_28106,N_10483,N_18233);
or U28107 (N_28107,N_19905,N_13314);
xor U28108 (N_28108,N_14674,N_16286);
and U28109 (N_28109,N_11257,N_18781);
nor U28110 (N_28110,N_19273,N_19653);
or U28111 (N_28111,N_10444,N_13228);
nor U28112 (N_28112,N_18358,N_11501);
or U28113 (N_28113,N_19831,N_12470);
nor U28114 (N_28114,N_11193,N_12541);
nor U28115 (N_28115,N_13497,N_19036);
and U28116 (N_28116,N_18008,N_15589);
nor U28117 (N_28117,N_13552,N_19121);
nor U28118 (N_28118,N_15357,N_15310);
nand U28119 (N_28119,N_13059,N_18665);
and U28120 (N_28120,N_18490,N_12780);
nand U28121 (N_28121,N_13365,N_10800);
nand U28122 (N_28122,N_19004,N_12215);
nor U28123 (N_28123,N_15892,N_13468);
or U28124 (N_28124,N_16813,N_14600);
and U28125 (N_28125,N_14755,N_13945);
nor U28126 (N_28126,N_17399,N_13417);
nand U28127 (N_28127,N_10918,N_14332);
nand U28128 (N_28128,N_18805,N_10690);
nor U28129 (N_28129,N_13774,N_15221);
nor U28130 (N_28130,N_12921,N_11825);
nand U28131 (N_28131,N_11437,N_14272);
nand U28132 (N_28132,N_15942,N_15372);
and U28133 (N_28133,N_12151,N_16924);
and U28134 (N_28134,N_16565,N_19398);
nand U28135 (N_28135,N_11272,N_12545);
nand U28136 (N_28136,N_18916,N_13948);
and U28137 (N_28137,N_14865,N_17759);
nor U28138 (N_28138,N_18875,N_19789);
and U28139 (N_28139,N_17732,N_16299);
nand U28140 (N_28140,N_10607,N_11451);
or U28141 (N_28141,N_18238,N_16480);
or U28142 (N_28142,N_19695,N_16237);
nand U28143 (N_28143,N_17185,N_19174);
nor U28144 (N_28144,N_16508,N_10250);
and U28145 (N_28145,N_13546,N_12099);
nand U28146 (N_28146,N_15517,N_17648);
nand U28147 (N_28147,N_18902,N_12601);
or U28148 (N_28148,N_16159,N_10142);
nor U28149 (N_28149,N_11831,N_10685);
nand U28150 (N_28150,N_14658,N_15596);
and U28151 (N_28151,N_15811,N_12611);
or U28152 (N_28152,N_17579,N_18920);
nand U28153 (N_28153,N_13460,N_14546);
or U28154 (N_28154,N_18180,N_18035);
or U28155 (N_28155,N_16103,N_17691);
and U28156 (N_28156,N_19735,N_11453);
nand U28157 (N_28157,N_17532,N_12999);
and U28158 (N_28158,N_14732,N_14498);
nand U28159 (N_28159,N_19750,N_15410);
nand U28160 (N_28160,N_16930,N_12749);
nor U28161 (N_28161,N_15862,N_17342);
and U28162 (N_28162,N_10406,N_18092);
nand U28163 (N_28163,N_11784,N_13218);
nor U28164 (N_28164,N_13844,N_15432);
nor U28165 (N_28165,N_16948,N_12559);
nand U28166 (N_28166,N_18266,N_13231);
and U28167 (N_28167,N_10171,N_16785);
or U28168 (N_28168,N_17156,N_12734);
and U28169 (N_28169,N_14662,N_14256);
nand U28170 (N_28170,N_18776,N_10945);
and U28171 (N_28171,N_11419,N_11787);
nor U28172 (N_28172,N_10468,N_13631);
or U28173 (N_28173,N_10900,N_10992);
and U28174 (N_28174,N_16227,N_19443);
and U28175 (N_28175,N_11034,N_16429);
nand U28176 (N_28176,N_13367,N_17723);
nand U28177 (N_28177,N_15404,N_17384);
xnor U28178 (N_28178,N_18871,N_17347);
nor U28179 (N_28179,N_17365,N_12443);
xor U28180 (N_28180,N_11236,N_11560);
or U28181 (N_28181,N_19154,N_17726);
and U28182 (N_28182,N_10341,N_13915);
nor U28183 (N_28183,N_14809,N_18445);
nor U28184 (N_28184,N_13405,N_18315);
nand U28185 (N_28185,N_19474,N_12169);
xnor U28186 (N_28186,N_15919,N_19588);
nand U28187 (N_28187,N_19406,N_12618);
xnor U28188 (N_28188,N_14590,N_10467);
nor U28189 (N_28189,N_13221,N_15389);
nor U28190 (N_28190,N_10762,N_17113);
nor U28191 (N_28191,N_16205,N_13086);
nand U28192 (N_28192,N_12718,N_19152);
and U28193 (N_28193,N_11673,N_13228);
and U28194 (N_28194,N_17159,N_12703);
xor U28195 (N_28195,N_19613,N_13573);
or U28196 (N_28196,N_19977,N_18405);
and U28197 (N_28197,N_16130,N_16463);
nor U28198 (N_28198,N_10627,N_11641);
nand U28199 (N_28199,N_11365,N_15597);
xor U28200 (N_28200,N_16495,N_10695);
nor U28201 (N_28201,N_14751,N_12618);
nand U28202 (N_28202,N_17761,N_18463);
and U28203 (N_28203,N_14995,N_10633);
and U28204 (N_28204,N_13975,N_15287);
or U28205 (N_28205,N_16773,N_10668);
nor U28206 (N_28206,N_19188,N_11234);
nand U28207 (N_28207,N_12855,N_12903);
or U28208 (N_28208,N_14032,N_18321);
nand U28209 (N_28209,N_12980,N_11514);
nand U28210 (N_28210,N_15040,N_15001);
nand U28211 (N_28211,N_18592,N_14108);
nor U28212 (N_28212,N_11890,N_18807);
or U28213 (N_28213,N_10766,N_15883);
nand U28214 (N_28214,N_14533,N_19594);
and U28215 (N_28215,N_11032,N_13253);
and U28216 (N_28216,N_14643,N_18610);
nand U28217 (N_28217,N_19549,N_17465);
nand U28218 (N_28218,N_19586,N_14096);
xor U28219 (N_28219,N_19306,N_19884);
nor U28220 (N_28220,N_14776,N_19098);
nor U28221 (N_28221,N_16844,N_11141);
nor U28222 (N_28222,N_19982,N_13387);
and U28223 (N_28223,N_16786,N_19611);
nand U28224 (N_28224,N_15940,N_17925);
and U28225 (N_28225,N_15932,N_12895);
or U28226 (N_28226,N_12350,N_14273);
nor U28227 (N_28227,N_14582,N_13897);
nand U28228 (N_28228,N_17639,N_13369);
and U28229 (N_28229,N_18731,N_18126);
or U28230 (N_28230,N_12509,N_16105);
or U28231 (N_28231,N_10396,N_16465);
and U28232 (N_28232,N_12048,N_19447);
nor U28233 (N_28233,N_16654,N_12989);
or U28234 (N_28234,N_19309,N_12133);
and U28235 (N_28235,N_19414,N_11220);
and U28236 (N_28236,N_12924,N_12214);
and U28237 (N_28237,N_11941,N_17382);
or U28238 (N_28238,N_12659,N_10218);
nand U28239 (N_28239,N_17826,N_11617);
or U28240 (N_28240,N_17402,N_11815);
nand U28241 (N_28241,N_16588,N_18760);
and U28242 (N_28242,N_14009,N_15727);
or U28243 (N_28243,N_17487,N_12495);
nor U28244 (N_28244,N_16005,N_18451);
or U28245 (N_28245,N_12280,N_14310);
nor U28246 (N_28246,N_18504,N_12220);
nor U28247 (N_28247,N_10929,N_19993);
or U28248 (N_28248,N_13671,N_11405);
or U28249 (N_28249,N_18476,N_14429);
and U28250 (N_28250,N_12373,N_17878);
or U28251 (N_28251,N_15306,N_11088);
nor U28252 (N_28252,N_10811,N_15556);
or U28253 (N_28253,N_17467,N_19375);
xor U28254 (N_28254,N_19720,N_14911);
xor U28255 (N_28255,N_18834,N_17369);
xor U28256 (N_28256,N_12190,N_11080);
nand U28257 (N_28257,N_12897,N_11904);
or U28258 (N_28258,N_10381,N_19593);
or U28259 (N_28259,N_12067,N_15042);
nand U28260 (N_28260,N_14488,N_14951);
xor U28261 (N_28261,N_11231,N_10217);
nor U28262 (N_28262,N_16528,N_17804);
xnor U28263 (N_28263,N_15887,N_19337);
xnor U28264 (N_28264,N_14408,N_12306);
and U28265 (N_28265,N_15945,N_11200);
nor U28266 (N_28266,N_13443,N_18633);
and U28267 (N_28267,N_15142,N_16837);
nand U28268 (N_28268,N_19935,N_12547);
nand U28269 (N_28269,N_12145,N_12579);
and U28270 (N_28270,N_14460,N_13024);
or U28271 (N_28271,N_18765,N_10377);
or U28272 (N_28272,N_17482,N_18014);
nand U28273 (N_28273,N_15128,N_11394);
or U28274 (N_28274,N_11758,N_17751);
and U28275 (N_28275,N_17866,N_16356);
nand U28276 (N_28276,N_10233,N_10953);
or U28277 (N_28277,N_12734,N_18763);
or U28278 (N_28278,N_11710,N_14376);
xor U28279 (N_28279,N_15380,N_11434);
xor U28280 (N_28280,N_19973,N_16171);
nand U28281 (N_28281,N_12997,N_19228);
nand U28282 (N_28282,N_17572,N_18020);
or U28283 (N_28283,N_15841,N_10752);
or U28284 (N_28284,N_15057,N_16117);
nand U28285 (N_28285,N_12914,N_16453);
nand U28286 (N_28286,N_13660,N_14873);
or U28287 (N_28287,N_15524,N_16771);
and U28288 (N_28288,N_11770,N_12001);
nand U28289 (N_28289,N_15738,N_13893);
nand U28290 (N_28290,N_10283,N_16255);
nand U28291 (N_28291,N_13737,N_11253);
or U28292 (N_28292,N_16414,N_13452);
or U28293 (N_28293,N_10624,N_15219);
or U28294 (N_28294,N_16825,N_19248);
nand U28295 (N_28295,N_10761,N_16266);
or U28296 (N_28296,N_11819,N_19054);
and U28297 (N_28297,N_11426,N_16926);
or U28298 (N_28298,N_15744,N_13439);
nor U28299 (N_28299,N_13608,N_16427);
nand U28300 (N_28300,N_17074,N_10795);
nand U28301 (N_28301,N_13465,N_17996);
or U28302 (N_28302,N_14899,N_16678);
and U28303 (N_28303,N_10391,N_16376);
and U28304 (N_28304,N_10625,N_10574);
and U28305 (N_28305,N_13216,N_16600);
nand U28306 (N_28306,N_17139,N_14007);
nand U28307 (N_28307,N_17677,N_15229);
nand U28308 (N_28308,N_19734,N_19264);
and U28309 (N_28309,N_11532,N_15024);
or U28310 (N_28310,N_14017,N_16093);
or U28311 (N_28311,N_14641,N_17135);
and U28312 (N_28312,N_13016,N_10726);
nor U28313 (N_28313,N_18751,N_17371);
xnor U28314 (N_28314,N_12300,N_11322);
nand U28315 (N_28315,N_15542,N_16329);
nand U28316 (N_28316,N_12487,N_11430);
nor U28317 (N_28317,N_16095,N_19963);
nand U28318 (N_28318,N_16464,N_14844);
and U28319 (N_28319,N_12068,N_16558);
nor U28320 (N_28320,N_11912,N_15293);
nand U28321 (N_28321,N_13860,N_14979);
nor U28322 (N_28322,N_16260,N_17642);
and U28323 (N_28323,N_15172,N_14746);
xor U28324 (N_28324,N_18128,N_14560);
nor U28325 (N_28325,N_17529,N_17183);
and U28326 (N_28326,N_18027,N_13917);
xor U28327 (N_28327,N_15936,N_13251);
nand U28328 (N_28328,N_12904,N_11449);
nor U28329 (N_28329,N_14106,N_10691);
or U28330 (N_28330,N_10319,N_15318);
xnor U28331 (N_28331,N_18154,N_18582);
nor U28332 (N_28332,N_14792,N_18297);
or U28333 (N_28333,N_16028,N_17239);
or U28334 (N_28334,N_16628,N_19095);
nor U28335 (N_28335,N_11957,N_19555);
nand U28336 (N_28336,N_18662,N_15571);
nand U28337 (N_28337,N_12305,N_18726);
nand U28338 (N_28338,N_14957,N_10582);
nand U28339 (N_28339,N_12818,N_14254);
and U28340 (N_28340,N_17609,N_10384);
or U28341 (N_28341,N_17191,N_12941);
or U28342 (N_28342,N_19435,N_17987);
and U28343 (N_28343,N_16859,N_14585);
and U28344 (N_28344,N_14499,N_13954);
or U28345 (N_28345,N_11959,N_10720);
nor U28346 (N_28346,N_16618,N_14699);
and U28347 (N_28347,N_18379,N_10053);
or U28348 (N_28348,N_13985,N_19434);
or U28349 (N_28349,N_12528,N_10127);
xor U28350 (N_28350,N_16644,N_19973);
and U28351 (N_28351,N_16732,N_18710);
and U28352 (N_28352,N_12530,N_10634);
or U28353 (N_28353,N_10521,N_11450);
and U28354 (N_28354,N_17511,N_10267);
and U28355 (N_28355,N_11590,N_13640);
or U28356 (N_28356,N_17011,N_18291);
xor U28357 (N_28357,N_10107,N_18750);
and U28358 (N_28358,N_11522,N_12213);
nand U28359 (N_28359,N_15942,N_18482);
and U28360 (N_28360,N_16816,N_13527);
nand U28361 (N_28361,N_17690,N_10106);
or U28362 (N_28362,N_19390,N_16432);
or U28363 (N_28363,N_14621,N_14436);
or U28364 (N_28364,N_18460,N_14406);
nor U28365 (N_28365,N_13177,N_12649);
nand U28366 (N_28366,N_12296,N_14704);
or U28367 (N_28367,N_10964,N_10397);
and U28368 (N_28368,N_18833,N_12554);
or U28369 (N_28369,N_13739,N_12715);
and U28370 (N_28370,N_10222,N_17153);
nand U28371 (N_28371,N_17958,N_17407);
nand U28372 (N_28372,N_12385,N_13988);
and U28373 (N_28373,N_16443,N_17815);
nand U28374 (N_28374,N_10261,N_10596);
nor U28375 (N_28375,N_14141,N_15375);
xnor U28376 (N_28376,N_12679,N_16432);
or U28377 (N_28377,N_17646,N_15327);
or U28378 (N_28378,N_19238,N_13852);
or U28379 (N_28379,N_13377,N_16823);
nor U28380 (N_28380,N_15146,N_10171);
nor U28381 (N_28381,N_12403,N_18933);
xnor U28382 (N_28382,N_15909,N_19229);
nor U28383 (N_28383,N_13898,N_19449);
nor U28384 (N_28384,N_18030,N_13315);
or U28385 (N_28385,N_10708,N_18090);
or U28386 (N_28386,N_18852,N_15685);
or U28387 (N_28387,N_17057,N_11516);
xor U28388 (N_28388,N_16253,N_15031);
nor U28389 (N_28389,N_19315,N_11583);
nand U28390 (N_28390,N_18940,N_14472);
nor U28391 (N_28391,N_10687,N_18795);
nand U28392 (N_28392,N_17481,N_18642);
and U28393 (N_28393,N_17434,N_17850);
nand U28394 (N_28394,N_11399,N_11226);
and U28395 (N_28395,N_17681,N_15299);
nand U28396 (N_28396,N_19166,N_15918);
nand U28397 (N_28397,N_15549,N_16717);
nand U28398 (N_28398,N_12001,N_11479);
nand U28399 (N_28399,N_17858,N_14747);
or U28400 (N_28400,N_12495,N_19632);
xor U28401 (N_28401,N_18689,N_15611);
or U28402 (N_28402,N_12411,N_18986);
and U28403 (N_28403,N_15679,N_15408);
nand U28404 (N_28404,N_12173,N_19150);
xor U28405 (N_28405,N_17634,N_15632);
or U28406 (N_28406,N_10580,N_12108);
nor U28407 (N_28407,N_16584,N_17378);
and U28408 (N_28408,N_13375,N_11954);
nor U28409 (N_28409,N_10594,N_14979);
and U28410 (N_28410,N_12919,N_11432);
nand U28411 (N_28411,N_14589,N_18937);
nor U28412 (N_28412,N_10605,N_17030);
and U28413 (N_28413,N_15195,N_17651);
nor U28414 (N_28414,N_10481,N_10561);
nand U28415 (N_28415,N_12386,N_11025);
and U28416 (N_28416,N_10215,N_10786);
xor U28417 (N_28417,N_18578,N_18394);
and U28418 (N_28418,N_10098,N_10600);
nor U28419 (N_28419,N_11944,N_18948);
nor U28420 (N_28420,N_19160,N_14152);
nand U28421 (N_28421,N_16436,N_16231);
or U28422 (N_28422,N_10103,N_14654);
nor U28423 (N_28423,N_11469,N_19329);
nor U28424 (N_28424,N_17560,N_13600);
nand U28425 (N_28425,N_18450,N_11829);
nor U28426 (N_28426,N_12440,N_14919);
xor U28427 (N_28427,N_19543,N_19378);
nor U28428 (N_28428,N_10650,N_19499);
and U28429 (N_28429,N_17470,N_14774);
nor U28430 (N_28430,N_11734,N_12568);
nand U28431 (N_28431,N_11301,N_13132);
nand U28432 (N_28432,N_11046,N_12799);
nor U28433 (N_28433,N_13382,N_19835);
nor U28434 (N_28434,N_13509,N_16717);
and U28435 (N_28435,N_14032,N_10605);
and U28436 (N_28436,N_18391,N_17373);
nor U28437 (N_28437,N_16258,N_14174);
xnor U28438 (N_28438,N_16668,N_17118);
nand U28439 (N_28439,N_14242,N_11002);
xor U28440 (N_28440,N_17515,N_19427);
or U28441 (N_28441,N_12313,N_16811);
or U28442 (N_28442,N_12809,N_10453);
or U28443 (N_28443,N_17639,N_19896);
nor U28444 (N_28444,N_14690,N_19440);
nand U28445 (N_28445,N_18777,N_10797);
and U28446 (N_28446,N_15225,N_16798);
or U28447 (N_28447,N_13979,N_14374);
nand U28448 (N_28448,N_10554,N_10895);
or U28449 (N_28449,N_15768,N_10065);
or U28450 (N_28450,N_13971,N_14155);
or U28451 (N_28451,N_12145,N_10062);
nand U28452 (N_28452,N_12196,N_15521);
or U28453 (N_28453,N_16841,N_16203);
nor U28454 (N_28454,N_15347,N_19657);
and U28455 (N_28455,N_10503,N_19434);
or U28456 (N_28456,N_19215,N_14546);
or U28457 (N_28457,N_11009,N_12706);
or U28458 (N_28458,N_19147,N_19291);
nand U28459 (N_28459,N_14184,N_18558);
or U28460 (N_28460,N_19078,N_15518);
xor U28461 (N_28461,N_15582,N_10245);
nand U28462 (N_28462,N_11717,N_19519);
and U28463 (N_28463,N_13522,N_12511);
or U28464 (N_28464,N_10033,N_17700);
nor U28465 (N_28465,N_11779,N_18660);
nand U28466 (N_28466,N_10236,N_15761);
nor U28467 (N_28467,N_19618,N_17770);
nand U28468 (N_28468,N_11818,N_18148);
nand U28469 (N_28469,N_18108,N_16476);
xor U28470 (N_28470,N_12922,N_15915);
and U28471 (N_28471,N_12701,N_13401);
and U28472 (N_28472,N_13408,N_14647);
nand U28473 (N_28473,N_11099,N_17991);
nor U28474 (N_28474,N_10136,N_14270);
or U28475 (N_28475,N_10634,N_16454);
or U28476 (N_28476,N_18480,N_16722);
and U28477 (N_28477,N_18531,N_15554);
nand U28478 (N_28478,N_18220,N_16009);
and U28479 (N_28479,N_13925,N_19149);
nand U28480 (N_28480,N_11016,N_19372);
nand U28481 (N_28481,N_17823,N_11568);
nand U28482 (N_28482,N_12315,N_13616);
nor U28483 (N_28483,N_13765,N_10518);
or U28484 (N_28484,N_17030,N_11294);
nand U28485 (N_28485,N_17315,N_18317);
nand U28486 (N_28486,N_17822,N_12634);
and U28487 (N_28487,N_11189,N_16716);
and U28488 (N_28488,N_11247,N_17909);
and U28489 (N_28489,N_12019,N_12678);
or U28490 (N_28490,N_11346,N_11033);
or U28491 (N_28491,N_12623,N_10211);
nand U28492 (N_28492,N_12512,N_17631);
or U28493 (N_28493,N_16982,N_17452);
and U28494 (N_28494,N_19193,N_14078);
nand U28495 (N_28495,N_10239,N_18933);
nand U28496 (N_28496,N_11958,N_16539);
nor U28497 (N_28497,N_15848,N_14027);
nor U28498 (N_28498,N_14352,N_15357);
or U28499 (N_28499,N_12850,N_19508);
nor U28500 (N_28500,N_10795,N_17899);
or U28501 (N_28501,N_15201,N_19681);
nand U28502 (N_28502,N_12806,N_10196);
xnor U28503 (N_28503,N_12565,N_12495);
nand U28504 (N_28504,N_14577,N_12992);
xor U28505 (N_28505,N_11279,N_10379);
nor U28506 (N_28506,N_19206,N_18112);
nor U28507 (N_28507,N_11605,N_10982);
and U28508 (N_28508,N_17317,N_13164);
and U28509 (N_28509,N_19113,N_11256);
nand U28510 (N_28510,N_16460,N_11177);
nor U28511 (N_28511,N_19807,N_19406);
or U28512 (N_28512,N_13902,N_16483);
or U28513 (N_28513,N_15209,N_16966);
or U28514 (N_28514,N_12708,N_19301);
nor U28515 (N_28515,N_18107,N_11193);
or U28516 (N_28516,N_15266,N_19968);
and U28517 (N_28517,N_14296,N_19343);
nor U28518 (N_28518,N_18092,N_12610);
or U28519 (N_28519,N_15119,N_12265);
nor U28520 (N_28520,N_10550,N_14394);
and U28521 (N_28521,N_17417,N_16086);
xnor U28522 (N_28522,N_10653,N_16787);
xnor U28523 (N_28523,N_11597,N_16693);
nand U28524 (N_28524,N_11334,N_14552);
and U28525 (N_28525,N_19641,N_15125);
nor U28526 (N_28526,N_10652,N_19610);
and U28527 (N_28527,N_11770,N_12979);
or U28528 (N_28528,N_19593,N_11419);
nor U28529 (N_28529,N_18278,N_16375);
and U28530 (N_28530,N_14205,N_19889);
and U28531 (N_28531,N_11418,N_12088);
xor U28532 (N_28532,N_10411,N_18869);
nand U28533 (N_28533,N_12552,N_15675);
and U28534 (N_28534,N_16354,N_17018);
xor U28535 (N_28535,N_16578,N_17953);
nand U28536 (N_28536,N_12328,N_15898);
nand U28537 (N_28537,N_11763,N_11316);
nor U28538 (N_28538,N_15679,N_16349);
nand U28539 (N_28539,N_18780,N_11969);
nor U28540 (N_28540,N_10579,N_15788);
nor U28541 (N_28541,N_11202,N_11401);
or U28542 (N_28542,N_12057,N_12490);
nand U28543 (N_28543,N_17310,N_17182);
nand U28544 (N_28544,N_15781,N_16536);
or U28545 (N_28545,N_13139,N_15132);
nor U28546 (N_28546,N_13627,N_14238);
and U28547 (N_28547,N_10777,N_11631);
xnor U28548 (N_28548,N_19687,N_16360);
xnor U28549 (N_28549,N_16381,N_15756);
nand U28550 (N_28550,N_13927,N_17696);
nand U28551 (N_28551,N_13927,N_11807);
nor U28552 (N_28552,N_16834,N_19126);
or U28553 (N_28553,N_10992,N_16075);
or U28554 (N_28554,N_17888,N_17554);
and U28555 (N_28555,N_18256,N_11878);
or U28556 (N_28556,N_15431,N_19273);
xnor U28557 (N_28557,N_10798,N_18165);
nand U28558 (N_28558,N_19298,N_14951);
xor U28559 (N_28559,N_12537,N_13208);
nor U28560 (N_28560,N_13198,N_19640);
or U28561 (N_28561,N_12789,N_16954);
and U28562 (N_28562,N_15378,N_10487);
nor U28563 (N_28563,N_19838,N_10116);
xor U28564 (N_28564,N_19571,N_16852);
nor U28565 (N_28565,N_16155,N_10815);
nand U28566 (N_28566,N_12537,N_15117);
nand U28567 (N_28567,N_17211,N_19041);
and U28568 (N_28568,N_17626,N_16361);
nor U28569 (N_28569,N_12828,N_18552);
or U28570 (N_28570,N_19443,N_13969);
nand U28571 (N_28571,N_14201,N_11612);
and U28572 (N_28572,N_11949,N_10438);
or U28573 (N_28573,N_16544,N_13676);
and U28574 (N_28574,N_10626,N_17263);
and U28575 (N_28575,N_19032,N_12613);
nor U28576 (N_28576,N_11512,N_18517);
and U28577 (N_28577,N_16693,N_18162);
or U28578 (N_28578,N_17988,N_16656);
nor U28579 (N_28579,N_13819,N_17561);
nand U28580 (N_28580,N_13803,N_13173);
xor U28581 (N_28581,N_14846,N_14394);
nor U28582 (N_28582,N_17252,N_11516);
nand U28583 (N_28583,N_10472,N_17967);
and U28584 (N_28584,N_11496,N_16632);
or U28585 (N_28585,N_18653,N_16760);
and U28586 (N_28586,N_10527,N_18183);
nor U28587 (N_28587,N_16969,N_14928);
or U28588 (N_28588,N_18458,N_15733);
xor U28589 (N_28589,N_15293,N_13100);
xnor U28590 (N_28590,N_11970,N_12070);
nand U28591 (N_28591,N_10078,N_16404);
nand U28592 (N_28592,N_17811,N_13802);
and U28593 (N_28593,N_16266,N_18052);
and U28594 (N_28594,N_18462,N_17781);
nand U28595 (N_28595,N_15273,N_13806);
nor U28596 (N_28596,N_12796,N_18080);
or U28597 (N_28597,N_19281,N_11662);
nand U28598 (N_28598,N_17486,N_17324);
nand U28599 (N_28599,N_10616,N_11156);
or U28600 (N_28600,N_10690,N_17498);
nor U28601 (N_28601,N_18848,N_15259);
nor U28602 (N_28602,N_16183,N_14265);
nor U28603 (N_28603,N_19435,N_19327);
nor U28604 (N_28604,N_13581,N_18649);
nor U28605 (N_28605,N_17132,N_18657);
or U28606 (N_28606,N_10666,N_15238);
and U28607 (N_28607,N_11092,N_19846);
or U28608 (N_28608,N_11276,N_11507);
nand U28609 (N_28609,N_11961,N_19280);
xor U28610 (N_28610,N_13008,N_19236);
nor U28611 (N_28611,N_19830,N_14545);
nor U28612 (N_28612,N_18353,N_18773);
nor U28613 (N_28613,N_19732,N_13645);
nand U28614 (N_28614,N_18295,N_13015);
nand U28615 (N_28615,N_15366,N_12772);
nand U28616 (N_28616,N_11542,N_16729);
nor U28617 (N_28617,N_10251,N_10809);
and U28618 (N_28618,N_15288,N_15421);
and U28619 (N_28619,N_16507,N_19743);
and U28620 (N_28620,N_13329,N_10139);
or U28621 (N_28621,N_12879,N_10605);
nor U28622 (N_28622,N_18916,N_15414);
nand U28623 (N_28623,N_11252,N_15304);
xor U28624 (N_28624,N_11612,N_19986);
and U28625 (N_28625,N_12334,N_17853);
nor U28626 (N_28626,N_11063,N_17955);
nand U28627 (N_28627,N_12397,N_11275);
or U28628 (N_28628,N_11885,N_19854);
or U28629 (N_28629,N_18336,N_14026);
or U28630 (N_28630,N_13239,N_19657);
and U28631 (N_28631,N_12965,N_12803);
nor U28632 (N_28632,N_10607,N_17297);
nand U28633 (N_28633,N_10086,N_15552);
and U28634 (N_28634,N_12488,N_14204);
or U28635 (N_28635,N_14443,N_15504);
or U28636 (N_28636,N_14562,N_17746);
and U28637 (N_28637,N_12167,N_13140);
nor U28638 (N_28638,N_19287,N_11769);
nand U28639 (N_28639,N_18210,N_12258);
nand U28640 (N_28640,N_17417,N_13458);
or U28641 (N_28641,N_11088,N_19042);
and U28642 (N_28642,N_17334,N_13296);
nor U28643 (N_28643,N_16400,N_13775);
xnor U28644 (N_28644,N_13387,N_18605);
or U28645 (N_28645,N_13315,N_17105);
nor U28646 (N_28646,N_17195,N_19075);
nand U28647 (N_28647,N_17797,N_19497);
nor U28648 (N_28648,N_13932,N_12934);
nor U28649 (N_28649,N_14376,N_15596);
and U28650 (N_28650,N_16591,N_17568);
or U28651 (N_28651,N_19396,N_19630);
and U28652 (N_28652,N_19847,N_11734);
and U28653 (N_28653,N_19140,N_18488);
nor U28654 (N_28654,N_15636,N_11673);
and U28655 (N_28655,N_16419,N_13366);
and U28656 (N_28656,N_16145,N_11649);
and U28657 (N_28657,N_12634,N_18833);
or U28658 (N_28658,N_13999,N_18060);
nand U28659 (N_28659,N_16821,N_19307);
nand U28660 (N_28660,N_12779,N_19930);
and U28661 (N_28661,N_14184,N_10334);
nor U28662 (N_28662,N_11479,N_11456);
nand U28663 (N_28663,N_15987,N_16900);
and U28664 (N_28664,N_18203,N_10349);
nand U28665 (N_28665,N_15856,N_10743);
xnor U28666 (N_28666,N_11952,N_12584);
and U28667 (N_28667,N_13564,N_16907);
and U28668 (N_28668,N_18713,N_14777);
or U28669 (N_28669,N_18646,N_19872);
nor U28670 (N_28670,N_16998,N_17466);
or U28671 (N_28671,N_17307,N_18951);
nor U28672 (N_28672,N_11837,N_17005);
or U28673 (N_28673,N_16155,N_15236);
xor U28674 (N_28674,N_14318,N_16390);
xor U28675 (N_28675,N_14613,N_19629);
and U28676 (N_28676,N_11618,N_12390);
nor U28677 (N_28677,N_10601,N_13688);
nor U28678 (N_28678,N_10764,N_17293);
or U28679 (N_28679,N_13294,N_17795);
or U28680 (N_28680,N_16869,N_18452);
nand U28681 (N_28681,N_10317,N_10729);
nor U28682 (N_28682,N_12484,N_12301);
or U28683 (N_28683,N_16818,N_14967);
and U28684 (N_28684,N_13420,N_17585);
or U28685 (N_28685,N_14082,N_11244);
and U28686 (N_28686,N_15945,N_15804);
or U28687 (N_28687,N_14657,N_16854);
nor U28688 (N_28688,N_17668,N_17098);
nor U28689 (N_28689,N_12706,N_14458);
nand U28690 (N_28690,N_11053,N_14551);
and U28691 (N_28691,N_18818,N_13256);
nand U28692 (N_28692,N_15213,N_12267);
nor U28693 (N_28693,N_15884,N_14287);
nand U28694 (N_28694,N_15362,N_12679);
nor U28695 (N_28695,N_13473,N_13078);
or U28696 (N_28696,N_11035,N_19416);
or U28697 (N_28697,N_13011,N_16012);
and U28698 (N_28698,N_15939,N_13829);
nand U28699 (N_28699,N_15742,N_14860);
or U28700 (N_28700,N_17699,N_12624);
nor U28701 (N_28701,N_15564,N_17730);
nand U28702 (N_28702,N_18422,N_19809);
nor U28703 (N_28703,N_10214,N_16181);
and U28704 (N_28704,N_17416,N_17365);
or U28705 (N_28705,N_16744,N_19071);
nor U28706 (N_28706,N_10938,N_17219);
nor U28707 (N_28707,N_11513,N_19196);
nor U28708 (N_28708,N_17059,N_16477);
nor U28709 (N_28709,N_19458,N_17525);
nand U28710 (N_28710,N_13741,N_14101);
xor U28711 (N_28711,N_18423,N_18447);
nor U28712 (N_28712,N_13547,N_19008);
nand U28713 (N_28713,N_15476,N_10711);
and U28714 (N_28714,N_10410,N_12101);
nor U28715 (N_28715,N_14299,N_19753);
xnor U28716 (N_28716,N_19336,N_10236);
nor U28717 (N_28717,N_11991,N_17095);
nor U28718 (N_28718,N_17042,N_11494);
or U28719 (N_28719,N_12715,N_16757);
or U28720 (N_28720,N_17458,N_15346);
nand U28721 (N_28721,N_17210,N_10422);
and U28722 (N_28722,N_12460,N_10486);
or U28723 (N_28723,N_14194,N_18501);
nor U28724 (N_28724,N_18454,N_13270);
nand U28725 (N_28725,N_11390,N_19834);
xor U28726 (N_28726,N_17753,N_12686);
nand U28727 (N_28727,N_13056,N_13378);
nand U28728 (N_28728,N_14596,N_19342);
nand U28729 (N_28729,N_12426,N_14807);
nand U28730 (N_28730,N_10833,N_16513);
nor U28731 (N_28731,N_17263,N_19416);
xor U28732 (N_28732,N_13025,N_14921);
nand U28733 (N_28733,N_19013,N_19899);
and U28734 (N_28734,N_12304,N_15489);
nand U28735 (N_28735,N_12715,N_17764);
or U28736 (N_28736,N_12745,N_19836);
nand U28737 (N_28737,N_10441,N_10698);
and U28738 (N_28738,N_19473,N_10975);
nor U28739 (N_28739,N_17885,N_12460);
nor U28740 (N_28740,N_15476,N_10251);
nor U28741 (N_28741,N_12829,N_14771);
nand U28742 (N_28742,N_15490,N_14264);
xnor U28743 (N_28743,N_13137,N_19586);
nor U28744 (N_28744,N_14113,N_18576);
or U28745 (N_28745,N_11286,N_10610);
nand U28746 (N_28746,N_13608,N_15846);
nand U28747 (N_28747,N_16923,N_11170);
or U28748 (N_28748,N_15846,N_15461);
or U28749 (N_28749,N_17055,N_16113);
nand U28750 (N_28750,N_17415,N_18931);
nand U28751 (N_28751,N_17695,N_19943);
or U28752 (N_28752,N_13784,N_11809);
and U28753 (N_28753,N_19852,N_18638);
xnor U28754 (N_28754,N_15224,N_13046);
xor U28755 (N_28755,N_17799,N_18349);
or U28756 (N_28756,N_13648,N_11485);
or U28757 (N_28757,N_12789,N_15383);
or U28758 (N_28758,N_17401,N_15621);
xnor U28759 (N_28759,N_13712,N_10703);
nor U28760 (N_28760,N_14033,N_11710);
or U28761 (N_28761,N_19807,N_14530);
and U28762 (N_28762,N_17988,N_19637);
and U28763 (N_28763,N_19728,N_14220);
and U28764 (N_28764,N_19490,N_18963);
or U28765 (N_28765,N_16640,N_12555);
and U28766 (N_28766,N_12219,N_15714);
nor U28767 (N_28767,N_18442,N_11278);
nor U28768 (N_28768,N_14233,N_14608);
nand U28769 (N_28769,N_11065,N_17325);
or U28770 (N_28770,N_17675,N_12417);
nor U28771 (N_28771,N_13858,N_15018);
and U28772 (N_28772,N_15689,N_16423);
or U28773 (N_28773,N_12541,N_19152);
or U28774 (N_28774,N_16518,N_17930);
nand U28775 (N_28775,N_13504,N_17568);
or U28776 (N_28776,N_19973,N_14144);
nand U28777 (N_28777,N_14773,N_11275);
nor U28778 (N_28778,N_15535,N_11399);
and U28779 (N_28779,N_12244,N_14997);
nand U28780 (N_28780,N_17652,N_19985);
nand U28781 (N_28781,N_11033,N_11994);
nand U28782 (N_28782,N_15105,N_14339);
and U28783 (N_28783,N_10718,N_15600);
nor U28784 (N_28784,N_11340,N_11854);
or U28785 (N_28785,N_17177,N_17985);
or U28786 (N_28786,N_12632,N_14960);
nor U28787 (N_28787,N_19389,N_11632);
nand U28788 (N_28788,N_19720,N_18308);
and U28789 (N_28789,N_12820,N_15687);
nand U28790 (N_28790,N_14714,N_17200);
nand U28791 (N_28791,N_12308,N_19045);
or U28792 (N_28792,N_10189,N_17473);
xnor U28793 (N_28793,N_19351,N_14490);
nand U28794 (N_28794,N_11556,N_13951);
xnor U28795 (N_28795,N_13810,N_13256);
or U28796 (N_28796,N_18046,N_17215);
nor U28797 (N_28797,N_13348,N_15507);
and U28798 (N_28798,N_17396,N_16798);
nand U28799 (N_28799,N_11144,N_14469);
or U28800 (N_28800,N_19553,N_16891);
xnor U28801 (N_28801,N_19812,N_12879);
nand U28802 (N_28802,N_15726,N_12878);
or U28803 (N_28803,N_10300,N_19006);
or U28804 (N_28804,N_18095,N_19717);
nor U28805 (N_28805,N_14301,N_13104);
nand U28806 (N_28806,N_17779,N_14988);
nor U28807 (N_28807,N_17365,N_19299);
and U28808 (N_28808,N_11425,N_13192);
nand U28809 (N_28809,N_11538,N_14435);
nor U28810 (N_28810,N_12392,N_14668);
and U28811 (N_28811,N_12056,N_14205);
nor U28812 (N_28812,N_19988,N_13674);
or U28813 (N_28813,N_19459,N_17503);
nor U28814 (N_28814,N_14170,N_15461);
nand U28815 (N_28815,N_18507,N_16160);
or U28816 (N_28816,N_17140,N_10207);
or U28817 (N_28817,N_18898,N_19810);
nand U28818 (N_28818,N_15311,N_10192);
nand U28819 (N_28819,N_12943,N_18504);
xor U28820 (N_28820,N_17056,N_14271);
nand U28821 (N_28821,N_12833,N_19052);
nor U28822 (N_28822,N_13235,N_14061);
or U28823 (N_28823,N_12811,N_11223);
xnor U28824 (N_28824,N_12218,N_12506);
or U28825 (N_28825,N_19432,N_18225);
or U28826 (N_28826,N_19431,N_11733);
nand U28827 (N_28827,N_13869,N_15450);
nand U28828 (N_28828,N_18972,N_15107);
and U28829 (N_28829,N_19068,N_15475);
or U28830 (N_28830,N_15245,N_11076);
nand U28831 (N_28831,N_18773,N_18100);
or U28832 (N_28832,N_11253,N_19297);
and U28833 (N_28833,N_12372,N_10335);
nand U28834 (N_28834,N_15712,N_16989);
and U28835 (N_28835,N_11911,N_13565);
nand U28836 (N_28836,N_14337,N_10407);
or U28837 (N_28837,N_18527,N_19723);
nand U28838 (N_28838,N_18331,N_13606);
nand U28839 (N_28839,N_17408,N_11669);
or U28840 (N_28840,N_10136,N_10714);
nand U28841 (N_28841,N_13995,N_11405);
xor U28842 (N_28842,N_12783,N_13303);
and U28843 (N_28843,N_18262,N_15194);
or U28844 (N_28844,N_13146,N_10879);
or U28845 (N_28845,N_16303,N_11346);
nand U28846 (N_28846,N_17079,N_10278);
or U28847 (N_28847,N_13894,N_14946);
nand U28848 (N_28848,N_18579,N_17339);
nand U28849 (N_28849,N_19796,N_19634);
nand U28850 (N_28850,N_14974,N_15048);
xor U28851 (N_28851,N_14371,N_16475);
or U28852 (N_28852,N_15205,N_17784);
nor U28853 (N_28853,N_12417,N_18431);
nor U28854 (N_28854,N_14725,N_13803);
nand U28855 (N_28855,N_17681,N_11552);
and U28856 (N_28856,N_18936,N_17291);
nor U28857 (N_28857,N_14320,N_13993);
nand U28858 (N_28858,N_13500,N_14500);
xor U28859 (N_28859,N_11290,N_14686);
xor U28860 (N_28860,N_18304,N_16048);
nand U28861 (N_28861,N_19640,N_16278);
nand U28862 (N_28862,N_10404,N_14446);
xnor U28863 (N_28863,N_14663,N_12872);
nand U28864 (N_28864,N_19135,N_11513);
nand U28865 (N_28865,N_15898,N_19338);
or U28866 (N_28866,N_12031,N_11732);
nor U28867 (N_28867,N_15389,N_18657);
nand U28868 (N_28868,N_18089,N_10619);
nand U28869 (N_28869,N_17145,N_13869);
nand U28870 (N_28870,N_15283,N_18109);
or U28871 (N_28871,N_19500,N_13461);
nor U28872 (N_28872,N_14784,N_10696);
xnor U28873 (N_28873,N_18832,N_17331);
nand U28874 (N_28874,N_16201,N_13289);
and U28875 (N_28875,N_12118,N_18513);
and U28876 (N_28876,N_12342,N_16463);
or U28877 (N_28877,N_16733,N_13259);
nor U28878 (N_28878,N_15480,N_18870);
nand U28879 (N_28879,N_19240,N_10511);
nor U28880 (N_28880,N_13381,N_11925);
and U28881 (N_28881,N_17368,N_10452);
and U28882 (N_28882,N_16265,N_15304);
or U28883 (N_28883,N_15723,N_15847);
nor U28884 (N_28884,N_10430,N_13392);
or U28885 (N_28885,N_19142,N_18538);
nor U28886 (N_28886,N_12223,N_15763);
or U28887 (N_28887,N_18167,N_13882);
nor U28888 (N_28888,N_19254,N_12316);
xor U28889 (N_28889,N_15172,N_11683);
nor U28890 (N_28890,N_18260,N_10563);
xnor U28891 (N_28891,N_11059,N_12141);
nand U28892 (N_28892,N_18057,N_16230);
or U28893 (N_28893,N_15798,N_16709);
nor U28894 (N_28894,N_11043,N_10609);
nand U28895 (N_28895,N_11640,N_10074);
nor U28896 (N_28896,N_19785,N_10811);
and U28897 (N_28897,N_16496,N_12524);
or U28898 (N_28898,N_12169,N_19175);
nand U28899 (N_28899,N_15909,N_12450);
nor U28900 (N_28900,N_17175,N_14493);
nor U28901 (N_28901,N_19931,N_18634);
nor U28902 (N_28902,N_14071,N_10158);
xnor U28903 (N_28903,N_19149,N_11209);
nand U28904 (N_28904,N_15717,N_14946);
and U28905 (N_28905,N_16935,N_17966);
nand U28906 (N_28906,N_13398,N_13845);
nand U28907 (N_28907,N_15684,N_16193);
and U28908 (N_28908,N_10569,N_10224);
or U28909 (N_28909,N_13703,N_19716);
and U28910 (N_28910,N_15400,N_12945);
nor U28911 (N_28911,N_10492,N_15487);
and U28912 (N_28912,N_10913,N_14465);
and U28913 (N_28913,N_13926,N_18421);
nand U28914 (N_28914,N_16037,N_11656);
or U28915 (N_28915,N_17925,N_10435);
and U28916 (N_28916,N_17459,N_11090);
and U28917 (N_28917,N_15260,N_17770);
nand U28918 (N_28918,N_17542,N_14794);
or U28919 (N_28919,N_17036,N_19520);
nand U28920 (N_28920,N_15237,N_16754);
nand U28921 (N_28921,N_19346,N_16570);
xnor U28922 (N_28922,N_14669,N_12558);
nor U28923 (N_28923,N_10381,N_15001);
xor U28924 (N_28924,N_10617,N_14907);
xnor U28925 (N_28925,N_14712,N_13671);
nor U28926 (N_28926,N_12714,N_16829);
nor U28927 (N_28927,N_14840,N_16053);
and U28928 (N_28928,N_17025,N_19564);
and U28929 (N_28929,N_11196,N_18660);
nor U28930 (N_28930,N_10517,N_12897);
nor U28931 (N_28931,N_10309,N_19040);
nor U28932 (N_28932,N_12893,N_19095);
nor U28933 (N_28933,N_19847,N_15397);
and U28934 (N_28934,N_14659,N_12585);
xnor U28935 (N_28935,N_10861,N_14901);
or U28936 (N_28936,N_12790,N_18857);
and U28937 (N_28937,N_16741,N_19623);
nand U28938 (N_28938,N_15581,N_14271);
nand U28939 (N_28939,N_11218,N_12393);
and U28940 (N_28940,N_12476,N_11017);
xnor U28941 (N_28941,N_18184,N_12827);
xor U28942 (N_28942,N_13848,N_13329);
and U28943 (N_28943,N_16050,N_15205);
or U28944 (N_28944,N_13026,N_11547);
and U28945 (N_28945,N_10404,N_13489);
or U28946 (N_28946,N_12153,N_13318);
nand U28947 (N_28947,N_19377,N_16417);
or U28948 (N_28948,N_10185,N_12410);
nor U28949 (N_28949,N_13273,N_12337);
nand U28950 (N_28950,N_11036,N_13711);
nor U28951 (N_28951,N_19891,N_18197);
nand U28952 (N_28952,N_14445,N_12040);
xnor U28953 (N_28953,N_11569,N_19734);
nand U28954 (N_28954,N_13227,N_14200);
nand U28955 (N_28955,N_10649,N_19714);
nand U28956 (N_28956,N_15830,N_11455);
nand U28957 (N_28957,N_10288,N_17783);
nor U28958 (N_28958,N_13777,N_16094);
nor U28959 (N_28959,N_12197,N_13661);
or U28960 (N_28960,N_10434,N_18670);
xnor U28961 (N_28961,N_17334,N_10380);
nor U28962 (N_28962,N_15992,N_13039);
nor U28963 (N_28963,N_18691,N_13052);
and U28964 (N_28964,N_19239,N_10556);
nand U28965 (N_28965,N_15138,N_13244);
and U28966 (N_28966,N_12181,N_12309);
nand U28967 (N_28967,N_16676,N_17225);
nor U28968 (N_28968,N_15503,N_14449);
nand U28969 (N_28969,N_10985,N_18899);
and U28970 (N_28970,N_12552,N_12931);
or U28971 (N_28971,N_12396,N_19404);
nor U28972 (N_28972,N_16430,N_16598);
or U28973 (N_28973,N_12364,N_18423);
and U28974 (N_28974,N_19686,N_15192);
or U28975 (N_28975,N_12130,N_17827);
or U28976 (N_28976,N_13190,N_13571);
or U28977 (N_28977,N_13827,N_19177);
and U28978 (N_28978,N_17235,N_14569);
nor U28979 (N_28979,N_18693,N_12570);
nor U28980 (N_28980,N_14312,N_15152);
nand U28981 (N_28981,N_17382,N_12209);
nor U28982 (N_28982,N_15988,N_18393);
nand U28983 (N_28983,N_15112,N_11140);
xor U28984 (N_28984,N_11537,N_11626);
or U28985 (N_28985,N_15355,N_10764);
and U28986 (N_28986,N_17889,N_18568);
or U28987 (N_28987,N_12689,N_16854);
or U28988 (N_28988,N_15980,N_18028);
and U28989 (N_28989,N_17358,N_18723);
and U28990 (N_28990,N_18799,N_14180);
nor U28991 (N_28991,N_15445,N_14462);
or U28992 (N_28992,N_16962,N_15286);
nor U28993 (N_28993,N_13238,N_19494);
nor U28994 (N_28994,N_14026,N_12768);
nor U28995 (N_28995,N_15086,N_16294);
or U28996 (N_28996,N_19396,N_13092);
and U28997 (N_28997,N_17948,N_12490);
and U28998 (N_28998,N_15578,N_12269);
nor U28999 (N_28999,N_14777,N_15426);
nand U29000 (N_29000,N_10092,N_14245);
and U29001 (N_29001,N_15485,N_19732);
or U29002 (N_29002,N_11935,N_18347);
xor U29003 (N_29003,N_17628,N_18806);
or U29004 (N_29004,N_15390,N_10605);
nor U29005 (N_29005,N_19016,N_13308);
nor U29006 (N_29006,N_18352,N_18576);
or U29007 (N_29007,N_19545,N_17421);
nor U29008 (N_29008,N_15833,N_14729);
nand U29009 (N_29009,N_14968,N_10169);
xor U29010 (N_29010,N_17333,N_18923);
and U29011 (N_29011,N_16370,N_18844);
nand U29012 (N_29012,N_15576,N_15389);
nand U29013 (N_29013,N_14920,N_11692);
or U29014 (N_29014,N_13037,N_18176);
nor U29015 (N_29015,N_11511,N_13319);
or U29016 (N_29016,N_18730,N_16884);
or U29017 (N_29017,N_10032,N_15538);
nand U29018 (N_29018,N_19421,N_17810);
and U29019 (N_29019,N_19009,N_19029);
nor U29020 (N_29020,N_16137,N_10287);
and U29021 (N_29021,N_14298,N_12807);
or U29022 (N_29022,N_14949,N_18180);
and U29023 (N_29023,N_17587,N_12112);
nor U29024 (N_29024,N_18655,N_15641);
xnor U29025 (N_29025,N_17725,N_18229);
or U29026 (N_29026,N_11827,N_17863);
or U29027 (N_29027,N_10861,N_17913);
nand U29028 (N_29028,N_12690,N_13263);
nor U29029 (N_29029,N_10846,N_10189);
nand U29030 (N_29030,N_14252,N_15103);
nor U29031 (N_29031,N_15617,N_11752);
and U29032 (N_29032,N_11687,N_10201);
and U29033 (N_29033,N_16375,N_15951);
or U29034 (N_29034,N_13501,N_11557);
and U29035 (N_29035,N_10492,N_13445);
nor U29036 (N_29036,N_11157,N_11943);
nor U29037 (N_29037,N_12217,N_19703);
nor U29038 (N_29038,N_19342,N_16409);
or U29039 (N_29039,N_16940,N_16161);
or U29040 (N_29040,N_11085,N_14872);
nand U29041 (N_29041,N_14012,N_13240);
and U29042 (N_29042,N_13222,N_14555);
or U29043 (N_29043,N_19113,N_16750);
and U29044 (N_29044,N_12480,N_18383);
xnor U29045 (N_29045,N_12716,N_16222);
or U29046 (N_29046,N_11397,N_17549);
and U29047 (N_29047,N_10620,N_11549);
and U29048 (N_29048,N_11518,N_10516);
nor U29049 (N_29049,N_18144,N_18798);
or U29050 (N_29050,N_14739,N_17356);
or U29051 (N_29051,N_19748,N_12229);
or U29052 (N_29052,N_11834,N_13394);
nor U29053 (N_29053,N_15148,N_15257);
nand U29054 (N_29054,N_18276,N_13190);
or U29055 (N_29055,N_12260,N_11636);
nor U29056 (N_29056,N_12737,N_15680);
or U29057 (N_29057,N_18543,N_12284);
or U29058 (N_29058,N_16744,N_15780);
xnor U29059 (N_29059,N_10075,N_16574);
and U29060 (N_29060,N_15151,N_19528);
nand U29061 (N_29061,N_19053,N_12130);
nand U29062 (N_29062,N_19879,N_10663);
nand U29063 (N_29063,N_11376,N_16737);
xor U29064 (N_29064,N_19159,N_10876);
nand U29065 (N_29065,N_18483,N_10820);
nor U29066 (N_29066,N_16842,N_12561);
nand U29067 (N_29067,N_17333,N_17191);
or U29068 (N_29068,N_10671,N_11708);
or U29069 (N_29069,N_18509,N_10287);
nand U29070 (N_29070,N_18996,N_16721);
and U29071 (N_29071,N_15273,N_18341);
nand U29072 (N_29072,N_10550,N_12141);
nand U29073 (N_29073,N_14484,N_11295);
xor U29074 (N_29074,N_13072,N_14803);
nor U29075 (N_29075,N_13497,N_11466);
nor U29076 (N_29076,N_19021,N_18569);
and U29077 (N_29077,N_18072,N_13130);
xor U29078 (N_29078,N_15212,N_12691);
xor U29079 (N_29079,N_11589,N_18485);
or U29080 (N_29080,N_14863,N_17006);
and U29081 (N_29081,N_15717,N_17823);
or U29082 (N_29082,N_10969,N_18682);
nor U29083 (N_29083,N_17979,N_15212);
and U29084 (N_29084,N_15851,N_10614);
or U29085 (N_29085,N_15422,N_15602);
nor U29086 (N_29086,N_10513,N_19475);
nand U29087 (N_29087,N_12706,N_12687);
nor U29088 (N_29088,N_10417,N_10591);
nand U29089 (N_29089,N_13520,N_16696);
and U29090 (N_29090,N_14943,N_11504);
or U29091 (N_29091,N_14731,N_15424);
or U29092 (N_29092,N_12303,N_11681);
nor U29093 (N_29093,N_18615,N_17538);
nand U29094 (N_29094,N_10505,N_14207);
xor U29095 (N_29095,N_14893,N_13955);
or U29096 (N_29096,N_11596,N_11780);
and U29097 (N_29097,N_12798,N_16074);
nor U29098 (N_29098,N_14616,N_16865);
or U29099 (N_29099,N_15719,N_13964);
and U29100 (N_29100,N_12082,N_11181);
or U29101 (N_29101,N_12934,N_14985);
nor U29102 (N_29102,N_17874,N_10241);
nor U29103 (N_29103,N_19980,N_10651);
and U29104 (N_29104,N_12759,N_15560);
and U29105 (N_29105,N_13967,N_11437);
nand U29106 (N_29106,N_15299,N_11464);
nand U29107 (N_29107,N_13704,N_12513);
nor U29108 (N_29108,N_14210,N_18613);
nand U29109 (N_29109,N_19145,N_15401);
and U29110 (N_29110,N_19581,N_11261);
nand U29111 (N_29111,N_19847,N_10744);
and U29112 (N_29112,N_14919,N_11549);
and U29113 (N_29113,N_13584,N_16851);
nor U29114 (N_29114,N_14406,N_14111);
nor U29115 (N_29115,N_14664,N_16190);
nand U29116 (N_29116,N_12844,N_11754);
or U29117 (N_29117,N_18299,N_10080);
and U29118 (N_29118,N_11167,N_15266);
and U29119 (N_29119,N_12873,N_13650);
nor U29120 (N_29120,N_17141,N_14630);
and U29121 (N_29121,N_15232,N_19339);
and U29122 (N_29122,N_12907,N_17049);
or U29123 (N_29123,N_13099,N_12595);
nand U29124 (N_29124,N_14428,N_11184);
nor U29125 (N_29125,N_19410,N_10654);
xnor U29126 (N_29126,N_13676,N_11854);
and U29127 (N_29127,N_17459,N_17110);
nand U29128 (N_29128,N_14351,N_12981);
or U29129 (N_29129,N_10792,N_10558);
xnor U29130 (N_29130,N_19801,N_17232);
nand U29131 (N_29131,N_12242,N_13008);
or U29132 (N_29132,N_12007,N_10015);
xor U29133 (N_29133,N_14501,N_18542);
nor U29134 (N_29134,N_14799,N_16990);
and U29135 (N_29135,N_15705,N_10503);
or U29136 (N_29136,N_12622,N_16289);
nor U29137 (N_29137,N_17846,N_19462);
or U29138 (N_29138,N_19961,N_16714);
or U29139 (N_29139,N_14364,N_19705);
xor U29140 (N_29140,N_14452,N_11303);
or U29141 (N_29141,N_11919,N_19288);
xnor U29142 (N_29142,N_11441,N_11012);
and U29143 (N_29143,N_10745,N_14061);
or U29144 (N_29144,N_11049,N_11510);
xor U29145 (N_29145,N_19906,N_12977);
nand U29146 (N_29146,N_11021,N_13553);
nand U29147 (N_29147,N_17163,N_11973);
or U29148 (N_29148,N_16398,N_10491);
nor U29149 (N_29149,N_16646,N_13967);
and U29150 (N_29150,N_16741,N_17149);
or U29151 (N_29151,N_17686,N_11206);
or U29152 (N_29152,N_14072,N_13507);
and U29153 (N_29153,N_17674,N_13910);
nor U29154 (N_29154,N_19552,N_19913);
and U29155 (N_29155,N_18220,N_10466);
nand U29156 (N_29156,N_18595,N_12038);
or U29157 (N_29157,N_16375,N_19122);
or U29158 (N_29158,N_12203,N_17048);
and U29159 (N_29159,N_11638,N_11682);
nor U29160 (N_29160,N_15207,N_12081);
nand U29161 (N_29161,N_12988,N_15546);
xor U29162 (N_29162,N_12041,N_14889);
or U29163 (N_29163,N_15423,N_18621);
nand U29164 (N_29164,N_12515,N_16981);
and U29165 (N_29165,N_14700,N_16222);
nand U29166 (N_29166,N_17014,N_13833);
and U29167 (N_29167,N_18075,N_12683);
and U29168 (N_29168,N_19675,N_13244);
or U29169 (N_29169,N_17406,N_14402);
xor U29170 (N_29170,N_11892,N_12093);
nand U29171 (N_29171,N_17688,N_10212);
nand U29172 (N_29172,N_12606,N_16356);
nor U29173 (N_29173,N_12557,N_11711);
or U29174 (N_29174,N_14513,N_14529);
xnor U29175 (N_29175,N_15181,N_16644);
xor U29176 (N_29176,N_15395,N_15425);
xnor U29177 (N_29177,N_13129,N_15464);
and U29178 (N_29178,N_10689,N_15464);
nor U29179 (N_29179,N_10221,N_10809);
or U29180 (N_29180,N_12891,N_18658);
nand U29181 (N_29181,N_10456,N_16195);
nand U29182 (N_29182,N_18842,N_10445);
or U29183 (N_29183,N_15696,N_10212);
and U29184 (N_29184,N_16354,N_18193);
or U29185 (N_29185,N_11030,N_17411);
or U29186 (N_29186,N_10027,N_13090);
or U29187 (N_29187,N_18365,N_13267);
or U29188 (N_29188,N_15357,N_14585);
nor U29189 (N_29189,N_19493,N_14991);
nand U29190 (N_29190,N_16277,N_10098);
xor U29191 (N_29191,N_18864,N_10089);
nand U29192 (N_29192,N_12290,N_15536);
nand U29193 (N_29193,N_10673,N_17260);
nand U29194 (N_29194,N_17005,N_14417);
nand U29195 (N_29195,N_10944,N_10246);
or U29196 (N_29196,N_14598,N_12642);
xnor U29197 (N_29197,N_14928,N_19742);
or U29198 (N_29198,N_10191,N_11100);
and U29199 (N_29199,N_14842,N_11189);
or U29200 (N_29200,N_11880,N_11765);
or U29201 (N_29201,N_11613,N_18245);
nand U29202 (N_29202,N_18275,N_13507);
nand U29203 (N_29203,N_16329,N_19233);
nand U29204 (N_29204,N_18695,N_11764);
or U29205 (N_29205,N_10429,N_12400);
nand U29206 (N_29206,N_10116,N_12686);
xnor U29207 (N_29207,N_18497,N_11850);
or U29208 (N_29208,N_11824,N_15368);
nor U29209 (N_29209,N_12400,N_16816);
nand U29210 (N_29210,N_10663,N_16251);
and U29211 (N_29211,N_14896,N_12112);
nor U29212 (N_29212,N_10210,N_13097);
and U29213 (N_29213,N_11563,N_19937);
nand U29214 (N_29214,N_16488,N_11221);
nor U29215 (N_29215,N_10972,N_11388);
xnor U29216 (N_29216,N_11310,N_13356);
nor U29217 (N_29217,N_10737,N_11397);
nand U29218 (N_29218,N_10253,N_11277);
or U29219 (N_29219,N_16881,N_12002);
and U29220 (N_29220,N_10475,N_16854);
nor U29221 (N_29221,N_10240,N_18246);
and U29222 (N_29222,N_17413,N_17041);
nor U29223 (N_29223,N_10019,N_11591);
nor U29224 (N_29224,N_11182,N_13220);
and U29225 (N_29225,N_19691,N_10788);
or U29226 (N_29226,N_17491,N_17237);
and U29227 (N_29227,N_19126,N_17263);
xor U29228 (N_29228,N_19008,N_18786);
and U29229 (N_29229,N_18423,N_15196);
nor U29230 (N_29230,N_15670,N_10090);
or U29231 (N_29231,N_16216,N_10058);
nand U29232 (N_29232,N_11418,N_11541);
nor U29233 (N_29233,N_12132,N_16659);
xnor U29234 (N_29234,N_19358,N_19772);
nor U29235 (N_29235,N_13340,N_11617);
nor U29236 (N_29236,N_10694,N_15902);
nand U29237 (N_29237,N_15236,N_12024);
nand U29238 (N_29238,N_15444,N_11822);
or U29239 (N_29239,N_16451,N_13530);
nand U29240 (N_29240,N_12276,N_19541);
or U29241 (N_29241,N_16538,N_11374);
or U29242 (N_29242,N_10618,N_16780);
nor U29243 (N_29243,N_14798,N_15107);
and U29244 (N_29244,N_14545,N_14653);
nand U29245 (N_29245,N_16142,N_11616);
nor U29246 (N_29246,N_13587,N_10483);
xnor U29247 (N_29247,N_12161,N_18307);
nor U29248 (N_29248,N_19458,N_13313);
xnor U29249 (N_29249,N_12381,N_10913);
and U29250 (N_29250,N_19433,N_11379);
nor U29251 (N_29251,N_13180,N_10330);
or U29252 (N_29252,N_14516,N_17018);
nor U29253 (N_29253,N_13198,N_10969);
nand U29254 (N_29254,N_13638,N_15712);
nand U29255 (N_29255,N_18987,N_14058);
or U29256 (N_29256,N_12759,N_13871);
and U29257 (N_29257,N_18996,N_15771);
and U29258 (N_29258,N_19516,N_12858);
or U29259 (N_29259,N_18073,N_14490);
and U29260 (N_29260,N_12271,N_10811);
nor U29261 (N_29261,N_19651,N_15385);
or U29262 (N_29262,N_12753,N_13183);
nor U29263 (N_29263,N_19161,N_13386);
or U29264 (N_29264,N_10751,N_10961);
nor U29265 (N_29265,N_18927,N_12936);
nor U29266 (N_29266,N_18394,N_12702);
nor U29267 (N_29267,N_14135,N_17353);
nand U29268 (N_29268,N_10249,N_14337);
xnor U29269 (N_29269,N_18002,N_12178);
nand U29270 (N_29270,N_10195,N_19988);
nor U29271 (N_29271,N_19279,N_12756);
xor U29272 (N_29272,N_19433,N_14382);
and U29273 (N_29273,N_19817,N_16957);
nand U29274 (N_29274,N_17124,N_11532);
nand U29275 (N_29275,N_11028,N_17807);
and U29276 (N_29276,N_13609,N_13538);
and U29277 (N_29277,N_12753,N_13603);
or U29278 (N_29278,N_18835,N_18372);
and U29279 (N_29279,N_15017,N_10873);
and U29280 (N_29280,N_15858,N_12511);
or U29281 (N_29281,N_18262,N_19878);
and U29282 (N_29282,N_10996,N_18168);
or U29283 (N_29283,N_18218,N_13184);
nor U29284 (N_29284,N_15627,N_15477);
nand U29285 (N_29285,N_10744,N_18718);
nor U29286 (N_29286,N_11729,N_19070);
or U29287 (N_29287,N_14792,N_11140);
nand U29288 (N_29288,N_10616,N_17818);
nor U29289 (N_29289,N_15710,N_14742);
or U29290 (N_29290,N_18434,N_15628);
nand U29291 (N_29291,N_18473,N_19418);
nand U29292 (N_29292,N_13806,N_10839);
nor U29293 (N_29293,N_18577,N_11845);
xnor U29294 (N_29294,N_14662,N_17805);
or U29295 (N_29295,N_16461,N_19762);
and U29296 (N_29296,N_17356,N_18236);
and U29297 (N_29297,N_16430,N_15275);
xor U29298 (N_29298,N_13317,N_14299);
or U29299 (N_29299,N_11577,N_15105);
nand U29300 (N_29300,N_12668,N_19834);
or U29301 (N_29301,N_10103,N_10428);
nor U29302 (N_29302,N_13586,N_14233);
nor U29303 (N_29303,N_14940,N_18326);
nand U29304 (N_29304,N_12444,N_14139);
nand U29305 (N_29305,N_10504,N_12149);
and U29306 (N_29306,N_14222,N_17558);
and U29307 (N_29307,N_11626,N_15180);
nand U29308 (N_29308,N_17834,N_10741);
nor U29309 (N_29309,N_10812,N_14880);
xor U29310 (N_29310,N_14191,N_15320);
or U29311 (N_29311,N_19938,N_18972);
and U29312 (N_29312,N_10506,N_11205);
nor U29313 (N_29313,N_10131,N_15136);
or U29314 (N_29314,N_19430,N_11070);
and U29315 (N_29315,N_13331,N_12989);
or U29316 (N_29316,N_10944,N_11105);
nand U29317 (N_29317,N_19737,N_19487);
or U29318 (N_29318,N_17248,N_17294);
or U29319 (N_29319,N_17291,N_19529);
nand U29320 (N_29320,N_14195,N_15114);
nand U29321 (N_29321,N_13883,N_16773);
nor U29322 (N_29322,N_10705,N_14470);
nor U29323 (N_29323,N_13529,N_19637);
and U29324 (N_29324,N_10619,N_17237);
xnor U29325 (N_29325,N_17316,N_17420);
nor U29326 (N_29326,N_11493,N_12053);
nor U29327 (N_29327,N_16817,N_16709);
nand U29328 (N_29328,N_12948,N_18401);
nand U29329 (N_29329,N_13844,N_10722);
or U29330 (N_29330,N_19600,N_12019);
nand U29331 (N_29331,N_10348,N_10130);
nand U29332 (N_29332,N_17543,N_10982);
nor U29333 (N_29333,N_15641,N_15999);
nor U29334 (N_29334,N_12356,N_10398);
or U29335 (N_29335,N_16600,N_18610);
nand U29336 (N_29336,N_19213,N_14834);
xor U29337 (N_29337,N_17370,N_13596);
nand U29338 (N_29338,N_18422,N_14469);
or U29339 (N_29339,N_14403,N_14811);
or U29340 (N_29340,N_18129,N_18928);
nor U29341 (N_29341,N_16456,N_17061);
or U29342 (N_29342,N_15880,N_14710);
or U29343 (N_29343,N_19682,N_11046);
nor U29344 (N_29344,N_19682,N_15004);
and U29345 (N_29345,N_11613,N_14280);
nor U29346 (N_29346,N_13990,N_12542);
or U29347 (N_29347,N_18166,N_15089);
and U29348 (N_29348,N_17888,N_12718);
and U29349 (N_29349,N_15180,N_13726);
nor U29350 (N_29350,N_13320,N_15871);
and U29351 (N_29351,N_17388,N_14873);
and U29352 (N_29352,N_15015,N_15760);
nand U29353 (N_29353,N_19521,N_10681);
nor U29354 (N_29354,N_12393,N_15638);
nor U29355 (N_29355,N_13586,N_19805);
or U29356 (N_29356,N_16280,N_13544);
or U29357 (N_29357,N_14796,N_18845);
nor U29358 (N_29358,N_19939,N_10993);
xnor U29359 (N_29359,N_10593,N_17035);
and U29360 (N_29360,N_14402,N_12251);
nor U29361 (N_29361,N_11987,N_16813);
or U29362 (N_29362,N_19086,N_12068);
nor U29363 (N_29363,N_18240,N_14498);
nand U29364 (N_29364,N_19288,N_12465);
nor U29365 (N_29365,N_14697,N_16918);
nand U29366 (N_29366,N_16032,N_18127);
nand U29367 (N_29367,N_16714,N_18600);
xnor U29368 (N_29368,N_19881,N_16355);
xor U29369 (N_29369,N_16212,N_19107);
and U29370 (N_29370,N_16547,N_11986);
nand U29371 (N_29371,N_11144,N_14994);
nor U29372 (N_29372,N_17749,N_19369);
and U29373 (N_29373,N_12008,N_10486);
or U29374 (N_29374,N_13480,N_16781);
or U29375 (N_29375,N_19032,N_12980);
nand U29376 (N_29376,N_17845,N_15229);
nand U29377 (N_29377,N_15193,N_10796);
xnor U29378 (N_29378,N_17326,N_12940);
or U29379 (N_29379,N_11800,N_19208);
and U29380 (N_29380,N_19390,N_14162);
nand U29381 (N_29381,N_12961,N_11201);
nor U29382 (N_29382,N_13297,N_11839);
nor U29383 (N_29383,N_10374,N_19440);
nor U29384 (N_29384,N_16188,N_13026);
or U29385 (N_29385,N_14206,N_12848);
or U29386 (N_29386,N_16791,N_15846);
or U29387 (N_29387,N_11000,N_15485);
and U29388 (N_29388,N_11665,N_16446);
nor U29389 (N_29389,N_16867,N_11375);
nor U29390 (N_29390,N_19364,N_17990);
and U29391 (N_29391,N_13628,N_17495);
and U29392 (N_29392,N_11845,N_17865);
xor U29393 (N_29393,N_12568,N_16608);
and U29394 (N_29394,N_12094,N_13040);
nor U29395 (N_29395,N_18255,N_12508);
and U29396 (N_29396,N_11769,N_14163);
or U29397 (N_29397,N_10923,N_14453);
or U29398 (N_29398,N_11420,N_17551);
nor U29399 (N_29399,N_15075,N_16860);
and U29400 (N_29400,N_19335,N_12526);
or U29401 (N_29401,N_18698,N_10630);
and U29402 (N_29402,N_11519,N_11954);
nand U29403 (N_29403,N_19165,N_11168);
and U29404 (N_29404,N_16890,N_10488);
nand U29405 (N_29405,N_18467,N_17571);
xor U29406 (N_29406,N_19541,N_14220);
or U29407 (N_29407,N_13109,N_17888);
nand U29408 (N_29408,N_10781,N_11357);
nor U29409 (N_29409,N_18308,N_15343);
nor U29410 (N_29410,N_13247,N_12172);
nor U29411 (N_29411,N_12370,N_14770);
nand U29412 (N_29412,N_17039,N_15130);
nand U29413 (N_29413,N_17614,N_12075);
nor U29414 (N_29414,N_12035,N_14529);
nor U29415 (N_29415,N_16509,N_10140);
nand U29416 (N_29416,N_10384,N_10067);
nor U29417 (N_29417,N_18241,N_18056);
nand U29418 (N_29418,N_13472,N_14426);
nand U29419 (N_29419,N_16565,N_14471);
nor U29420 (N_29420,N_17454,N_19625);
and U29421 (N_29421,N_18950,N_17337);
nand U29422 (N_29422,N_17085,N_13954);
nor U29423 (N_29423,N_14249,N_17866);
and U29424 (N_29424,N_13574,N_17185);
and U29425 (N_29425,N_10256,N_11012);
nor U29426 (N_29426,N_16577,N_16082);
nor U29427 (N_29427,N_17020,N_12736);
and U29428 (N_29428,N_19741,N_18796);
nand U29429 (N_29429,N_10377,N_12965);
or U29430 (N_29430,N_16103,N_19258);
and U29431 (N_29431,N_14119,N_18523);
or U29432 (N_29432,N_14662,N_11535);
nand U29433 (N_29433,N_15776,N_16671);
nand U29434 (N_29434,N_11556,N_18848);
and U29435 (N_29435,N_11690,N_16290);
and U29436 (N_29436,N_14471,N_15657);
nand U29437 (N_29437,N_15116,N_12760);
nor U29438 (N_29438,N_11609,N_10878);
or U29439 (N_29439,N_15523,N_16989);
nand U29440 (N_29440,N_15040,N_18027);
nand U29441 (N_29441,N_19393,N_12227);
and U29442 (N_29442,N_17799,N_19806);
xor U29443 (N_29443,N_19834,N_16316);
and U29444 (N_29444,N_14245,N_18533);
and U29445 (N_29445,N_14047,N_11776);
xnor U29446 (N_29446,N_14704,N_12685);
nand U29447 (N_29447,N_16132,N_18051);
and U29448 (N_29448,N_11710,N_15408);
nand U29449 (N_29449,N_12332,N_19072);
or U29450 (N_29450,N_13234,N_10243);
or U29451 (N_29451,N_14472,N_15331);
or U29452 (N_29452,N_14253,N_10840);
and U29453 (N_29453,N_15344,N_17125);
and U29454 (N_29454,N_11778,N_11402);
xor U29455 (N_29455,N_16114,N_12701);
nand U29456 (N_29456,N_13997,N_13863);
and U29457 (N_29457,N_10337,N_12042);
and U29458 (N_29458,N_17066,N_14557);
nand U29459 (N_29459,N_13153,N_18585);
nand U29460 (N_29460,N_14899,N_15302);
and U29461 (N_29461,N_12806,N_13017);
and U29462 (N_29462,N_18956,N_19154);
or U29463 (N_29463,N_17446,N_16307);
nor U29464 (N_29464,N_19333,N_12688);
nand U29465 (N_29465,N_16092,N_11321);
nor U29466 (N_29466,N_19868,N_12370);
nor U29467 (N_29467,N_10386,N_17524);
nand U29468 (N_29468,N_12938,N_13067);
or U29469 (N_29469,N_10956,N_16006);
or U29470 (N_29470,N_15629,N_10255);
nand U29471 (N_29471,N_14154,N_15651);
nor U29472 (N_29472,N_13917,N_11358);
and U29473 (N_29473,N_13004,N_14789);
or U29474 (N_29474,N_13089,N_13448);
and U29475 (N_29475,N_11612,N_18238);
or U29476 (N_29476,N_16500,N_18567);
xor U29477 (N_29477,N_16620,N_11038);
nor U29478 (N_29478,N_14942,N_14813);
and U29479 (N_29479,N_17123,N_17871);
nand U29480 (N_29480,N_12988,N_16185);
nor U29481 (N_29481,N_10123,N_17954);
nor U29482 (N_29482,N_12303,N_12905);
and U29483 (N_29483,N_13895,N_17188);
nor U29484 (N_29484,N_18015,N_12176);
nand U29485 (N_29485,N_18072,N_14737);
or U29486 (N_29486,N_11351,N_14719);
nor U29487 (N_29487,N_14166,N_14684);
and U29488 (N_29488,N_18160,N_12639);
nand U29489 (N_29489,N_18052,N_14817);
or U29490 (N_29490,N_14138,N_13967);
nand U29491 (N_29491,N_19513,N_16468);
nor U29492 (N_29492,N_11641,N_19715);
xnor U29493 (N_29493,N_19794,N_11168);
or U29494 (N_29494,N_12788,N_10841);
nand U29495 (N_29495,N_12771,N_13793);
and U29496 (N_29496,N_12328,N_17987);
nand U29497 (N_29497,N_19131,N_10032);
nand U29498 (N_29498,N_11950,N_18114);
and U29499 (N_29499,N_15446,N_16885);
xnor U29500 (N_29500,N_16879,N_11843);
nor U29501 (N_29501,N_11394,N_11279);
xnor U29502 (N_29502,N_14290,N_15200);
or U29503 (N_29503,N_15381,N_14967);
or U29504 (N_29504,N_18245,N_11236);
nor U29505 (N_29505,N_15883,N_13826);
or U29506 (N_29506,N_14098,N_16556);
or U29507 (N_29507,N_18571,N_11627);
nor U29508 (N_29508,N_15181,N_10375);
nand U29509 (N_29509,N_19023,N_11710);
nor U29510 (N_29510,N_16669,N_18530);
nand U29511 (N_29511,N_16706,N_10608);
and U29512 (N_29512,N_14764,N_17910);
xnor U29513 (N_29513,N_12837,N_18868);
or U29514 (N_29514,N_11355,N_11244);
and U29515 (N_29515,N_14628,N_11972);
and U29516 (N_29516,N_11207,N_19156);
nand U29517 (N_29517,N_11018,N_13596);
nor U29518 (N_29518,N_18654,N_10988);
or U29519 (N_29519,N_11964,N_14981);
nand U29520 (N_29520,N_16118,N_11278);
nor U29521 (N_29521,N_14476,N_13796);
or U29522 (N_29522,N_10022,N_11765);
nor U29523 (N_29523,N_12386,N_16261);
nand U29524 (N_29524,N_19647,N_14512);
and U29525 (N_29525,N_10482,N_17085);
and U29526 (N_29526,N_11888,N_12724);
and U29527 (N_29527,N_17202,N_15642);
or U29528 (N_29528,N_16453,N_12377);
nor U29529 (N_29529,N_16601,N_10069);
xnor U29530 (N_29530,N_18558,N_14354);
nor U29531 (N_29531,N_12748,N_18010);
and U29532 (N_29532,N_10975,N_14817);
nand U29533 (N_29533,N_10672,N_14756);
nor U29534 (N_29534,N_11459,N_11353);
or U29535 (N_29535,N_10455,N_17190);
or U29536 (N_29536,N_16966,N_19039);
and U29537 (N_29537,N_19532,N_12993);
nor U29538 (N_29538,N_17358,N_19512);
nor U29539 (N_29539,N_13765,N_11465);
and U29540 (N_29540,N_16799,N_14347);
xor U29541 (N_29541,N_13346,N_18931);
nor U29542 (N_29542,N_15471,N_16453);
and U29543 (N_29543,N_12980,N_19320);
nor U29544 (N_29544,N_12410,N_12334);
nand U29545 (N_29545,N_14707,N_11421);
nor U29546 (N_29546,N_12526,N_11165);
xnor U29547 (N_29547,N_10214,N_14611);
nor U29548 (N_29548,N_14373,N_14367);
and U29549 (N_29549,N_14052,N_18746);
or U29550 (N_29550,N_16614,N_13813);
or U29551 (N_29551,N_18834,N_13706);
nand U29552 (N_29552,N_15690,N_18578);
nand U29553 (N_29553,N_18782,N_12381);
nand U29554 (N_29554,N_14546,N_14145);
nor U29555 (N_29555,N_13836,N_16661);
or U29556 (N_29556,N_18587,N_15063);
xor U29557 (N_29557,N_19749,N_17851);
nand U29558 (N_29558,N_18292,N_17184);
and U29559 (N_29559,N_12173,N_16821);
xnor U29560 (N_29560,N_14233,N_14990);
nor U29561 (N_29561,N_14462,N_10904);
nor U29562 (N_29562,N_12833,N_15720);
nor U29563 (N_29563,N_18186,N_11889);
and U29564 (N_29564,N_13927,N_13017);
and U29565 (N_29565,N_14875,N_13081);
nor U29566 (N_29566,N_12875,N_19893);
and U29567 (N_29567,N_15583,N_14844);
nand U29568 (N_29568,N_15505,N_17954);
or U29569 (N_29569,N_16218,N_15811);
nand U29570 (N_29570,N_13307,N_14393);
nor U29571 (N_29571,N_10662,N_15730);
nor U29572 (N_29572,N_15869,N_17962);
nor U29573 (N_29573,N_15953,N_11487);
and U29574 (N_29574,N_14626,N_13089);
nor U29575 (N_29575,N_17631,N_15123);
nand U29576 (N_29576,N_13485,N_11916);
or U29577 (N_29577,N_10998,N_16059);
nor U29578 (N_29578,N_13678,N_19938);
or U29579 (N_29579,N_16511,N_12695);
and U29580 (N_29580,N_11590,N_18116);
and U29581 (N_29581,N_17755,N_10971);
xor U29582 (N_29582,N_19644,N_16508);
nor U29583 (N_29583,N_13688,N_11058);
and U29584 (N_29584,N_11633,N_11086);
nand U29585 (N_29585,N_13486,N_11744);
nand U29586 (N_29586,N_15677,N_15705);
or U29587 (N_29587,N_10835,N_14152);
and U29588 (N_29588,N_18925,N_18866);
xor U29589 (N_29589,N_10622,N_12257);
nor U29590 (N_29590,N_17139,N_19065);
and U29591 (N_29591,N_16166,N_16125);
and U29592 (N_29592,N_15986,N_12680);
or U29593 (N_29593,N_17468,N_18745);
xnor U29594 (N_29594,N_15761,N_12820);
or U29595 (N_29595,N_19303,N_10761);
or U29596 (N_29596,N_17998,N_11917);
or U29597 (N_29597,N_14682,N_18934);
nand U29598 (N_29598,N_17952,N_10695);
xnor U29599 (N_29599,N_10052,N_13718);
nand U29600 (N_29600,N_19080,N_14113);
or U29601 (N_29601,N_16511,N_15090);
and U29602 (N_29602,N_19864,N_12001);
nand U29603 (N_29603,N_19137,N_19925);
and U29604 (N_29604,N_11413,N_17195);
and U29605 (N_29605,N_10456,N_16504);
nand U29606 (N_29606,N_19275,N_15165);
or U29607 (N_29607,N_16539,N_15849);
nor U29608 (N_29608,N_16431,N_19980);
xor U29609 (N_29609,N_16385,N_12004);
or U29610 (N_29610,N_19770,N_16663);
nor U29611 (N_29611,N_10887,N_10419);
or U29612 (N_29612,N_18517,N_17776);
nor U29613 (N_29613,N_12705,N_14863);
xor U29614 (N_29614,N_17560,N_12350);
or U29615 (N_29615,N_13374,N_13373);
nor U29616 (N_29616,N_12398,N_10523);
nand U29617 (N_29617,N_10743,N_17357);
nor U29618 (N_29618,N_18452,N_18330);
nor U29619 (N_29619,N_16980,N_11379);
nand U29620 (N_29620,N_19418,N_12872);
nor U29621 (N_29621,N_14532,N_13653);
nand U29622 (N_29622,N_17657,N_10082);
or U29623 (N_29623,N_19237,N_13715);
or U29624 (N_29624,N_11577,N_14044);
nor U29625 (N_29625,N_16059,N_14018);
nand U29626 (N_29626,N_14752,N_18187);
nor U29627 (N_29627,N_19576,N_14162);
and U29628 (N_29628,N_19270,N_18475);
and U29629 (N_29629,N_18850,N_19753);
nor U29630 (N_29630,N_14522,N_11704);
nor U29631 (N_29631,N_14830,N_10468);
or U29632 (N_29632,N_12829,N_10441);
xor U29633 (N_29633,N_13404,N_19931);
xor U29634 (N_29634,N_16895,N_14795);
or U29635 (N_29635,N_16532,N_19170);
and U29636 (N_29636,N_19407,N_11258);
nor U29637 (N_29637,N_12655,N_16072);
nand U29638 (N_29638,N_19177,N_17148);
nand U29639 (N_29639,N_19957,N_15262);
nand U29640 (N_29640,N_19949,N_11994);
and U29641 (N_29641,N_19871,N_15119);
nor U29642 (N_29642,N_13944,N_19001);
and U29643 (N_29643,N_10341,N_14867);
nor U29644 (N_29644,N_16760,N_16991);
or U29645 (N_29645,N_12214,N_12113);
nand U29646 (N_29646,N_18955,N_17769);
or U29647 (N_29647,N_18511,N_11800);
or U29648 (N_29648,N_18618,N_13370);
nand U29649 (N_29649,N_13390,N_18818);
or U29650 (N_29650,N_13624,N_14401);
nor U29651 (N_29651,N_13920,N_18620);
nor U29652 (N_29652,N_10204,N_16188);
or U29653 (N_29653,N_19662,N_19717);
or U29654 (N_29654,N_11539,N_15593);
nor U29655 (N_29655,N_10084,N_13009);
or U29656 (N_29656,N_14082,N_16018);
nor U29657 (N_29657,N_17016,N_10003);
nor U29658 (N_29658,N_11563,N_16594);
nor U29659 (N_29659,N_12172,N_12351);
or U29660 (N_29660,N_19764,N_11495);
or U29661 (N_29661,N_12621,N_19808);
or U29662 (N_29662,N_16656,N_19363);
nand U29663 (N_29663,N_19774,N_16289);
or U29664 (N_29664,N_10622,N_16163);
and U29665 (N_29665,N_15957,N_15582);
or U29666 (N_29666,N_15540,N_18741);
or U29667 (N_29667,N_15789,N_12807);
and U29668 (N_29668,N_13828,N_14503);
nand U29669 (N_29669,N_11082,N_12513);
nor U29670 (N_29670,N_10154,N_12800);
xnor U29671 (N_29671,N_18790,N_15268);
nor U29672 (N_29672,N_15935,N_17965);
or U29673 (N_29673,N_18957,N_12438);
and U29674 (N_29674,N_18700,N_10685);
or U29675 (N_29675,N_17241,N_14532);
nor U29676 (N_29676,N_17407,N_13173);
nor U29677 (N_29677,N_18391,N_16098);
nand U29678 (N_29678,N_13469,N_15281);
nand U29679 (N_29679,N_17951,N_12783);
or U29680 (N_29680,N_14304,N_10415);
nor U29681 (N_29681,N_16880,N_14267);
nand U29682 (N_29682,N_10154,N_11901);
nor U29683 (N_29683,N_17532,N_11383);
nor U29684 (N_29684,N_10432,N_10918);
nor U29685 (N_29685,N_11371,N_12200);
or U29686 (N_29686,N_19568,N_10516);
nand U29687 (N_29687,N_12146,N_10662);
nand U29688 (N_29688,N_18557,N_16642);
and U29689 (N_29689,N_17440,N_16532);
nand U29690 (N_29690,N_17799,N_19706);
nor U29691 (N_29691,N_18350,N_13810);
nand U29692 (N_29692,N_13971,N_16213);
nand U29693 (N_29693,N_15614,N_18108);
nor U29694 (N_29694,N_10288,N_13927);
and U29695 (N_29695,N_13535,N_17308);
xnor U29696 (N_29696,N_19292,N_12489);
or U29697 (N_29697,N_13370,N_18655);
xnor U29698 (N_29698,N_11342,N_16729);
or U29699 (N_29699,N_18585,N_16299);
or U29700 (N_29700,N_14458,N_15537);
or U29701 (N_29701,N_15512,N_14601);
nand U29702 (N_29702,N_10936,N_19111);
nor U29703 (N_29703,N_14329,N_15712);
nor U29704 (N_29704,N_18505,N_17148);
or U29705 (N_29705,N_12269,N_14592);
and U29706 (N_29706,N_13247,N_19076);
and U29707 (N_29707,N_15313,N_10964);
nor U29708 (N_29708,N_13368,N_17573);
and U29709 (N_29709,N_17786,N_12395);
and U29710 (N_29710,N_18895,N_18117);
nor U29711 (N_29711,N_19326,N_18624);
or U29712 (N_29712,N_14994,N_17050);
nand U29713 (N_29713,N_10678,N_15558);
xnor U29714 (N_29714,N_11633,N_17211);
nand U29715 (N_29715,N_18376,N_15700);
and U29716 (N_29716,N_19052,N_19287);
xnor U29717 (N_29717,N_13738,N_17981);
or U29718 (N_29718,N_11787,N_14720);
nor U29719 (N_29719,N_13320,N_19464);
or U29720 (N_29720,N_14405,N_11014);
xnor U29721 (N_29721,N_14647,N_19213);
or U29722 (N_29722,N_11700,N_16998);
and U29723 (N_29723,N_17236,N_14936);
or U29724 (N_29724,N_15447,N_14308);
nand U29725 (N_29725,N_13117,N_14315);
nor U29726 (N_29726,N_18297,N_14772);
nor U29727 (N_29727,N_11108,N_14309);
nor U29728 (N_29728,N_16133,N_17338);
and U29729 (N_29729,N_16100,N_12927);
nor U29730 (N_29730,N_14301,N_18900);
nand U29731 (N_29731,N_10134,N_11422);
or U29732 (N_29732,N_13370,N_12604);
or U29733 (N_29733,N_15835,N_12209);
or U29734 (N_29734,N_10270,N_10606);
or U29735 (N_29735,N_15454,N_15442);
nor U29736 (N_29736,N_15810,N_15594);
nor U29737 (N_29737,N_19469,N_13834);
and U29738 (N_29738,N_10270,N_16410);
nand U29739 (N_29739,N_14801,N_18833);
nand U29740 (N_29740,N_19435,N_17792);
or U29741 (N_29741,N_12119,N_17775);
nand U29742 (N_29742,N_13806,N_16397);
nor U29743 (N_29743,N_17377,N_18115);
and U29744 (N_29744,N_19339,N_18540);
or U29745 (N_29745,N_14205,N_18990);
or U29746 (N_29746,N_14531,N_11031);
nor U29747 (N_29747,N_14831,N_12796);
nand U29748 (N_29748,N_15102,N_10519);
nand U29749 (N_29749,N_13367,N_18227);
nor U29750 (N_29750,N_15868,N_14338);
nand U29751 (N_29751,N_19167,N_13092);
or U29752 (N_29752,N_15775,N_18232);
or U29753 (N_29753,N_18433,N_12351);
nand U29754 (N_29754,N_15519,N_14352);
and U29755 (N_29755,N_12541,N_11244);
and U29756 (N_29756,N_14566,N_14545);
or U29757 (N_29757,N_17921,N_16986);
and U29758 (N_29758,N_10634,N_13216);
xor U29759 (N_29759,N_19480,N_15239);
nor U29760 (N_29760,N_12328,N_17274);
nand U29761 (N_29761,N_11694,N_19839);
nor U29762 (N_29762,N_15941,N_10910);
or U29763 (N_29763,N_19538,N_17412);
nand U29764 (N_29764,N_17756,N_16079);
xor U29765 (N_29765,N_11670,N_10573);
nand U29766 (N_29766,N_12205,N_16942);
or U29767 (N_29767,N_16706,N_11556);
nor U29768 (N_29768,N_12808,N_15211);
and U29769 (N_29769,N_19813,N_13980);
nor U29770 (N_29770,N_17512,N_11606);
nand U29771 (N_29771,N_13182,N_11279);
nor U29772 (N_29772,N_14282,N_11762);
or U29773 (N_29773,N_15074,N_14031);
nand U29774 (N_29774,N_16086,N_14998);
or U29775 (N_29775,N_17025,N_14153);
or U29776 (N_29776,N_13125,N_15670);
nor U29777 (N_29777,N_12567,N_15464);
and U29778 (N_29778,N_13278,N_10837);
xnor U29779 (N_29779,N_15420,N_19429);
nand U29780 (N_29780,N_12575,N_19681);
nor U29781 (N_29781,N_10712,N_16485);
xor U29782 (N_29782,N_11340,N_10620);
or U29783 (N_29783,N_15964,N_16785);
or U29784 (N_29784,N_11119,N_15044);
nand U29785 (N_29785,N_18070,N_16051);
nor U29786 (N_29786,N_15725,N_12590);
and U29787 (N_29787,N_18187,N_11093);
nand U29788 (N_29788,N_13310,N_19798);
nor U29789 (N_29789,N_14339,N_11106);
nand U29790 (N_29790,N_12467,N_19126);
and U29791 (N_29791,N_13356,N_18332);
nor U29792 (N_29792,N_13983,N_16832);
or U29793 (N_29793,N_17975,N_19727);
nor U29794 (N_29794,N_19718,N_10313);
or U29795 (N_29795,N_17863,N_14336);
and U29796 (N_29796,N_13571,N_10774);
nand U29797 (N_29797,N_10445,N_15888);
or U29798 (N_29798,N_13890,N_15442);
nand U29799 (N_29799,N_15978,N_11691);
nand U29800 (N_29800,N_14004,N_18086);
nor U29801 (N_29801,N_12002,N_12418);
nor U29802 (N_29802,N_11450,N_19997);
nand U29803 (N_29803,N_11894,N_17781);
or U29804 (N_29804,N_12152,N_17334);
and U29805 (N_29805,N_12264,N_14315);
nor U29806 (N_29806,N_11325,N_13839);
nand U29807 (N_29807,N_14922,N_11904);
nand U29808 (N_29808,N_11328,N_11820);
and U29809 (N_29809,N_11252,N_19891);
or U29810 (N_29810,N_18179,N_10274);
nand U29811 (N_29811,N_11438,N_17347);
xor U29812 (N_29812,N_14377,N_12265);
nor U29813 (N_29813,N_12742,N_18265);
nor U29814 (N_29814,N_11502,N_16070);
nor U29815 (N_29815,N_11182,N_18368);
xnor U29816 (N_29816,N_14081,N_18273);
xnor U29817 (N_29817,N_13413,N_11990);
nand U29818 (N_29818,N_19457,N_16411);
and U29819 (N_29819,N_13577,N_11164);
and U29820 (N_29820,N_16533,N_17861);
or U29821 (N_29821,N_12440,N_19324);
and U29822 (N_29822,N_19584,N_13370);
nor U29823 (N_29823,N_17245,N_11862);
xnor U29824 (N_29824,N_11967,N_10098);
nor U29825 (N_29825,N_19668,N_12537);
or U29826 (N_29826,N_12010,N_11083);
xnor U29827 (N_29827,N_13922,N_12444);
nor U29828 (N_29828,N_11307,N_19004);
xor U29829 (N_29829,N_10729,N_12316);
and U29830 (N_29830,N_15073,N_19845);
nand U29831 (N_29831,N_15233,N_10528);
or U29832 (N_29832,N_17885,N_13129);
or U29833 (N_29833,N_12045,N_12116);
nand U29834 (N_29834,N_14322,N_17599);
nand U29835 (N_29835,N_11340,N_13011);
nor U29836 (N_29836,N_17680,N_13988);
or U29837 (N_29837,N_16105,N_16636);
xor U29838 (N_29838,N_15173,N_11485);
nor U29839 (N_29839,N_17807,N_13361);
nand U29840 (N_29840,N_11081,N_17554);
xor U29841 (N_29841,N_13791,N_17397);
and U29842 (N_29842,N_17649,N_19037);
and U29843 (N_29843,N_16168,N_11499);
nand U29844 (N_29844,N_15698,N_19757);
nor U29845 (N_29845,N_14455,N_16898);
or U29846 (N_29846,N_15977,N_15373);
xnor U29847 (N_29847,N_18471,N_17281);
or U29848 (N_29848,N_15836,N_16885);
and U29849 (N_29849,N_11451,N_18569);
and U29850 (N_29850,N_18216,N_15043);
or U29851 (N_29851,N_18619,N_17161);
nor U29852 (N_29852,N_13184,N_10371);
nand U29853 (N_29853,N_15208,N_19129);
or U29854 (N_29854,N_15943,N_13914);
nor U29855 (N_29855,N_18254,N_10156);
and U29856 (N_29856,N_14088,N_19731);
or U29857 (N_29857,N_14799,N_19684);
nor U29858 (N_29858,N_19665,N_12466);
xnor U29859 (N_29859,N_12631,N_14577);
nor U29860 (N_29860,N_19936,N_15997);
and U29861 (N_29861,N_15677,N_19105);
or U29862 (N_29862,N_19561,N_15871);
nand U29863 (N_29863,N_10230,N_11045);
nand U29864 (N_29864,N_12133,N_15147);
nand U29865 (N_29865,N_13744,N_14004);
xor U29866 (N_29866,N_11463,N_12814);
nand U29867 (N_29867,N_10534,N_18725);
nor U29868 (N_29868,N_10313,N_15303);
and U29869 (N_29869,N_13022,N_16416);
xor U29870 (N_29870,N_13651,N_17730);
nor U29871 (N_29871,N_11251,N_14562);
nand U29872 (N_29872,N_15113,N_19138);
nor U29873 (N_29873,N_13047,N_17463);
and U29874 (N_29874,N_14926,N_18357);
nand U29875 (N_29875,N_12489,N_11492);
or U29876 (N_29876,N_16977,N_18244);
nand U29877 (N_29877,N_15152,N_19578);
or U29878 (N_29878,N_11475,N_11556);
or U29879 (N_29879,N_10726,N_16519);
xor U29880 (N_29880,N_10949,N_14122);
and U29881 (N_29881,N_19027,N_18665);
nor U29882 (N_29882,N_19563,N_15905);
nor U29883 (N_29883,N_14853,N_10305);
or U29884 (N_29884,N_18856,N_14908);
or U29885 (N_29885,N_19797,N_17342);
nand U29886 (N_29886,N_16354,N_16892);
and U29887 (N_29887,N_18516,N_15503);
or U29888 (N_29888,N_15842,N_11281);
nand U29889 (N_29889,N_15039,N_17009);
or U29890 (N_29890,N_19767,N_15162);
or U29891 (N_29891,N_13431,N_15741);
nor U29892 (N_29892,N_15218,N_17379);
and U29893 (N_29893,N_13902,N_17041);
xor U29894 (N_29894,N_16639,N_16701);
nand U29895 (N_29895,N_15016,N_16931);
and U29896 (N_29896,N_14980,N_18004);
and U29897 (N_29897,N_18260,N_12646);
nand U29898 (N_29898,N_19984,N_17273);
nand U29899 (N_29899,N_14211,N_10665);
or U29900 (N_29900,N_18424,N_19667);
and U29901 (N_29901,N_15670,N_16965);
or U29902 (N_29902,N_18996,N_15356);
nor U29903 (N_29903,N_14304,N_19612);
nand U29904 (N_29904,N_18692,N_18148);
or U29905 (N_29905,N_16167,N_17092);
and U29906 (N_29906,N_17523,N_11015);
nor U29907 (N_29907,N_10154,N_13620);
or U29908 (N_29908,N_11081,N_12424);
and U29909 (N_29909,N_11181,N_18231);
xor U29910 (N_29910,N_13488,N_10339);
nor U29911 (N_29911,N_15925,N_17445);
nand U29912 (N_29912,N_13842,N_15230);
xnor U29913 (N_29913,N_14907,N_10862);
xnor U29914 (N_29914,N_17129,N_14569);
xnor U29915 (N_29915,N_10719,N_16253);
or U29916 (N_29916,N_11723,N_17105);
nor U29917 (N_29917,N_15394,N_18398);
or U29918 (N_29918,N_11148,N_17316);
nand U29919 (N_29919,N_18316,N_16561);
nor U29920 (N_29920,N_12073,N_12449);
nor U29921 (N_29921,N_11028,N_14815);
or U29922 (N_29922,N_10949,N_18558);
nand U29923 (N_29923,N_13976,N_16260);
nor U29924 (N_29924,N_11077,N_18142);
nand U29925 (N_29925,N_19142,N_19430);
xnor U29926 (N_29926,N_12382,N_18138);
or U29927 (N_29927,N_14283,N_11334);
nor U29928 (N_29928,N_12664,N_14442);
nor U29929 (N_29929,N_13524,N_16614);
or U29930 (N_29930,N_11257,N_18339);
xnor U29931 (N_29931,N_15951,N_18901);
xnor U29932 (N_29932,N_15085,N_14211);
nor U29933 (N_29933,N_19234,N_12937);
xor U29934 (N_29934,N_18739,N_16414);
nand U29935 (N_29935,N_19775,N_15393);
nor U29936 (N_29936,N_16312,N_14789);
or U29937 (N_29937,N_13935,N_10546);
nand U29938 (N_29938,N_16218,N_12428);
xor U29939 (N_29939,N_17780,N_10965);
or U29940 (N_29940,N_13548,N_12160);
or U29941 (N_29941,N_11366,N_11281);
and U29942 (N_29942,N_15311,N_14637);
xnor U29943 (N_29943,N_12194,N_14966);
and U29944 (N_29944,N_17072,N_15992);
and U29945 (N_29945,N_13124,N_12027);
nand U29946 (N_29946,N_15364,N_11421);
or U29947 (N_29947,N_11366,N_16914);
and U29948 (N_29948,N_16783,N_12522);
and U29949 (N_29949,N_10688,N_16426);
and U29950 (N_29950,N_10481,N_17565);
nor U29951 (N_29951,N_11699,N_11703);
or U29952 (N_29952,N_10586,N_13071);
or U29953 (N_29953,N_16227,N_12422);
nand U29954 (N_29954,N_10861,N_14979);
nand U29955 (N_29955,N_14305,N_18261);
and U29956 (N_29956,N_14929,N_14390);
nor U29957 (N_29957,N_17340,N_19160);
nor U29958 (N_29958,N_10019,N_10605);
nand U29959 (N_29959,N_16885,N_14519);
or U29960 (N_29960,N_17163,N_15073);
or U29961 (N_29961,N_10807,N_11605);
nand U29962 (N_29962,N_16711,N_11074);
or U29963 (N_29963,N_10077,N_17187);
nand U29964 (N_29964,N_19490,N_10231);
and U29965 (N_29965,N_11013,N_13764);
and U29966 (N_29966,N_11375,N_19971);
nand U29967 (N_29967,N_16959,N_17382);
nor U29968 (N_29968,N_16879,N_11949);
nor U29969 (N_29969,N_15246,N_14710);
and U29970 (N_29970,N_16653,N_15371);
nand U29971 (N_29971,N_14987,N_19905);
nor U29972 (N_29972,N_18525,N_16050);
nand U29973 (N_29973,N_16529,N_19997);
and U29974 (N_29974,N_13205,N_13780);
and U29975 (N_29975,N_18038,N_18780);
and U29976 (N_29976,N_10122,N_11702);
or U29977 (N_29977,N_14836,N_19452);
and U29978 (N_29978,N_15737,N_19755);
and U29979 (N_29979,N_10255,N_17016);
nand U29980 (N_29980,N_16496,N_12931);
nor U29981 (N_29981,N_10135,N_13388);
nand U29982 (N_29982,N_17420,N_14903);
nor U29983 (N_29983,N_11195,N_10113);
or U29984 (N_29984,N_11614,N_19816);
nor U29985 (N_29985,N_19848,N_13233);
nor U29986 (N_29986,N_18126,N_10678);
nor U29987 (N_29987,N_16477,N_12408);
nand U29988 (N_29988,N_18101,N_18685);
and U29989 (N_29989,N_13319,N_19021);
or U29990 (N_29990,N_12515,N_15443);
and U29991 (N_29991,N_15372,N_18540);
nand U29992 (N_29992,N_12872,N_10871);
xnor U29993 (N_29993,N_11119,N_14268);
xor U29994 (N_29994,N_16958,N_16212);
xnor U29995 (N_29995,N_17989,N_17868);
xnor U29996 (N_29996,N_11451,N_17732);
nor U29997 (N_29997,N_11998,N_10762);
xor U29998 (N_29998,N_18851,N_16552);
nand U29999 (N_29999,N_15646,N_14940);
and UO_0 (O_0,N_26107,N_24293);
nand UO_1 (O_1,N_22871,N_29474);
nor UO_2 (O_2,N_21478,N_25368);
or UO_3 (O_3,N_26173,N_25754);
nand UO_4 (O_4,N_27605,N_26731);
or UO_5 (O_5,N_23459,N_24770);
or UO_6 (O_6,N_28663,N_21988);
and UO_7 (O_7,N_29163,N_24553);
nand UO_8 (O_8,N_22239,N_29964);
or UO_9 (O_9,N_21571,N_29411);
nor UO_10 (O_10,N_26405,N_26588);
or UO_11 (O_11,N_29462,N_29919);
or UO_12 (O_12,N_21687,N_28500);
nor UO_13 (O_13,N_26411,N_24581);
nor UO_14 (O_14,N_23263,N_27531);
or UO_15 (O_15,N_21313,N_27763);
nand UO_16 (O_16,N_23642,N_24592);
nor UO_17 (O_17,N_22024,N_24137);
nor UO_18 (O_18,N_27472,N_23118);
nand UO_19 (O_19,N_23984,N_27959);
nand UO_20 (O_20,N_22387,N_22579);
or UO_21 (O_21,N_25703,N_24507);
and UO_22 (O_22,N_21881,N_26468);
nor UO_23 (O_23,N_25071,N_26289);
or UO_24 (O_24,N_27366,N_25866);
and UO_25 (O_25,N_24971,N_22960);
nor UO_26 (O_26,N_28953,N_20859);
or UO_27 (O_27,N_27999,N_24746);
and UO_28 (O_28,N_23963,N_22134);
nand UO_29 (O_29,N_22536,N_27830);
or UO_30 (O_30,N_29172,N_29368);
nor UO_31 (O_31,N_21286,N_23374);
and UO_32 (O_32,N_23148,N_26524);
or UO_33 (O_33,N_28900,N_28177);
nor UO_34 (O_34,N_22009,N_29062);
nand UO_35 (O_35,N_22447,N_22659);
nor UO_36 (O_36,N_28085,N_23705);
nor UO_37 (O_37,N_28383,N_23946);
nor UO_38 (O_38,N_25561,N_20582);
or UO_39 (O_39,N_24346,N_22096);
nand UO_40 (O_40,N_25461,N_20598);
nor UO_41 (O_41,N_21936,N_22230);
and UO_42 (O_42,N_28939,N_28906);
or UO_43 (O_43,N_25138,N_29714);
nand UO_44 (O_44,N_23463,N_27945);
and UO_45 (O_45,N_20565,N_27343);
nor UO_46 (O_46,N_24183,N_20111);
nand UO_47 (O_47,N_27777,N_29820);
xor UO_48 (O_48,N_28898,N_22876);
and UO_49 (O_49,N_21346,N_29180);
nand UO_50 (O_50,N_22461,N_20971);
nand UO_51 (O_51,N_25521,N_20169);
nand UO_52 (O_52,N_29870,N_29115);
or UO_53 (O_53,N_23590,N_28676);
nor UO_54 (O_54,N_23874,N_29252);
xnor UO_55 (O_55,N_20611,N_22188);
xnor UO_56 (O_56,N_23494,N_29161);
nand UO_57 (O_57,N_20133,N_27938);
nand UO_58 (O_58,N_20746,N_21354);
and UO_59 (O_59,N_25331,N_26084);
nor UO_60 (O_60,N_24966,N_26057);
nand UO_61 (O_61,N_23959,N_22887);
and UO_62 (O_62,N_24376,N_29050);
nor UO_63 (O_63,N_22611,N_21087);
nor UO_64 (O_64,N_20455,N_27622);
nand UO_65 (O_65,N_22028,N_28076);
nand UO_66 (O_66,N_27878,N_23773);
or UO_67 (O_67,N_21444,N_27943);
and UO_68 (O_68,N_20340,N_24875);
nand UO_69 (O_69,N_23023,N_23681);
nand UO_70 (O_70,N_26056,N_29518);
or UO_71 (O_71,N_21254,N_27602);
nand UO_72 (O_72,N_24421,N_29405);
or UO_73 (O_73,N_23304,N_22768);
nand UO_74 (O_74,N_24445,N_27417);
and UO_75 (O_75,N_25335,N_23175);
and UO_76 (O_76,N_21797,N_29188);
or UO_77 (O_77,N_21191,N_29699);
xor UO_78 (O_78,N_20013,N_28783);
and UO_79 (O_79,N_27801,N_21579);
nor UO_80 (O_80,N_29196,N_26387);
and UO_81 (O_81,N_29855,N_23438);
nand UO_82 (O_82,N_24928,N_23534);
nor UO_83 (O_83,N_28265,N_23126);
and UO_84 (O_84,N_25601,N_23356);
nand UO_85 (O_85,N_27655,N_25574);
or UO_86 (O_86,N_21063,N_20538);
nand UO_87 (O_87,N_21641,N_24528);
and UO_88 (O_88,N_28253,N_29843);
and UO_89 (O_89,N_29361,N_23844);
nand UO_90 (O_90,N_22229,N_29294);
or UO_91 (O_91,N_23246,N_24378);
nand UO_92 (O_92,N_28461,N_28516);
xor UO_93 (O_93,N_29935,N_23317);
or UO_94 (O_94,N_25733,N_23911);
or UO_95 (O_95,N_21592,N_24814);
xor UO_96 (O_96,N_27312,N_24898);
and UO_97 (O_97,N_22026,N_23557);
and UO_98 (O_98,N_21074,N_24893);
nor UO_99 (O_99,N_25051,N_28107);
and UO_100 (O_100,N_20329,N_21955);
and UO_101 (O_101,N_29787,N_24843);
and UO_102 (O_102,N_21850,N_28689);
and UO_103 (O_103,N_24428,N_28029);
and UO_104 (O_104,N_23472,N_20448);
and UO_105 (O_105,N_21047,N_27058);
nor UO_106 (O_106,N_26479,N_26578);
nand UO_107 (O_107,N_25847,N_28039);
nand UO_108 (O_108,N_24361,N_24709);
and UO_109 (O_109,N_21075,N_21239);
xnor UO_110 (O_110,N_25549,N_28169);
nor UO_111 (O_111,N_20588,N_26043);
nand UO_112 (O_112,N_27235,N_23301);
and UO_113 (O_113,N_21767,N_25027);
nand UO_114 (O_114,N_26406,N_29463);
and UO_115 (O_115,N_25036,N_22295);
or UO_116 (O_116,N_27245,N_20862);
nor UO_117 (O_117,N_26424,N_26502);
nor UO_118 (O_118,N_21498,N_23528);
xnor UO_119 (O_119,N_22888,N_25390);
and UO_120 (O_120,N_24591,N_26817);
and UO_121 (O_121,N_26637,N_28140);
nor UO_122 (O_122,N_22300,N_24383);
xor UO_123 (O_123,N_23566,N_26865);
nand UO_124 (O_124,N_23955,N_25102);
or UO_125 (O_125,N_21602,N_29961);
nand UO_126 (O_126,N_26307,N_26660);
and UO_127 (O_127,N_23555,N_25179);
and UO_128 (O_128,N_23057,N_27179);
nor UO_129 (O_129,N_27671,N_27505);
or UO_130 (O_130,N_28644,N_26852);
xor UO_131 (O_131,N_23992,N_26400);
nand UO_132 (O_132,N_27126,N_28712);
xor UO_133 (O_133,N_20733,N_20550);
or UO_134 (O_134,N_21624,N_27285);
nand UO_135 (O_135,N_24233,N_26167);
nor UO_136 (O_136,N_26685,N_27786);
nor UO_137 (O_137,N_21553,N_28701);
nand UO_138 (O_138,N_24610,N_26415);
nor UO_139 (O_139,N_23303,N_20066);
or UO_140 (O_140,N_27627,N_27917);
nand UO_141 (O_141,N_22878,N_21344);
nand UO_142 (O_142,N_20210,N_24622);
or UO_143 (O_143,N_23313,N_23025);
or UO_144 (O_144,N_24640,N_22775);
nand UO_145 (O_145,N_23114,N_28459);
and UO_146 (O_146,N_20176,N_28010);
nand UO_147 (O_147,N_29493,N_23991);
and UO_148 (O_148,N_21860,N_21323);
and UO_149 (O_149,N_25202,N_24940);
nand UO_150 (O_150,N_23961,N_26977);
nor UO_151 (O_151,N_24853,N_26379);
or UO_152 (O_152,N_23347,N_27883);
nand UO_153 (O_153,N_26035,N_21422);
and UO_154 (O_154,N_21655,N_24290);
and UO_155 (O_155,N_29176,N_24391);
nand UO_156 (O_156,N_28601,N_24865);
nand UO_157 (O_157,N_27135,N_22151);
or UO_158 (O_158,N_24562,N_23189);
and UO_159 (O_159,N_27411,N_28470);
nor UO_160 (O_160,N_22110,N_23388);
and UO_161 (O_161,N_20316,N_26794);
or UO_162 (O_162,N_27708,N_28454);
nor UO_163 (O_163,N_25572,N_22748);
or UO_164 (O_164,N_27517,N_21015);
and UO_165 (O_165,N_23142,N_20090);
nor UO_166 (O_166,N_24094,N_29619);
or UO_167 (O_167,N_27132,N_28831);
and UO_168 (O_168,N_24168,N_20843);
nand UO_169 (O_169,N_28674,N_24552);
nand UO_170 (O_170,N_24599,N_29721);
nor UO_171 (O_171,N_23503,N_20494);
and UO_172 (O_172,N_24969,N_27735);
and UO_173 (O_173,N_22422,N_24232);
nand UO_174 (O_174,N_28067,N_28003);
and UO_175 (O_175,N_28284,N_23651);
or UO_176 (O_176,N_24159,N_27566);
nand UO_177 (O_177,N_24309,N_23731);
nor UO_178 (O_178,N_28023,N_22388);
nor UO_179 (O_179,N_24054,N_24783);
nand UO_180 (O_180,N_25990,N_21798);
nand UO_181 (O_181,N_20955,N_21390);
nor UO_182 (O_182,N_23351,N_29974);
nor UO_183 (O_183,N_29969,N_23713);
or UO_184 (O_184,N_24896,N_24467);
nand UO_185 (O_185,N_22564,N_20374);
nor UO_186 (O_186,N_20431,N_23781);
and UO_187 (O_187,N_23353,N_29891);
or UO_188 (O_188,N_23738,N_28445);
and UO_189 (O_189,N_26220,N_26929);
xnor UO_190 (O_190,N_26197,N_27662);
nor UO_191 (O_191,N_22493,N_22515);
or UO_192 (O_192,N_25174,N_25756);
or UO_193 (O_193,N_28315,N_21493);
and UO_194 (O_194,N_25357,N_22732);
nand UO_195 (O_195,N_29972,N_26603);
or UO_196 (O_196,N_20154,N_21205);
and UO_197 (O_197,N_23149,N_24555);
nand UO_198 (O_198,N_25412,N_25736);
xor UO_199 (O_199,N_29984,N_25177);
xor UO_200 (O_200,N_24827,N_25049);
or UO_201 (O_201,N_27346,N_24460);
and UO_202 (O_202,N_23883,N_28804);
or UO_203 (O_203,N_24052,N_28343);
nand UO_204 (O_204,N_23450,N_20742);
or UO_205 (O_205,N_26887,N_24604);
or UO_206 (O_206,N_27975,N_29562);
or UO_207 (O_207,N_21227,N_22770);
nand UO_208 (O_208,N_29554,N_25951);
or UO_209 (O_209,N_29773,N_28020);
nor UO_210 (O_210,N_25158,N_27184);
or UO_211 (O_211,N_20098,N_22345);
or UO_212 (O_212,N_27008,N_29053);
and UO_213 (O_213,N_21653,N_24835);
nand UO_214 (O_214,N_29668,N_26932);
and UO_215 (O_215,N_22988,N_21685);
nand UO_216 (O_216,N_26413,N_23838);
nor UO_217 (O_217,N_20776,N_23646);
nor UO_218 (O_218,N_27757,N_25740);
and UO_219 (O_219,N_24164,N_25950);
nor UO_220 (O_220,N_28376,N_24509);
nor UO_221 (O_221,N_27133,N_27431);
or UO_222 (O_222,N_22218,N_23457);
nor UO_223 (O_223,N_20863,N_29996);
and UO_224 (O_224,N_20123,N_23306);
nor UO_225 (O_225,N_26276,N_25047);
or UO_226 (O_226,N_27846,N_20819);
and UO_227 (O_227,N_22806,N_20332);
nand UO_228 (O_228,N_24007,N_24485);
and UO_229 (O_229,N_27679,N_22513);
and UO_230 (O_230,N_24154,N_29929);
or UO_231 (O_231,N_27254,N_23093);
or UO_232 (O_232,N_29741,N_24613);
or UO_233 (O_233,N_23897,N_25594);
or UO_234 (O_234,N_28536,N_20422);
and UO_235 (O_235,N_24768,N_26873);
and UO_236 (O_236,N_27901,N_29846);
nor UO_237 (O_237,N_24093,N_28669);
nand UO_238 (O_238,N_29685,N_20314);
nor UO_239 (O_239,N_26708,N_27717);
nand UO_240 (O_240,N_23501,N_27150);
or UO_241 (O_241,N_21870,N_24654);
and UO_242 (O_242,N_22969,N_22546);
nor UO_243 (O_243,N_28219,N_22487);
or UO_244 (O_244,N_26678,N_26296);
xnor UO_245 (O_245,N_25189,N_26861);
or UO_246 (O_246,N_22642,N_23711);
nor UO_247 (O_247,N_28427,N_21795);
nand UO_248 (O_248,N_20773,N_28522);
nand UO_249 (O_249,N_25217,N_22533);
nor UO_250 (O_250,N_27116,N_23033);
and UO_251 (O_251,N_21186,N_26211);
nand UO_252 (O_252,N_28242,N_26571);
nand UO_253 (O_253,N_24988,N_26665);
or UO_254 (O_254,N_26349,N_28282);
nand UO_255 (O_255,N_27389,N_29234);
and UO_256 (O_256,N_27212,N_28204);
nand UO_257 (O_257,N_28263,N_25725);
or UO_258 (O_258,N_24194,N_27042);
nor UO_259 (O_259,N_24579,N_26357);
xor UO_260 (O_260,N_21983,N_29231);
nand UO_261 (O_261,N_22905,N_21089);
nor UO_262 (O_262,N_28374,N_22675);
and UO_263 (O_263,N_27654,N_28588);
nand UO_264 (O_264,N_21397,N_24250);
nand UO_265 (O_265,N_27643,N_27205);
nand UO_266 (O_266,N_28336,N_27140);
nor UO_267 (O_267,N_24689,N_22799);
or UO_268 (O_268,N_27282,N_27376);
nand UO_269 (O_269,N_26111,N_26554);
xor UO_270 (O_270,N_23725,N_27070);
nor UO_271 (O_271,N_20269,N_28303);
nand UO_272 (O_272,N_21891,N_26066);
nor UO_273 (O_273,N_25583,N_20673);
xnor UO_274 (O_274,N_28050,N_24515);
xnor UO_275 (O_275,N_24678,N_25713);
and UO_276 (O_276,N_21985,N_24932);
xor UO_277 (O_277,N_24994,N_29153);
nor UO_278 (O_278,N_20909,N_21182);
or UO_279 (O_279,N_28979,N_27762);
and UO_280 (O_280,N_20680,N_20998);
nor UO_281 (O_281,N_29697,N_29317);
nand UO_282 (O_282,N_20921,N_22179);
nor UO_283 (O_283,N_21359,N_27626);
xor UO_284 (O_284,N_21698,N_20001);
or UO_285 (O_285,N_24750,N_20871);
xnor UO_286 (O_286,N_23066,N_25487);
and UO_287 (O_287,N_23389,N_24894);
or UO_288 (O_288,N_22049,N_24112);
or UO_289 (O_289,N_28962,N_20032);
or UO_290 (O_290,N_29406,N_20814);
nand UO_291 (O_291,N_24518,N_27911);
and UO_292 (O_292,N_29858,N_28838);
xnor UO_293 (O_293,N_20250,N_22814);
nor UO_294 (O_294,N_28879,N_24602);
or UO_295 (O_295,N_26015,N_27395);
or UO_296 (O_296,N_21278,N_21011);
and UO_297 (O_297,N_24121,N_20046);
and UO_298 (O_298,N_26223,N_27853);
nor UO_299 (O_299,N_28069,N_29928);
nor UO_300 (O_300,N_29500,N_21805);
and UO_301 (O_301,N_25396,N_28869);
or UO_302 (O_302,N_29456,N_25037);
nand UO_303 (O_303,N_22130,N_26103);
nand UO_304 (O_304,N_22530,N_25527);
nor UO_305 (O_305,N_29922,N_20805);
nand UO_306 (O_306,N_25744,N_24379);
xnor UO_307 (O_307,N_24393,N_20913);
and UO_308 (O_308,N_29370,N_29949);
nand UO_309 (O_309,N_23538,N_23947);
and UO_310 (O_310,N_29340,N_23591);
nand UO_311 (O_311,N_23721,N_24645);
nor UO_312 (O_312,N_27737,N_29635);
nand UO_313 (O_313,N_20626,N_25118);
or UO_314 (O_314,N_26684,N_29383);
nand UO_315 (O_315,N_25826,N_23486);
and UO_316 (O_316,N_29558,N_20248);
or UO_317 (O_317,N_27418,N_26607);
xor UO_318 (O_318,N_24521,N_26694);
xor UO_319 (O_319,N_24976,N_21841);
nor UO_320 (O_320,N_23633,N_26585);
nand UO_321 (O_321,N_27991,N_21258);
and UO_322 (O_322,N_28326,N_21762);
nor UO_323 (O_323,N_27913,N_20362);
nor UO_324 (O_324,N_20305,N_29446);
and UO_325 (O_325,N_22901,N_22697);
and UO_326 (O_326,N_26958,N_29139);
xnor UO_327 (O_327,N_21546,N_29098);
or UO_328 (O_328,N_26631,N_27244);
and UO_329 (O_329,N_24899,N_28774);
or UO_330 (O_330,N_28785,N_20681);
and UO_331 (O_331,N_24696,N_21051);
nor UO_332 (O_332,N_29630,N_21532);
and UO_333 (O_333,N_22846,N_20902);
or UO_334 (O_334,N_23321,N_27903);
and UO_335 (O_335,N_20655,N_26813);
nand UO_336 (O_336,N_29519,N_22918);
and UO_337 (O_337,N_27102,N_26770);
or UO_338 (O_338,N_28892,N_27512);
nand UO_339 (O_339,N_27355,N_26425);
xnor UO_340 (O_340,N_21410,N_23007);
nor UO_341 (O_341,N_27894,N_21709);
and UO_342 (O_342,N_25290,N_21833);
nand UO_343 (O_343,N_24661,N_20472);
or UO_344 (O_344,N_29228,N_27380);
and UO_345 (O_345,N_27340,N_29162);
and UO_346 (O_346,N_29016,N_27297);
xor UO_347 (O_347,N_20286,N_23592);
nor UO_348 (O_348,N_22650,N_29142);
or UO_349 (O_349,N_24401,N_26615);
and UO_350 (O_350,N_23585,N_21459);
and UO_351 (O_351,N_29117,N_29344);
nand UO_352 (O_352,N_28727,N_26931);
or UO_353 (O_353,N_26561,N_20497);
and UO_354 (O_354,N_28197,N_23256);
nand UO_355 (O_355,N_21362,N_20864);
nand UO_356 (O_356,N_28566,N_22524);
or UO_357 (O_357,N_26267,N_20205);
or UO_358 (O_358,N_29695,N_25213);
nand UO_359 (O_359,N_25278,N_23858);
xor UO_360 (O_360,N_24425,N_21465);
and UO_361 (O_361,N_24717,N_22469);
nand UO_362 (O_362,N_29743,N_25885);
nor UO_363 (O_363,N_27902,N_20058);
nand UO_364 (O_364,N_26146,N_28686);
nand UO_365 (O_365,N_27549,N_20635);
and UO_366 (O_366,N_27251,N_26506);
and UO_367 (O_367,N_20504,N_25336);
nor UO_368 (O_368,N_22604,N_22115);
and UO_369 (O_369,N_29548,N_20558);
or UO_370 (O_370,N_28557,N_22303);
and UO_371 (O_371,N_22448,N_22754);
or UO_372 (O_372,N_20231,N_21490);
or UO_373 (O_373,N_25135,N_28255);
and UO_374 (O_374,N_20226,N_20424);
nand UO_375 (O_375,N_24813,N_28846);
and UO_376 (O_376,N_21462,N_28772);
and UO_377 (O_377,N_26516,N_26341);
or UO_378 (O_378,N_20643,N_29242);
and UO_379 (O_379,N_26291,N_28796);
nor UO_380 (O_380,N_28233,N_20170);
and UO_381 (O_381,N_27947,N_23782);
nor UO_382 (O_382,N_29782,N_21842);
or UO_383 (O_383,N_21432,N_29539);
xor UO_384 (O_384,N_21071,N_22165);
and UO_385 (O_385,N_22817,N_22571);
nand UO_386 (O_386,N_23582,N_20918);
nor UO_387 (O_387,N_24122,N_27397);
nor UO_388 (O_388,N_26201,N_27906);
xnor UO_389 (O_389,N_24432,N_22706);
nor UO_390 (O_390,N_25587,N_22607);
nand UO_391 (O_391,N_28867,N_28092);
and UO_392 (O_392,N_22951,N_28407);
and UO_393 (O_393,N_24506,N_29760);
xnor UO_394 (O_394,N_28043,N_26208);
and UO_395 (O_395,N_29097,N_22099);
nand UO_396 (O_396,N_21666,N_21965);
nand UO_397 (O_397,N_25356,N_28745);
nor UO_398 (O_398,N_23084,N_28604);
nand UO_399 (O_399,N_28697,N_29997);
or UO_400 (O_400,N_24979,N_25681);
nor UO_401 (O_401,N_21215,N_27681);
nor UO_402 (O_402,N_29193,N_20945);
or UO_403 (O_403,N_22037,N_24322);
and UO_404 (O_404,N_26001,N_21489);
nand UO_405 (O_405,N_20542,N_29573);
and UO_406 (O_406,N_26002,N_24484);
nand UO_407 (O_407,N_25663,N_29236);
and UO_408 (O_408,N_23371,N_24905);
or UO_409 (O_409,N_28858,N_27493);
nand UO_410 (O_410,N_22291,N_22109);
nand UO_411 (O_411,N_23045,N_25595);
nor UO_412 (O_412,N_23843,N_22298);
and UO_413 (O_413,N_25887,N_27394);
nor UO_414 (O_414,N_21406,N_29947);
and UO_415 (O_415,N_28593,N_22153);
nor UO_416 (O_416,N_21809,N_26414);
or UO_417 (O_417,N_22260,N_29037);
nor UO_418 (O_418,N_26740,N_21564);
or UO_419 (O_419,N_22522,N_21807);
nor UO_420 (O_420,N_20988,N_28024);
nor UO_421 (O_421,N_27214,N_26681);
nor UO_422 (O_422,N_28749,N_23678);
nand UO_423 (O_423,N_24152,N_26488);
and UO_424 (O_424,N_22600,N_29376);
nor UO_425 (O_425,N_21427,N_20320);
and UO_426 (O_426,N_26819,N_25645);
nand UO_427 (O_427,N_25706,N_27513);
nor UO_428 (O_428,N_20095,N_28058);
or UO_429 (O_429,N_21567,N_23153);
nand UO_430 (O_430,N_26947,N_29679);
and UO_431 (O_431,N_22972,N_25930);
and UO_432 (O_432,N_26616,N_25326);
nor UO_433 (O_433,N_22790,N_26150);
and UO_434 (O_434,N_25058,N_28853);
nand UO_435 (O_435,N_25072,N_25763);
and UO_436 (O_436,N_20406,N_24206);
nor UO_437 (O_437,N_20670,N_27667);
and UO_438 (O_438,N_25809,N_25545);
or UO_439 (O_439,N_25010,N_24160);
or UO_440 (O_440,N_25157,N_29826);
nand UO_441 (O_441,N_29149,N_28565);
or UO_442 (O_442,N_20729,N_24590);
and UO_443 (O_443,N_20115,N_26247);
nor UO_444 (O_444,N_22625,N_28080);
or UO_445 (O_445,N_25091,N_29305);
and UO_446 (O_446,N_24742,N_22082);
and UO_447 (O_447,N_20888,N_26364);
and UO_448 (O_448,N_23821,N_25526);
and UO_449 (O_449,N_28090,N_29588);
nand UO_450 (O_450,N_27561,N_28964);
nor UO_451 (O_451,N_26541,N_25710);
xnor UO_452 (O_452,N_28331,N_25178);
or UO_453 (O_453,N_24043,N_26936);
and UO_454 (O_454,N_25044,N_20545);
and UO_455 (O_455,N_26998,N_21606);
or UO_456 (O_456,N_22678,N_28532);
nor UO_457 (O_457,N_25244,N_22312);
nand UO_458 (O_458,N_28668,N_25610);
xnor UO_459 (O_459,N_29363,N_26657);
and UO_460 (O_460,N_21621,N_28424);
nand UO_461 (O_461,N_25176,N_22392);
nor UO_462 (O_462,N_26012,N_29219);
and UO_463 (O_463,N_23088,N_25730);
nor UO_464 (O_464,N_21552,N_23512);
and UO_465 (O_465,N_28030,N_21322);
nand UO_466 (O_466,N_22302,N_23030);
and UO_467 (O_467,N_23654,N_23701);
or UO_468 (O_468,N_22902,N_23842);
nand UO_469 (O_469,N_26097,N_21487);
xor UO_470 (O_470,N_21725,N_24086);
xor UO_471 (O_471,N_21578,N_21481);
and UO_472 (O_472,N_27769,N_28720);
nand UO_473 (O_473,N_25359,N_25657);
nand UO_474 (O_474,N_28885,N_25170);
nor UO_475 (O_475,N_27939,N_20136);
nand UO_476 (O_476,N_25766,N_22631);
nand UO_477 (O_477,N_23390,N_25555);
nand UO_478 (O_478,N_21178,N_27462);
or UO_479 (O_479,N_22480,N_26255);
and UO_480 (O_480,N_27748,N_21961);
xor UO_481 (O_481,N_24469,N_22764);
or UO_482 (O_482,N_22508,N_25022);
nand UO_483 (O_483,N_21442,N_25670);
xnor UO_484 (O_484,N_29624,N_26149);
and UO_485 (O_485,N_24849,N_29747);
and UO_486 (O_486,N_20941,N_26445);
nand UO_487 (O_487,N_24576,N_27159);
nor UO_488 (O_488,N_20311,N_20505);
nor UO_489 (O_489,N_22680,N_23466);
and UO_490 (O_490,N_22286,N_25862);
or UO_491 (O_491,N_29030,N_29621);
xor UO_492 (O_492,N_26126,N_21528);
nor UO_493 (O_493,N_22470,N_27555);
xnor UO_494 (O_494,N_28583,N_21598);
and UO_495 (O_495,N_23456,N_27071);
xor UO_496 (O_496,N_23914,N_24177);
or UO_497 (O_497,N_22358,N_29414);
nand UO_498 (O_498,N_28737,N_26741);
xor UO_499 (O_499,N_22145,N_21347);
nor UO_500 (O_500,N_21266,N_26353);
or UO_501 (O_501,N_20278,N_29878);
or UO_502 (O_502,N_20323,N_26920);
nand UO_503 (O_503,N_20200,N_28534);
nor UO_504 (O_504,N_23990,N_21557);
and UO_505 (O_505,N_28012,N_24762);
and UO_506 (O_506,N_23483,N_28175);
nor UO_507 (O_507,N_26964,N_21828);
nor UO_508 (O_508,N_20881,N_26017);
nand UO_509 (O_509,N_23630,N_28491);
nor UO_510 (O_510,N_29315,N_29703);
xnor UO_511 (O_511,N_27253,N_25120);
nor UO_512 (O_512,N_29479,N_25519);
or UO_513 (O_513,N_25287,N_25458);
and UO_514 (O_514,N_24626,N_21190);
nand UO_515 (O_515,N_22870,N_24221);
nand UO_516 (O_516,N_24105,N_25061);
and UO_517 (O_517,N_24657,N_27776);
or UO_518 (O_518,N_27303,N_24193);
nand UO_519 (O_519,N_22336,N_25949);
nand UO_520 (O_520,N_20232,N_23136);
nand UO_521 (O_521,N_21240,N_28834);
nand UO_522 (O_522,N_23146,N_25112);
or UO_523 (O_523,N_20844,N_28401);
and UO_524 (O_524,N_20801,N_26070);
and UO_525 (O_525,N_26980,N_25737);
nor UO_526 (O_526,N_29642,N_24439);
nor UO_527 (O_527,N_21907,N_26923);
or UO_528 (O_528,N_20656,N_23953);
or UO_529 (O_529,N_24572,N_26326);
nand UO_530 (O_530,N_23709,N_22190);
nor UO_531 (O_531,N_27379,N_29357);
and UO_532 (O_532,N_21591,N_24990);
or UO_533 (O_533,N_26855,N_27641);
nand UO_534 (O_534,N_21992,N_24731);
or UO_535 (O_535,N_26117,N_26297);
and UO_536 (O_536,N_26675,N_28444);
nor UO_537 (O_537,N_21932,N_29401);
xor UO_538 (O_538,N_22520,N_28009);
nand UO_539 (O_539,N_23794,N_21249);
and UO_540 (O_540,N_21315,N_21111);
nand UO_541 (O_541,N_21041,N_24323);
nand UO_542 (O_542,N_20457,N_20308);
and UO_543 (O_543,N_22360,N_25919);
nand UO_544 (O_544,N_20524,N_26841);
nand UO_545 (O_545,N_20996,N_23227);
xnor UO_546 (O_546,N_23212,N_23272);
nand UO_547 (O_547,N_25108,N_23169);
nand UO_548 (O_548,N_28488,N_24129);
nor UO_549 (O_549,N_20114,N_24303);
xnor UO_550 (O_550,N_23116,N_23765);
nor UO_551 (O_551,N_27115,N_22417);
and UO_552 (O_552,N_27004,N_22877);
xnor UO_553 (O_553,N_22002,N_29890);
and UO_554 (O_554,N_28591,N_28648);
nor UO_555 (O_555,N_22630,N_27577);
xnor UO_556 (O_556,N_29689,N_26672);
and UO_557 (O_557,N_20031,N_20573);
or UO_558 (O_558,N_24695,N_29329);
and UO_559 (O_559,N_28104,N_26369);
nor UO_560 (O_560,N_20694,N_28116);
and UO_561 (O_561,N_24146,N_25160);
nor UO_562 (O_562,N_27357,N_28456);
and UO_563 (O_563,N_29122,N_24385);
nand UO_564 (O_564,N_26367,N_20521);
nor UO_565 (O_565,N_26441,N_29603);
and UO_566 (O_566,N_24329,N_26181);
nor UO_567 (O_567,N_22069,N_28258);
nor UO_568 (O_568,N_23972,N_23158);
or UO_569 (O_569,N_28753,N_26788);
nor UO_570 (O_570,N_21729,N_28695);
or UO_571 (O_571,N_26751,N_21233);
and UO_572 (O_572,N_28943,N_22328);
and UO_573 (O_573,N_24575,N_27600);
and UO_574 (O_574,N_27572,N_23832);
nand UO_575 (O_575,N_29508,N_29048);
nor UO_576 (O_576,N_21456,N_20936);
nor UO_577 (O_577,N_22735,N_26839);
nor UO_578 (O_578,N_27078,N_24118);
and UO_579 (O_579,N_25499,N_25580);
nand UO_580 (O_580,N_25739,N_28447);
and UO_581 (O_581,N_21863,N_27713);
or UO_582 (O_582,N_28888,N_27588);
and UO_583 (O_583,N_26921,N_22289);
and UO_584 (O_584,N_24204,N_24627);
xor UO_585 (O_585,N_24065,N_23194);
nor UO_586 (O_586,N_25232,N_21674);
and UO_587 (O_587,N_28716,N_29765);
nand UO_588 (O_588,N_22350,N_28997);
and UO_589 (O_589,N_20107,N_24948);
or UO_590 (O_590,N_26328,N_27112);
xnor UO_591 (O_591,N_27226,N_28742);
xor UO_592 (O_592,N_22999,N_23589);
and UO_593 (O_593,N_27305,N_26040);
xnor UO_594 (O_594,N_23100,N_20360);
or UO_595 (O_595,N_25655,N_29672);
or UO_596 (O_596,N_24114,N_26919);
or UO_597 (O_597,N_21689,N_24733);
or UO_598 (O_598,N_25283,N_25789);
nand UO_599 (O_599,N_22976,N_21980);
or UO_600 (O_600,N_26895,N_21825);
nand UO_601 (O_601,N_25258,N_24808);
and UO_602 (O_602,N_21670,N_23629);
nand UO_603 (O_603,N_23710,N_23516);
nand UO_604 (O_604,N_28539,N_25635);
or UO_605 (O_605,N_29019,N_22225);
or UO_606 (O_606,N_24842,N_25607);
or UO_607 (O_607,N_28118,N_28225);
and UO_608 (O_608,N_22994,N_24345);
nand UO_609 (O_609,N_27536,N_23739);
or UO_610 (O_610,N_20659,N_22504);
nor UO_611 (O_611,N_25184,N_23597);
or UO_612 (O_612,N_21915,N_25531);
nand UO_613 (O_613,N_20958,N_20564);
nor UO_614 (O_614,N_24855,N_24652);
or UO_615 (O_615,N_25416,N_22811);
nand UO_616 (O_616,N_21873,N_26274);
and UO_617 (O_617,N_29484,N_25402);
or UO_618 (O_618,N_27817,N_28493);
and UO_619 (O_619,N_20962,N_27316);
nor UO_620 (O_620,N_22856,N_26950);
or UO_621 (O_621,N_20830,N_29303);
nand UO_622 (O_622,N_21811,N_20999);
and UO_623 (O_623,N_26240,N_26707);
nor UO_624 (O_624,N_22468,N_29136);
xnor UO_625 (O_625,N_21683,N_23508);
or UO_626 (O_626,N_27647,N_22597);
or UO_627 (O_627,N_24777,N_22281);
nor UO_628 (O_628,N_22462,N_20185);
nor UO_629 (O_629,N_24880,N_25362);
and UO_630 (O_630,N_29107,N_29164);
nand UO_631 (O_631,N_20744,N_22052);
xnor UO_632 (O_632,N_23117,N_29031);
nor UO_633 (O_633,N_27217,N_24254);
nor UO_634 (O_634,N_27401,N_26500);
and UO_635 (O_635,N_21435,N_20914);
nor UO_636 (O_636,N_25796,N_29485);
and UO_637 (O_637,N_21010,N_23915);
xnor UO_638 (O_638,N_25050,N_25528);
nor UO_639 (O_639,N_28385,N_26799);
and UO_640 (O_640,N_22534,N_22047);
xor UO_641 (O_641,N_27542,N_23319);
nor UO_642 (O_642,N_25182,N_28497);
and UO_643 (O_643,N_25475,N_20810);
nand UO_644 (O_644,N_25849,N_29475);
nor UO_645 (O_645,N_26995,N_20097);
nor UO_646 (O_646,N_28054,N_22752);
or UO_647 (O_647,N_23541,N_29937);
nand UO_648 (O_648,N_23124,N_22700);
nor UO_649 (O_649,N_24530,N_26044);
nand UO_650 (O_650,N_25541,N_22416);
xnor UO_651 (O_651,N_26654,N_24660);
nand UO_652 (O_652,N_24143,N_27501);
and UO_653 (O_653,N_22689,N_25448);
and UO_654 (O_654,N_27031,N_24027);
nand UO_655 (O_655,N_20212,N_23537);
nor UO_656 (O_656,N_29124,N_20930);
nor UO_657 (O_657,N_28037,N_27359);
xnor UO_658 (O_658,N_27367,N_24815);
nand UO_659 (O_659,N_27231,N_27569);
nand UO_660 (O_660,N_24534,N_21389);
nor UO_661 (O_661,N_29780,N_24596);
or UO_662 (O_662,N_22653,N_25620);
and UO_663 (O_663,N_24051,N_23465);
xor UO_664 (O_664,N_21243,N_28517);
nand UO_665 (O_665,N_20462,N_21309);
nand UO_666 (O_666,N_26714,N_28670);
and UO_667 (O_667,N_20004,N_29786);
nor UO_668 (O_668,N_24897,N_24266);
nor UO_669 (O_669,N_29589,N_22760);
nor UO_670 (O_670,N_25409,N_21402);
or UO_671 (O_671,N_27994,N_22429);
nand UO_672 (O_672,N_22124,N_26090);
and UO_673 (O_673,N_23565,N_27683);
and UO_674 (O_674,N_24687,N_22593);
nand UO_675 (O_675,N_28525,N_23853);
or UO_676 (O_676,N_20857,N_23443);
nor UO_677 (O_677,N_28211,N_26469);
and UO_678 (O_678,N_20400,N_22418);
xnor UO_679 (O_679,N_25612,N_26354);
nand UO_680 (O_680,N_25103,N_26582);
and UO_681 (O_681,N_21211,N_26658);
nor UO_682 (O_682,N_27839,N_22712);
and UO_683 (O_683,N_23147,N_29837);
nand UO_684 (O_684,N_27117,N_27870);
xnor UO_685 (O_685,N_20866,N_21361);
or UO_686 (O_686,N_20042,N_28923);
xor UO_687 (O_687,N_20041,N_27318);
and UO_688 (O_688,N_24965,N_20957);
and UO_689 (O_689,N_27034,N_22326);
or UO_690 (O_690,N_21281,N_29884);
xnor UO_691 (O_691,N_28847,N_24357);
or UO_692 (O_692,N_24840,N_21576);
nand UO_693 (O_693,N_20233,N_26937);
nor UO_694 (O_694,N_27241,N_20282);
or UO_695 (O_695,N_27097,N_23498);
or UO_696 (O_696,N_27611,N_24045);
nor UO_697 (O_697,N_23650,N_21536);
nand UO_698 (O_698,N_29260,N_23619);
and UO_699 (O_699,N_21993,N_20633);
nand UO_700 (O_700,N_21492,N_25679);
or UO_701 (O_701,N_25026,N_25300);
or UO_702 (O_702,N_20561,N_24109);
nand UO_703 (O_703,N_29407,N_23288);
or UO_704 (O_704,N_29254,N_24917);
or UO_705 (O_705,N_20932,N_29960);
xnor UO_706 (O_706,N_29904,N_23477);
nor UO_707 (O_707,N_24273,N_24310);
and UO_708 (O_708,N_22354,N_29111);
nand UO_709 (O_709,N_21069,N_22914);
nor UO_710 (O_710,N_24725,N_29267);
nor UO_711 (O_711,N_20087,N_22139);
xnor UO_712 (O_712,N_25195,N_29976);
nor UO_713 (O_713,N_25097,N_29087);
nand UO_714 (O_714,N_29585,N_23395);
and UO_715 (O_715,N_21953,N_20034);
or UO_716 (O_716,N_21469,N_28325);
and UO_717 (O_717,N_24113,N_22103);
or UO_718 (O_718,N_29223,N_21803);
and UO_719 (O_719,N_23223,N_26161);
or UO_720 (O_720,N_20823,N_27040);
nor UO_721 (O_721,N_28227,N_24088);
and UO_722 (O_722,N_29885,N_21539);
nor UO_723 (O_723,N_27745,N_22922);
nand UO_724 (O_724,N_24062,N_28934);
xor UO_725 (O_725,N_23644,N_24058);
or UO_726 (O_726,N_25812,N_27729);
nand UO_727 (O_727,N_27773,N_21800);
xor UO_728 (O_728,N_20021,N_27405);
and UO_729 (O_729,N_21701,N_28222);
and UO_730 (O_730,N_23283,N_24745);
nor UO_731 (O_731,N_24718,N_21381);
nand UO_732 (O_732,N_22247,N_25738);
or UO_733 (O_733,N_27584,N_24487);
or UO_734 (O_734,N_27966,N_26471);
nor UO_735 (O_735,N_23890,N_29596);
nor UO_736 (O_736,N_28283,N_28344);
nand UO_737 (O_737,N_21950,N_21008);
and UO_738 (O_738,N_22849,N_21061);
and UO_739 (O_739,N_20893,N_23808);
and UO_740 (O_740,N_23325,N_22222);
nor UO_741 (O_741,N_27852,N_25523);
and UO_742 (O_742,N_28631,N_26184);
and UO_743 (O_743,N_26885,N_26147);
nand UO_744 (O_744,N_24796,N_23723);
nand UO_745 (O_745,N_24402,N_26403);
nand UO_746 (O_746,N_24205,N_29032);
or UO_747 (O_747,N_20488,N_24798);
nor UO_748 (O_748,N_24153,N_23692);
or UO_749 (O_749,N_21196,N_24225);
nand UO_750 (O_750,N_21816,N_24671);
or UO_751 (O_751,N_23815,N_26851);
nand UO_752 (O_752,N_25391,N_28224);
nor UO_753 (O_753,N_25935,N_20217);
or UO_754 (O_754,N_20162,N_24336);
nor UO_755 (O_755,N_23468,N_25619);
or UO_756 (O_756,N_23933,N_26670);
or UO_757 (O_757,N_27436,N_29502);
or UO_758 (O_758,N_28684,N_25654);
or UO_759 (O_759,N_24751,N_22851);
or UO_760 (O_760,N_27292,N_29594);
and UO_761 (O_761,N_28157,N_25508);
or UO_762 (O_762,N_25857,N_29191);
or UO_763 (O_763,N_20089,N_24819);
and UO_764 (O_764,N_28238,N_24307);
xor UO_765 (O_765,N_21236,N_22926);
or UO_766 (O_766,N_28795,N_24806);
nand UO_767 (O_767,N_22080,N_21457);
nand UO_768 (O_768,N_20403,N_22989);
nand UO_769 (O_769,N_26483,N_29517);
nor UO_770 (O_770,N_29209,N_24501);
and UO_771 (O_771,N_29473,N_23674);
and UO_772 (O_772,N_29749,N_27232);
nor UO_773 (O_773,N_29195,N_28519);
nand UO_774 (O_774,N_22051,N_21844);
and UO_775 (O_775,N_26597,N_20622);
or UO_776 (O_776,N_22828,N_22125);
nand UO_777 (O_777,N_22968,N_20458);
nor UO_778 (O_778,N_28764,N_20533);
nand UO_779 (O_779,N_20092,N_25239);
or UO_780 (O_780,N_20085,N_24003);
nand UO_781 (O_781,N_28971,N_28108);
or UO_782 (O_782,N_26832,N_27836);
nand UO_783 (O_783,N_22471,N_28622);
or UO_784 (O_784,N_26372,N_29505);
xor UO_785 (O_785,N_20731,N_22646);
nand UO_786 (O_786,N_26437,N_27813);
and UO_787 (O_787,N_20997,N_20043);
and UO_788 (O_788,N_27326,N_28339);
nor UO_789 (O_789,N_29616,N_29450);
and UO_790 (O_790,N_25879,N_25059);
and UO_791 (O_791,N_26257,N_25197);
or UO_792 (O_792,N_25484,N_29975);
nor UO_793 (O_793,N_21073,N_24429);
and UO_794 (O_794,N_24395,N_26628);
or UO_795 (O_795,N_22170,N_29512);
or UO_796 (O_796,N_22331,N_27384);
xnor UO_797 (O_797,N_20350,N_25711);
or UO_798 (O_798,N_27541,N_21981);
and UO_799 (O_799,N_24333,N_24406);
and UO_800 (O_800,N_21219,N_21255);
nor UO_801 (O_801,N_26775,N_23847);
or UO_802 (O_802,N_29182,N_20952);
or UO_803 (O_803,N_23574,N_20771);
or UO_804 (O_804,N_21398,N_23975);
nand UO_805 (O_805,N_23595,N_24851);
nor UO_806 (O_806,N_27344,N_23003);
nand UO_807 (O_807,N_25693,N_27222);
and UO_808 (O_808,N_29873,N_20865);
nand UO_809 (O_809,N_26762,N_24715);
nand UO_810 (O_810,N_21209,N_22150);
nor UO_811 (O_811,N_27506,N_25551);
or UO_812 (O_812,N_20758,N_27272);
xor UO_813 (O_813,N_22017,N_29348);
nor UO_814 (O_814,N_25734,N_27791);
and UO_815 (O_815,N_20453,N_20723);
or UO_816 (O_816,N_20597,N_24292);
nor UO_817 (O_817,N_22305,N_26774);
nand UO_818 (O_818,N_28773,N_21118);
and UO_819 (O_819,N_26722,N_29279);
nand UO_820 (O_820,N_24340,N_21352);
nor UO_821 (O_821,N_24244,N_20601);
and UO_822 (O_822,N_26848,N_24187);
nand UO_823 (O_823,N_26390,N_28802);
xnor UO_824 (O_824,N_28335,N_29150);
or UO_825 (O_825,N_25110,N_27993);
nand UO_826 (O_826,N_21386,N_25131);
nor UO_827 (O_827,N_24190,N_26933);
or UO_828 (O_828,N_22815,N_28205);
nand UO_829 (O_829,N_29039,N_20426);
and UO_830 (O_830,N_27752,N_27686);
nand UO_831 (O_831,N_23499,N_25637);
and UO_832 (O_832,N_23679,N_20238);
or UO_833 (O_833,N_21110,N_29690);
nor UO_834 (O_834,N_25716,N_24694);
and UO_835 (O_835,N_23187,N_28235);
and UO_836 (O_836,N_23011,N_25621);
nand UO_837 (O_837,N_26472,N_21078);
or UO_838 (O_838,N_27905,N_26399);
nand UO_839 (O_839,N_22774,N_26456);
nand UO_840 (O_840,N_22507,N_20848);
nor UO_841 (O_841,N_28635,N_28578);
xnor UO_842 (O_842,N_20832,N_20719);
xnor UO_843 (O_843,N_29864,N_21711);
and UO_844 (O_844,N_25969,N_22979);
nand UO_845 (O_845,N_29116,N_27747);
nor UO_846 (O_846,N_27551,N_29764);
nor UO_847 (O_847,N_20356,N_24539);
and UO_848 (O_848,N_23892,N_26221);
nor UO_849 (O_849,N_25085,N_24264);
xnor UO_850 (O_850,N_27682,N_26736);
and UO_851 (O_851,N_26109,N_27891);
nor UO_852 (O_852,N_26960,N_28174);
or UO_853 (O_853,N_24703,N_20926);
nor UO_854 (O_854,N_20140,N_25004);
and UO_855 (O_855,N_28696,N_22085);
nor UO_856 (O_856,N_23594,N_24120);
nand UO_857 (O_857,N_23816,N_21697);
nor UO_858 (O_858,N_23790,N_24211);
nor UO_859 (O_859,N_20718,N_22692);
and UO_860 (O_860,N_27940,N_23097);
nand UO_861 (O_861,N_26230,N_24356);
or UO_862 (O_862,N_28439,N_24235);
nand UO_863 (O_863,N_29882,N_26099);
nor UO_864 (O_864,N_26941,N_23962);
nor UO_865 (O_865,N_27915,N_21785);
nor UO_866 (O_866,N_25094,N_23604);
and UO_867 (O_867,N_28597,N_22670);
and UO_868 (O_868,N_26018,N_24584);
nor UO_869 (O_869,N_25425,N_26983);
nand UO_870 (O_870,N_29666,N_29090);
nand UO_871 (O_871,N_27141,N_27522);
and UO_872 (O_872,N_27562,N_26375);
and UO_873 (O_873,N_28504,N_28932);
nand UO_874 (O_874,N_22798,N_26309);
nand UO_875 (O_875,N_20906,N_26930);
nor UO_876 (O_876,N_23180,N_20346);
nand UO_877 (O_877,N_27822,N_23755);
nand UO_878 (O_878,N_27617,N_28495);
or UO_879 (O_879,N_24741,N_24918);
nor UO_880 (O_880,N_28630,N_28931);
nor UO_881 (O_881,N_26648,N_25310);
nand UO_882 (O_882,N_27778,N_25342);
and UO_883 (O_883,N_28678,N_24227);
nand UO_884 (O_884,N_21941,N_22282);
nor UO_885 (O_885,N_20847,N_24646);
xnor UO_886 (O_886,N_22961,N_25084);
or UO_887 (O_887,N_26259,N_21140);
nor UO_888 (O_888,N_26574,N_23047);
nor UO_889 (O_889,N_27125,N_24107);
nand UO_890 (O_890,N_21512,N_21142);
or UO_891 (O_891,N_28158,N_26519);
nor UO_892 (O_892,N_26778,N_24556);
nor UO_893 (O_893,N_23683,N_24066);
nor UO_894 (O_894,N_29394,N_21911);
nand UO_895 (O_895,N_28976,N_26130);
and UO_896 (O_896,N_23602,N_23835);
nor UO_897 (O_897,N_23458,N_29024);
nor UO_898 (O_898,N_20427,N_24423);
xor UO_899 (O_899,N_26677,N_26689);
nand UO_900 (O_900,N_28702,N_27702);
nor UO_901 (O_901,N_26939,N_29877);
nand UO_902 (O_902,N_25973,N_24669);
or UO_903 (O_903,N_24504,N_22545);
or UO_904 (O_904,N_25633,N_26888);
or UO_905 (O_905,N_20619,N_28217);
or UO_906 (O_906,N_23840,N_26460);
nand UO_907 (O_907,N_23228,N_27515);
nor UO_908 (O_908,N_21802,N_28342);
or UO_909 (O_909,N_23247,N_23487);
and UO_910 (O_910,N_24267,N_26767);
or UO_911 (O_911,N_29566,N_21148);
or UO_912 (O_912,N_27821,N_26434);
and UO_913 (O_913,N_20509,N_29134);
or UO_914 (O_914,N_29145,N_26725);
or UO_915 (O_915,N_21770,N_25345);
nor UO_916 (O_916,N_28918,N_20082);
and UO_917 (O_917,N_24906,N_21101);
and UO_918 (O_918,N_22996,N_22269);
or UO_919 (O_919,N_22261,N_28546);
or UO_920 (O_920,N_23139,N_29409);
and UO_921 (O_921,N_26567,N_23479);
or UO_922 (O_922,N_20118,N_20748);
and UO_923 (O_923,N_24970,N_26508);
nor UO_924 (O_924,N_21784,N_22568);
nand UO_925 (O_925,N_20782,N_22813);
xnor UO_926 (O_926,N_20500,N_20772);
nand UO_927 (O_927,N_20954,N_20256);
and UO_928 (O_928,N_25891,N_29268);
or UO_929 (O_929,N_20809,N_25579);
or UO_930 (O_930,N_27403,N_27468);
and UO_931 (O_931,N_20285,N_23653);
or UO_932 (O_932,N_26721,N_24436);
or UO_933 (O_933,N_22574,N_25971);
or UO_934 (O_934,N_28166,N_28647);
nand UO_935 (O_935,N_21105,N_22831);
nor UO_936 (O_936,N_27658,N_28129);
nor UO_937 (O_937,N_27332,N_20541);
nor UO_938 (O_938,N_25873,N_20125);
nor UO_939 (O_939,N_26872,N_27674);
or UO_940 (O_940,N_21971,N_25757);
and UO_941 (O_941,N_24480,N_24442);
and UO_942 (O_942,N_26729,N_29615);
and UO_943 (O_943,N_29841,N_25101);
nand UO_944 (O_944,N_24850,N_24838);
or UO_945 (O_945,N_23199,N_25125);
xor UO_946 (O_946,N_27443,N_24306);
nor UO_947 (O_947,N_25277,N_25443);
nand UO_948 (O_948,N_27167,N_26060);
xor UO_949 (O_949,N_23408,N_28105);
nor UO_950 (O_950,N_22057,N_23942);
xor UO_951 (O_951,N_27044,N_23060);
nand UO_952 (O_952,N_29444,N_22511);
nor UO_953 (O_953,N_23193,N_20479);
nand UO_954 (O_954,N_23488,N_26458);
or UO_955 (O_955,N_22402,N_21019);
or UO_956 (O_956,N_22561,N_27689);
or UO_957 (O_957,N_26287,N_23156);
nand UO_958 (O_958,N_21143,N_27457);
nor UO_959 (O_959,N_22081,N_23943);
nand UO_960 (O_960,N_22695,N_27614);
nor UO_961 (O_961,N_26065,N_27893);
xnor UO_962 (O_962,N_23005,N_25578);
nor UO_963 (O_963,N_25570,N_25772);
nor UO_964 (O_964,N_23409,N_23230);
nor UO_965 (O_965,N_24123,N_27884);
nand UO_966 (O_966,N_28094,N_24001);
and UO_967 (O_967,N_22256,N_22393);
or UO_968 (O_968,N_26419,N_28352);
nor UO_969 (O_969,N_26000,N_29670);
or UO_970 (O_970,N_20293,N_23793);
or UO_971 (O_971,N_26791,N_25001);
and UO_972 (O_972,N_29809,N_22895);
or UO_973 (O_973,N_21287,N_20969);
nand UO_974 (O_974,N_29571,N_26389);
and UO_975 (O_975,N_25916,N_23511);
nand UO_976 (O_976,N_24956,N_27345);
or UO_977 (O_977,N_27848,N_22737);
nor UO_978 (O_978,N_28089,N_20328);
nand UO_979 (O_979,N_27624,N_25205);
or UO_980 (O_980,N_23208,N_29157);
and UO_981 (O_981,N_22537,N_20518);
xor UO_982 (O_982,N_22845,N_29448);
or UO_983 (O_983,N_25346,N_25000);
or UO_984 (O_984,N_29696,N_27151);
nand UO_985 (O_985,N_25628,N_29380);
and UO_986 (O_986,N_23111,N_21330);
and UO_987 (O_987,N_22086,N_26281);
nor UO_988 (O_988,N_24908,N_23020);
nand UO_989 (O_989,N_21060,N_21064);
nand UO_990 (O_990,N_28378,N_27172);
and UO_991 (O_991,N_27278,N_29871);
and UO_992 (O_992,N_23041,N_21238);
nor UO_993 (O_993,N_28787,N_22590);
and UO_994 (O_994,N_21145,N_23018);
nor UO_995 (O_995,N_29052,N_27725);
nand UO_996 (O_996,N_29273,N_29089);
and UO_997 (O_997,N_20587,N_27806);
xnor UO_998 (O_998,N_25136,N_29076);
nor UO_999 (O_999,N_25420,N_28758);
nand UO_1000 (O_1000,N_22213,N_22352);
and UO_1001 (O_1001,N_26433,N_21547);
or UO_1002 (O_1002,N_28201,N_29040);
nor UO_1003 (O_1003,N_24795,N_20077);
or UO_1004 (O_1004,N_28288,N_25151);
and UO_1005 (O_1005,N_23067,N_23201);
nor UO_1006 (O_1006,N_21162,N_25422);
and UO_1007 (O_1007,N_22473,N_21460);
or UO_1008 (O_1008,N_25662,N_27953);
nor UO_1009 (O_1009,N_21377,N_27781);
xnor UO_1010 (O_1010,N_20124,N_20956);
nand UO_1011 (O_1011,N_22011,N_22019);
or UO_1012 (O_1012,N_27038,N_27698);
nor UO_1013 (O_1013,N_26837,N_29437);
and UO_1014 (O_1014,N_24262,N_21813);
and UO_1015 (O_1015,N_21234,N_21780);
and UO_1016 (O_1016,N_24417,N_26655);
nand UO_1017 (O_1017,N_20753,N_29565);
nand UO_1018 (O_1018,N_23803,N_26343);
or UO_1019 (O_1019,N_25188,N_27833);
or UO_1020 (O_1020,N_27320,N_22992);
nor UO_1021 (O_1021,N_29568,N_28610);
or UO_1022 (O_1022,N_28819,N_26024);
nor UO_1023 (O_1023,N_21385,N_21304);
or UO_1024 (O_1024,N_27743,N_26165);
and UO_1025 (O_1025,N_25718,N_21664);
and UO_1026 (O_1026,N_27000,N_24279);
xnor UO_1027 (O_1027,N_23750,N_25701);
or UO_1028 (O_1028,N_28659,N_20732);
or UO_1029 (O_1029,N_23531,N_25867);
and UO_1030 (O_1030,N_27056,N_20761);
nand UO_1031 (O_1031,N_24202,N_24497);
nand UO_1032 (O_1032,N_26917,N_23172);
nor UO_1033 (O_1033,N_27061,N_29824);
or UO_1034 (O_1034,N_26860,N_20702);
nor UO_1035 (O_1035,N_20388,N_24440);
nor UO_1036 (O_1036,N_24135,N_26131);
and UO_1037 (O_1037,N_24077,N_21156);
and UO_1038 (O_1038,N_23042,N_26338);
and UO_1039 (O_1039,N_20152,N_23616);
or UO_1040 (O_1040,N_23936,N_28852);
and UO_1041 (O_1041,N_25584,N_27799);
or UO_1042 (O_1042,N_22532,N_21348);
nand UO_1043 (O_1043,N_23764,N_20836);
and UO_1044 (O_1044,N_22714,N_25721);
and UO_1045 (O_1045,N_27216,N_26031);
xor UO_1046 (O_1046,N_25841,N_26717);
or UO_1047 (O_1047,N_29026,N_29214);
xor UO_1048 (O_1048,N_21869,N_27337);
or UO_1049 (O_1049,N_24136,N_23530);
or UO_1050 (O_1050,N_28261,N_20228);
or UO_1051 (O_1051,N_23608,N_20589);
or UO_1052 (O_1052,N_25782,N_23393);
and UO_1053 (O_1053,N_26323,N_21338);
and UO_1054 (O_1054,N_21779,N_25810);
and UO_1055 (O_1055,N_22639,N_20009);
xnor UO_1056 (O_1056,N_23864,N_23647);
nand UO_1057 (O_1057,N_24603,N_28545);
and UO_1058 (O_1058,N_23717,N_20047);
and UO_1059 (O_1059,N_28778,N_23497);
and UO_1060 (O_1060,N_28081,N_28685);
and UO_1061 (O_1061,N_22494,N_29438);
and UO_1062 (O_1062,N_25005,N_24195);
and UO_1063 (O_1063,N_26112,N_21409);
or UO_1064 (O_1064,N_26713,N_29525);
nor UO_1065 (O_1065,N_24415,N_20641);
or UO_1066 (O_1066,N_25765,N_26674);
xor UO_1067 (O_1067,N_24859,N_29439);
nor UO_1068 (O_1068,N_23165,N_27545);
nand UO_1069 (O_1069,N_28395,N_22531);
nor UO_1070 (O_1070,N_22292,N_22991);
and UO_1071 (O_1071,N_28143,N_27864);
nand UO_1072 (O_1072,N_27302,N_22349);
nand UO_1073 (O_1073,N_22397,N_27556);
or UO_1074 (O_1074,N_26025,N_23880);
nor UO_1075 (O_1075,N_23248,N_22583);
nor UO_1076 (O_1076,N_27371,N_27630);
or UO_1077 (O_1077,N_24644,N_28220);
xor UO_1078 (O_1078,N_26611,N_27528);
nor UO_1079 (O_1079,N_22610,N_25618);
nor UO_1080 (O_1080,N_27459,N_21480);
nor UO_1081 (O_1081,N_25028,N_27433);
nor UO_1082 (O_1082,N_26752,N_26520);
or UO_1083 (O_1083,N_21045,N_25363);
xnor UO_1084 (O_1084,N_24420,N_22250);
nand UO_1085 (O_1085,N_23983,N_24833);
and UO_1086 (O_1086,N_29452,N_25495);
or UO_1087 (O_1087,N_29408,N_20148);
nor UO_1088 (O_1088,N_21994,N_20934);
nor UO_1089 (O_1089,N_20695,N_25626);
nand UO_1090 (O_1090,N_22198,N_24704);
nor UO_1091 (O_1091,N_25522,N_22053);
or UO_1092 (O_1092,N_20419,N_29712);
and UO_1093 (O_1093,N_25095,N_22788);
nand UO_1094 (O_1094,N_29477,N_23398);
nand UO_1095 (O_1095,N_25870,N_27489);
and UO_1096 (O_1096,N_22375,N_29639);
and UO_1097 (O_1097,N_27750,N_29158);
or UO_1098 (O_1098,N_26647,N_27492);
nor UO_1099 (O_1099,N_20334,N_24489);
nor UO_1100 (O_1100,N_29058,N_24268);
and UO_1101 (O_1101,N_29746,N_21968);
nor UO_1102 (O_1102,N_20236,N_20677);
or UO_1103 (O_1103,N_28942,N_27575);
and UO_1104 (O_1104,N_29626,N_24013);
or UO_1105 (O_1105,N_28538,N_25430);
and UO_1106 (O_1106,N_24836,N_23791);
or UO_1107 (O_1107,N_28132,N_20357);
and UO_1108 (O_1108,N_28193,N_21307);
nor UO_1109 (O_1109,N_24245,N_24433);
nand UO_1110 (O_1110,N_27197,N_26759);
nand UO_1111 (O_1111,N_23403,N_21270);
xnor UO_1112 (O_1112,N_28600,N_27919);
nor UO_1113 (O_1113,N_21188,N_26757);
and UO_1114 (O_1114,N_28981,N_22821);
and UO_1115 (O_1115,N_20781,N_28599);
or UO_1116 (O_1116,N_20951,N_24377);
nor UO_1117 (O_1117,N_23211,N_26234);
and UO_1118 (O_1118,N_25685,N_27956);
nor UO_1119 (O_1119,N_23415,N_20079);
or UO_1120 (O_1120,N_25275,N_27390);
nand UO_1121 (O_1121,N_27181,N_26892);
and UO_1122 (O_1122,N_27609,N_26693);
and UO_1123 (O_1123,N_26642,N_27009);
nand UO_1124 (O_1124,N_22757,N_20556);
nor UO_1125 (O_1125,N_29229,N_24830);
nand UO_1126 (O_1126,N_22592,N_22894);
and UO_1127 (O_1127,N_28929,N_25333);
or UO_1128 (O_1128,N_23806,N_22364);
nor UO_1129 (O_1129,N_22523,N_25052);
nand UO_1130 (O_1130,N_22407,N_28341);
xor UO_1131 (O_1131,N_27243,N_23397);
and UO_1132 (O_1132,N_21096,N_24559);
nand UO_1133 (O_1133,N_28462,N_28730);
nor UO_1134 (O_1134,N_22589,N_27741);
nor UO_1135 (O_1135,N_24400,N_20591);
xor UO_1136 (O_1136,N_26288,N_28607);
and UO_1137 (O_1137,N_28880,N_29154);
or UO_1138 (O_1138,N_29283,N_25907);
and UO_1139 (O_1139,N_26733,N_21001);
and UO_1140 (O_1140,N_25745,N_26308);
nand UO_1141 (O_1141,N_29569,N_27719);
or UO_1142 (O_1142,N_23584,N_20608);
nor UO_1143 (O_1143,N_29923,N_22636);
or UO_1144 (O_1144,N_24874,N_22394);
nand UO_1145 (O_1145,N_21617,N_25271);
and UO_1146 (O_1146,N_24101,N_29794);
and UO_1147 (O_1147,N_23026,N_24710);
and UO_1148 (O_1148,N_23504,N_21900);
and UO_1149 (O_1149,N_20186,N_27842);
or UO_1150 (O_1150,N_20491,N_21124);
nor UO_1151 (O_1151,N_20828,N_29807);
and UO_1152 (O_1152,N_29816,N_24490);
and UO_1153 (O_1153,N_27193,N_21171);
or UO_1154 (O_1154,N_27208,N_23121);
nor UO_1155 (O_1155,N_25525,N_25163);
nor UO_1156 (O_1156,N_24623,N_22785);
nand UO_1157 (O_1157,N_25921,N_21765);
nor UO_1158 (O_1158,N_29436,N_22320);
or UO_1159 (O_1159,N_23363,N_21099);
and UO_1160 (O_1160,N_28063,N_28814);
xnor UO_1161 (O_1161,N_28883,N_20149);
nand UO_1162 (O_1162,N_21159,N_21715);
nor UO_1163 (O_1163,N_25915,N_23523);
xor UO_1164 (O_1164,N_25735,N_28180);
nor UO_1165 (O_1165,N_26593,N_22444);
nand UO_1166 (O_1166,N_23960,N_28798);
nand UO_1167 (O_1167,N_25159,N_29341);
and UO_1168 (O_1168,N_28062,N_29610);
nor UO_1169 (O_1169,N_29489,N_20876);
nor UO_1170 (O_1170,N_20853,N_28734);
nor UO_1171 (O_1171,N_22656,N_21013);
or UO_1172 (O_1172,N_27325,N_25819);
nand UO_1173 (O_1173,N_25510,N_27645);
nand UO_1174 (O_1174,N_23945,N_29285);
and UO_1175 (O_1175,N_26264,N_21808);
nor UO_1176 (O_1176,N_24117,N_25132);
nand UO_1177 (O_1177,N_29766,N_21424);
or UO_1178 (O_1178,N_20413,N_24021);
nand UO_1179 (O_1179,N_24947,N_25354);
nor UO_1180 (O_1180,N_21091,N_23242);
nor UO_1181 (O_1181,N_26313,N_25424);
nand UO_1182 (O_1182,N_22844,N_20783);
nand UO_1183 (O_1183,N_28887,N_22936);
nor UO_1184 (O_1184,N_22353,N_27051);
nand UO_1185 (O_1185,N_23733,N_24275);
nor UO_1186 (O_1186,N_24951,N_29224);
nand UO_1187 (O_1187,N_26152,N_26037);
and UO_1188 (O_1188,N_23899,N_29166);
and UO_1189 (O_1189,N_24341,N_28055);
and UO_1190 (O_1190,N_27845,N_20821);
or UO_1191 (O_1191,N_25168,N_26371);
nand UO_1192 (O_1192,N_26183,N_24473);
nor UO_1193 (O_1193,N_27766,N_28621);
nor UO_1194 (O_1194,N_22141,N_25469);
or UO_1195 (O_1195,N_21501,N_28586);
xnor UO_1196 (O_1196,N_26253,N_23980);
or UO_1197 (O_1197,N_24611,N_27880);
xor UO_1198 (O_1198,N_22169,N_24456);
nor UO_1199 (O_1199,N_22665,N_23471);
nand UO_1200 (O_1200,N_23820,N_26719);
and UO_1201 (O_1201,N_22420,N_29068);
nor UO_1202 (O_1202,N_29486,N_26962);
or UO_1203 (O_1203,N_26049,N_23298);
nand UO_1204 (O_1204,N_21508,N_26342);
nor UO_1205 (O_1205,N_26540,N_21914);
or UO_1206 (O_1206,N_28982,N_27347);
nand UO_1207 (O_1207,N_20666,N_20110);
xor UO_1208 (O_1208,N_20933,N_24508);
nor UO_1209 (O_1209,N_26745,N_23266);
and UO_1210 (O_1210,N_26273,N_28388);
or UO_1211 (O_1211,N_27854,N_29723);
nor UO_1212 (O_1212,N_24413,N_20679);
nand UO_1213 (O_1213,N_20192,N_28337);
xor UO_1214 (O_1214,N_20576,N_29065);
or UO_1215 (O_1215,N_21678,N_22971);
nand UO_1216 (O_1216,N_20924,N_20908);
nand UO_1217 (O_1217,N_24597,N_21283);
nand UO_1218 (O_1218,N_28983,N_20172);
xor UO_1219 (O_1219,N_22904,N_28809);
or UO_1220 (O_1220,N_28627,N_28891);
nor UO_1221 (O_1221,N_24952,N_20751);
or UO_1222 (O_1222,N_20532,N_23159);
and UO_1223 (O_1223,N_22254,N_24252);
and UO_1224 (O_1224,N_28301,N_26748);
nand UO_1225 (O_1225,N_25544,N_24587);
or UO_1226 (O_1226,N_23763,N_28747);
xnor UO_1227 (O_1227,N_28392,N_26638);
nand UO_1228 (O_1228,N_26595,N_20020);
nor UO_1229 (O_1229,N_23150,N_21082);
or UO_1230 (O_1230,N_28944,N_26312);
nand UO_1231 (O_1231,N_23405,N_29034);
and UO_1232 (O_1232,N_27548,N_29379);
nand UO_1233 (O_1233,N_23378,N_20414);
nor UO_1234 (O_1234,N_26692,N_24009);
nor UO_1235 (O_1235,N_20964,N_22014);
or UO_1236 (O_1236,N_23596,N_25967);
or UO_1237 (O_1237,N_24902,N_29347);
and UO_1238 (O_1238,N_20786,N_25581);
and UO_1239 (O_1239,N_20104,N_27452);
nor UO_1240 (O_1240,N_23807,N_26753);
xor UO_1241 (O_1241,N_24320,N_21684);
xnor UO_1242 (O_1242,N_22959,N_27524);
nand UO_1243 (O_1243,N_28324,N_29595);
and UO_1244 (O_1244,N_29168,N_27113);
nor UO_1245 (O_1245,N_27100,N_23324);
and UO_1246 (O_1246,N_25379,N_20173);
and UO_1247 (O_1247,N_20454,N_24422);
or UO_1248 (O_1248,N_23505,N_21335);
nor UO_1249 (O_1249,N_23893,N_25220);
and UO_1250 (O_1250,N_26034,N_28851);
nor UO_1251 (O_1251,N_24238,N_24359);
xnor UO_1252 (O_1252,N_21594,N_29722);
nand UO_1253 (O_1253,N_20061,N_27886);
nor UO_1254 (O_1254,N_27185,N_27413);
nor UO_1255 (O_1255,N_22481,N_27053);
and UO_1256 (O_1256,N_29278,N_23081);
nor UO_1257 (O_1257,N_29802,N_25046);
nand UO_1258 (O_1258,N_22465,N_21103);
or UO_1259 (O_1259,N_21497,N_25497);
xor UO_1260 (O_1260,N_27849,N_26360);
nand UO_1261 (O_1261,N_22803,N_26160);
and UO_1262 (O_1262,N_21288,N_28618);
nand UO_1263 (O_1263,N_28016,N_29141);
nor UO_1264 (O_1264,N_28434,N_22874);
xnor UO_1265 (O_1265,N_20965,N_25625);
nand UO_1266 (O_1266,N_21350,N_22497);
xor UO_1267 (O_1267,N_25650,N_25261);
xor UO_1268 (O_1268,N_26350,N_28498);
nor UO_1269 (O_1269,N_22661,N_21530);
or UO_1270 (O_1270,N_24166,N_20987);
nand UO_1271 (O_1271,N_24512,N_29324);
and UO_1272 (O_1272,N_27942,N_23358);
xor UO_1273 (O_1273,N_22759,N_22506);
and UO_1274 (O_1274,N_29143,N_26189);
or UO_1275 (O_1275,N_26282,N_26068);
nand UO_1276 (O_1276,N_27469,N_26537);
nand UO_1277 (O_1277,N_22747,N_22679);
nor UO_1278 (O_1278,N_27668,N_20692);
and UO_1279 (O_1279,N_25111,N_28285);
and UO_1280 (O_1280,N_23309,N_21294);
or UO_1281 (O_1281,N_20722,N_25223);
nand UO_1282 (O_1282,N_20911,N_28423);
nand UO_1283 (O_1283,N_29707,N_29353);
and UO_1284 (O_1284,N_20937,N_22251);
nand UO_1285 (O_1285,N_20726,N_21526);
and UO_1286 (O_1286,N_21251,N_25385);
nor UO_1287 (O_1287,N_29509,N_28347);
and UO_1288 (O_1288,N_29784,N_20204);
and UO_1289 (O_1289,N_23338,N_22867);
nand UO_1290 (O_1290,N_29869,N_20358);
and UO_1291 (O_1291,N_21610,N_25898);
or UO_1292 (O_1292,N_22542,N_28980);
nor UO_1293 (O_1293,N_27944,N_22424);
nor UO_1294 (O_1294,N_20604,N_26188);
and UO_1295 (O_1295,N_28786,N_21328);
nor UO_1296 (O_1296,N_25423,N_20385);
and UO_1297 (O_1297,N_24811,N_27107);
nand UO_1298 (O_1298,N_29790,N_23059);
nand UO_1299 (O_1299,N_28501,N_24989);
and UO_1300 (O_1300,N_29761,N_29515);
nand UO_1301 (O_1301,N_29128,N_25090);
nor UO_1302 (O_1302,N_26735,N_26594);
xor UO_1303 (O_1303,N_22476,N_22467);
and UO_1304 (O_1304,N_26901,N_20167);
xnor UO_1305 (O_1305,N_29968,N_20363);
and UO_1306 (O_1306,N_27646,N_28234);
and UO_1307 (O_1307,N_25939,N_21031);
or UO_1308 (O_1308,N_22720,N_29856);
and UO_1309 (O_1309,N_20685,N_26874);
nand UO_1310 (O_1310,N_24255,N_23618);
nor UO_1311 (O_1311,N_24825,N_24085);
nor UO_1312 (O_1312,N_20421,N_27152);
nand UO_1313 (O_1313,N_20706,N_29177);
or UO_1314 (O_1314,N_22217,N_22721);
nand UO_1315 (O_1315,N_20487,N_25494);
nor UO_1316 (O_1316,N_23928,N_27962);
xor UO_1317 (O_1317,N_23394,N_25934);
xor UO_1318 (O_1318,N_28231,N_28452);
nor UO_1319 (O_1319,N_21889,N_28229);
nand UO_1320 (O_1320,N_25421,N_22910);
and UO_1321 (O_1321,N_22935,N_20254);
or UO_1322 (O_1322,N_29318,N_26166);
xnor UO_1323 (O_1323,N_22056,N_25762);
nor UO_1324 (O_1324,N_28482,N_27215);
nand UO_1325 (O_1325,N_28548,N_23226);
nand UO_1326 (O_1326,N_20468,N_20445);
and UO_1327 (O_1327,N_23702,N_23016);
or UO_1328 (O_1328,N_27967,N_29836);
nor UO_1329 (O_1329,N_26327,N_21301);
nand UO_1330 (O_1330,N_25634,N_29197);
nor UO_1331 (O_1331,N_21719,N_25743);
nand UO_1332 (O_1332,N_27322,N_21723);
nor UO_1333 (O_1333,N_28995,N_27560);
and UO_1334 (O_1334,N_25651,N_27449);
and UO_1335 (O_1335,N_21721,N_25760);
nand UO_1336 (O_1336,N_26179,N_22705);
xnor UO_1337 (O_1337,N_27685,N_20271);
nand UO_1338 (O_1338,N_23178,N_29025);
nor UO_1339 (O_1339,N_20779,N_27356);
nand UO_1340 (O_1340,N_22731,N_21901);
and UO_1341 (O_1341,N_26806,N_21155);
nand UO_1342 (O_1342,N_27527,N_27733);
xor UO_1343 (O_1343,N_28605,N_28490);
or UO_1344 (O_1344,N_28875,N_26418);
nor UO_1345 (O_1345,N_20833,N_21036);
nand UO_1346 (O_1346,N_23952,N_25603);
and UO_1347 (O_1347,N_21413,N_20780);
xnor UO_1348 (O_1348,N_23740,N_20253);
nand UO_1349 (O_1349,N_26191,N_21017);
and UO_1350 (O_1350,N_24127,N_28380);
or UO_1351 (O_1351,N_21007,N_24614);
or UO_1352 (O_1352,N_24222,N_23006);
nand UO_1353 (O_1353,N_24258,N_21938);
nand UO_1354 (O_1354,N_29028,N_21416);
or UO_1355 (O_1355,N_29792,N_28743);
nand UO_1356 (O_1356,N_29326,N_25880);
nand UO_1357 (O_1357,N_26709,N_20463);
nor UO_1358 (O_1358,N_24780,N_27109);
nand UO_1359 (O_1359,N_22724,N_27896);
and UO_1360 (O_1360,N_22100,N_25234);
and UO_1361 (O_1361,N_23280,N_22567);
nand UO_1362 (O_1362,N_22236,N_27895);
or UO_1363 (O_1363,N_27730,N_23884);
nor UO_1364 (O_1364,N_27767,N_22539);
nand UO_1365 (O_1365,N_26795,N_28429);
nor UO_1366 (O_1366,N_25860,N_27204);
nand UO_1367 (O_1367,N_23275,N_27249);
nand UO_1368 (O_1368,N_26700,N_25161);
and UO_1369 (O_1369,N_27550,N_21995);
and UO_1370 (O_1370,N_29842,N_21764);
and UO_1371 (O_1371,N_23091,N_27073);
xnor UO_1372 (O_1372,N_27011,N_23906);
nor UO_1373 (O_1373,N_26206,N_21732);
nor UO_1374 (O_1374,N_29987,N_28681);
or UO_1375 (O_1375,N_24128,N_28993);
nor UO_1376 (O_1376,N_25478,N_21042);
nand UO_1377 (O_1377,N_23202,N_21650);
and UO_1378 (O_1378,N_29605,N_23185);
nor UO_1379 (O_1379,N_23873,N_29664);
and UO_1380 (O_1380,N_23110,N_29894);
and UO_1381 (O_1381,N_23168,N_20331);
and UO_1382 (O_1382,N_23525,N_22215);
nand UO_1383 (O_1383,N_23220,N_23968);
nand UO_1384 (O_1384,N_29832,N_25779);
nand UO_1385 (O_1385,N_28102,N_23424);
nand UO_1386 (O_1386,N_25431,N_26820);
and UO_1387 (O_1387,N_23070,N_26779);
nor UO_1388 (O_1388,N_23290,N_25035);
and UO_1389 (O_1389,N_28683,N_26330);
and UO_1390 (O_1390,N_23308,N_24561);
nor UO_1391 (O_1391,N_22645,N_28248);
and UO_1392 (O_1392,N_24447,N_29675);
nor UO_1393 (O_1393,N_25582,N_25427);
or UO_1394 (O_1394,N_23688,N_27219);
or UO_1395 (O_1395,N_23839,N_29652);
nor UO_1396 (O_1396,N_24938,N_24360);
and UO_1397 (O_1397,N_28933,N_24691);
or UO_1398 (O_1398,N_26376,N_20868);
and UO_1399 (O_1399,N_29102,N_24817);
nand UO_1400 (O_1400,N_20096,N_21749);
or UO_1401 (O_1401,N_27266,N_29175);
or UO_1402 (O_1402,N_26381,N_21886);
or UO_1403 (O_1403,N_26430,N_24708);
nor UO_1404 (O_1404,N_21366,N_21067);
and UO_1405 (O_1405,N_25720,N_21384);
nor UO_1406 (O_1406,N_20769,N_29010);
xor UO_1407 (O_1407,N_20580,N_24207);
nand UO_1408 (O_1408,N_29389,N_27236);
nor UO_1409 (O_1409,N_29421,N_22883);
and UO_1410 (O_1410,N_28182,N_23867);
nor UO_1411 (O_1411,N_27925,N_20275);
and UO_1412 (O_1412,N_20980,N_26059);
and UO_1413 (O_1413,N_25240,N_24674);
and UO_1414 (O_1414,N_24701,N_29332);
or UO_1415 (O_1415,N_23685,N_26092);
nand UO_1416 (O_1416,N_27727,N_28437);
nor UO_1417 (O_1417,N_28160,N_28713);
and UO_1418 (O_1418,N_23769,N_26485);
nor UO_1419 (O_1419,N_21479,N_20883);
and UO_1420 (O_1420,N_28328,N_28125);
nand UO_1421 (O_1421,N_21342,N_25286);
nand UO_1422 (O_1422,N_25613,N_20897);
and UO_1423 (O_1423,N_28820,N_26278);
nor UO_1424 (O_1424,N_22609,N_26536);
xnor UO_1425 (O_1425,N_23062,N_20973);
nor UO_1426 (O_1426,N_23077,N_24217);
xnor UO_1427 (O_1427,N_26318,N_27640);
nor UO_1428 (O_1428,N_25014,N_22740);
nor UO_1429 (O_1429,N_29617,N_22949);
and UO_1430 (O_1430,N_24716,N_25340);
or UO_1431 (O_1431,N_25802,N_29498);
or UO_1432 (O_1432,N_28741,N_21922);
and UO_1433 (O_1433,N_25235,N_26756);
or UO_1434 (O_1434,N_20372,N_25210);
and UO_1435 (O_1435,N_26581,N_29901);
nand UO_1436 (O_1436,N_21791,N_28321);
or UO_1437 (O_1437,N_29495,N_27756);
and UO_1438 (O_1438,N_23645,N_24807);
or UO_1439 (O_1439,N_24289,N_24324);
or UO_1440 (O_1440,N_21198,N_22196);
nor UO_1441 (O_1441,N_28334,N_21874);
nor UO_1442 (O_1442,N_20131,N_25133);
and UO_1443 (O_1443,N_25648,N_26750);
nor UO_1444 (O_1444,N_24020,N_28159);
or UO_1445 (O_1445,N_22729,N_26737);
xnor UO_1446 (O_1446,N_28127,N_28881);
and UO_1447 (O_1447,N_25683,N_22565);
and UO_1448 (O_1448,N_29004,N_21772);
nand UO_1449 (O_1449,N_20482,N_26509);
and UO_1450 (O_1450,N_22766,N_27625);
nor UO_1451 (O_1451,N_21748,N_20838);
and UO_1452 (O_1452,N_26209,N_23522);
nor UO_1453 (O_1453,N_24200,N_28430);
and UO_1454 (O_1454,N_28637,N_21123);
or UO_1455 (O_1455,N_21648,N_26720);
nand UO_1456 (O_1456,N_23216,N_20741);
nand UO_1457 (O_1457,N_20646,N_24739);
nor UO_1458 (O_1458,N_23542,N_24496);
nor UO_1459 (O_1459,N_28826,N_29649);
and UO_1460 (O_1460,N_21369,N_29750);
or UO_1461 (O_1461,N_24810,N_29788);
or UO_1462 (O_1462,N_21114,N_22226);
nand UO_1463 (O_1463,N_26224,N_21128);
xor UO_1464 (O_1464,N_23521,N_21599);
and UO_1465 (O_1465,N_28850,N_29282);
nand UO_1466 (O_1466,N_29713,N_28032);
or UO_1467 (O_1467,N_25428,N_28571);
xor UO_1468 (O_1468,N_23186,N_27829);
nor UO_1469 (O_1469,N_20103,N_20371);
nor UO_1470 (O_1470,N_22634,N_28789);
nor UO_1471 (O_1471,N_20016,N_29194);
or UO_1472 (O_1472,N_27754,N_23783);
nand UO_1473 (O_1473,N_27013,N_26207);
or UO_1474 (O_1474,N_22690,N_24409);
xor UO_1475 (O_1475,N_20563,N_22796);
xor UO_1476 (O_1476,N_29418,N_29185);
and UO_1477 (O_1477,N_21514,N_23320);
nor UO_1478 (O_1478,N_26336,N_27083);
xor UO_1479 (O_1479,N_21531,N_28874);
nand UO_1480 (O_1480,N_20808,N_21626);
nand UO_1481 (O_1481,N_20220,N_25251);
nand UO_1482 (O_1482,N_22745,N_21540);
and UO_1483 (O_1483,N_22483,N_23719);
or UO_1484 (O_1484,N_29783,N_26589);
nor UO_1485 (O_1485,N_26564,N_26683);
or UO_1486 (O_1486,N_28450,N_24111);
nor UO_1487 (O_1487,N_21274,N_20586);
and UO_1488 (O_1488,N_26083,N_28137);
and UO_1489 (O_1489,N_26551,N_27746);
nand UO_1490 (O_1490,N_23418,N_26724);
and UO_1491 (O_1491,N_29314,N_28040);
nand UO_1492 (O_1492,N_26286,N_29857);
nand UO_1493 (O_1493,N_25632,N_28988);
or UO_1494 (O_1494,N_25198,N_26549);
nor UO_1495 (O_1495,N_23535,N_20802);
nor UO_1496 (O_1496,N_28411,N_21401);
nor UO_1497 (O_1497,N_27525,N_27706);
nand UO_1498 (O_1498,N_24236,N_29420);
xor UO_1499 (O_1499,N_28139,N_27142);
or UO_1500 (O_1500,N_26755,N_28199);
nand UO_1501 (O_1501,N_25324,N_29426);
and UO_1502 (O_1502,N_22104,N_24162);
xnor UO_1503 (O_1503,N_21280,N_24856);
nand UO_1504 (O_1504,N_22135,N_24163);
or UO_1505 (O_1505,N_28736,N_25726);
nand UO_1506 (O_1506,N_29683,N_24925);
or UO_1507 (O_1507,N_24450,N_26644);
and UO_1508 (O_1508,N_24997,N_28658);
nand UO_1509 (O_1509,N_25291,N_28594);
or UO_1510 (O_1510,N_29205,N_27257);
nor UO_1511 (O_1511,N_26798,N_27889);
or UO_1512 (O_1512,N_23540,N_22857);
or UO_1513 (O_1513,N_24036,N_23857);
and UO_1514 (O_1514,N_25811,N_24583);
or UO_1515 (O_1515,N_21644,N_29226);
nor UO_1516 (O_1516,N_27793,N_23145);
xor UO_1517 (O_1517,N_20459,N_29216);
and UO_1518 (O_1518,N_23179,N_27327);
and UO_1519 (O_1519,N_25998,N_26159);
nand UO_1520 (O_1520,N_24463,N_23238);
and UO_1521 (O_1521,N_28950,N_28473);
and UO_1522 (O_1522,N_29284,N_25850);
xor UO_1523 (O_1523,N_28001,N_22699);
and UO_1524 (O_1524,N_27820,N_25859);
or UO_1525 (O_1525,N_25045,N_29943);
xor UO_1526 (O_1526,N_25914,N_27175);
nor UO_1527 (O_1527,N_28362,N_23727);
or UO_1528 (O_1528,N_26277,N_26227);
nor UO_1529 (O_1529,N_24863,N_29227);
and UO_1530 (O_1530,N_22673,N_20735);
or UO_1531 (O_1531,N_24769,N_27284);
or UO_1532 (O_1532,N_20763,N_21261);
xnor UO_1533 (O_1533,N_27731,N_22558);
nand UO_1534 (O_1534,N_29126,N_24115);
nand UO_1535 (O_1535,N_28723,N_25747);
and UO_1536 (O_1536,N_26967,N_29069);
nor UO_1537 (O_1537,N_27012,N_26987);
or UO_1538 (O_1538,N_23252,N_28292);
nor UO_1539 (O_1539,N_29078,N_23273);
nand UO_1540 (O_1540,N_25203,N_22963);
nand UO_1541 (O_1541,N_25183,N_26401);
and UO_1542 (O_1542,N_22931,N_25533);
nor UO_1543 (O_1543,N_27001,N_27599);
or UO_1544 (O_1544,N_29351,N_27559);
and UO_1545 (O_1545,N_21327,N_20026);
xnor UO_1546 (O_1546,N_29358,N_26535);
nor UO_1547 (O_1547,N_22892,N_29388);
and UO_1548 (O_1548,N_26701,N_21374);
and UO_1549 (O_1549,N_21673,N_27415);
or UO_1550 (O_1550,N_24474,N_29410);
and UO_1551 (O_1551,N_24388,N_21618);
xnor UO_1552 (O_1552,N_27761,N_20668);
nor UO_1553 (O_1553,N_26074,N_24805);
and UO_1554 (O_1554,N_22189,N_21522);
nor UO_1555 (O_1555,N_28196,N_25717);
xnor UO_1556 (O_1556,N_25462,N_27851);
xnor UO_1557 (O_1557,N_29550,N_23617);
xnor UO_1558 (O_1558,N_26486,N_21158);
nor UO_1559 (O_1559,N_22018,N_29003);
or UO_1560 (O_1560,N_27897,N_29499);
or UO_1561 (O_1561,N_28296,N_23559);
nand UO_1562 (O_1562,N_21224,N_20466);
nand UO_1563 (O_1563,N_29333,N_27471);
nor UO_1564 (O_1564,N_21009,N_24366);
or UO_1565 (O_1565,N_20225,N_27779);
xnor UO_1566 (O_1566,N_28624,N_23287);
and UO_1567 (O_1567,N_24492,N_24934);
xnor UO_1568 (O_1568,N_20059,N_28198);
or UO_1569 (O_1569,N_25813,N_20224);
nand UO_1570 (O_1570,N_27035,N_25282);
or UO_1571 (O_1571,N_21388,N_24545);
nor UO_1572 (O_1572,N_20553,N_25653);
and UO_1573 (O_1573,N_24015,N_23279);
or UO_1574 (O_1574,N_23420,N_20867);
nor UO_1575 (O_1575,N_26912,N_22182);
or UO_1576 (O_1576,N_29991,N_29718);
and UO_1577 (O_1577,N_22684,N_22552);
nor UO_1578 (O_1578,N_26972,N_20721);
and UO_1579 (O_1579,N_22346,N_26904);
and UO_1580 (O_1580,N_28951,N_26139);
xnor UO_1581 (O_1581,N_21524,N_27594);
nor UO_1582 (O_1582,N_29398,N_26169);
or UO_1583 (O_1583,N_26760,N_20852);
or UO_1584 (O_1584,N_20370,N_20317);
xnor UO_1585 (O_1585,N_29244,N_29021);
nor UO_1586 (O_1586,N_26063,N_29859);
and UO_1587 (O_1587,N_28359,N_27446);
nand UO_1588 (O_1588,N_26366,N_29883);
nor UO_1589 (O_1589,N_28188,N_20188);
nor UO_1590 (O_1590,N_22008,N_24097);
nor UO_1591 (O_1591,N_24318,N_28554);
or UO_1592 (O_1592,N_29867,N_27788);
or UO_1593 (O_1593,N_23262,N_28004);
or UO_1594 (O_1594,N_21783,N_26417);
and UO_1595 (O_1595,N_21275,N_23786);
nor UO_1596 (O_1596,N_26408,N_22562);
nor UO_1597 (O_1597,N_22756,N_22620);
xor UO_1598 (O_1598,N_21818,N_22514);
nand UO_1599 (O_1599,N_23850,N_25029);
or UO_1600 (O_1600,N_29698,N_22245);
or UO_1601 (O_1601,N_22330,N_27022);
xor UO_1602 (O_1602,N_20062,N_23797);
or UO_1603 (O_1603,N_20886,N_27621);
nand UO_1604 (O_1604,N_20577,N_24304);
and UO_1605 (O_1605,N_28784,N_24213);
xnor UO_1606 (O_1606,N_25643,N_29059);
nand UO_1607 (O_1607,N_21308,N_25814);
nand UO_1608 (O_1608,N_22276,N_27595);
or UO_1609 (O_1609,N_27315,N_29657);
or UO_1610 (O_1610,N_20147,N_25304);
nand UO_1611 (O_1611,N_23772,N_25874);
and UO_1612 (O_1612,N_27670,N_22943);
or UO_1613 (O_1613,N_21454,N_21647);
xnor UO_1614 (O_1614,N_27275,N_27029);
nor UO_1615 (O_1615,N_28365,N_20605);
nand UO_1616 (O_1616,N_28561,N_28623);
nand UO_1617 (O_1617,N_29393,N_27705);
or UO_1618 (O_1618,N_25673,N_25076);
nand UO_1619 (O_1619,N_26602,N_22496);
nor UO_1620 (O_1620,N_23411,N_29360);
and UO_1621 (O_1621,N_25697,N_20380);
or UO_1622 (O_1622,N_20599,N_22886);
nor UO_1623 (O_1623,N_20484,N_21904);
and UO_1624 (O_1624,N_20623,N_28735);
nand UO_1625 (O_1625,N_22339,N_21337);
nor UO_1626 (O_1626,N_23467,N_27723);
nor UO_1627 (O_1627,N_20961,N_23345);
nor UO_1628 (O_1628,N_20036,N_24551);
nor UO_1629 (O_1629,N_29402,N_24219);
nor UO_1630 (O_1630,N_25500,N_25351);
nand UO_1631 (O_1631,N_26556,N_24764);
or UO_1632 (O_1632,N_25631,N_26067);
or UO_1633 (O_1633,N_24792,N_21282);
or UO_1634 (O_1634,N_24580,N_20201);
nand UO_1635 (O_1635,N_22343,N_21686);
or UO_1636 (O_1636,N_21946,N_22413);
and UO_1637 (O_1637,N_21812,N_24775);
or UO_1638 (O_1638,N_24727,N_24041);
and UO_1639 (O_1639,N_25274,N_28523);
nand UO_1640 (O_1640,N_20130,N_23426);
nor UO_1641 (O_1641,N_23675,N_24676);
nand UO_1642 (O_1642,N_26513,N_26467);
nand UO_1643 (O_1643,N_27124,N_23379);
or UO_1644 (O_1644,N_20052,N_29264);
nor UO_1645 (O_1645,N_25418,N_27797);
nor UO_1646 (O_1646,N_24313,N_26426);
nor UO_1647 (O_1647,N_22006,N_29148);
nand UO_1648 (O_1648,N_20770,N_25215);
or UO_1649 (O_1649,N_24910,N_28293);
or UO_1650 (O_1650,N_28913,N_22500);
nor UO_1651 (O_1651,N_22013,N_28642);
nand UO_1652 (O_1652,N_25350,N_26739);
nor UO_1653 (O_1653,N_20309,N_25100);
and UO_1654 (O_1654,N_28371,N_24296);
nor UO_1655 (O_1655,N_29913,N_23161);
nor UO_1656 (O_1656,N_21829,N_23514);
nor UO_1657 (O_1657,N_26528,N_25064);
and UO_1658 (O_1658,N_23265,N_21634);
or UO_1659 (O_1659,N_22074,N_20522);
nand UO_1660 (O_1660,N_25698,N_21728);
or UO_1661 (O_1661,N_23871,N_24276);
nand UO_1662 (O_1662,N_27467,N_24786);
xnor UO_1663 (O_1663,N_25116,N_27059);
and UO_1664 (O_1664,N_25459,N_23311);
or UO_1665 (O_1665,N_25270,N_29537);
and UO_1666 (O_1666,N_20993,N_27104);
xnor UO_1667 (O_1667,N_23106,N_29213);
nand UO_1668 (O_1668,N_25433,N_28738);
nor UO_1669 (O_1669,N_28446,N_24637);
or UO_1670 (O_1670,N_22113,N_25315);
nor UO_1671 (O_1671,N_23732,N_20653);
and UO_1672 (O_1672,N_22884,N_28639);
and UO_1673 (O_1673,N_20121,N_22484);
nor UO_1674 (O_1674,N_27690,N_23833);
and UO_1675 (O_1675,N_21782,N_21651);
nand UO_1676 (O_1676,N_24647,N_25688);
nand UO_1677 (O_1677,N_23518,N_26796);
nor UO_1678 (O_1678,N_20390,N_27792);
or UO_1679 (O_1679,N_20523,N_20737);
nor UO_1680 (O_1680,N_29979,N_22915);
nand UO_1681 (O_1681,N_25672,N_25473);
nand UO_1682 (O_1682,N_24821,N_28709);
nand UO_1683 (O_1683,N_23663,N_29938);
or UO_1684 (O_1684,N_25468,N_29492);
nand UO_1685 (O_1685,N_21225,N_22881);
nand UO_1686 (O_1686,N_29520,N_24926);
and UO_1687 (O_1687,N_26814,N_28390);
and UO_1688 (O_1688,N_25573,N_28478);
and UO_1689 (O_1689,N_27930,N_22322);
and UO_1690 (O_1690,N_25532,N_24737);
nand UO_1691 (O_1691,N_21751,N_29432);
or UO_1692 (O_1692,N_20799,N_24134);
or UO_1693 (O_1693,N_24363,N_25608);
nor UO_1694 (O_1694,N_24618,N_29501);
nand UO_1695 (O_1695,N_26999,N_26172);
or UO_1696 (O_1696,N_24023,N_25032);
nor UO_1697 (O_1697,N_25056,N_24541);
or UO_1698 (O_1698,N_22355,N_20817);
nand UO_1699 (O_1699,N_25384,N_24912);
nor UO_1700 (O_1700,N_27484,N_28305);
nor UO_1701 (O_1701,N_24301,N_21098);
nand UO_1702 (O_1702,N_23553,N_27455);
xor UO_1703 (O_1703,N_24008,N_29762);
xnor UO_1704 (O_1704,N_27310,N_20736);
or UO_1705 (O_1705,N_26293,N_22015);
nor UO_1706 (O_1706,N_28329,N_20470);
nand UO_1707 (O_1707,N_21021,N_26011);
nor UO_1708 (O_1708,N_29241,N_26843);
nor UO_1709 (O_1709,N_27700,N_24936);
nor UO_1710 (O_1710,N_23115,N_29631);
xnor UO_1711 (O_1711,N_29572,N_27875);
nor UO_1712 (O_1712,N_23289,N_24191);
or UO_1713 (O_1713,N_21555,N_21761);
nor UO_1714 (O_1714,N_22038,N_21367);
nor UO_1715 (O_1715,N_24749,N_25843);
or UO_1716 (O_1716,N_22203,N_26743);
nand UO_1717 (O_1717,N_24571,N_21453);
nand UO_1718 (O_1718,N_24398,N_27823);
nor UO_1719 (O_1719,N_20299,N_26489);
nand UO_1720 (O_1720,N_21349,N_26464);
xnor UO_1721 (O_1721,N_21169,N_25691);
nor UO_1722 (O_1722,N_23029,N_26606);
nor UO_1723 (O_1723,N_26027,N_27388);
or UO_1724 (O_1724,N_28916,N_22970);
xnor UO_1725 (O_1725,N_29217,N_28366);
and UO_1726 (O_1726,N_25048,N_24543);
or UO_1727 (O_1727,N_24375,N_22076);
or UO_1728 (O_1728,N_23355,N_26164);
nor UO_1729 (O_1729,N_28937,N_27518);
nand UO_1730 (O_1730,N_23698,N_23234);
nor UO_1731 (O_1731,N_29879,N_24334);
nand UO_1732 (O_1732,N_24767,N_25307);
xnor UO_1733 (O_1733,N_21693,N_28109);
nand UO_1734 (O_1734,N_25675,N_25767);
nor UO_1735 (O_1735,N_20312,N_20451);
and UO_1736 (O_1736,N_27410,N_22430);
and UO_1737 (O_1737,N_22569,N_26004);
and UO_1738 (O_1738,N_28115,N_24011);
xnor UO_1739 (O_1739,N_20469,N_27795);
and UO_1740 (O_1740,N_27055,N_26769);
nand UO_1741 (O_1741,N_28396,N_26974);
nand UO_1742 (O_1742,N_21284,N_24747);
xnor UO_1743 (O_1743,N_28629,N_24502);
and UO_1744 (O_1744,N_28457,N_24110);
nor UO_1745 (O_1745,N_26599,N_26859);
and UO_1746 (O_1746,N_24312,N_28817);
xor UO_1747 (O_1747,N_26869,N_21201);
xnor UO_1748 (O_1748,N_25142,N_20885);
nor UO_1749 (O_1749,N_26847,N_27770);
and UO_1750 (O_1750,N_29924,N_28810);
nor UO_1751 (O_1751,N_28369,N_25375);
nand UO_1752 (O_1752,N_20672,N_26952);
nand UO_1753 (O_1753,N_26945,N_29715);
nand UO_1754 (O_1754,N_23656,N_29246);
or UO_1755 (O_1755,N_22316,N_27971);
and UO_1756 (O_1756,N_24957,N_29002);
or UO_1757 (O_1757,N_27280,N_23105);
nand UO_1758 (O_1758,N_29835,N_28718);
and UO_1759 (O_1759,N_27378,N_23745);
and UO_1760 (O_1760,N_29751,N_27018);
nand UO_1761 (O_1761,N_21161,N_29889);
nand UO_1762 (O_1762,N_28002,N_22284);
nand UO_1763 (O_1763,N_21975,N_23233);
nor UO_1764 (O_1764,N_26036,N_24019);
nor UO_1765 (O_1765,N_29327,N_21677);
nor UO_1766 (O_1766,N_24881,N_26412);
or UO_1767 (O_1767,N_22023,N_29545);
nand UO_1768 (O_1768,N_24939,N_22297);
nor UO_1769 (O_1769,N_24692,N_28350);
and UO_1770 (O_1770,N_23369,N_23099);
and UO_1771 (O_1771,N_24818,N_20221);
or UO_1772 (O_1772,N_25567,N_24405);
xnor UO_1773 (O_1773,N_23587,N_26879);
or UO_1774 (O_1774,N_24862,N_26132);
nand UO_1775 (O_1775,N_20534,N_26407);
and UO_1776 (O_1776,N_29827,N_21868);
and UO_1777 (O_1777,N_22107,N_26022);
or UO_1778 (O_1778,N_21405,N_26030);
nand UO_1779 (O_1779,N_28998,N_26271);
nor UO_1780 (O_1780,N_24799,N_23563);
nor UO_1781 (O_1781,N_28925,N_23668);
or UO_1782 (O_1782,N_20574,N_26256);
and UO_1783 (O_1783,N_22259,N_21157);
and UO_1784 (O_1784,N_24040,N_24141);
nor UO_1785 (O_1785,N_22357,N_20974);
xor UO_1786 (O_1786,N_26928,N_27338);
nand UO_1787 (O_1787,N_28313,N_28653);
nor UO_1788 (O_1788,N_23404,N_28269);
xnor UO_1789 (O_1789,N_24348,N_20910);
xor UO_1790 (O_1790,N_22311,N_29757);
xor UO_1791 (O_1791,N_28320,N_20284);
nor UO_1792 (O_1792,N_26938,N_27482);
nand UO_1793 (O_1793,N_22719,N_22662);
nor UO_1794 (O_1794,N_24315,N_25883);
or UO_1795 (O_1795,N_22386,N_27843);
or UO_1796 (O_1796,N_25954,N_28330);
nor UO_1797 (O_1797,N_20289,N_27091);
or UO_1798 (O_1798,N_23948,N_26522);
nor UO_1799 (O_1799,N_29921,N_25190);
nand UO_1800 (O_1800,N_27961,N_27300);
or UO_1801 (O_1801,N_29447,N_25272);
nand UO_1802 (O_1802,N_25122,N_21184);
nor UO_1803 (O_1803,N_21084,N_22937);
nor UO_1804 (O_1804,N_21300,N_22030);
nor UO_1805 (O_1805,N_21899,N_25586);
nand UO_1806 (O_1806,N_25961,N_28245);
xnor UO_1807 (O_1807,N_25977,N_26355);
nand UO_1808 (O_1808,N_20684,N_29905);
or UO_1809 (O_1809,N_23917,N_25313);
xnor UO_1810 (O_1810,N_25991,N_26552);
nand UO_1811 (O_1811,N_20637,N_25851);
and UO_1812 (O_1812,N_20664,N_22891);
or UO_1813 (O_1813,N_23970,N_26261);
and UO_1814 (O_1814,N_22990,N_28123);
nor UO_1815 (O_1815,N_25535,N_25800);
xor UO_1816 (O_1816,N_29830,N_23294);
nor UO_1817 (O_1817,N_22965,N_24170);
or UO_1818 (O_1818,N_26435,N_29269);
nor UO_1819 (O_1819,N_21502,N_26992);
xnor UO_1820 (O_1820,N_29898,N_24130);
nor UO_1821 (O_1821,N_27652,N_28859);
nor UO_1822 (O_1822,N_22861,N_24773);
nand UO_1823 (O_1823,N_20632,N_20142);
and UO_1824 (O_1824,N_22231,N_29349);
and UO_1825 (O_1825,N_27648,N_23441);
nor UO_1826 (O_1826,N_21048,N_25568);
nand UO_1827 (O_1827,N_23448,N_21608);
xnor UO_1828 (O_1828,N_21014,N_24288);
and UO_1829 (O_1829,N_22278,N_20803);
xnor UO_1830 (O_1830,N_23449,N_25509);
and UO_1831 (O_1831,N_25854,N_22039);
xnor UO_1832 (O_1832,N_26584,N_29201);
nor UO_1833 (O_1833,N_27632,N_24454);
or UO_1834 (O_1834,N_20355,N_21412);
or UO_1835 (O_1835,N_22022,N_22527);
or UO_1836 (O_1836,N_27148,N_27844);
xor UO_1837 (O_1837,N_23539,N_21351);
or UO_1838 (O_1838,N_28025,N_27573);
xor UO_1839 (O_1839,N_27509,N_26440);
nand UO_1840 (O_1840,N_27319,N_23401);
nand UO_1841 (O_1841,N_28426,N_23716);
or UO_1842 (O_1842,N_22472,N_22617);
nand UO_1843 (O_1843,N_28803,N_23771);
nand UO_1844 (O_1844,N_25419,N_23151);
or UO_1845 (O_1845,N_29538,N_20241);
or UO_1846 (O_1846,N_20392,N_26496);
or UO_1847 (O_1847,N_28096,N_24427);
nand UO_1848 (O_1848,N_24650,N_21628);
or UO_1849 (O_1849,N_25209,N_24828);
or UO_1850 (O_1850,N_26305,N_26154);
xor UO_1851 (O_1851,N_22366,N_28837);
and UO_1852 (O_1852,N_26953,N_22324);
and UO_1853 (O_1853,N_24566,N_28214);
nor UO_1854 (O_1854,N_24089,N_23903);
and UO_1855 (O_1855,N_28592,N_22985);
nor UO_1856 (O_1856,N_23724,N_23533);
nor UO_1857 (O_1857,N_24338,N_26532);
or UO_1858 (O_1858,N_24758,N_29528);
or UO_1859 (O_1859,N_23607,N_22751);
nand UO_1860 (O_1860,N_26890,N_27258);
or UO_1861 (O_1861,N_25856,N_23666);
nand UO_1862 (O_1862,N_28512,N_28677);
nand UO_1863 (O_1863,N_29653,N_24510);
nand UO_1864 (O_1864,N_20525,N_29839);
or UO_1865 (O_1865,N_28363,N_23749);
and UO_1866 (O_1866,N_20178,N_22551);
or UO_1867 (O_1867,N_21070,N_28049);
nand UO_1868 (O_1868,N_29613,N_20270);
nand UO_1869 (O_1869,N_20755,N_28860);
or UO_1870 (O_1870,N_23891,N_28904);
xnor UO_1871 (O_1871,N_28999,N_27408);
and UO_1872 (O_1872,N_24210,N_26370);
and UO_1873 (O_1873,N_22547,N_22351);
and UO_1874 (O_1874,N_22945,N_28316);
and UO_1875 (O_1875,N_20712,N_25387);
or UO_1876 (O_1876,N_20777,N_28840);
or UO_1877 (O_1877,N_27984,N_28902);
or UO_1878 (O_1878,N_24380,N_20827);
and UO_1879 (O_1879,N_27825,N_25250);
nand UO_1880 (O_1880,N_29834,N_26436);
or UO_1881 (O_1881,N_27426,N_21206);
and UO_1882 (O_1882,N_22853,N_20631);
and UO_1883 (O_1883,N_26055,N_20983);
nor UO_1884 (O_1884,N_29535,N_24347);
or UO_1885 (O_1885,N_27422,N_26510);
nand UO_1886 (O_1886,N_26455,N_29001);
nand UO_1887 (O_1887,N_22274,N_20341);
and UO_1888 (O_1888,N_29271,N_21948);
nand UO_1889 (O_1889,N_20076,N_28186);
nand UO_1890 (O_1890,N_27909,N_24964);
nor UO_1891 (O_1891,N_25024,N_21147);
nand UO_1892 (O_1892,N_22359,N_25616);
nand UO_1893 (O_1893,N_21537,N_20182);
nor UO_1894 (O_1894,N_26557,N_29795);
xnor UO_1895 (O_1895,N_20116,N_26123);
nand UO_1896 (O_1896,N_21029,N_20411);
nand UO_1897 (O_1897,N_27106,N_22187);
xor UO_1898 (O_1898,N_24330,N_23526);
or UO_1899 (O_1899,N_29339,N_28420);
and UO_1900 (O_1900,N_22795,N_24407);
or UO_1901 (O_1901,N_20337,N_21392);
nand UO_1902 (O_1902,N_27865,N_27444);
and UO_1903 (O_1903,N_28960,N_21000);
nand UO_1904 (O_1904,N_22956,N_28638);
or UO_1905 (O_1905,N_25501,N_29990);
and UO_1906 (O_1906,N_20056,N_26176);
nand UO_1907 (O_1907,N_22863,N_21778);
and UO_1908 (O_1908,N_20112,N_28574);
nor UO_1909 (O_1909,N_27067,N_22434);
nor UO_1910 (O_1910,N_29443,N_29119);
and UO_1911 (O_1911,N_27077,N_27869);
and UO_1912 (O_1912,N_25152,N_25355);
and UO_1913 (O_1913,N_27016,N_28739);
nand UO_1914 (O_1914,N_25822,N_23249);
nand UO_1915 (O_1915,N_27289,N_25993);
or UO_1916 (O_1916,N_20793,N_26145);
nand UO_1917 (O_1917,N_21034,N_22632);
or UO_1918 (O_1918,N_21888,N_22978);
or UO_1919 (O_1919,N_22896,N_29230);
and UO_1920 (O_1920,N_27997,N_20211);
and UO_1921 (O_1921,N_29304,N_22577);
nor UO_1922 (O_1922,N_23312,N_22021);
and UO_1923 (O_1923,N_28765,N_24000);
and UO_1924 (O_1924,N_28399,N_29085);
nor UO_1925 (O_1925,N_23191,N_26652);
nor UO_1926 (O_1926,N_23022,N_23550);
nor UO_1927 (O_1927,N_27263,N_22615);
and UO_1928 (O_1928,N_24064,N_29206);
and UO_1929 (O_1929,N_25055,N_23478);
or UO_1930 (O_1930,N_27635,N_27157);
or UO_1931 (O_1931,N_23901,N_27985);
and UO_1932 (O_1932,N_21977,N_25600);
or UO_1933 (O_1933,N_29681,N_24639);
or UO_1934 (O_1934,N_21570,N_25041);
and UO_1935 (O_1935,N_28479,N_22668);
or UO_1936 (O_1936,N_23454,N_25976);
nor UO_1937 (O_1937,N_27354,N_28027);
nor UO_1938 (O_1938,N_22055,N_23951);
nor UO_1939 (O_1939,N_22451,N_21411);
nand UO_1940 (O_1940,N_28208,N_22658);
or UO_1941 (O_1941,N_22599,N_21831);
nor UO_1942 (O_1942,N_26517,N_28762);
nor UO_1943 (O_1943,N_20242,N_26512);
or UO_1944 (O_1944,N_27290,N_21638);
and UO_1945 (O_1945,N_27755,N_21276);
nand UO_1946 (O_1946,N_21086,N_21793);
xor UO_1947 (O_1947,N_29397,N_28451);
or UO_1948 (O_1948,N_26531,N_26186);
nand UO_1949 (O_1949,N_26746,N_29377);
and UO_1950 (O_1950,N_27177,N_24883);
and UO_1951 (O_1951,N_21760,N_21353);
or UO_1952 (O_1952,N_23562,N_23780);
nor UO_1953 (O_1953,N_21885,N_21141);
or UO_1954 (O_1954,N_21058,N_20728);
nor UO_1955 (O_1955,N_21913,N_23354);
xnor UO_1956 (O_1956,N_29184,N_20990);
nor UO_1957 (O_1957,N_26667,N_26515);
or UO_1958 (O_1958,N_28698,N_23580);
nand UO_1959 (O_1959,N_28841,N_24760);
nand UO_1960 (O_1960,N_24809,N_22818);
nand UO_1961 (O_1961,N_29599,N_29736);
nor UO_1962 (O_1962,N_24537,N_29629);
or UO_1963 (O_1963,N_28632,N_25877);
xor UO_1964 (O_1964,N_28908,N_21404);
or UO_1965 (O_1965,N_28652,N_28018);
nand UO_1966 (O_1966,N_25844,N_23087);
xor UO_1967 (O_1967,N_20260,N_21343);
and UO_1968 (O_1968,N_26514,N_20057);
nand UO_1969 (O_1969,N_29999,N_20797);
and UO_1970 (O_1970,N_29096,N_24468);
nor UO_1971 (O_1971,N_28884,N_22855);
and UO_1972 (O_1972,N_21616,N_25401);
nand UO_1973 (O_1973,N_28117,N_23919);
or UO_1974 (O_1974,N_21926,N_25371);
nor UO_1975 (O_1975,N_28168,N_29049);
nor UO_1976 (O_1976,N_26673,N_29151);
and UO_1977 (O_1977,N_25417,N_22550);
nor UO_1978 (O_1978,N_21228,N_29074);
and UO_1979 (O_1979,N_23658,N_26946);
nor UO_1980 (O_1980,N_28189,N_29931);
or UO_1981 (O_1981,N_23795,N_21305);
xor UO_1982 (O_1982,N_28813,N_24864);
nand UO_1983 (O_1983,N_27283,N_20839);
and UO_1984 (O_1984,N_21909,N_29321);
nand UO_1985 (O_1985,N_25769,N_20562);
or UO_1986 (O_1986,N_23648,N_22649);
and UO_1987 (O_1987,N_23577,N_25381);
nor UO_1988 (O_1988,N_21586,N_24987);
nand UO_1989 (O_1989,N_27794,N_21920);
and UO_1990 (O_1990,N_22045,N_20880);
and UO_1991 (O_1991,N_21440,N_21068);
nand UO_1992 (O_1992,N_28207,N_28710);
and UO_1993 (O_1993,N_22713,N_27520);
or UO_1994 (O_1994,N_26566,N_22172);
and UO_1995 (O_1995,N_29293,N_23622);
nand UO_1996 (O_1996,N_21551,N_28172);
and UO_1997 (O_1997,N_26633,N_24824);
nand UO_1998 (O_1998,N_20663,N_21700);
or UO_1999 (O_1999,N_21866,N_24547);
or UO_2000 (O_2000,N_23554,N_25732);
or UO_2001 (O_2001,N_20651,N_26385);
nor UO_2002 (O_2002,N_28518,N_25074);
or UO_2003 (O_2003,N_24308,N_29908);
nand UO_2004 (O_2004,N_27920,N_20995);
xor UO_2005 (O_2005,N_20166,N_22398);
nand UO_2006 (O_2006,N_21470,N_29899);
xnor UO_2007 (O_2007,N_24295,N_22043);
nor UO_2008 (O_2008,N_23561,N_20088);
or UO_2009 (O_2009,N_29567,N_20307);
or UO_2010 (O_2010,N_25817,N_24659);
or UO_2011 (O_2011,N_25834,N_27304);
nor UO_2012 (O_2012,N_27642,N_22663);
nor UO_2013 (O_2013,N_20105,N_21636);
nand UO_2014 (O_2014,N_24072,N_28021);
nor UO_2015 (O_2015,N_22805,N_25445);
nand UO_2016 (O_2016,N_21210,N_24542);
nand UO_2017 (O_2017,N_26475,N_24656);
or UO_2018 (O_2018,N_22084,N_20939);
nor UO_2019 (O_2019,N_29810,N_22341);
nor UO_2020 (O_2020,N_27739,N_25719);
or UO_2021 (O_2021,N_23300,N_21216);
or UO_2022 (O_2022,N_24246,N_20086);
nand UO_2023 (O_2023,N_21607,N_26867);
and UO_2024 (O_2024,N_29730,N_20638);
nand UO_2025 (O_2025,N_29973,N_27877);
nor UO_2026 (O_2026,N_22488,N_27201);
nand UO_2027 (O_2027,N_25181,N_29371);
and UO_2028 (O_2028,N_27321,N_29356);
and UO_2029 (O_2029,N_24538,N_28882);
or UO_2030 (O_2030,N_20343,N_24712);
and UO_2031 (O_2031,N_23829,N_22850);
and UO_2032 (O_2032,N_27165,N_29378);
nor UO_2033 (O_2033,N_27170,N_28986);
and UO_2034 (O_2034,N_27074,N_26835);
nor UO_2035 (O_2035,N_20202,N_29957);
and UO_2036 (O_2036,N_20447,N_27406);
xor UO_2037 (O_2037,N_28275,N_28587);
or UO_2038 (O_2038,N_25314,N_24286);
and UO_2039 (O_2039,N_25093,N_20650);
nand UO_2040 (O_2040,N_22580,N_29950);
nor UO_2041 (O_2041,N_23762,N_20379);
nand UO_2042 (O_2042,N_28968,N_26643);
xnor UO_2043 (O_2043,N_20796,N_27192);
or UO_2044 (O_2044,N_22241,N_20368);
nor UO_2045 (O_2045,N_20223,N_25590);
nor UO_2046 (O_2046,N_28357,N_20391);
nor UO_2047 (O_2047,N_25878,N_26577);
or UO_2048 (O_2048,N_22958,N_25562);
or UO_2049 (O_2049,N_28271,N_24536);
nor UO_2050 (O_2050,N_20165,N_29114);
nor UO_2051 (O_2051,N_22068,N_22907);
and UO_2052 (O_2052,N_22211,N_24679);
nor UO_2053 (O_2053,N_24524,N_25687);
xor UO_2054 (O_2054,N_23130,N_26905);
or UO_2055 (O_2055,N_26883,N_22390);
nor UO_2056 (O_2056,N_28144,N_27447);
nor UO_2057 (O_2057,N_29112,N_20443);
and UO_2058 (O_2058,N_25659,N_26135);
or UO_2059 (O_2059,N_29302,N_26959);
or UO_2060 (O_2060,N_29469,N_27017);
nor UO_2061 (O_2061,N_26039,N_21151);
nand UO_2062 (O_2062,N_22778,N_26963);
nor UO_2063 (O_2063,N_20007,N_22964);
or UO_2064 (O_2064,N_24720,N_21963);
and UO_2065 (O_2065,N_20774,N_24982);
and UO_2066 (O_2066,N_21556,N_28825);
nand UO_2067 (O_2067,N_27789,N_26663);
nor UO_2068 (O_2068,N_25196,N_29018);
and UO_2069 (O_2069,N_20634,N_20335);
and UO_2070 (O_2070,N_24208,N_22885);
or UO_2071 (O_2071,N_29309,N_20697);
nor UO_2072 (O_2072,N_20870,N_21517);
nand UO_2073 (O_2073,N_22373,N_28612);
and UO_2074 (O_2074,N_27262,N_20000);
nor UO_2075 (O_2075,N_24074,N_23204);
and UO_2076 (O_2076,N_25208,N_25636);
or UO_2077 (O_2077,N_26078,N_24464);
or UO_2078 (O_2078,N_22941,N_29541);
and UO_2079 (O_2079,N_25966,N_20216);
nand UO_2080 (O_2080,N_29524,N_20811);
and UO_2081 (O_2081,N_26494,N_28443);
xor UO_2082 (O_2082,N_29423,N_21474);
or UO_2083 (O_2083,N_23430,N_21794);
nand UO_2084 (O_2084,N_23707,N_23380);
nand UO_2085 (O_2085,N_29738,N_26934);
xor UO_2086 (O_2086,N_21221,N_22591);
and UO_2087 (O_2087,N_20113,N_25306);
and UO_2088 (O_2088,N_26462,N_23894);
nor UO_2089 (O_2089,N_20519,N_26970);
and UO_2090 (O_2090,N_24868,N_21587);
nand UO_2091 (O_2091,N_25398,N_20846);
nor UO_2092 (O_2092,N_29338,N_29993);
and UO_2093 (O_2093,N_20099,N_25020);
nand UO_2094 (O_2094,N_21894,N_26050);
nand UO_2095 (O_2095,N_28767,N_22438);
nand UO_2096 (O_2096,N_29311,N_25803);
nand UO_2097 (O_2097,N_28857,N_28876);
and UO_2098 (O_2098,N_26636,N_29472);
nor UO_2099 (O_2099,N_24784,N_24608);
and UO_2100 (O_2100,N_28893,N_20887);
and UO_2101 (O_2101,N_22266,N_21970);
xnor UO_2102 (O_2102,N_26219,N_24321);
and UO_2103 (O_2103,N_25759,N_27586);
xor UO_2104 (O_2104,N_25827,N_25089);
or UO_2105 (O_2105,N_22517,N_28691);
and UO_2106 (O_2106,N_24156,N_22118);
nand UO_2107 (O_2107,N_22822,N_21445);
or UO_2108 (O_2108,N_27223,N_24239);
nor UO_2109 (O_2109,N_23819,N_24930);
nand UO_2110 (O_2110,N_26570,N_25382);
or UO_2111 (O_2111,N_24034,N_22816);
nor UO_2112 (O_2112,N_29109,N_26525);
and UO_2113 (O_2113,N_26765,N_24119);
nor UO_2114 (O_2114,N_20959,N_20657);
and UO_2115 (O_2115,N_20054,N_29739);
or UO_2116 (O_2116,N_20630,N_25964);
nor UO_2117 (O_2117,N_23908,N_29369);
nor UO_2118 (O_2118,N_29433,N_28750);
or UO_2119 (O_2119,N_22717,N_22627);
nor UO_2120 (O_2120,N_28210,N_24677);
nand UO_2121 (O_2121,N_23183,N_26052);
and UO_2122 (O_2122,N_28823,N_25211);
and UO_2123 (O_2123,N_24975,N_25429);
or UO_2124 (O_2124,N_23432,N_23966);
nor UO_2125 (O_2125,N_23613,N_23200);
nand UO_2126 (O_2126,N_28073,N_25925);
and UO_2127 (O_2127,N_25369,N_28984);
nor UO_2128 (O_2128,N_25472,N_20158);
nand UO_2129 (O_2129,N_29093,N_27694);
or UO_2130 (O_2130,N_29460,N_23412);
or UO_2131 (O_2131,N_24251,N_22585);
or UO_2132 (O_2132,N_24871,N_29207);
nor UO_2133 (O_2133,N_23877,N_22128);
nand UO_2134 (O_2134,N_20276,N_29310);
nand UO_2135 (O_2135,N_29483,N_27023);
xor UO_2136 (O_2136,N_28410,N_20435);
or UO_2137 (O_2137,N_25530,N_25709);
and UO_2138 (O_2138,N_24390,N_23285);
nor UO_2139 (O_2139,N_20890,N_24434);
nor UO_2140 (O_2140,N_20189,N_28381);
xor UO_2141 (O_2141,N_22060,N_23704);
or UO_2142 (O_2142,N_24670,N_22207);
and UO_2143 (O_2143,N_23268,N_28361);
and UO_2144 (O_2144,N_24684,N_24035);
or UO_2145 (O_2145,N_21892,N_21919);
or UO_2146 (O_2146,N_21024,N_21468);
or UO_2147 (O_2147,N_23896,N_24680);
and UO_2148 (O_2148,N_22458,N_27032);
and UO_2149 (O_2149,N_25792,N_26266);
and UO_2150 (O_2150,N_24452,N_22161);
nor UO_2151 (O_2151,N_21119,N_28667);
nand UO_2152 (O_2152,N_29275,N_28145);
nand UO_2153 (O_2153,N_23981,N_25705);
and UO_2154 (O_2154,N_20749,N_20373);
nor UO_2155 (O_2155,N_29043,N_26635);
or UO_2156 (O_2156,N_21906,N_23909);
and UO_2157 (O_2157,N_20310,N_28035);
and UO_2158 (O_2158,N_26792,N_29218);
xnor UO_2159 (O_2159,N_24185,N_25480);
xor UO_2160 (O_2160,N_20850,N_28864);
or UO_2161 (O_2161,N_29523,N_25690);
nor UO_2162 (O_2162,N_28699,N_22138);
nand UO_2163 (O_2163,N_28005,N_20048);
nor UO_2164 (O_2164,N_24184,N_26984);
nand UO_2165 (O_2165,N_20981,N_29077);
xor UO_2166 (O_2166,N_29295,N_23722);
or UO_2167 (O_2167,N_25216,N_29135);
nand UO_2168 (O_2168,N_21095,N_29261);
or UO_2169 (O_2169,N_22376,N_25956);
or UO_2170 (O_2170,N_23302,N_28075);
nand UO_2171 (O_2171,N_25298,N_28486);
or UO_2172 (O_2172,N_25038,N_25837);
and UO_2173 (O_2173,N_29658,N_23012);
nand UO_2174 (O_2174,N_23197,N_29592);
or UO_2175 (O_2175,N_28270,N_27814);
nor UO_2176 (O_2176,N_25109,N_23655);
and UO_2177 (O_2177,N_23751,N_27521);
and UO_2178 (O_2178,N_25997,N_25265);
nor UO_2179 (O_2179,N_25790,N_22723);
and UO_2180 (O_2180,N_28608,N_21690);
and UO_2181 (O_2181,N_28634,N_27499);
nand UO_2182 (O_2182,N_26818,N_23510);
or UO_2183 (O_2183,N_24612,N_26526);
or UO_2184 (O_2184,N_29717,N_29692);
nand UO_2185 (O_2185,N_22243,N_20474);
or UO_2186 (O_2186,N_29449,N_23239);
nand UO_2187 (O_2187,N_28973,N_27876);
and UO_2188 (O_2188,N_27025,N_28112);
xor UO_2189 (O_2189,N_28556,N_28581);
or UO_2190 (O_2190,N_22581,N_29769);
nor UO_2191 (O_2191,N_24913,N_26612);
nand UO_2192 (O_2192,N_24698,N_25614);
xor UO_2193 (O_2193,N_22441,N_27435);
nor UO_2194 (O_2194,N_25441,N_24574);
nor UO_2195 (O_2195,N_29129,N_24482);
or UO_2196 (O_2196,N_22321,N_25884);
nand UO_2197 (O_2197,N_25658,N_24628);
or UO_2198 (O_2198,N_25006,N_22572);
nor UO_2199 (O_2199,N_24700,N_29167);
or UO_2200 (O_2200,N_26927,N_23610);
or UO_2201 (O_2201,N_27045,N_23357);
nor UO_2202 (O_2202,N_24367,N_28360);
nor UO_2203 (O_2203,N_20520,N_21373);
or UO_2204 (O_2204,N_26252,N_25986);
or UO_2205 (O_2205,N_25171,N_28031);
and UO_2206 (O_2206,N_29620,N_22923);
nand UO_2207 (O_2207,N_29574,N_24387);
or UO_2208 (O_2208,N_23307,N_23543);
or UO_2209 (O_2209,N_26101,N_25788);
nor UO_2210 (O_2210,N_28977,N_28782);
xor UO_2211 (O_2211,N_25276,N_25344);
nor UO_2212 (O_2212,N_25115,N_29532);
and UO_2213 (O_2213,N_22342,N_22131);
and UO_2214 (O_2214,N_22025,N_29480);
or UO_2215 (O_2215,N_23969,N_27982);
nand UO_2216 (O_2216,N_23621,N_25781);
and UO_2217 (O_2217,N_22637,N_26442);
nand UO_2218 (O_2218,N_28458,N_26108);
and UO_2219 (O_2219,N_21846,N_24284);
nor UO_2220 (O_2220,N_21898,N_28564);
nand UO_2221 (O_2221,N_26481,N_20384);
and UO_2222 (O_2222,N_29165,N_25727);
nor UO_2223 (O_2223,N_23318,N_29006);
or UO_2224 (O_2224,N_20928,N_21485);
nand UO_2225 (O_2225,N_26831,N_23251);
and UO_2226 (O_2226,N_24826,N_27237);
nand UO_2227 (O_2227,N_28135,N_24915);
nand UO_2228 (O_2228,N_25498,N_27565);
nor UO_2229 (O_2229,N_29081,N_25538);
nor UO_2230 (O_2230,N_28480,N_29934);
nor UO_2231 (O_2231,N_24916,N_21917);
nand UO_2232 (O_2232,N_24438,N_21325);
and UO_2233 (O_2233,N_20585,N_24992);
and UO_2234 (O_2234,N_28921,N_20917);
or UO_2235 (O_2235,N_20636,N_20649);
and UO_2236 (O_2236,N_27663,N_20093);
xor UO_2237 (O_2237,N_24455,N_22459);
and UO_2238 (O_2238,N_21958,N_25186);
nand UO_2239 (O_2239,N_27002,N_22648);
or UO_2240 (O_2240,N_20040,N_22967);
nand UO_2241 (O_2241,N_21408,N_26922);
and UO_2242 (O_2242,N_28106,N_28379);
nor UO_2243 (O_2243,N_28790,N_23095);
or UO_2244 (O_2244,N_29962,N_26659);
or UO_2245 (O_2245,N_22075,N_20300);
nand UO_2246 (O_2246,N_26590,N_25928);
nor UO_2247 (O_2247,N_20826,N_28570);
nor UO_2248 (O_2248,N_29881,N_23997);
or UO_2249 (O_2249,N_23297,N_26451);
nor UO_2250 (O_2250,N_26703,N_27014);
or UO_2251 (O_2251,N_22606,N_29818);
nand UO_2252 (O_2252,N_28259,N_29978);
and UO_2253 (O_2253,N_22306,N_21302);
and UO_2254 (O_2254,N_21954,N_29663);
and UO_2255 (O_2255,N_24648,N_23292);
nor UO_2256 (O_2256,N_23792,N_23419);
and UO_2257 (O_2257,N_22000,N_20790);
nor UO_2258 (O_2258,N_26764,N_28161);
nor UO_2259 (O_2259,N_22277,N_29138);
xnor UO_2260 (O_2260,N_20164,N_23278);
nand UO_2261 (O_2261,N_25003,N_27250);
or UO_2262 (O_2262,N_27510,N_21376);
xnor UO_2263 (O_2263,N_21365,N_24155);
nand UO_2264 (O_2264,N_28289,N_22309);
and UO_2265 (O_2265,N_26459,N_23641);
or UO_2266 (O_2266,N_26284,N_20381);
nand UO_2267 (O_2267,N_20243,N_20354);
and UO_2268 (O_2268,N_26009,N_22993);
nand UO_2269 (O_2269,N_24368,N_26275);
or UO_2270 (O_2270,N_28131,N_22070);
nor UO_2271 (O_2271,N_20596,N_28408);
and UO_2272 (O_2272,N_21403,N_25957);
nor UO_2273 (O_2273,N_22119,N_29897);
and UO_2274 (O_2274,N_25546,N_20720);
nor UO_2275 (O_2275,N_27502,N_29733);
nand UO_2276 (O_2276,N_21065,N_23827);
or UO_2277 (O_2277,N_29110,N_28946);
nand UO_2278 (O_2278,N_21212,N_27478);
nor UO_2279 (O_2279,N_25449,N_22749);
and UO_2280 (O_2280,N_28625,N_28620);
nor UO_2281 (O_2281,N_24996,N_29298);
or UO_2282 (O_2282,N_22601,N_29812);
xnor UO_2283 (O_2283,N_28746,N_22711);
or UO_2284 (O_2284,N_28184,N_20044);
nor UO_2285 (O_2285,N_24476,N_22092);
and UO_2286 (O_2286,N_20709,N_26438);
and UO_2287 (O_2287,N_27228,N_29980);
nor UO_2288 (O_2288,N_27437,N_28714);
nand UO_2289 (O_2289,N_29131,N_20244);
nor UO_2290 (O_2290,N_25328,N_25248);
nor UO_2291 (O_2291,N_23452,N_29442);
and UO_2292 (O_2292,N_22050,N_27570);
nor UO_2293 (O_2293,N_28645,N_23882);
nor UO_2294 (O_2294,N_22184,N_22733);
nor UO_2295 (O_2295,N_27716,N_28515);
nor UO_2296 (O_2296,N_21429,N_28046);
and UO_2297 (O_2297,N_25869,N_28725);
nand UO_2298 (O_2298,N_22802,N_29560);
or UO_2299 (O_2299,N_25173,N_24016);
nor UO_2300 (O_2300,N_20433,N_24004);
nor UO_2301 (O_2301,N_26120,N_23509);
or UO_2302 (O_2302,N_23295,N_21423);
nand UO_2303 (O_2303,N_28141,N_21370);
nand UO_2304 (O_2304,N_22957,N_26981);
xnor UO_2305 (O_2305,N_29985,N_28351);
nor UO_2306 (O_2306,N_28513,N_22836);
nor UO_2307 (O_2307,N_29199,N_20119);
nor UO_2308 (O_2308,N_24793,N_26910);
and UO_2309 (O_2309,N_23691,N_28404);
nand UO_2310 (O_2310,N_24624,N_22521);
or UO_2311 (O_2311,N_21790,N_29015);
nand UO_2312 (O_2312,N_28059,N_21120);
nor UO_2313 (O_2313,N_21996,N_20982);
nor UO_2314 (O_2314,N_26321,N_21436);
xnor UO_2315 (O_2315,N_24337,N_23898);
nand UO_2316 (O_2316,N_21558,N_27815);
and UO_2317 (O_2317,N_22063,N_24223);
nand UO_2318 (O_2318,N_23174,N_27960);
nand UO_2319 (O_2319,N_20296,N_20549);
nor UO_2320 (O_2320,N_29354,N_23492);
and UO_2321 (O_2321,N_23988,N_24544);
or UO_2322 (O_2322,N_28671,N_25515);
nand UO_2323 (O_2323,N_22973,N_25301);
and UO_2324 (O_2324,N_20701,N_24586);
or UO_2325 (O_2325,N_28066,N_24215);
and UO_2326 (O_2326,N_26116,N_20060);
and UO_2327 (O_2327,N_25560,N_23024);
nor UO_2328 (O_2328,N_23994,N_28873);
nor UO_2329 (O_2329,N_27693,N_20575);
xnor UO_2330 (O_2330,N_20800,N_24371);
or UO_2331 (O_2331,N_26238,N_25361);
and UO_2332 (O_2332,N_22986,N_29598);
nand UO_2333 (O_2333,N_20747,N_26142);
xor UO_2334 (O_2334,N_25807,N_27372);
nor UO_2335 (O_2335,N_20450,N_24765);
and UO_2336 (O_2336,N_24458,N_29981);
and UO_2337 (O_2337,N_23112,N_20126);
or UO_2338 (O_2338,N_24520,N_25865);
nor UO_2339 (O_2339,N_22725,N_24369);
nand UO_2340 (O_2340,N_20517,N_28448);
and UO_2341 (O_2341,N_22939,N_21438);
nor UO_2342 (O_2342,N_21703,N_24776);
nor UO_2343 (O_2343,N_20069,N_26175);
nor UO_2344 (O_2344,N_26171,N_20199);
nand UO_2345 (O_2345,N_20544,N_28136);
nor UO_2346 (O_2346,N_23407,N_21375);
and UO_2347 (O_2347,N_22526,N_28297);
and UO_2348 (O_2348,N_20264,N_21028);
and UO_2349 (O_2349,N_22681,N_24270);
nand UO_2350 (O_2350,N_21964,N_23400);
nand UO_2351 (O_2351,N_21630,N_28471);
nor UO_2352 (O_2352,N_25279,N_21484);
and UO_2353 (O_2353,N_22065,N_24642);
xnor UO_2354 (O_2354,N_25801,N_22034);
or UO_2355 (O_2355,N_28469,N_29453);
or UO_2356 (O_2356,N_23188,N_20429);
or UO_2357 (O_2357,N_26877,N_25699);
or UO_2358 (O_2358,N_26237,N_24144);
and UO_2359 (O_2359,N_21394,N_24151);
and UO_2360 (O_2360,N_28812,N_26562);
and UO_2361 (O_2361,N_26265,N_29251);
nand UO_2362 (O_2362,N_24658,N_27760);
and UO_2363 (O_2363,N_29570,N_28808);
nor UO_2364 (O_2364,N_28250,N_22629);
xor UO_2365 (O_2365,N_29918,N_23708);
xor UO_2366 (O_2366,N_27637,N_28776);
nor UO_2367 (O_2367,N_21612,N_20101);
nand UO_2368 (O_2368,N_22262,N_26868);
nor UO_2369 (O_2369,N_25285,N_23620);
nor UO_2370 (O_2370,N_21037,N_24370);
and UO_2371 (O_2371,N_24995,N_21379);
or UO_2372 (O_2372,N_28994,N_22750);
and UO_2373 (O_2373,N_21223,N_24399);
xnor UO_2374 (O_2374,N_22035,N_28797);
nand UO_2375 (O_2375,N_23976,N_27785);
and UO_2376 (O_2376,N_29956,N_22966);
nand UO_2377 (O_2377,N_21022,N_21202);
or UO_2378 (O_2378,N_29054,N_22669);
and UO_2379 (O_2379,N_20555,N_25909);
and UO_2380 (O_2380,N_23985,N_22433);
and UO_2381 (O_2381,N_28302,N_22379);
and UO_2382 (O_2382,N_27156,N_24522);
or UO_2383 (O_2383,N_24498,N_26352);
nor UO_2384 (O_2384,N_22862,N_26187);
or UO_2385 (O_2385,N_22163,N_28091);
xnor UO_2386 (O_2386,N_20927,N_20446);
nor UO_2387 (O_2387,N_27784,N_23934);
and UO_2388 (O_2388,N_24224,N_27453);
xor UO_2389 (O_2389,N_29677,N_29735);
nand UO_2390 (O_2390,N_23255,N_26236);
or UO_2391 (O_2391,N_23677,N_21183);
xor UO_2392 (O_2392,N_29343,N_26373);
or UO_2393 (O_2393,N_29200,N_26651);
and UO_2394 (O_2394,N_29886,N_29255);
and UO_2395 (O_2395,N_24060,N_20647);
nor UO_2396 (O_2396,N_23614,N_29464);
nor UO_2397 (O_2397,N_25154,N_27697);
nand UO_2398 (O_2398,N_26666,N_23455);
nor UO_2399 (O_2399,N_21714,N_27221);
nand UO_2400 (O_2400,N_25404,N_28187);
xor UO_2401 (O_2401,N_21194,N_20280);
nor UO_2402 (O_2402,N_23776,N_21043);
xnor UO_2403 (O_2403,N_27676,N_20986);
or UO_2404 (O_2404,N_29513,N_24430);
and UO_2405 (O_2405,N_25395,N_21012);
nand UO_2406 (O_2406,N_28800,N_25297);
nand UO_2407 (O_2407,N_28393,N_20707);
or UO_2408 (O_2408,N_21199,N_20513);
nor UO_2409 (O_2409,N_26573,N_21569);
nor UO_2410 (O_2410,N_28431,N_29711);
and UO_2411 (O_2411,N_25435,N_29963);
or UO_2412 (O_2412,N_25771,N_24673);
xnor UO_2413 (O_2413,N_24339,N_28835);
and UO_2414 (O_2414,N_29700,N_22167);
nor UO_2415 (O_2415,N_23373,N_22858);
xor UO_2416 (O_2416,N_24212,N_24834);
and UO_2417 (O_2417,N_26432,N_21787);
or UO_2418 (O_2418,N_21633,N_24068);
nand UO_2419 (O_2419,N_20351,N_22555);
and UO_2420 (O_2420,N_23314,N_27348);
nor UO_2421 (O_2421,N_28553,N_26006);
or UO_2422 (O_2422,N_20393,N_28728);
or UO_2423 (O_2423,N_21832,N_20146);
nor UO_2424 (O_2424,N_25896,N_21312);
and UO_2425 (O_2425,N_29724,N_20972);
nand UO_2426 (O_2426,N_28955,N_23669);
nand UO_2427 (O_2427,N_23137,N_24588);
nand UO_2428 (O_2428,N_26279,N_21949);
nand UO_2429 (O_2429,N_26222,N_22117);
and UO_2430 (O_2430,N_21450,N_23862);
and UO_2431 (O_2431,N_20869,N_26096);
nor UO_2432 (O_2432,N_29152,N_25975);
xnor UO_2433 (O_2433,N_21297,N_23261);
and UO_2434 (O_2434,N_22329,N_20740);
nor UO_2435 (O_2435,N_28340,N_22338);
or UO_2436 (O_2436,N_21152,N_22029);
nand UO_2437 (O_2437,N_24126,N_25374);
nor UO_2438 (O_2438,N_21420,N_29986);
nand UO_2439 (O_2439,N_23775,N_29688);
nor UO_2440 (O_2440,N_23695,N_20916);
nand UO_2441 (O_2441,N_22185,N_28391);
nor UO_2442 (O_2442,N_25104,N_25823);
or UO_2443 (O_2443,N_28654,N_28114);
and UO_2444 (O_2444,N_25520,N_28113);
xnor UO_2445 (O_2445,N_23570,N_25712);
and UO_2446 (O_2446,N_25666,N_22208);
or UO_2447 (O_2447,N_27383,N_25269);
and UO_2448 (O_2448,N_28416,N_27060);
or UO_2449 (O_2449,N_20155,N_22367);
and UO_2450 (O_2450,N_23429,N_20298);
and UO_2451 (O_2451,N_20778,N_27264);
nor UO_2452 (O_2452,N_29155,N_20027);
or UO_2453 (O_2453,N_29374,N_23907);
nand UO_2454 (O_2454,N_24643,N_20067);
xor UO_2455 (O_2455,N_22194,N_22823);
nand UO_2456 (O_2456,N_26691,N_23460);
xnor UO_2457 (O_2457,N_23737,N_24150);
or UO_2458 (O_2458,N_27585,N_28179);
nand UO_2459 (O_2459,N_29092,N_20730);
xnor UO_2460 (O_2460,N_27047,N_20081);
nand UO_2461 (O_2461,N_20612,N_24665);
nand UO_2462 (O_2462,N_28306,N_26699);
nor UO_2463 (O_2463,N_20425,N_26087);
nand UO_2464 (O_2464,N_28924,N_24872);
nor UO_2465 (O_2465,N_27707,N_21434);
nor UO_2466 (O_2466,N_27440,N_25836);
nor UO_2467 (O_2467,N_25937,N_21320);
nand UO_2468 (O_2468,N_24499,N_26744);
nor UO_2469 (O_2469,N_21499,N_28719);
nand UO_2470 (O_2470,N_22573,N_22492);
nand UO_2471 (O_2471,N_29982,N_22847);
or UO_2472 (O_2472,N_20190,N_26881);
nor UO_2473 (O_2473,N_27644,N_24209);
nor UO_2474 (O_2474,N_20083,N_20438);
and UO_2475 (O_2475,N_26362,N_25900);
and UO_2476 (O_2476,N_21660,N_21426);
nand UO_2477 (O_2477,N_29814,N_21025);
or UO_2478 (O_2478,N_22683,N_20812);
xor UO_2479 (O_2479,N_28223,N_22776);
and UO_2480 (O_2480,N_21175,N_29880);
nor UO_2481 (O_2481,N_27307,N_27030);
or UO_2482 (O_2482,N_20014,N_20600);
nor UO_2483 (O_2483,N_25799,N_28138);
or UO_2484 (O_2484,N_29183,N_29416);
nor UO_2485 (O_2485,N_23870,N_24567);
and UO_2486 (O_2486,N_23881,N_28499);
nand UO_2487 (O_2487,N_22793,N_28413);
and UO_2488 (O_2488,N_22908,N_28722);
nor UO_2489 (O_2489,N_25141,N_25187);
nor UO_2490 (O_2490,N_25563,N_24048);
nor UO_2491 (O_2491,N_23001,N_26639);
and UO_2492 (O_2492,N_24037,N_28575);
or UO_2493 (O_2493,N_26680,N_22746);
nor UO_2494 (O_2494,N_27986,N_26246);
nand UO_2495 (O_2495,N_28957,N_25507);
and UO_2496 (O_2496,N_26396,N_29702);
xor UO_2497 (O_2497,N_28966,N_29328);
and UO_2498 (O_2498,N_24092,N_24635);
and UO_2499 (O_2499,N_28563,N_24186);
nand UO_2500 (O_2500,N_22716,N_21299);
or UO_2501 (O_2501,N_25941,N_27972);
or UO_2502 (O_2502,N_26605,N_25015);
nand UO_2503 (O_2503,N_27039,N_26866);
or UO_2504 (O_2504,N_23600,N_22635);
nor UO_2505 (O_2505,N_25994,N_25783);
nor UO_2506 (O_2506,N_24595,N_28744);
nor UO_2507 (O_2507,N_20237,N_23235);
or UO_2508 (O_2508,N_23236,N_23342);
nor UO_2509 (O_2509,N_23209,N_23639);
nand UO_2510 (O_2510,N_23680,N_27194);
and UO_2511 (O_2511,N_23779,N_26404);
or UO_2512 (O_2512,N_27861,N_20301);
or UO_2513 (O_2513,N_20920,N_26978);
nor UO_2514 (O_2514,N_20326,N_22676);
and UO_2515 (O_2515,N_29676,N_26402);
nor UO_2516 (O_2516,N_22540,N_20960);
nor UO_2517 (O_2517,N_25953,N_23323);
nand UO_2518 (O_2518,N_28262,N_21694);
nand UO_2519 (O_2519,N_29607,N_25804);
nand UO_2520 (O_2520,N_25113,N_26805);
nor UO_2521 (O_2521,N_22140,N_28543);
xnor UO_2522 (O_2522,N_25067,N_22335);
or UO_2523 (O_2523,N_23361,N_26118);
nand UO_2524 (O_2524,N_29778,N_25039);
and UO_2525 (O_2525,N_27619,N_26521);
nand UO_2526 (O_2526,N_24734,N_22940);
or UO_2527 (O_2527,N_23439,N_20503);
nand UO_2528 (O_2528,N_26858,N_27554);
nor UO_2529 (O_2529,N_22621,N_29872);
nand UO_2530 (O_2530,N_29204,N_27333);
or UO_2531 (O_2531,N_23978,N_23138);
or UO_2532 (O_2532,N_24831,N_21935);
nor UO_2533 (O_2533,N_21214,N_21643);
and UO_2534 (O_2534,N_23128,N_20977);
or UO_2535 (O_2535,N_21896,N_21840);
and UO_2536 (O_2536,N_28294,N_29618);
nand UO_2537 (O_2537,N_23532,N_25227);
or UO_2538 (O_2538,N_25615,N_28213);
nor UO_2539 (O_2539,N_28756,N_20569);
or UO_2540 (O_2540,N_29178,N_27526);
or UO_2541 (O_2541,N_21121,N_28072);
nand UO_2542 (O_2542,N_29334,N_24513);
nand UO_2543 (O_2543,N_28609,N_21989);
nand UO_2544 (O_2544,N_24832,N_29801);
or UO_2545 (O_2545,N_27634,N_29047);
and UO_2546 (O_2546,N_25829,N_25411);
nor UO_2547 (O_2547,N_26900,N_21268);
and UO_2548 (O_2548,N_24404,N_28400);
or UO_2549 (O_2549,N_22385,N_25529);
or UO_2550 (O_2550,N_22205,N_21631);
nand UO_2551 (O_2551,N_23113,N_21527);
nand UO_2552 (O_2552,N_24049,N_21814);
xnor UO_2553 (O_2553,N_27267,N_22837);
nor UO_2554 (O_2554,N_22041,N_21250);
nand UO_2555 (O_2555,N_20976,N_24167);
nor UO_2556 (O_2556,N_26789,N_26243);
or UO_2557 (O_2557,N_23564,N_23078);
and UO_2558 (O_2558,N_29239,N_26064);
or UO_2559 (O_2559,N_29046,N_22535);
or UO_2560 (O_2560,N_29623,N_27311);
and UO_2561 (O_2561,N_21222,N_24533);
nand UO_2562 (O_2562,N_21016,N_28264);
or UO_2563 (O_2563,N_28015,N_27699);
and UO_2564 (O_2564,N_22122,N_25962);
and UO_2565 (O_2565,N_21923,N_24350);
nor UO_2566 (O_2566,N_28122,N_28788);
or UO_2567 (O_2567,N_27020,N_29249);
and UO_2568 (O_2568,N_26973,N_25918);
or UO_2569 (O_2569,N_28617,N_21471);
xor UO_2570 (O_2570,N_27563,N_25995);
nor UO_2571 (O_2571,N_22427,N_25457);
xor UO_2572 (O_2572,N_20938,N_25165);
and UO_2573 (O_2573,N_26629,N_21507);
and UO_2574 (O_2574,N_29813,N_21050);
or UO_2575 (O_2575,N_20108,N_29169);
xor UO_2576 (O_2576,N_28780,N_24131);
nor UO_2577 (O_2577,N_29106,N_24178);
nand UO_2578 (O_2578,N_20219,N_27187);
nor UO_2579 (O_2579,N_22175,N_20024);
nand UO_2580 (O_2580,N_28690,N_25558);
or UO_2581 (O_2581,N_28274,N_23935);
and UO_2582 (O_2582,N_29277,N_28811);
or UO_2583 (O_2583,N_21727,N_23291);
xor UO_2584 (O_2584,N_29243,N_21872);
and UO_2585 (O_2585,N_21003,N_20849);
nand UO_2586 (O_2586,N_24852,N_26591);
and UO_2587 (O_2587,N_28715,N_29504);
nand UO_2588 (O_2588,N_28870,N_27358);
and UO_2589 (O_2589,N_21279,N_20705);
xnor UO_2590 (O_2590,N_22651,N_20658);
and UO_2591 (O_2591,N_21750,N_26544);
xnor UO_2592 (O_2592,N_23687,N_22237);
and UO_2593 (O_2593,N_29726,N_27122);
xor UO_2594 (O_2594,N_28440,N_25325);
nand UO_2595 (O_2595,N_22952,N_29208);
and UO_2596 (O_2596,N_23941,N_21046);
xnor UO_2597 (O_2597,N_26986,N_25245);
nand UO_2598 (O_2598,N_26143,N_22566);
or UO_2599 (O_2599,N_24095,N_21966);
xnor UO_2600 (O_2600,N_23841,N_21271);
nand UO_2601 (O_2601,N_29238,N_27155);
or UO_2602 (O_2602,N_25311,N_29014);
xor UO_2603 (O_2603,N_27601,N_26216);
or UO_2604 (O_2604,N_23387,N_20407);
and UO_2605 (O_2605,N_23916,N_27062);
or UO_2606 (O_2606,N_27432,N_26849);
or UO_2607 (O_2607,N_25889,N_22869);
nor UO_2608 (O_2608,N_26966,N_26641);
and UO_2609 (O_2609,N_22136,N_21173);
nor UO_2610 (O_2610,N_28855,N_29632);
xnor UO_2611 (O_2611,N_26913,N_25996);
nand UO_2612 (O_2612,N_23869,N_23517);
xnor UO_2613 (O_2613,N_25008,N_24523);
nor UO_2614 (O_2614,N_20313,N_20294);
nor UO_2615 (O_2615,N_23182,N_27095);
and UO_2616 (O_2616,N_23885,N_29415);
nor UO_2617 (O_2617,N_24980,N_25674);
xor UO_2618 (O_2618,N_20344,N_21269);
or UO_2619 (O_2619,N_29667,N_25761);
xor UO_2620 (O_2620,N_27274,N_29419);
nand UO_2621 (O_2621,N_24257,N_25753);
or UO_2622 (O_2622,N_22560,N_27775);
nand UO_2623 (O_2623,N_22463,N_22147);
or UO_2624 (O_2624,N_21852,N_29503);
xnor UO_2625 (O_2625,N_27659,N_22975);
nand UO_2626 (O_2626,N_28195,N_27259);
and UO_2627 (O_2627,N_20716,N_26182);
nor UO_2628 (O_2628,N_22613,N_25543);
nor UO_2629 (O_2629,N_24231,N_22980);
or UO_2630 (O_2630,N_28680,N_23127);
and UO_2631 (O_2631,N_22094,N_21195);
xnor UO_2632 (O_2632,N_24025,N_27618);
nand UO_2633 (O_2633,N_25083,N_24179);
and UO_2634 (O_2634,N_24753,N_26454);
and UO_2635 (O_2635,N_25453,N_26008);
nor UO_2636 (O_2636,N_21545,N_28051);
or UO_2637 (O_2637,N_25167,N_22784);
and UO_2638 (O_2638,N_24294,N_20978);
and UO_2639 (O_2639,N_29272,N_21109);
or UO_2640 (O_2640,N_23863,N_29017);
nand UO_2641 (O_2641,N_23886,N_24858);
nand UO_2642 (O_2642,N_25886,N_21038);
nor UO_2643 (O_2643,N_21865,N_22906);
nand UO_2644 (O_2644,N_25774,N_20325);
or UO_2645 (O_2645,N_20891,N_23825);
nor UO_2646 (O_2646,N_25389,N_27089);
and UO_2647 (O_2647,N_22123,N_23258);
or UO_2648 (O_2648,N_29611,N_28000);
nor UO_2649 (O_2649,N_28221,N_27990);
xnor UO_2650 (O_2650,N_23546,N_25214);
and UO_2651 (O_2651,N_26880,N_21246);
or UO_2652 (O_2652,N_27899,N_22490);
or UO_2653 (O_2653,N_25019,N_25087);
nand UO_2654 (O_2654,N_22718,N_28164);
and UO_2655 (O_2655,N_28317,N_26447);
xor UO_2656 (O_2656,N_25236,N_25929);
xnor UO_2657 (O_2657,N_29637,N_23002);
and UO_2658 (O_2658,N_29127,N_27099);
and UO_2659 (O_2659,N_25642,N_25162);
or UO_2660 (O_2660,N_22466,N_27391);
and UO_2661 (O_2661,N_29350,N_27935);
and UO_2662 (O_2662,N_22841,N_20274);
nor UO_2663 (O_2663,N_23715,N_28185);
xnor UO_2664 (O_2664,N_29825,N_27169);
nand UO_2665 (O_2665,N_20404,N_28662);
nand UO_2666 (O_2666,N_29036,N_28781);
and UO_2667 (O_2667,N_26586,N_25322);
nand UO_2668 (O_2668,N_26125,N_29130);
or UO_2669 (O_2669,N_25624,N_29994);
nand UO_2670 (O_2670,N_29817,N_24699);
nand UO_2671 (O_2671,N_22840,N_23435);
nor UO_2672 (O_2672,N_21681,N_27546);
nor UO_2673 (O_2673,N_28215,N_29038);
and UO_2674 (O_2674,N_29771,N_21387);
and UO_2675 (O_2675,N_25242,N_21473);
or UO_2676 (O_2676,N_21509,N_23667);
or UO_2677 (O_2677,N_25262,N_23598);
nor UO_2678 (O_2678,N_29640,N_27271);
nand UO_2679 (O_2679,N_27265,N_21208);
or UO_2680 (O_2680,N_21554,N_26807);
and UO_2681 (O_2681,N_21943,N_25968);
nor UO_2682 (O_2682,N_27368,N_26539);
or UO_2683 (O_2683,N_21921,N_28466);
xnor UO_2684 (O_2684,N_22890,N_24563);
nor UO_2685 (O_2685,N_29833,N_23796);
and UO_2686 (O_2686,N_28485,N_23495);
nand UO_2687 (O_2687,N_27574,N_26303);
xnor UO_2688 (O_2688,N_26870,N_22556);
nand UO_2689 (O_2689,N_27650,N_28087);
or UO_2690 (O_2690,N_22832,N_26862);
nor UO_2691 (O_2691,N_23089,N_29316);
nand UO_2692 (O_2692,N_23474,N_26202);
and UO_2693 (O_2693,N_28901,N_27592);
xnor UO_2694 (O_2694,N_21248,N_23004);
nand UO_2695 (O_2695,N_20304,N_24942);
nor UO_2696 (O_2696,N_28441,N_26976);
nor UO_2697 (O_2697,N_29967,N_20303);
nor UO_2698 (O_2698,N_28844,N_22586);
nor UO_2699 (O_2699,N_27373,N_25933);
and UO_2700 (O_2700,N_29636,N_23231);
nand UO_2701 (O_2701,N_26392,N_21174);
or UO_2702 (O_2702,N_28510,N_27996);
or UO_2703 (O_2703,N_23125,N_22509);
or UO_2704 (O_2704,N_26337,N_28494);
nand UO_2705 (O_2705,N_25980,N_20507);
or UO_2706 (O_2706,N_27703,N_21496);
nor UO_2707 (O_2707,N_22510,N_23924);
nor UO_2708 (O_2708,N_21559,N_21245);
xnor UO_2709 (O_2709,N_20415,N_27424);
xor UO_2710 (O_2710,N_28278,N_24984);
and UO_2711 (O_2711,N_29534,N_24102);
or UO_2712 (O_2712,N_26133,N_24174);
nand UO_2713 (O_2713,N_26726,N_24517);
nor UO_2714 (O_2714,N_24104,N_25622);
and UO_2715 (O_2715,N_26949,N_25454);
nor UO_2716 (O_2716,N_29373,N_22827);
or UO_2717 (O_2717,N_27072,N_20417);
xor UO_2718 (O_2718,N_24055,N_25296);
nand UO_2719 (O_2719,N_24214,N_22707);
nor UO_2720 (O_2720,N_21959,N_20878);
or UO_2721 (O_2721,N_20102,N_24147);
nand UO_2722 (O_2722,N_21834,N_24944);
xnor UO_2723 (O_2723,N_20073,N_20410);
and UO_2724 (O_2724,N_27615,N_23044);
xor UO_2725 (O_2725,N_20627,N_27339);
or UO_2726 (O_2726,N_27239,N_26864);
and UO_2727 (O_2727,N_29120,N_23905);
nand UO_2728 (O_2728,N_22304,N_21810);
and UO_2729 (O_2729,N_28436,N_25212);
nor UO_2730 (O_2730,N_29752,N_21695);
nor UO_2731 (O_2731,N_21544,N_26781);
nand UO_2732 (O_2732,N_25838,N_29510);
nand UO_2733 (O_2733,N_24274,N_29590);
and UO_2734 (O_2734,N_20144,N_21931);
xnor UO_2735 (O_2735,N_28126,N_23921);
and UO_2736 (O_2736,N_29365,N_21861);
or UO_2737 (O_2737,N_20557,N_25012);
xnor UO_2738 (O_2738,N_25386,N_20349);
or UO_2739 (O_2739,N_26420,N_23336);
and UO_2740 (O_2740,N_26969,N_23316);
nor UO_2741 (O_2741,N_28367,N_21951);
nand UO_2742 (O_2742,N_21080,N_24636);
nor UO_2743 (O_2743,N_27119,N_23741);
xor UO_2744 (O_2744,N_21477,N_24693);
xor UO_2745 (O_2745,N_26100,N_24558);
nor UO_2746 (O_2746,N_29256,N_29266);
or UO_2747 (O_2747,N_20055,N_21675);
xor UO_2748 (O_2748,N_22879,N_24081);
nor UO_2749 (O_2749,N_26233,N_25550);
or UO_2750 (O_2750,N_21856,N_22368);
or UO_2751 (O_2751,N_20436,N_23104);
nand UO_2752 (O_2752,N_20489,N_25741);
and UO_2753 (O_2753,N_22088,N_29774);
or UO_2754 (O_2754,N_27807,N_26272);
or UO_2755 (O_2755,N_24744,N_20675);
nand UO_2756 (O_2756,N_29125,N_21235);
nor UO_2757 (O_2757,N_25746,N_21032);
nor UO_2758 (O_2758,N_28531,N_25784);
nor UO_2759 (O_2759,N_21862,N_23855);
and UO_2760 (O_2760,N_20787,N_28914);
or UO_2761 (O_2761,N_27234,N_28322);
and UO_2762 (O_2762,N_21197,N_24929);
nor UO_2763 (O_2763,N_22880,N_23068);
or UO_2764 (O_2764,N_24073,N_27936);
nor UO_2765 (O_2765,N_20181,N_28878);
and UO_2766 (O_2766,N_27656,N_28508);
nor UO_2767 (O_2767,N_20756,N_24548);
nor UO_2768 (O_2768,N_27086,N_24771);
and UO_2769 (O_2769,N_27782,N_20156);
nand UO_2770 (O_2770,N_23672,N_23210);
and UO_2771 (O_2771,N_26046,N_26723);
or UO_2772 (O_2772,N_29557,N_20872);
or UO_2773 (O_2773,N_26490,N_22612);
and UO_2774 (O_2774,N_28509,N_28070);
nor UO_2775 (O_2775,N_23052,N_24392);
or UO_2776 (O_2776,N_24954,N_23383);
or UO_2777 (O_2777,N_25238,N_27749);
and UO_2778 (O_2778,N_26170,N_26926);
xor UO_2779 (O_2779,N_22641,N_28967);
xnor UO_2780 (O_2780,N_24847,N_22436);
and UO_2781 (O_2781,N_21393,N_20261);
nand UO_2782 (O_2782,N_29323,N_26803);
and UO_2783 (O_2783,N_21077,N_24188);
nand UO_2784 (O_2784,N_26339,N_28176);
nand UO_2785 (O_2785,N_24047,N_28535);
nand UO_2786 (O_2786,N_23756,N_24593);
or UO_2787 (O_2787,N_21905,N_23579);
or UO_2788 (O_2788,N_26491,N_21720);
nor UO_2789 (O_2789,N_21960,N_27498);
and UO_2790 (O_2790,N_24397,N_23083);
and UO_2791 (O_2791,N_27381,N_26410);
xnor UO_2792 (O_2792,N_27065,N_21620);
nor UO_2793 (O_2793,N_26138,N_20439);
nor UO_2794 (O_2794,N_29804,N_27246);
and UO_2795 (O_2795,N_23637,N_24535);
and UO_2796 (O_2796,N_23856,N_22576);
xnor UO_2797 (O_2797,N_26062,N_29533);
and UO_2798 (O_2798,N_20683,N_27834);
nand UO_2799 (O_2799,N_20725,N_20595);
nand UO_2800 (O_2800,N_23676,N_29478);
or UO_2801 (O_2801,N_29428,N_29853);
xor UO_2802 (O_2802,N_21488,N_27838);
xor UO_2803 (O_2803,N_22426,N_21745);
or UO_2804 (O_2804,N_24943,N_21611);
nor UO_2805 (O_2805,N_28183,N_26306);
xor UO_2806 (O_2806,N_25931,N_27533);
nor UO_2807 (O_2807,N_27396,N_22238);
and UO_2808 (O_2808,N_25758,N_26427);
or UO_2809 (O_2809,N_22212,N_22787);
nand UO_2810 (O_2810,N_22624,N_27751);
xor UO_2811 (O_2811,N_22900,N_26461);
or UO_2812 (O_2812,N_27954,N_21671);
or UO_2813 (O_2813,N_27827,N_27929);
nand UO_2814 (O_2814,N_21649,N_27977);
and UO_2815 (O_2815,N_23927,N_21566);
and UO_2816 (O_2816,N_29796,N_24280);
or UO_2817 (O_2817,N_23879,N_24803);
nor UO_2818 (O_2818,N_22983,N_27363);
nor UO_2819 (O_2819,N_24998,N_21560);
or UO_2820 (O_2820,N_28732,N_22932);
nand UO_2821 (O_2821,N_25542,N_22095);
xnor UO_2822 (O_2822,N_28987,N_21957);
or UO_2823 (O_2823,N_22158,N_26550);
nand UO_2824 (O_2824,N_20903,N_22825);
nor UO_2825 (O_2825,N_24759,N_22046);
nor UO_2826 (O_2826,N_25153,N_22762);
nand UO_2827 (O_2827,N_22200,N_22272);
and UO_2828 (O_2828,N_21057,N_22265);
nand UO_2829 (O_2829,N_28290,N_29602);
or UO_2830 (O_2830,N_21333,N_21679);
xnor UO_2831 (O_2831,N_24967,N_26121);
or UO_2832 (O_2832,N_23349,N_27874);
and UO_2833 (O_2833,N_23386,N_27114);
or UO_2834 (O_2834,N_26482,N_21774);
and UO_2835 (O_2835,N_24779,N_27255);
nor UO_2836 (O_2836,N_22623,N_24557);
and UO_2837 (O_2837,N_25146,N_24681);
or UO_2838 (O_2838,N_27487,N_22439);
nor UO_2839 (O_2839,N_26127,N_28149);
or UO_2840 (O_2840,N_27458,N_27382);
nand UO_2841 (O_2841,N_28682,N_23536);
or UO_2842 (O_2842,N_21976,N_28665);
xor UO_2843 (O_2843,N_29791,N_21590);
xnor UO_2844 (O_2844,N_23552,N_25855);
and UO_2845 (O_2845,N_29719,N_29644);
nand UO_2846 (O_2846,N_21295,N_28822);
nand UO_2847 (O_2847,N_21838,N_26793);
or UO_2848 (O_2848,N_20738,N_24781);
nand UO_2849 (O_2849,N_22771,N_24889);
nor UO_2850 (O_2850,N_23049,N_27064);
nand UO_2851 (O_2851,N_28865,N_24516);
or UO_2852 (O_2852,N_25339,N_24719);
and UO_2853 (O_2853,N_21433,N_26538);
or UO_2854 (O_2854,N_26114,N_25128);
and UO_2855 (O_2855,N_20590,N_23931);
or UO_2856 (O_2856,N_22830,N_20252);
xor UO_2857 (O_2857,N_23889,N_20184);
or UO_2858 (O_2858,N_21839,N_21040);
and UO_2859 (O_2859,N_25073,N_25863);
or UO_2860 (O_2860,N_22156,N_24192);
nor UO_2861 (O_2861,N_22859,N_23229);
nand UO_2862 (O_2862,N_29245,N_25749);
or UO_2863 (O_2863,N_26925,N_25924);
nor UO_2864 (O_2864,N_20145,N_24978);
nor UO_2865 (O_2865,N_24099,N_21758);
and UO_2866 (O_2866,N_21998,N_21819);
and UO_2867 (O_2867,N_27048,N_27567);
or UO_2868 (O_2868,N_25815,N_20493);
nor UO_2869 (O_2869,N_28243,N_28938);
or UO_2870 (O_2870,N_25476,N_23196);
nand UO_2871 (O_2871,N_20257,N_22193);
nand UO_2872 (O_2872,N_26073,N_29296);
and UO_2873 (O_2873,N_23801,N_20246);
or UO_2874 (O_2874,N_27050,N_27675);
xor UO_2875 (O_2875,N_29917,N_26783);
or UO_2876 (O_2876,N_24877,N_25119);
nor UO_2877 (O_2877,N_24974,N_28827);
or UO_2878 (O_2878,N_25820,N_24218);
nand UO_2879 (O_2879,N_20900,N_27046);
or UO_2880 (O_2880,N_24860,N_24090);
nor UO_2881 (O_2881,N_22528,N_21400);
nor UO_2882 (O_2882,N_20222,N_22220);
and UO_2883 (O_2883,N_26944,N_20287);
or UO_2884 (O_2884,N_20895,N_29650);
and UO_2885 (O_2885,N_29497,N_25222);
nor UO_2886 (O_2886,N_20159,N_29430);
xor UO_2887 (O_2887,N_29094,N_27057);
nand UO_2888 (O_2888,N_28872,N_23861);
nand UO_2889 (O_2889,N_20367,N_22348);
and UO_2890 (O_2890,N_27921,N_21726);
and UO_2891 (O_2891,N_20473,N_21464);
nand UO_2892 (O_2892,N_25092,N_27519);
or UO_2893 (O_2893,N_27288,N_26416);
nand UO_2894 (O_2894,N_23699,N_21189);
and UO_2895 (O_2895,N_20292,N_24702);
nor UO_2896 (O_2896,N_23682,N_28216);
nor UO_2897 (O_2897,N_28708,N_24598);
nand UO_2898 (O_2898,N_27593,N_28755);
and UO_2899 (O_2899,N_28661,N_20288);
and UO_2900 (O_2900,N_27094,N_22820);
and UO_2901 (O_2901,N_21100,N_21167);
and UO_2902 (O_2902,N_20648,N_22554);
nand UO_2903 (O_2903,N_29866,N_25241);
and UO_2904 (O_2904,N_23217,N_24364);
nor UO_2905 (O_2905,N_28527,N_27692);
nand UO_2906 (O_2906,N_24059,N_21052);
nand UO_2907 (O_2907,N_24449,N_20784);
nor UO_2908 (O_2908,N_20970,N_24148);
nand UO_2909 (O_2909,N_25266,N_29777);
or UO_2910 (O_2910,N_26156,N_26377);
nand UO_2911 (O_2911,N_29840,N_26924);
or UO_2912 (O_2912,N_20529,N_26822);
or UO_2913 (O_2913,N_25677,N_21277);
nor UO_2914 (O_2914,N_29646,N_29045);
or UO_2915 (O_2915,N_26383,N_22313);
or UO_2916 (O_2916,N_28576,N_25185);
xor UO_2917 (O_2917,N_23205,N_24785);
nor UO_2918 (O_2918,N_22064,N_27335);
nor UO_2919 (O_2919,N_24242,N_21637);
nand UO_2920 (O_2920,N_23162,N_23872);
and UO_2921 (O_2921,N_26332,N_22608);
nor UO_2922 (O_2922,N_22396,N_26443);
or UO_2923 (O_2923,N_24017,N_21849);
xor UO_2924 (O_2924,N_22098,N_21030);
or UO_2925 (O_2925,N_21072,N_24962);
or UO_2926 (O_2926,N_24886,N_22177);
nand UO_2927 (O_2927,N_21134,N_26583);
nor UO_2928 (O_2928,N_27425,N_25288);
and UO_2929 (O_2929,N_22685,N_27386);
nor UO_2930 (O_2930,N_21585,N_22938);
nand UO_2931 (O_2931,N_26876,N_25623);
or UO_2932 (O_2932,N_25708,N_26882);
xnor UO_2933 (O_2933,N_27101,N_27597);
and UO_2934 (O_2934,N_23814,N_22518);
nand UO_2935 (O_2935,N_26596,N_29451);
xnor UO_2936 (O_2936,N_20440,N_27428);
nor UO_2937 (O_2937,N_26609,N_23096);
or UO_2938 (O_2938,N_23119,N_28333);
nand UO_2939 (O_2939,N_21738,N_24861);
nand UO_2940 (O_2940,N_20698,N_22694);
nand UO_2941 (O_2941,N_25597,N_26530);
xor UO_2942 (O_2942,N_20053,N_23902);
and UO_2943 (O_2943,N_21903,N_29808);
nand UO_2944 (O_2944,N_21956,N_29023);
nand UO_2945 (O_2945,N_20593,N_22384);
and UO_2946 (O_2946,N_22792,N_25366);
and UO_2947 (O_2947,N_24419,N_27857);
or UO_2948 (O_2948,N_29300,N_22405);
and UO_2949 (O_2949,N_23274,N_23090);
nor UO_2950 (O_2950,N_21864,N_25392);
nor UO_2951 (O_2951,N_25664,N_20251);
nand UO_2952 (O_2952,N_25327,N_28077);
nand UO_2953 (O_2953,N_25318,N_20342);
nor UO_2954 (O_2954,N_26622,N_23572);
nand UO_2955 (O_2955,N_20546,N_23854);
nand UO_2956 (O_2956,N_27539,N_29785);
nor UO_2957 (O_2957,N_23778,N_22553);
nand UO_2958 (O_2958,N_20006,N_27805);
and UO_2959 (O_2959,N_25534,N_24180);
nand UO_2960 (O_2960,N_24311,N_20306);
or UO_2961 (O_2961,N_25148,N_23799);
and UO_2962 (O_2962,N_20688,N_29609);
nor UO_2963 (O_2963,N_25081,N_28170);
nand UO_2964 (O_2964,N_26498,N_22440);
nor UO_2965 (O_2965,N_27196,N_24414);
and UO_2966 (O_2966,N_21475,N_27974);
xor UO_2967 (O_2967,N_22753,N_22093);
and UO_2968 (O_2968,N_21619,N_25068);
and UO_2969 (O_2969,N_25764,N_28348);
nand UO_2970 (O_2970,N_26935,N_24931);
nor UO_2971 (O_2971,N_22197,N_25207);
or UO_2972 (O_2972,N_26021,N_27162);
and UO_2973 (O_2973,N_20084,N_28203);
and UO_2974 (O_2974,N_22995,N_24625);
and UO_2975 (O_2975,N_25481,N_25145);
and UO_2976 (O_2976,N_22001,N_28679);
nand UO_2977 (O_2977,N_22410,N_21942);
nand UO_2978 (O_2978,N_20141,N_26782);
nand UO_2979 (O_2979,N_28763,N_25775);
nand UO_2980 (O_2980,N_26690,N_25156);
nand UO_2981 (O_2981,N_22512,N_20132);
xor UO_2982 (O_2982,N_23484,N_29936);
and UO_2983 (O_2983,N_26645,N_21614);
nor UO_2984 (O_2984,N_23352,N_22704);
and UO_2985 (O_2985,N_29604,N_20263);
and UO_2986 (O_2986,N_29729,N_20187);
and UO_2987 (O_2987,N_22114,N_21549);
or UO_2988 (O_2988,N_21672,N_26439);
or UO_2989 (O_2989,N_21461,N_28863);
and UO_2990 (O_2990,N_29306,N_26072);
nor UO_2991 (O_2991,N_25489,N_21680);
nor UO_2992 (O_2992,N_26816,N_26771);
nor UO_2993 (O_2993,N_24569,N_25021);
nand UO_2994 (O_2994,N_23141,N_21122);
nand UO_2995 (O_2995,N_25797,N_23817);
xnor UO_2996 (O_2996,N_29507,N_26891);
nand UO_2997 (O_2997,N_21421,N_26842);
or UO_2998 (O_2998,N_21383,N_29977);
and UO_2999 (O_2999,N_27464,N_27054);
nor UO_3000 (O_3000,N_28821,N_24638);
or UO_3001 (O_3001,N_27638,N_28911);
nor UO_3002 (O_3002,N_23269,N_21107);
nor UO_3003 (O_3003,N_28660,N_29684);
nor UO_3004 (O_3004,N_28711,N_23787);
nor UO_3005 (O_3005,N_22372,N_26854);
or UO_3006 (O_3006,N_25805,N_25018);
nand UO_3007 (O_3007,N_29071,N_26780);
nor UO_3008 (O_3008,N_24342,N_26290);
nand UO_3009 (O_3009,N_21172,N_27922);
nand UO_3010 (O_3010,N_21166,N_26627);
and UO_3011 (O_3011,N_27892,N_24435);
xnor UO_3012 (O_3012,N_26283,N_25652);
xnor UO_3013 (O_3013,N_25219,N_21890);
and UO_3014 (O_3014,N_20071,N_22835);
xnor UO_3015 (O_3015,N_26423,N_25780);
nor UO_3016 (O_3016,N_28477,N_22477);
nor UO_3017 (O_3017,N_28549,N_21625);
nor UO_3018 (O_3018,N_29895,N_26205);
and UO_3019 (O_3019,N_29680,N_29829);
or UO_3020 (O_3020,N_24662,N_27912);
nor UO_3021 (O_3021,N_21584,N_28754);
and UO_3022 (O_3022,N_24922,N_26195);
nor UO_3023 (O_3023,N_22486,N_21601);
nor UO_3024 (O_3024,N_25467,N_24876);
or UO_3025 (O_3025,N_23826,N_28008);
nor UO_3026 (O_3026,N_29457,N_29336);
and UO_3027 (O_3027,N_28120,N_22666);
xnor UO_3028 (O_3028,N_26374,N_27168);
or UO_3029 (O_3029,N_21691,N_21947);
nor UO_3030 (O_3030,N_23888,N_28124);
or UO_3031 (O_3031,N_29005,N_26180);
or UO_3032 (O_3032,N_22144,N_28171);
or UO_3033 (O_3033,N_27317,N_29705);
or UO_3034 (O_3034,N_28148,N_28389);
or UO_3035 (O_3035,N_29221,N_23527);
or UO_3036 (O_3036,N_23331,N_20946);
xnor UO_3037 (O_3037,N_23576,N_27696);
or UO_3038 (O_3038,N_27336,N_23427);
and UO_3039 (O_3039,N_23987,N_28300);
nand UO_3040 (O_3040,N_25791,N_23958);
nor UO_3041 (O_3041,N_20640,N_26626);
or UO_3042 (O_3042,N_29725,N_26361);
nand UO_3043 (O_3043,N_22120,N_21692);
and UO_3044 (O_3044,N_21676,N_27015);
or UO_3045 (O_3045,N_28098,N_21439);
or UO_3046 (O_3046,N_29488,N_27907);
nor UO_3047 (O_3047,N_28449,N_24904);
or UO_3048 (O_3048,N_27465,N_29819);
nand UO_3049 (O_3049,N_22739,N_23322);
nor UO_3050 (O_3050,N_27006,N_28097);
xnor UO_3051 (O_3051,N_25504,N_28947);
nor UO_3052 (O_3052,N_21991,N_22866);
or UO_3053 (O_3053,N_24873,N_24884);
nand UO_3054 (O_3054,N_26811,N_28110);
or UO_3055 (O_3055,N_23568,N_28806);
and UO_3056 (O_3056,N_22728,N_23766);
nor UO_3057 (O_3057,N_29022,N_25511);
and UO_3058 (O_3058,N_21516,N_27420);
nand UO_3059 (O_3059,N_27098,N_25660);
and UO_3060 (O_3060,N_20739,N_27500);
xor UO_3061 (O_3061,N_26533,N_26113);
xor UO_3062 (O_3062,N_28045,N_29391);
xor UO_3063 (O_3063,N_24721,N_20161);
and UO_3064 (O_3064,N_23222,N_26604);
and UO_3065 (O_3065,N_22559,N_26889);
nor UO_3066 (O_3066,N_20690,N_25641);
and UO_3067 (O_3067,N_22054,N_25646);
and UO_3068 (O_3068,N_25075,N_20642);
or UO_3069 (O_3069,N_25927,N_23822);
xor UO_3070 (O_3070,N_29716,N_23237);
nand UO_3071 (O_3071,N_20347,N_23241);
nand UO_3072 (O_3072,N_23109,N_23135);
nor UO_3073 (O_3073,N_29755,N_24667);
or UO_3074 (O_3074,N_20138,N_28355);
and UO_3075 (O_3075,N_22273,N_22132);
and UO_3076 (O_3076,N_22181,N_28673);
or UO_3077 (O_3077,N_22797,N_25237);
nand UO_3078 (O_3078,N_29070,N_26587);
and UO_3079 (O_3079,N_24462,N_23520);
or UO_3080 (O_3080,N_22563,N_20432);
xor UO_3081 (O_3081,N_29481,N_22327);
nor UO_3082 (O_3082,N_27027,N_24278);
nand UO_3083 (O_3083,N_28551,N_25539);
nor UO_3084 (O_3084,N_29235,N_28433);
and UO_3085 (O_3085,N_29942,N_20949);
nand UO_3086 (O_3086,N_27580,N_21836);
or UO_3087 (O_3087,N_22404,N_22083);
xor UO_3088 (O_3088,N_22920,N_29440);
nor UO_3089 (O_3089,N_24937,N_20687);
xnor UO_3090 (O_3090,N_28128,N_28619);
nand UO_3091 (O_3091,N_24220,N_22929);
or UO_3092 (O_3092,N_25557,N_29959);
nor UO_3093 (O_3093,N_23760,N_24589);
nand UO_3094 (O_3094,N_24475,N_20511);
and UO_3095 (O_3095,N_26990,N_21768);
nand UO_3096 (O_3096,N_27195,N_25107);
or UO_3097 (O_3097,N_26548,N_22176);
nand UO_3098 (O_3098,N_23431,N_29556);
and UO_3099 (O_3099,N_28165,N_23736);
or UO_3100 (O_3100,N_23305,N_21734);
nand UO_3101 (O_3101,N_26193,N_20063);
nand UO_3102 (O_3102,N_24787,N_27598);
and UO_3103 (O_3103,N_29366,N_22852);
and UO_3104 (O_3104,N_27276,N_20855);
and UO_3105 (O_3105,N_29118,N_22412);
nand UO_3106 (O_3106,N_26559,N_28799);
xor UO_3107 (O_3107,N_23140,N_20273);
nor UO_3108 (O_3108,N_20572,N_23865);
nor UO_3109 (O_3109,N_23937,N_22061);
or UO_3110 (O_3110,N_26821,N_21135);
or UO_3111 (O_3111,N_27768,N_28614);
nand UO_3112 (O_3112,N_29854,N_24621);
or UO_3113 (O_3113,N_27931,N_20840);
nand UO_3114 (O_3114,N_25979,N_25054);
and UO_3115 (O_3115,N_26310,N_20502);
nand UO_3116 (O_3116,N_26495,N_21752);
and UO_3117 (O_3117,N_26918,N_23362);
nor UO_3118 (O_3118,N_27153,N_28146);
or UO_3119 (O_3119,N_23276,N_28717);
and UO_3120 (O_3120,N_25066,N_22730);
xnor UO_3121 (O_3121,N_27918,N_28839);
and UO_3122 (O_3122,N_25353,N_24230);
and UO_3123 (O_3123,N_26026,N_23804);
and UO_3124 (O_3124,N_24076,N_23624);
nand UO_3125 (O_3125,N_23131,N_27965);
or UO_3126 (O_3126,N_21878,N_28956);
nand UO_3127 (O_3127,N_25785,N_25451);
and UO_3128 (O_3128,N_20818,N_24139);
nor UO_3129 (O_3129,N_23661,N_23859);
nand UO_3130 (O_3130,N_27233,N_21160);
nand UO_3131 (O_3131,N_20789,N_21596);
nor UO_3132 (O_3132,N_26844,N_21837);
nor UO_3133 (O_3133,N_26269,N_29798);
nand UO_3134 (O_3134,N_20629,N_22807);
nand UO_3135 (O_3135,N_24349,N_25715);
or UO_3136 (O_3136,N_29000,N_27277);
and UO_3137 (O_3137,N_29140,N_25566);
nor UO_3138 (O_3138,N_26398,N_27587);
nand UO_3139 (O_3139,N_22727,N_22255);
xor UO_3140 (O_3140,N_24615,N_21741);
and UO_3141 (O_3141,N_21293,N_25598);
nand UO_3142 (O_3142,N_23434,N_22741);
and UO_3143 (O_3143,N_29559,N_29061);
and UO_3144 (O_3144,N_25777,N_22308);
nand UO_3145 (O_3145,N_28455,N_27772);
nand UO_3146 (O_3146,N_29553,N_29915);
or UO_3147 (O_3147,N_28134,N_26715);
nand UO_3148 (O_3148,N_21563,N_28052);
nor UO_3149 (O_3149,N_27826,N_23414);
or UO_3150 (O_3150,N_22332,N_25611);
nand UO_3151 (O_3151,N_23878,N_21311);
xnor UO_3152 (O_3152,N_23690,N_20259);
nor UO_3153 (O_3153,N_20382,N_26840);
and UO_3154 (O_3154,N_27837,N_27923);
nor UO_3155 (O_3155,N_21229,N_29720);
or UO_3156 (O_3156,N_26262,N_21193);
or UO_3157 (O_3157,N_20584,N_27613);
nor UO_3158 (O_3158,N_22769,N_29799);
nor UO_3159 (O_3159,N_22575,N_23551);
or UO_3160 (O_3160,N_26251,N_20460);
nor UO_3161 (O_3161,N_28861,N_22012);
nand UO_3162 (O_3162,N_22005,N_27281);
xnor UO_3163 (O_3163,N_20791,N_21446);
nor UO_3164 (O_3164,N_21910,N_23206);
and UO_3165 (O_3165,N_27438,N_26042);
nand UO_3166 (O_3166,N_28487,N_22942);
xnor UO_3167 (O_3167,N_23652,N_26391);
and UO_3168 (O_3168,N_28152,N_20526);
xor UO_3169 (O_3169,N_24351,N_25194);
or UO_3170 (O_3170,N_27691,N_28641);
nand UO_3171 (O_3171,N_27753,N_21575);
nor UO_3172 (O_3172,N_21329,N_24327);
and UO_3173 (O_3173,N_27530,N_21505);
nor UO_3174 (O_3174,N_26014,N_26507);
nor UO_3175 (O_3175,N_21656,N_21130);
nor UO_3176 (O_3176,N_25684,N_27331);
xnor UO_3177 (O_3177,N_20235,N_22325);
nor UO_3178 (O_3178,N_26356,N_24396);
or UO_3179 (O_3179,N_27535,N_22121);
nor UO_3180 (O_3180,N_23134,N_28007);
nor UO_3181 (O_3181,N_27309,N_24822);
nand UO_3182 (O_3182,N_23686,N_27576);
nor UO_3183 (O_3183,N_28256,N_21272);
nand UO_3184 (O_3184,N_22502,N_22264);
xnor UO_3185 (O_3185,N_22924,N_22460);
or UO_3186 (O_3186,N_29606,N_22925);
nand UO_3187 (O_3187,N_20947,N_22947);
or UO_3188 (O_3188,N_22584,N_23606);
nor UO_3189 (O_3189,N_22974,N_20704);
xnor UO_3190 (O_3190,N_28273,N_26875);
and UO_3191 (O_3191,N_29121,N_21360);
or UO_3192 (O_3192,N_20137,N_25293);
and UO_3193 (O_3193,N_21428,N_23343);
nand UO_3194 (O_3194,N_26898,N_25070);
or UO_3195 (O_3195,N_29768,N_21740);
and UO_3196 (O_3196,N_22314,N_29916);
and UO_3197 (O_3197,N_27969,N_29848);
nand UO_3198 (O_3198,N_21593,N_28156);
and UO_3199 (O_3199,N_27299,N_20485);
and UO_3200 (O_3200,N_20713,N_27803);
and UO_3201 (O_3201,N_25305,N_20461);
nor UO_3202 (O_3202,N_29536,N_27491);
and UO_3203 (O_3203,N_26331,N_23493);
nand UO_3204 (O_3204,N_21170,N_20017);
nor UO_3205 (O_3205,N_28064,N_26105);
and UO_3206 (O_3206,N_22442,N_21589);
or UO_3207 (O_3207,N_20327,N_26446);
nand UO_3208 (O_3208,N_21090,N_29971);
nand UO_3209 (O_3209,N_29404,N_23053);
xnor UO_3210 (O_3210,N_23491,N_25013);
nor UO_3211 (O_3211,N_21658,N_29822);
or UO_3212 (O_3212,N_21027,N_20395);
nand UO_3213 (O_3213,N_21533,N_25604);
nand UO_3214 (O_3214,N_26893,N_20177);
nor UO_3215 (O_3215,N_26386,N_23218);
nor UO_3216 (O_3216,N_21079,N_27684);
xor UO_3217 (O_3217,N_22004,N_24527);
or UO_3218 (O_3218,N_28121,N_24526);
nand UO_3219 (O_3219,N_22216,N_28666);
or UO_3220 (O_3220,N_28167,N_20074);
or UO_3221 (O_3221,N_28975,N_21763);
and UO_3222 (O_3222,N_26993,N_25982);
nand UO_3223 (O_3223,N_25821,N_28917);
nand UO_3224 (O_3224,N_23744,N_29280);
and UO_3225 (O_3225,N_23490,N_21668);
and UO_3226 (O_3226,N_28577,N_28573);
and UO_3227 (O_3227,N_21396,N_24018);
nor UO_3228 (O_3228,N_29308,N_25252);
and UO_3229 (O_3229,N_28533,N_27473);
and UO_3230 (O_3230,N_29203,N_23428);
or UO_3231 (O_3231,N_25959,N_27296);
nand UO_3232 (O_3232,N_20247,N_23636);
nor UO_3233 (O_3233,N_26951,N_24053);
nor UO_3234 (O_3234,N_20174,N_21094);
or UO_3235 (O_3235,N_24249,N_20127);
nand UO_3236 (O_3236,N_21125,N_21875);
nor UO_3237 (O_3237,N_26344,N_25432);
and UO_3238 (O_3238,N_22909,N_21318);
or UO_3239 (O_3239,N_20923,N_25917);
and UO_3240 (O_3240,N_25748,N_28589);
xor UO_3241 (O_3241,N_29645,N_20547);
nor UO_3242 (O_3242,N_25123,N_24697);
or UO_3243 (O_3243,N_23368,N_28585);
or UO_3244 (O_3244,N_25965,N_27230);
or UO_3245 (O_3245,N_25317,N_22186);
or UO_3246 (O_3246,N_23103,N_22516);
nor UO_3247 (O_3247,N_25256,N_29307);
or UO_3248 (O_3248,N_26311,N_20592);
and UO_3249 (O_3249,N_27330,N_25825);
nor UO_3250 (O_3250,N_25714,N_27937);
nand UO_3251 (O_3251,N_20369,N_22594);
nor UO_3252 (O_3252,N_21289,N_20662);
and UO_3253 (O_3253,N_21613,N_29095);
xnor UO_3254 (O_3254,N_27603,N_29865);
nand UO_3255 (O_3255,N_28212,N_28251);
xor UO_3256 (O_3256,N_24493,N_22174);
and UO_3257 (O_3257,N_29491,N_28200);
xor UO_3258 (O_3258,N_27661,N_21296);
and UO_3259 (O_3259,N_29531,N_28042);
xnor UO_3260 (O_3260,N_21635,N_21930);
or UO_3261 (O_3261,N_23413,N_21769);
or UO_3262 (O_3262,N_21066,N_28567);
nor UO_3263 (O_3263,N_28026,N_25329);
and UO_3264 (O_3264,N_24344,N_20481);
nand UO_3265 (O_3265,N_24755,N_29189);
nor UO_3266 (O_3266,N_24335,N_21290);
and UO_3267 (O_3267,N_27916,N_26856);
xor UO_3268 (O_3268,N_28596,N_23689);
nor UO_3269 (O_3269,N_24991,N_26838);
and UO_3270 (O_3270,N_29542,N_23171);
nand UO_3271 (O_3271,N_26975,N_27441);
or UO_3272 (O_3272,N_20734,N_22917);
nor UO_3273 (O_3273,N_26163,N_20531);
and UO_3274 (O_3274,N_21707,N_25638);
nor UO_3275 (O_3275,N_28866,N_22479);
nand UO_3276 (O_3276,N_21542,N_24483);
and UO_3277 (O_3277,N_29082,N_21753);
nor UO_3278 (O_3278,N_22808,N_21146);
nor UO_3279 (O_3279,N_21595,N_20339);
or UO_3280 (O_3280,N_26210,N_26477);
nor UO_3281 (O_3281,N_25149,N_25446);
and UO_3282 (O_3282,N_22317,N_26334);
or UO_3283 (O_3283,N_27688,N_22950);
xnor UO_3284 (O_3284,N_28909,N_20171);
and UO_3285 (O_3285,N_22108,N_27607);
nand UO_3286 (O_3286,N_27007,N_20194);
nor UO_3287 (O_3287,N_28643,N_21139);
and UO_3288 (O_3288,N_28181,N_26200);
nor UO_3289 (O_3289,N_25513,N_20258);
or UO_3290 (O_3290,N_29386,N_23271);
and UO_3291 (O_3291,N_20948,N_21200);
or UO_3292 (O_3292,N_22921,N_25901);
nor UO_3293 (O_3293,N_21319,N_21952);
or UO_3294 (O_3294,N_28082,N_22587);
and UO_3295 (O_3295,N_20714,N_20760);
nor UO_3296 (O_3296,N_23177,N_25722);
nand UO_3297 (O_3297,N_22860,N_20183);
nor UO_3298 (O_3298,N_23442,N_23069);
xor UO_3299 (O_3299,N_24031,N_21605);
or UO_3300 (O_3300,N_29815,N_29851);
and UO_3301 (O_3301,N_23031,N_25144);
nor UO_3302 (O_3302,N_24686,N_20035);
xor UO_3303 (O_3303,N_20606,N_23758);
nor UO_3304 (O_3304,N_21044,N_20798);
and UO_3305 (O_3305,N_25316,N_29458);
or UO_3306 (O_3306,N_29156,N_25842);
or UO_3307 (O_3307,N_27651,N_27718);
or UO_3308 (O_3308,N_29331,N_24823);
and UO_3309 (O_3309,N_20297,N_20639);
nor UO_3310 (O_3310,N_27092,N_21292);
xnor UO_3311 (O_3311,N_28703,N_20570);
and UO_3312 (O_3312,N_25503,N_28048);
or UO_3313 (O_3313,N_24529,N_25372);
and UO_3314 (O_3314,N_25247,N_23219);
nand UO_3315 (O_3315,N_28266,N_21822);
nand UO_3316 (O_3316,N_28704,N_29655);
or UO_3317 (O_3317,N_29063,N_27127);
nor UO_3318 (O_3318,N_24672,N_22159);
or UO_3319 (O_3319,N_29876,N_24594);
nand UO_3320 (O_3320,N_25150,N_21380);
nor UO_3321 (O_3321,N_22801,N_28503);
and UO_3322 (O_3322,N_26174,N_26823);
or UO_3323 (O_3323,N_20579,N_26790);
or UO_3324 (O_3324,N_20153,N_23662);
nand UO_3325 (O_3325,N_21054,N_21665);
xnor UO_3326 (O_3326,N_28252,N_25455);
or UO_3327 (O_3327,N_29337,N_27932);
and UO_3328 (O_3328,N_28555,N_28267);
or UO_3329 (O_3329,N_22478,N_20267);
or UO_3330 (O_3330,N_24466,N_25388);
xor UO_3331 (O_3331,N_29775,N_24816);
nand UO_3332 (O_3332,N_27421,N_28687);
xnor UO_3333 (O_3333,N_22736,N_29029);
or UO_3334 (O_3334,N_28969,N_29496);
and UO_3335 (O_3335,N_25692,N_21574);
or UO_3336 (O_3336,N_23632,N_28047);
or UO_3337 (O_3337,N_28163,N_26102);
or UO_3338 (O_3338,N_26754,N_25452);
nand UO_3339 (O_3339,N_23830,N_20602);
nor UO_3340 (O_3340,N_20049,N_20896);
nand UO_3341 (O_3341,N_20764,N_21395);
and UO_3342 (O_3342,N_26232,N_24891);
nand UO_3343 (O_3343,N_23476,N_27758);
nor UO_3344 (O_3344,N_23481,N_26085);
or UO_3345 (O_3345,N_20464,N_27564);
nand UO_3346 (O_3346,N_21876,N_29682);
xor UO_3347 (O_3347,N_28281,N_25486);
or UO_3348 (O_3348,N_27202,N_20012);
and UO_3349 (O_3349,N_25617,N_26894);
xor UO_3350 (O_3350,N_26098,N_24907);
xor UO_3351 (O_3351,N_29893,N_25731);
nor UO_3352 (O_3352,N_25669,N_23260);
nor UO_3353 (O_3353,N_20693,N_29647);
nand UO_3354 (O_3354,N_22242,N_28761);
xnor UO_3355 (O_3355,N_25033,N_22127);
nand UO_3356 (O_3356,N_23284,N_23270);
or UO_3357 (O_3357,N_29067,N_26212);
and UO_3358 (O_3358,N_25832,N_29909);
xor UO_3359 (O_3359,N_27160,N_23485);
or UO_3360 (O_3360,N_23277,N_29259);
nand UO_3361 (O_3361,N_23470,N_25295);
nor UO_3362 (O_3362,N_28312,N_25893);
nor UO_3363 (O_3363,N_21020,N_29925);
nor UO_3364 (O_3364,N_26069,N_20874);
and UO_3365 (O_3365,N_28428,N_21731);
and UO_3366 (O_3366,N_20628,N_21781);
nand UO_3367 (O_3367,N_20621,N_21754);
nand UO_3368 (O_3368,N_27581,N_24634);
and UO_3369 (O_3369,N_21247,N_24885);
or UO_3370 (O_3370,N_27036,N_27665);
and UO_3371 (O_3371,N_21717,N_29487);
or UO_3372 (O_3372,N_23094,N_20892);
and UO_3373 (O_3373,N_26501,N_27612);
and UO_3374 (O_3374,N_26380,N_24260);
nand UO_3375 (O_3375,N_23625,N_22059);
nor UO_3376 (O_3376,N_25377,N_25134);
or UO_3377 (O_3377,N_26916,N_21163);
nor UO_3378 (O_3378,N_29529,N_26329);
nor UO_3379 (O_3379,N_29133,N_22399);
and UO_3380 (O_3380,N_20129,N_23244);
nor UO_3381 (O_3381,N_23034,N_26619);
nand UO_3382 (O_3382,N_27850,N_25695);
or UO_3383 (O_3383,N_20676,N_28572);
or UO_3384 (O_3384,N_22246,N_28526);
nand UO_3385 (O_3385,N_26110,N_22228);
and UO_3386 (O_3386,N_26047,N_28206);
or UO_3387 (O_3387,N_20272,N_23605);
nand UO_3388 (O_3388,N_23573,N_26809);
nand UO_3389 (O_3389,N_29320,N_28559);
xor UO_3390 (O_3390,N_29933,N_27149);
nand UO_3391 (O_3391,N_25778,N_29342);
or UO_3392 (O_3392,N_24578,N_27726);
and UO_3393 (O_3393,N_29989,N_26239);
nand UO_3394 (O_3394,N_21525,N_24138);
or UO_3395 (O_3395,N_28930,N_24149);
nor UO_3396 (O_3396,N_27831,N_28562);
nor UO_3397 (O_3397,N_28752,N_25899);
and UO_3398 (O_3398,N_28595,N_20197);
and UO_3399 (O_3399,N_22287,N_27154);
or UO_3400 (O_3400,N_23327,N_20661);
nand UO_3401 (O_3401,N_24172,N_22301);
and UO_3402 (O_3402,N_27404,N_23524);
nand UO_3403 (O_3403,N_21733,N_21788);
nor UO_3404 (O_3404,N_27759,N_27451);
and UO_3405 (O_3405,N_25474,N_25397);
nor UO_3406 (O_3406,N_21137,N_20536);
or UO_3407 (O_3407,N_21340,N_25913);
or UO_3408 (O_3408,N_27238,N_22734);
and UO_3409 (O_3409,N_24605,N_26601);
nor UO_3410 (O_3410,N_21667,N_28489);
and UO_3411 (O_3411,N_27957,N_27904);
nand UO_3412 (O_3412,N_28101,N_23154);
nand UO_3413 (O_3413,N_24228,N_21724);
nand UO_3414 (O_3414,N_23451,N_24038);
nand UO_3415 (O_3415,N_29424,N_20203);
nor UO_3416 (O_3416,N_26320,N_29844);
xnor UO_3417 (O_3417,N_29582,N_29758);
nor UO_3418 (O_3418,N_24199,N_29132);
nand UO_3419 (O_3419,N_24243,N_23382);
nand UO_3420 (O_3420,N_28895,N_24968);
nor UO_3421 (O_3421,N_20227,N_20143);
xor UO_3422 (O_3422,N_27532,N_29345);
nor UO_3423 (O_3423,N_26322,N_25787);
nand UO_3424 (O_3424,N_23017,N_28726);
nand UO_3425 (O_3425,N_26712,N_24914);
and UO_3426 (O_3426,N_23967,N_25062);
and UO_3427 (O_3427,N_20315,N_24790);
and UO_3428 (O_3428,N_27672,N_21324);
xnor UO_3429 (O_3429,N_23659,N_24766);
and UO_3430 (O_3430,N_26634,N_22984);
nor UO_3431 (O_3431,N_20377,N_29910);
nor UO_3432 (O_3432,N_25588,N_29906);
or UO_3433 (O_3433,N_21939,N_22224);
nor UO_3434 (O_3434,N_28398,N_22783);
nor UO_3435 (O_3435,N_27268,N_25321);
nand UO_3436 (O_3436,N_29352,N_23638);
or UO_3437 (O_3437,N_27871,N_27143);
and UO_3438 (O_3438,N_26429,N_22233);
or UO_3439 (O_3439,N_21511,N_20837);
nand UO_3440 (O_3440,N_25752,N_24010);
nand UO_3441 (O_3441,N_27496,N_25589);
and UO_3442 (O_3442,N_21321,N_27722);
or UO_3443 (O_3443,N_24514,N_22779);
and UO_3444 (O_3444,N_29101,N_22688);
nand UO_3445 (O_3445,N_29955,N_22529);
and UO_3446 (O_3446,N_22897,N_28130);
and UO_3447 (O_3447,N_27213,N_26845);
xor UO_3448 (O_3448,N_26656,N_23473);
or UO_3449 (O_3449,N_21663,N_24983);
or UO_3450 (O_3450,N_24263,N_23364);
xnor UO_3451 (O_3451,N_23157,N_26971);
nand UO_3452 (O_3452,N_25117,N_26560);
xor UO_3453 (O_3453,N_24096,N_27855);
or UO_3454 (O_3454,N_21927,N_22455);
and UO_3455 (O_3455,N_20122,N_29091);
nand UO_3456 (O_3456,N_28287,N_22767);
or UO_3457 (O_3457,N_25987,N_20072);
or UO_3458 (O_3458,N_20815,N_20571);
nand UO_3459 (O_3459,N_21023,N_25537);
nand UO_3460 (O_3460,N_28672,N_22223);
and UO_3461 (O_3461,N_28832,N_29709);
nor UO_3462 (O_3462,N_27710,N_29763);
and UO_3463 (O_3463,N_20134,N_21773);
or UO_3464 (O_3464,N_28280,N_29325);
nor UO_3465 (O_3465,N_20539,N_24949);
xnor UO_3466 (O_3466,N_25294,N_26319);
xor UO_3467 (O_3467,N_26421,N_21604);
nor UO_3468 (O_3468,N_21669,N_29847);
and UO_3469 (O_3469,N_20552,N_22285);
nor UO_3470 (O_3470,N_26632,N_20644);
xnor UO_3471 (O_3471,N_27981,N_23583);
and UO_3472 (O_3472,N_20568,N_20560);
or UO_3473 (O_3473,N_23932,N_29381);
nor UO_3474 (O_3474,N_24063,N_23010);
or UO_3475 (O_3475,N_23122,N_21775);
and UO_3476 (O_3476,N_25639,N_23464);
and UO_3477 (O_3477,N_23729,N_27819);
nand UO_3478 (O_3478,N_27992,N_25352);
nor UO_3479 (O_3479,N_21127,N_20230);
or UO_3480 (O_3480,N_20157,N_23120);
nor UO_3481 (O_3481,N_24314,N_21642);
and UO_3482 (O_3482,N_22962,N_28086);
and UO_3483 (O_3483,N_25249,N_20291);
and UO_3484 (O_3484,N_23376,N_29797);
or UO_3485 (O_3485,N_24247,N_28777);
nor UO_3486 (O_3486,N_22192,N_20543);
nand UO_3487 (O_3487,N_24854,N_21092);
or UO_3488 (O_3488,N_22409,N_23144);
and UO_3489 (O_3489,N_24169,N_20434);
and UO_3490 (O_3490,N_23446,N_23293);
nand UO_3491 (O_3491,N_27137,N_23575);
or UO_3492 (O_3492,N_21704,N_27494);
nand UO_3493 (O_3493,N_24846,N_29137);
nand UO_3494 (O_3494,N_27804,N_26902);
or UO_3495 (O_3495,N_24973,N_21972);
and UO_3496 (O_3496,N_20762,N_24617);
nor UO_3497 (O_3497,N_29737,N_28733);
or UO_3498 (O_3498,N_23767,N_22977);
and UO_3499 (O_3499,N_20825,N_27863);
endmodule