module basic_2000_20000_2500_5_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1228,In_1349);
nor U1 (N_1,In_868,In_397);
or U2 (N_2,In_1823,In_1852);
xnor U3 (N_3,In_508,In_684);
nand U4 (N_4,In_332,In_1570);
nor U5 (N_5,In_399,In_254);
nand U6 (N_6,In_1583,In_143);
xor U7 (N_7,In_1865,In_1704);
and U8 (N_8,In_1328,In_1857);
nor U9 (N_9,In_639,In_1694);
and U10 (N_10,In_1761,In_1038);
nor U11 (N_11,In_609,In_1166);
xor U12 (N_12,In_1628,In_590);
or U13 (N_13,In_553,In_530);
nor U14 (N_14,In_1483,In_1279);
and U15 (N_15,In_1635,In_346);
and U16 (N_16,In_1611,In_1095);
and U17 (N_17,In_966,In_1954);
xor U18 (N_18,In_1990,In_662);
or U19 (N_19,In_1042,In_1579);
nand U20 (N_20,In_1090,In_1170);
or U21 (N_21,In_488,In_221);
or U22 (N_22,In_805,In_39);
or U23 (N_23,In_574,In_294);
nor U24 (N_24,In_1837,In_1630);
nand U25 (N_25,In_53,In_1451);
and U26 (N_26,In_555,In_533);
or U27 (N_27,In_260,In_991);
or U28 (N_28,In_1624,In_1571);
nand U29 (N_29,In_699,In_1353);
nor U30 (N_30,In_281,In_1608);
nand U31 (N_31,In_121,In_1358);
nor U32 (N_32,In_1400,In_237);
nand U33 (N_33,In_1475,In_944);
xor U34 (N_34,In_350,In_416);
nand U35 (N_35,In_901,In_1469);
and U36 (N_36,In_1677,In_165);
nand U37 (N_37,In_768,In_69);
and U38 (N_38,In_1866,In_1953);
nor U39 (N_39,In_1562,In_1736);
and U40 (N_40,In_931,In_536);
or U41 (N_41,In_947,In_560);
or U42 (N_42,In_1526,In_1266);
or U43 (N_43,In_686,In_504);
nand U44 (N_44,In_631,In_1537);
xnor U45 (N_45,In_235,In_849);
xnor U46 (N_46,In_109,In_740);
and U47 (N_47,In_541,In_1669);
xor U48 (N_48,In_1871,In_1177);
xnor U49 (N_49,In_640,In_1629);
and U50 (N_50,In_1899,In_614);
or U51 (N_51,In_879,In_93);
nor U52 (N_52,In_851,In_604);
or U53 (N_53,In_1334,In_1165);
nor U54 (N_54,In_232,In_1278);
or U55 (N_55,In_712,In_1352);
or U56 (N_56,In_1930,In_637);
nand U57 (N_57,In_714,In_1119);
nand U58 (N_58,In_316,In_510);
and U59 (N_59,In_1726,In_565);
and U60 (N_60,In_1113,In_199);
and U61 (N_61,In_1815,In_86);
and U62 (N_62,In_468,In_1981);
and U63 (N_63,In_1111,In_683);
or U64 (N_64,In_1644,In_1344);
and U65 (N_65,In_1587,In_726);
and U66 (N_66,In_999,In_941);
nand U67 (N_67,In_1060,In_695);
and U68 (N_68,In_1816,In_617);
nand U69 (N_69,In_1124,In_172);
and U70 (N_70,In_1584,In_1895);
nor U71 (N_71,In_1196,In_3);
nor U72 (N_72,In_1500,In_778);
nor U73 (N_73,In_278,In_520);
or U74 (N_74,In_148,In_1337);
nand U75 (N_75,In_538,In_423);
and U76 (N_76,In_1455,In_1620);
nor U77 (N_77,In_1189,In_1153);
and U78 (N_78,In_1006,In_1592);
and U79 (N_79,In_597,In_892);
nor U80 (N_80,In_471,In_1938);
or U81 (N_81,In_1986,In_1420);
xnor U82 (N_82,In_1133,In_1903);
or U83 (N_83,In_516,In_1925);
nand U84 (N_84,In_9,In_487);
and U85 (N_85,In_1181,In_1361);
nor U86 (N_86,In_700,In_13);
or U87 (N_87,In_542,In_1586);
nor U88 (N_88,In_460,In_1947);
nor U89 (N_89,In_1398,In_479);
xnor U90 (N_90,In_1351,In_1504);
nor U91 (N_91,In_255,In_1803);
nand U92 (N_92,In_1224,In_343);
nor U93 (N_93,In_502,In_222);
and U94 (N_94,In_677,In_1538);
and U95 (N_95,In_983,In_353);
and U96 (N_96,In_1506,In_251);
nand U97 (N_97,In_1286,In_665);
nand U98 (N_98,In_540,In_757);
and U99 (N_99,In_464,In_1879);
or U100 (N_100,In_1663,In_1952);
xor U101 (N_101,In_1988,In_10);
or U102 (N_102,In_1945,In_845);
xor U103 (N_103,In_1796,In_1589);
or U104 (N_104,In_70,In_996);
xnor U105 (N_105,In_1687,In_641);
and U106 (N_106,In_385,In_959);
and U107 (N_107,In_698,In_454);
and U108 (N_108,In_1164,In_1012);
and U109 (N_109,In_383,In_128);
nor U110 (N_110,In_155,In_681);
or U111 (N_111,In_1627,In_1969);
nor U112 (N_112,In_1000,In_1484);
nand U113 (N_113,In_1901,In_1147);
and U114 (N_114,In_1122,In_1854);
nor U115 (N_115,In_1826,In_779);
nor U116 (N_116,In_776,In_351);
xnor U117 (N_117,In_76,In_167);
and U118 (N_118,In_1924,In_356);
nand U119 (N_119,In_382,In_880);
or U120 (N_120,In_1632,In_706);
and U121 (N_121,In_1371,In_719);
and U122 (N_122,In_1757,In_421);
xor U123 (N_123,In_888,In_1313);
or U124 (N_124,In_1780,In_751);
and U125 (N_125,In_1450,In_156);
and U126 (N_126,In_670,In_1789);
and U127 (N_127,In_887,In_1432);
and U128 (N_128,In_1192,In_742);
and U129 (N_129,In_929,In_1199);
and U130 (N_130,In_274,In_654);
xor U131 (N_131,In_787,In_485);
or U132 (N_132,In_82,In_348);
or U133 (N_133,In_1876,In_934);
or U134 (N_134,In_1399,In_687);
or U135 (N_135,In_1972,In_335);
nor U136 (N_136,In_276,In_284);
nor U137 (N_137,In_928,In_1270);
and U138 (N_138,In_1786,In_169);
nand U139 (N_139,In_767,In_1473);
or U140 (N_140,In_679,In_63);
xor U141 (N_141,In_1116,In_1017);
nor U142 (N_142,In_1712,In_1673);
xnor U143 (N_143,In_1827,In_1835);
nand U144 (N_144,In_444,In_64);
nand U145 (N_145,In_1206,In_937);
nor U146 (N_146,In_478,In_418);
nor U147 (N_147,In_1856,In_1581);
nor U148 (N_148,In_1029,In_1832);
and U149 (N_149,In_1552,In_1249);
nand U150 (N_150,In_975,In_1312);
or U151 (N_151,In_1120,In_660);
and U152 (N_152,In_241,In_1531);
xor U153 (N_153,In_666,In_1653);
nand U154 (N_154,In_1014,In_1243);
and U155 (N_155,In_1516,In_414);
and U156 (N_156,In_210,In_1281);
and U157 (N_157,In_1906,In_170);
xnor U158 (N_158,In_1777,In_1652);
nand U159 (N_159,In_132,In_784);
or U160 (N_160,In_1428,In_15);
nand U161 (N_161,In_793,In_797);
xor U162 (N_162,In_1023,In_1887);
or U163 (N_163,In_858,In_0);
nor U164 (N_164,In_90,In_1867);
nor U165 (N_165,In_1998,In_1480);
nand U166 (N_166,In_1028,In_323);
and U167 (N_167,In_1752,In_832);
nand U168 (N_168,In_126,In_451);
nor U169 (N_169,In_442,In_6);
and U170 (N_170,In_543,In_386);
nor U171 (N_171,In_517,In_362);
or U172 (N_172,In_1067,In_1394);
nor U173 (N_173,In_1997,In_1907);
or U174 (N_174,In_737,In_1942);
nor U175 (N_175,In_790,In_864);
and U176 (N_176,In_754,In_994);
nand U177 (N_177,In_1773,In_1191);
and U178 (N_178,In_1853,In_850);
nand U179 (N_179,In_819,In_189);
or U180 (N_180,In_1244,In_905);
xnor U181 (N_181,In_1276,In_1639);
and U182 (N_182,In_1379,In_799);
xor U183 (N_183,In_734,In_1710);
and U184 (N_184,In_85,In_924);
and U185 (N_185,In_91,In_214);
nand U186 (N_186,In_127,In_680);
or U187 (N_187,In_979,In_1173);
and U188 (N_188,In_1146,In_441);
and U189 (N_189,In_919,In_1005);
or U190 (N_190,In_922,In_1707);
nand U191 (N_191,In_1878,In_572);
nor U192 (N_192,In_174,In_1190);
nor U193 (N_193,In_509,In_716);
nand U194 (N_194,In_1785,In_1975);
nand U195 (N_195,In_1214,In_1555);
nor U196 (N_196,In_181,In_300);
and U197 (N_197,In_347,In_582);
nand U198 (N_198,In_1343,In_373);
nand U199 (N_199,In_473,In_1102);
and U200 (N_200,In_1053,In_424);
xnor U201 (N_201,In_549,In_659);
or U202 (N_202,In_1631,In_157);
nor U203 (N_203,In_1955,In_1962);
and U204 (N_204,In_669,In_548);
nand U205 (N_205,In_1395,In_325);
and U206 (N_206,In_245,In_789);
or U207 (N_207,In_285,In_591);
and U208 (N_208,In_1658,In_1819);
nor U209 (N_209,In_1967,In_306);
nand U210 (N_210,In_1126,In_775);
and U211 (N_211,In_81,In_465);
or U212 (N_212,In_1864,In_1123);
nor U213 (N_213,In_1999,In_1472);
or U214 (N_214,In_1063,In_1933);
nor U215 (N_215,In_1117,In_1642);
nand U216 (N_216,In_1869,In_515);
nand U217 (N_217,In_932,In_1580);
and U218 (N_218,In_606,In_1292);
or U219 (N_219,In_1366,In_448);
nor U220 (N_220,In_438,In_1690);
nand U221 (N_221,In_1223,In_619);
nor U222 (N_222,In_404,In_462);
or U223 (N_223,In_627,In_1062);
xor U224 (N_224,In_1833,In_1657);
or U225 (N_225,In_1168,In_1222);
or U226 (N_226,In_1659,In_14);
and U227 (N_227,In_1521,In_925);
nor U228 (N_228,In_1476,In_372);
xor U229 (N_229,In_1265,In_1944);
nor U230 (N_230,In_1740,In_697);
nor U231 (N_231,In_1209,In_1460);
and U232 (N_232,In_763,In_1756);
or U233 (N_233,In_1474,In_927);
and U234 (N_234,In_1964,In_1599);
xor U235 (N_235,In_1817,In_1965);
or U236 (N_236,In_1084,In_173);
or U237 (N_237,In_1479,In_129);
and U238 (N_238,In_1109,In_1308);
nand U239 (N_239,In_611,In_1129);
or U240 (N_240,In_731,In_376);
nand U241 (N_241,In_739,In_1596);
and U242 (N_242,In_164,In_1702);
or U243 (N_243,In_113,In_301);
or U244 (N_244,In_546,In_1503);
nand U245 (N_245,In_769,In_914);
nand U246 (N_246,In_1417,In_958);
or U247 (N_247,In_897,In_656);
and U248 (N_248,In_1547,In_962);
nand U249 (N_249,In_37,In_1215);
nor U250 (N_250,In_1490,In_94);
or U251 (N_251,In_554,In_1057);
nand U252 (N_252,In_432,In_1543);
nor U253 (N_253,In_1549,In_1448);
or U254 (N_254,In_1296,In_721);
nand U255 (N_255,In_1753,In_1155);
nand U256 (N_256,In_1163,In_1254);
or U257 (N_257,In_60,In_1435);
or U258 (N_258,In_357,In_162);
and U259 (N_259,In_956,In_1442);
xor U260 (N_260,In_31,In_1180);
or U261 (N_261,In_1297,In_252);
nand U262 (N_262,In_783,In_1850);
nor U263 (N_263,In_1405,In_302);
or U264 (N_264,In_989,In_1825);
and U265 (N_265,In_98,In_494);
and U266 (N_266,In_1686,In_995);
nand U267 (N_267,In_1783,In_1982);
and U268 (N_268,In_1750,In_1309);
nand U269 (N_269,In_1618,In_87);
or U270 (N_270,In_567,In_1843);
nor U271 (N_271,In_985,In_981);
nand U272 (N_272,In_653,In_800);
and U273 (N_273,In_758,In_1735);
nor U274 (N_274,In_387,In_1572);
or U275 (N_275,In_1805,In_728);
xnor U276 (N_276,In_238,In_190);
or U277 (N_277,In_430,In_146);
nor U278 (N_278,In_1948,In_638);
xnor U279 (N_279,In_19,In_435);
and U280 (N_280,In_1623,In_99);
nand U281 (N_281,In_1365,In_227);
and U282 (N_282,In_1691,In_1920);
and U283 (N_283,In_1251,In_1518);
xor U284 (N_284,In_1136,In_176);
nor U285 (N_285,In_1489,In_311);
nor U286 (N_286,In_1421,In_1323);
nor U287 (N_287,In_326,In_1205);
nand U288 (N_288,In_1762,In_144);
or U289 (N_289,In_1212,In_1041);
nand U290 (N_290,In_1022,In_771);
and U291 (N_291,In_961,In_29);
nor U292 (N_292,In_630,In_102);
nor U293 (N_293,In_643,In_1454);
or U294 (N_294,In_770,In_1654);
nand U295 (N_295,In_140,In_1648);
nand U296 (N_296,In_163,In_184);
nand U297 (N_297,In_592,In_1557);
and U298 (N_298,In_410,In_1427);
nand U299 (N_299,In_1935,In_1992);
nor U300 (N_300,In_18,In_987);
and U301 (N_301,In_1493,In_1385);
nand U302 (N_302,In_1429,In_1809);
nand U303 (N_303,In_1995,In_1025);
or U304 (N_304,In_26,In_1104);
and U305 (N_305,In_579,In_1892);
nand U306 (N_306,In_25,In_512);
nand U307 (N_307,In_1847,In_1923);
nor U308 (N_308,In_142,In_1675);
nor U309 (N_309,In_513,In_1647);
and U310 (N_310,In_405,In_196);
and U311 (N_311,In_672,In_263);
nand U312 (N_312,In_893,In_842);
nand U313 (N_313,In_1889,In_1340);
and U314 (N_314,In_183,In_378);
or U315 (N_315,In_545,In_1021);
or U316 (N_316,In_965,In_205);
nand U317 (N_317,In_1069,In_878);
nor U318 (N_318,In_218,In_561);
or U319 (N_319,In_792,In_65);
xor U320 (N_320,In_625,In_1985);
or U321 (N_321,In_1729,In_1403);
or U322 (N_322,In_1533,In_1966);
nor U323 (N_323,In_1464,In_702);
nand U324 (N_324,In_380,In_598);
xnor U325 (N_325,In_997,In_1711);
nor U326 (N_326,In_1510,In_1723);
or U327 (N_327,In_1179,In_309);
or U328 (N_328,In_484,In_1101);
or U329 (N_329,In_1877,In_1068);
or U330 (N_330,In_859,In_963);
and U331 (N_331,In_1207,In_433);
nand U332 (N_332,In_360,In_259);
nor U333 (N_333,In_1453,In_133);
nand U334 (N_334,In_288,In_1364);
xor U335 (N_335,In_587,In_809);
and U336 (N_336,In_1315,In_506);
nor U337 (N_337,In_1708,In_1775);
and U338 (N_338,In_491,In_1664);
xnor U339 (N_339,In_159,In_1305);
nand U340 (N_340,In_612,In_1078);
and U341 (N_341,In_1529,In_661);
and U342 (N_342,In_1217,In_853);
nand U343 (N_343,In_187,In_945);
and U344 (N_344,In_1044,In_1422);
nor U345 (N_345,In_580,In_459);
nor U346 (N_346,In_1839,In_158);
or U347 (N_347,In_1951,In_1092);
nor U348 (N_348,In_896,In_601);
xnor U349 (N_349,In_525,In_624);
nor U350 (N_350,In_179,In_1787);
nor U351 (N_351,In_1193,In_828);
nand U352 (N_352,In_599,In_733);
and U353 (N_353,In_367,In_1280);
nand U354 (N_354,In_379,In_1551);
and U355 (N_355,In_440,In_812);
and U356 (N_356,In_766,In_1693);
nor U357 (N_357,In_1517,In_171);
nor U358 (N_358,In_1043,In_588);
nor U359 (N_359,In_762,In_1380);
or U360 (N_360,In_613,In_1739);
and U361 (N_361,In_1713,In_1605);
and U362 (N_362,In_1227,In_1175);
or U363 (N_363,In_1868,In_1900);
nor U364 (N_364,In_1134,In_1316);
and U365 (N_365,In_824,In_1667);
nor U366 (N_366,In_1471,In_752);
or U367 (N_367,In_1758,In_1443);
nand U368 (N_368,In_523,In_890);
nand U369 (N_369,In_1643,In_1246);
nor U370 (N_370,In_547,In_1650);
or U371 (N_371,In_715,In_717);
or U372 (N_372,In_110,In_514);
nor U373 (N_373,In_365,In_138);
nand U374 (N_374,In_648,In_36);
nand U375 (N_375,In_396,In_229);
nor U376 (N_376,In_1625,In_452);
nand U377 (N_377,In_1367,In_1883);
and U378 (N_378,In_920,In_271);
nor U379 (N_379,In_247,In_96);
and U380 (N_380,In_486,In_898);
nand U381 (N_381,In_1426,In_1372);
xnor U382 (N_382,In_1715,In_275);
nor U383 (N_383,In_651,In_1311);
nand U384 (N_384,In_1829,In_823);
and U385 (N_385,In_705,In_1848);
nand U386 (N_386,In_701,In_1588);
and U387 (N_387,In_984,In_1376);
or U388 (N_388,In_32,In_759);
nand U389 (N_389,In_948,In_1003);
nand U390 (N_390,In_1974,In_577);
nor U391 (N_391,In_1325,In_1219);
and U392 (N_392,In_224,In_1719);
nand U393 (N_393,In_470,In_1797);
xor U394 (N_394,In_35,In_1247);
nand U395 (N_395,In_1671,In_363);
and U396 (N_396,In_1162,In_1083);
and U397 (N_397,In_1545,In_1978);
xnor U398 (N_398,In_1668,In_231);
nand U399 (N_399,In_1054,In_415);
nor U400 (N_400,In_282,In_1884);
and U401 (N_401,In_295,In_104);
or U402 (N_402,In_220,In_1804);
nor U403 (N_403,In_233,In_1106);
nor U404 (N_404,In_1130,In_248);
and U405 (N_405,In_258,In_95);
nand U406 (N_406,In_1345,In_1751);
or U407 (N_407,In_246,In_437);
xor U408 (N_408,In_1891,In_557);
nor U409 (N_409,In_1461,In_1438);
nand U410 (N_410,In_1968,In_1597);
nor U411 (N_411,In_1468,In_389);
and U412 (N_412,In_457,In_860);
xnor U413 (N_413,In_1174,In_1097);
nor U414 (N_414,In_650,In_1263);
nor U415 (N_415,In_1556,In_345);
or U416 (N_416,In_1019,In_1875);
or U417 (N_417,In_957,In_1178);
or U418 (N_418,In_180,In_149);
nand U419 (N_419,In_1110,In_1148);
nor U420 (N_420,In_483,In_671);
and U421 (N_421,In_375,In_1061);
and U422 (N_422,In_907,In_814);
or U423 (N_423,In_629,In_1703);
and U424 (N_424,In_28,In_349);
nand U425 (N_425,In_333,In_1695);
nand U426 (N_426,In_1984,In_1431);
xor U427 (N_427,In_1226,In_49);
nor U428 (N_428,In_1844,In_1040);
or U429 (N_429,In_1306,In_455);
nor U430 (N_430,In_1210,In_571);
and U431 (N_431,In_1501,In_1956);
and U432 (N_432,In_12,In_1058);
nor U433 (N_433,In_881,In_198);
and U434 (N_434,In_303,In_1622);
or U435 (N_435,In_1389,In_1811);
xor U436 (N_436,In_889,In_1798);
nand U437 (N_437,In_201,In_1011);
or U438 (N_438,In_213,In_1718);
nand U439 (N_439,In_1259,In_1100);
and U440 (N_440,In_1156,In_1784);
and U441 (N_441,In_392,In_1885);
xnor U442 (N_442,In_339,In_1274);
nand U443 (N_443,In_1689,In_1527);
nor U444 (N_444,In_844,In_1682);
nor U445 (N_445,In_1145,In_265);
nor U446 (N_446,In_1076,In_911);
or U447 (N_447,In_1347,In_1649);
nor U448 (N_448,In_244,In_1722);
nand U449 (N_449,In_1674,In_875);
xor U450 (N_450,In_802,In_11);
nand U451 (N_451,In_111,In_857);
or U452 (N_452,In_1742,In_943);
and U453 (N_453,In_1233,In_735);
or U454 (N_454,In_1154,In_891);
or U455 (N_455,In_1466,In_1559);
and U456 (N_456,In_935,In_1494);
and U457 (N_457,In_135,In_1356);
nand U458 (N_458,In_990,In_658);
or U459 (N_459,In_1374,In_1160);
nor U460 (N_460,In_1931,In_960);
nor U461 (N_461,In_1035,In_822);
nand U462 (N_462,In_331,In_1958);
and U463 (N_463,In_723,In_810);
nand U464 (N_464,In_1724,In_202);
xor U465 (N_465,In_1560,In_355);
and U466 (N_466,In_1615,In_1821);
nor U467 (N_467,In_1324,In_324);
or U468 (N_468,In_1338,In_1013);
nor U469 (N_469,In_1220,In_1055);
and U470 (N_470,In_50,In_1121);
and U471 (N_471,In_175,In_420);
and U472 (N_472,In_101,In_108);
nand U473 (N_473,In_1331,In_338);
nand U474 (N_474,In_528,In_100);
or U475 (N_475,In_1402,In_336);
and U476 (N_476,In_593,In_1514);
nand U477 (N_477,In_1327,In_1943);
or U478 (N_478,In_839,In_1872);
and U479 (N_479,In_556,In_1354);
or U480 (N_480,In_1941,In_431);
nor U481 (N_481,In_1094,In_1577);
nand U482 (N_482,In_1187,In_689);
or U483 (N_483,In_75,In_1370);
and U484 (N_484,In_1709,In_703);
and U485 (N_485,In_1937,In_1200);
nand U486 (N_486,In_1524,In_1996);
or U487 (N_487,In_429,In_492);
nor U488 (N_488,In_458,In_16);
and U489 (N_489,In_308,In_1738);
or U490 (N_490,In_1778,In_1194);
or U491 (N_491,In_1140,In_1457);
or U492 (N_492,In_1375,In_1834);
nand U493 (N_493,In_1582,In_250);
or U494 (N_494,In_1066,In_1262);
or U495 (N_495,In_334,In_1563);
xor U496 (N_496,In_782,In_474);
nand U497 (N_497,In_305,In_566);
or U498 (N_498,In_1275,In_1234);
or U499 (N_499,In_449,In_57);
nand U500 (N_500,In_381,In_391);
and U501 (N_501,In_1378,In_655);
or U502 (N_502,In_707,In_1911);
nor U503 (N_503,In_1575,In_884);
and U504 (N_504,In_1820,In_1488);
and U505 (N_505,In_54,In_1108);
nor U506 (N_506,In_48,In_1481);
and U507 (N_507,In_1651,In_72);
and U508 (N_508,In_2,In_1755);
nor U509 (N_509,In_1633,In_522);
nand U510 (N_510,In_634,In_1444);
nor U511 (N_511,In_453,In_1018);
xor U512 (N_512,In_1391,In_342);
and U513 (N_513,In_970,In_710);
nand U514 (N_514,In_708,In_837);
nand U515 (N_515,In_277,In_20);
or U516 (N_516,In_916,In_1082);
and U517 (N_517,In_967,In_1310);
or U518 (N_518,In_369,In_772);
and U519 (N_519,In_765,In_1030);
xor U520 (N_520,In_209,In_1922);
or U521 (N_521,In_633,In_532);
nor U522 (N_522,In_1152,In_1861);
nand U523 (N_523,In_761,In_243);
or U524 (N_524,In_1478,In_569);
xor U525 (N_525,In_481,In_835);
or U526 (N_526,In_1801,In_256);
nor U527 (N_527,In_657,In_1072);
nor U528 (N_528,In_527,In_297);
or U529 (N_529,In_826,In_66);
nor U530 (N_530,In_804,In_1073);
xor U531 (N_531,In_1137,In_1045);
nand U532 (N_532,In_124,In_1157);
and U533 (N_533,In_817,In_1253);
nor U534 (N_534,In_1957,In_1446);
or U535 (N_535,In_477,In_103);
nand U536 (N_536,In_1897,In_366);
and U537 (N_537,In_1499,In_1322);
xnor U538 (N_538,In_1734,In_745);
nor U539 (N_539,In_1052,In_535);
xor U540 (N_540,In_1766,In_1135);
nor U541 (N_541,In_861,In_570);
xnor U542 (N_542,In_622,In_992);
or U543 (N_543,In_1606,In_647);
and U544 (N_544,In_621,In_1230);
nor U545 (N_545,In_820,In_821);
nor U546 (N_546,In_1027,In_217);
and U547 (N_547,In_1568,In_341);
and U548 (N_548,In_668,In_873);
xor U549 (N_549,In_685,In_1383);
and U550 (N_550,In_785,In_1242);
and U551 (N_551,In_1085,In_692);
xor U552 (N_552,In_718,In_1637);
nand U553 (N_553,In_1335,In_1950);
or U554 (N_554,In_242,In_652);
nor U555 (N_555,In_1882,In_1720);
nand U556 (N_556,In_1046,In_551);
nor U557 (N_557,In_412,In_1684);
nand U558 (N_558,In_408,In_971);
nor U559 (N_559,In_1749,In_1321);
nor U560 (N_560,In_1634,In_1036);
and U561 (N_561,In_1363,In_434);
and U562 (N_562,In_1613,In_939);
nand U563 (N_563,In_1239,In_1714);
and U564 (N_564,In_178,In_1828);
xor U565 (N_565,In_730,In_136);
and U566 (N_566,In_848,In_207);
nand U567 (N_567,In_393,In_436);
and U568 (N_568,In_41,In_973);
nand U569 (N_569,In_1699,In_1416);
nor U570 (N_570,In_489,In_503);
or U571 (N_571,In_1357,In_280);
or U572 (N_572,In_1617,In_673);
and U573 (N_573,In_1240,In_480);
and U574 (N_574,In_777,In_1768);
nor U575 (N_575,In_204,In_83);
nand U576 (N_576,In_1373,In_674);
or U577 (N_577,In_1171,In_1467);
nor U578 (N_578,In_1976,In_986);
nor U579 (N_579,In_1728,In_1293);
xor U580 (N_580,In_1330,In_289);
nand U581 (N_581,In_1849,In_1301);
or U582 (N_582,In_1567,In_836);
or U583 (N_583,In_1886,In_568);
nor U584 (N_584,In_940,In_1112);
nor U585 (N_585,In_1115,In_371);
and U586 (N_586,In_402,In_1346);
nor U587 (N_587,In_1683,In_626);
xor U588 (N_588,In_1788,In_1603);
and U589 (N_589,In_1158,In_1812);
and U590 (N_590,In_56,In_1970);
and U591 (N_591,In_1824,In_846);
and U592 (N_592,In_526,In_328);
nor U593 (N_593,In_1544,In_909);
and U594 (N_594,In_223,In_511);
or U595 (N_595,In_1727,In_84);
and U596 (N_596,In_1881,In_1273);
nand U597 (N_597,In_1002,In_160);
nand U598 (N_598,In_1138,In_1238);
and U599 (N_599,In_829,In_713);
or U600 (N_600,In_1929,In_293);
xor U601 (N_601,In_1341,In_1646);
nand U602 (N_602,In_134,In_322);
nand U603 (N_603,In_1680,In_38);
nor U604 (N_604,In_827,In_1142);
nor U605 (N_605,In_1382,In_736);
nand U606 (N_606,In_1492,In_374);
or U607 (N_607,In_1511,In_1218);
nor U608 (N_608,In_262,In_1285);
and U609 (N_609,In_895,In_445);
or U610 (N_610,In_114,In_539);
or U611 (N_611,In_17,In_1991);
nand U612 (N_612,In_1267,In_186);
nand U613 (N_613,In_320,In_46);
nor U614 (N_614,In_1791,In_1621);
and U615 (N_615,In_1496,In_1236);
and U616 (N_616,In_1176,In_1088);
or U617 (N_617,In_1477,In_1841);
nand U618 (N_618,In_950,In_1607);
or U619 (N_619,In_1961,In_1600);
nor U620 (N_620,In_270,In_1411);
and U621 (N_621,In_788,In_1548);
nand U622 (N_622,In_1831,In_704);
and U623 (N_623,In_1792,In_521);
and U624 (N_624,In_30,In_693);
nor U625 (N_625,In_290,In_1934);
xor U626 (N_626,In_321,In_855);
and U627 (N_627,In_272,In_773);
nor U628 (N_628,In_1591,In_915);
or U629 (N_629,In_1128,In_1260);
or U630 (N_630,In_1554,In_1932);
nand U631 (N_631,In_1188,In_403);
or U632 (N_632,In_1692,In_1079);
nor U633 (N_633,In_1105,In_1401);
and U634 (N_634,In_413,In_1359);
nor U635 (N_635,In_1721,In_1415);
and U636 (N_636,In_1509,In_1048);
and U637 (N_637,In_211,In_906);
or U638 (N_638,In_107,In_1874);
or U639 (N_639,In_62,In_1523);
nand U640 (N_640,In_1842,In_1830);
and U641 (N_641,In_422,In_92);
nand U642 (N_642,In_664,In_1977);
nor U643 (N_643,In_1730,In_498);
and U644 (N_644,In_603,In_1681);
xnor U645 (N_645,In_188,In_1660);
xnor U646 (N_646,In_1896,In_1182);
nand U647 (N_647,In_1419,In_748);
and U648 (N_648,In_1495,In_267);
nand U649 (N_649,In_623,In_1541);
nor U650 (N_650,In_946,In_507);
or U651 (N_651,In_1732,In_1594);
and U652 (N_652,In_867,In_1915);
or U653 (N_653,In_1034,In_781);
xnor U654 (N_654,In_1486,In_1656);
xnor U655 (N_655,In_327,In_1598);
nand U656 (N_656,In_646,In_1590);
nand U657 (N_657,In_894,In_1733);
nor U658 (N_658,In_1908,In_1221);
nor U659 (N_659,In_1342,In_125);
xor U660 (N_660,In_1771,In_1150);
nand U661 (N_661,In_257,In_1745);
nand U662 (N_662,In_151,In_1360);
nand U663 (N_663,In_1118,In_602);
nand U664 (N_664,In_1498,In_1909);
xnor U665 (N_665,In_1141,In_1528);
nor U666 (N_666,In_1269,In_409);
and U667 (N_667,In_732,In_236);
nand U668 (N_668,In_524,In_1257);
nor U669 (N_669,In_1845,In_364);
and U670 (N_670,In_645,In_1008);
and U671 (N_671,In_1913,In_1747);
nor U672 (N_672,In_1065,In_818);
and U673 (N_673,In_1184,In_807);
nor U674 (N_674,In_446,In_1350);
or U675 (N_675,In_249,In_21);
and U676 (N_676,In_1566,In_1449);
and U677 (N_677,In_682,In_1298);
nor U678 (N_678,In_803,In_1198);
or U679 (N_679,In_595,In_368);
nand U680 (N_680,In_1880,In_44);
and U681 (N_681,In_1336,In_1211);
nand U682 (N_682,In_1638,In_1470);
or U683 (N_683,In_1989,In_1007);
and U684 (N_684,In_988,In_1277);
or U685 (N_685,In_688,In_161);
nand U686 (N_686,In_921,In_1697);
nor U687 (N_687,In_1979,In_678);
and U688 (N_688,In_1512,In_1696);
nor U689 (N_689,In_1093,In_1339);
xor U690 (N_690,In_663,In_1522);
and U691 (N_691,In_1802,In_869);
xnor U692 (N_692,In_1075,In_840);
xnor U693 (N_693,In_283,In_1700);
and U694 (N_694,In_760,In_1050);
nor U695 (N_695,In_1818,In_496);
nor U696 (N_696,In_722,In_1939);
xor U697 (N_697,In_1229,In_1368);
or U698 (N_698,In_475,In_1390);
nor U699 (N_699,In_1231,In_1741);
and U700 (N_700,In_1388,In_203);
and U701 (N_701,In_750,In_1917);
xnor U702 (N_702,In_1326,In_1392);
nor U703 (N_703,In_1256,In_493);
and U704 (N_704,In_97,In_1074);
xor U705 (N_705,In_261,In_384);
or U706 (N_706,In_34,In_1539);
or U707 (N_707,In_900,In_1814);
xnor U708 (N_708,In_727,In_1414);
nor U709 (N_709,In_1424,In_1799);
and U710 (N_710,In_1107,In_863);
and U711 (N_711,In_813,In_1225);
or U712 (N_712,In_52,In_1299);
nor U713 (N_713,In_1497,In_1381);
or U714 (N_714,In_808,In_1010);
and U715 (N_715,In_1525,In_1595);
and U716 (N_716,In_388,In_1558);
nand U717 (N_717,In_1425,In_1487);
nor U718 (N_718,In_1051,In_1081);
xnor U719 (N_719,In_1410,In_1167);
nand U720 (N_720,In_780,In_862);
xnor U721 (N_721,In_575,In_61);
and U722 (N_722,In_1926,In_191);
or U723 (N_723,In_977,In_825);
and U724 (N_724,In_675,In_1208);
nor U725 (N_725,In_1377,In_417);
nand U726 (N_726,In_709,In_1670);
nor U727 (N_727,In_1569,In_377);
xnor U728 (N_728,In_628,In_1836);
and U729 (N_729,In_89,In_1666);
and U730 (N_730,In_1790,In_615);
nand U731 (N_731,In_495,In_1250);
and U732 (N_732,In_1031,In_1255);
or U733 (N_733,In_1172,In_1641);
nor U734 (N_734,In_406,In_1776);
nor U735 (N_735,In_505,In_1404);
nand U736 (N_736,In_1959,In_208);
nor U737 (N_737,In_476,In_1546);
and U738 (N_738,In_1725,In_1439);
nor U739 (N_739,In_1574,In_1037);
xnor U740 (N_740,In_1928,In_291);
and U741 (N_741,In_838,In_594);
nand U742 (N_742,In_1807,In_352);
nor U743 (N_743,In_834,In_1406);
or U744 (N_744,In_978,In_816);
nand U745 (N_745,In_1091,In_4);
or U746 (N_746,In_1282,In_1905);
or U747 (N_747,In_870,In_1851);
nor U748 (N_748,In_1186,In_969);
nand U749 (N_749,In_1610,In_1759);
nand U750 (N_750,In_912,In_1125);
or U751 (N_751,In_936,In_620);
nor U752 (N_752,In_1767,In_193);
nor U753 (N_753,In_1774,In_74);
nor U754 (N_754,In_815,In_71);
and U755 (N_755,In_910,In_1946);
and U756 (N_756,In_1447,In_531);
and U757 (N_757,In_1731,In_1744);
nand U758 (N_758,In_871,In_1283);
nor U759 (N_759,In_1860,In_1232);
or U760 (N_760,In_304,In_266);
nor U761 (N_761,In_27,In_1362);
nand U762 (N_762,In_1127,In_490);
and U763 (N_763,In_518,In_1320);
nor U764 (N_764,In_1304,In_1604);
and U765 (N_765,In_856,In_725);
and U766 (N_766,In_1245,In_1185);
xor U767 (N_767,In_1769,In_753);
or U768 (N_768,In_696,In_443);
and U769 (N_769,In_852,In_400);
xnor U770 (N_770,In_1898,In_177);
or U771 (N_771,In_313,In_273);
nand U772 (N_772,In_1463,In_1386);
and U773 (N_773,In_1765,In_876);
nor U774 (N_774,In_904,In_1973);
and U775 (N_775,In_1994,In_1890);
nor U776 (N_776,In_117,In_1936);
or U777 (N_777,In_1532,In_1077);
nand U778 (N_778,In_573,In_1071);
nor U779 (N_779,In_1149,In_1348);
nor U780 (N_780,In_1396,In_192);
xnor U781 (N_781,In_1258,In_1502);
and U782 (N_782,In_185,In_1912);
and U783 (N_783,In_607,In_115);
or U784 (N_784,In_1840,In_563);
xnor U785 (N_785,In_253,In_296);
nor U786 (N_786,In_43,In_562);
and U787 (N_787,In_1307,In_550);
nor U788 (N_788,In_1910,In_1585);
nor U789 (N_789,In_1902,In_951);
nor U790 (N_790,In_1114,In_954);
or U791 (N_791,In_1565,In_854);
nor U792 (N_792,In_1676,In_1333);
nor U793 (N_793,In_1015,In_642);
nand U794 (N_794,In_497,In_1300);
xnor U795 (N_795,In_131,In_1601);
or U796 (N_796,In_993,In_312);
xor U797 (N_797,In_5,In_795);
nand U798 (N_798,In_286,In_51);
nor U799 (N_799,In_930,In_287);
nor U800 (N_800,In_885,In_1004);
or U801 (N_801,In_450,In_315);
or U802 (N_802,In_40,In_425);
and U803 (N_803,In_1519,In_1578);
or U804 (N_804,In_584,In_644);
nor U805 (N_805,In_1151,In_329);
nand U806 (N_806,In_340,In_1781);
and U807 (N_807,In_632,In_1319);
and U808 (N_808,In_116,In_139);
nand U809 (N_809,In_938,In_1550);
or U810 (N_810,In_168,In_1748);
nand U811 (N_811,In_667,In_596);
nand U812 (N_812,In_1561,In_1195);
nand U813 (N_813,In_953,In_1070);
and U814 (N_814,In_1716,In_1870);
nor U815 (N_815,In_206,In_1303);
nor U816 (N_816,In_1858,In_1838);
nor U817 (N_817,In_519,In_738);
nand U818 (N_818,In_145,In_427);
nand U819 (N_819,In_883,In_872);
and U820 (N_820,In_886,In_1237);
or U821 (N_821,In_1927,In_798);
or U822 (N_822,In_1536,In_1271);
or U823 (N_823,In_1318,In_1033);
nand U824 (N_824,In_310,In_314);
nand U825 (N_825,In_1024,In_439);
and U826 (N_826,In_581,In_1640);
nor U827 (N_827,In_307,In_123);
nor U828 (N_828,In_649,In_1678);
nor U829 (N_829,In_463,In_1564);
nand U830 (N_830,In_130,In_67);
nand U831 (N_831,In_1893,In_1131);
nor U832 (N_832,In_1863,In_219);
or U833 (N_833,In_976,In_230);
or U834 (N_834,In_1540,In_694);
or U835 (N_835,In_841,In_359);
nand U836 (N_836,In_1515,In_68);
nor U837 (N_837,In_1782,In_150);
and U838 (N_838,In_1423,In_552);
or U839 (N_839,In_724,In_1553);
nor U840 (N_840,In_831,In_1701);
nor U841 (N_841,In_1314,In_1505);
nand U842 (N_842,In_1020,In_1369);
nor U843 (N_843,In_1412,In_1264);
xor U844 (N_844,In_756,In_1413);
and U845 (N_845,In_1434,In_24);
or U846 (N_846,In_1144,In_830);
nor U847 (N_847,In_1949,In_917);
and U848 (N_848,In_1779,In_398);
nand U849 (N_849,In_1772,In_1302);
nand U850 (N_850,In_882,In_903);
xor U851 (N_851,In_106,In_358);
nand U852 (N_852,In_216,In_1513);
nor U853 (N_853,In_228,In_1159);
xnor U854 (N_854,In_1916,In_1202);
and U855 (N_855,In_1009,In_949);
and U856 (N_856,In_112,In_33);
nand U857 (N_857,In_1795,In_1593);
nand U858 (N_858,In_720,In_1754);
nor U859 (N_859,In_317,In_1859);
or U860 (N_860,In_877,In_1846);
xor U861 (N_861,In_47,In_578);
nand U862 (N_862,In_1272,In_80);
and U863 (N_863,In_447,In_1203);
nand U864 (N_864,In_1655,In_1626);
nand U865 (N_865,In_1197,In_746);
nand U866 (N_866,In_1332,In_968);
nand U867 (N_867,In_791,In_22);
nand U868 (N_868,In_1047,In_902);
nand U869 (N_869,In_1143,In_239);
nand U870 (N_870,In_182,In_1800);
xor U871 (N_871,In_1418,In_1387);
nor U872 (N_872,In_918,In_1520);
and U873 (N_873,In_1822,In_618);
nor U874 (N_874,In_833,In_1268);
xnor U875 (N_875,In_73,In_1183);
nand U876 (N_876,In_691,In_147);
nand U877 (N_877,In_1614,In_1284);
or U878 (N_878,In_401,In_1290);
nor U879 (N_879,In_1919,In_1001);
xor U880 (N_880,In_1662,In_1534);
and U881 (N_881,In_212,In_749);
or U882 (N_882,In_472,In_500);
and U883 (N_883,In_137,In_1491);
xor U884 (N_884,In_955,In_589);
and U885 (N_885,In_1,In_461);
and U886 (N_886,In_564,In_743);
or U887 (N_887,In_1288,In_501);
xnor U888 (N_888,In_225,In_395);
or U889 (N_889,In_1665,In_1980);
or U890 (N_890,In_1252,In_1408);
and U891 (N_891,In_88,In_1602);
nand U892 (N_892,In_42,In_337);
nor U893 (N_893,In_1169,In_1616);
nor U894 (N_894,In_7,In_786);
and U895 (N_895,In_998,In_1216);
and U896 (N_896,In_152,In_118);
nand U897 (N_897,In_166,In_847);
and U898 (N_898,In_843,In_269);
nor U899 (N_899,In_1987,In_1436);
xor U900 (N_900,In_1888,In_1813);
nand U901 (N_901,In_1971,In_1397);
nor U902 (N_902,In_1261,In_1894);
or U903 (N_903,In_1430,In_1576);
nor U904 (N_904,In_1289,In_1904);
nand U905 (N_905,In_467,In_774);
nor U906 (N_906,In_330,In_1441);
and U907 (N_907,In_411,In_1535);
nand U908 (N_908,In_299,In_585);
or U909 (N_909,In_428,In_1862);
nor U910 (N_910,In_1688,In_1459);
nor U911 (N_911,In_534,In_1161);
or U912 (N_912,In_1241,In_926);
or U913 (N_913,In_1698,In_874);
xor U914 (N_914,In_1291,In_794);
xnor U915 (N_915,In_1609,In_1213);
nor U916 (N_916,In_1465,In_529);
or U917 (N_917,In_407,In_1706);
or U918 (N_918,In_1636,In_899);
and U919 (N_919,In_1612,In_908);
nand U920 (N_920,In_1016,In_122);
or U921 (N_921,In_1737,In_344);
and U922 (N_922,In_1793,In_120);
nor U923 (N_923,In_77,In_964);
and U924 (N_924,In_1080,In_105);
nor U925 (N_925,In_1508,In_1089);
and U926 (N_926,In_676,In_811);
nor U927 (N_927,In_1407,In_78);
or U928 (N_928,In_744,In_354);
or U929 (N_929,In_1201,In_79);
nor U930 (N_930,In_1810,In_482);
nor U931 (N_931,In_866,In_153);
and U932 (N_932,In_1914,In_1456);
and U933 (N_933,In_913,In_319);
and U934 (N_934,In_318,In_1132);
nor U935 (N_935,In_974,In_499);
and U936 (N_936,In_1940,In_1026);
and U937 (N_937,In_1086,In_59);
nor U938 (N_938,In_1098,In_1573);
nand U939 (N_939,In_55,In_1452);
and U940 (N_940,In_390,In_1746);
nand U941 (N_941,In_200,In_466);
and U942 (N_942,In_583,In_1437);
and U943 (N_943,In_58,In_1921);
nor U944 (N_944,In_195,In_741);
xnor U945 (N_945,In_394,In_1542);
nand U946 (N_946,In_194,In_1087);
and U947 (N_947,In_1806,In_1485);
and U948 (N_948,In_1059,In_982);
nand U949 (N_949,In_1743,In_796);
nor U950 (N_950,In_729,In_610);
nand U951 (N_951,In_370,In_1717);
and U952 (N_952,In_1855,In_1672);
nor U953 (N_953,In_197,In_558);
and U954 (N_954,In_1993,In_1963);
nand U955 (N_955,In_1204,In_298);
nor U956 (N_956,In_1139,In_215);
nor U957 (N_957,In_1235,In_154);
or U958 (N_958,In_1409,In_1507);
and U959 (N_959,In_576,In_456);
and U960 (N_960,In_426,In_636);
and U961 (N_961,In_933,In_923);
nor U962 (N_962,In_1445,In_1619);
nand U963 (N_963,In_119,In_544);
or U964 (N_964,In_1039,In_952);
nor U965 (N_965,In_8,In_469);
and U966 (N_966,In_1049,In_764);
nor U967 (N_967,In_1679,In_586);
or U968 (N_968,In_1103,In_1462);
xnor U969 (N_969,In_1705,In_1248);
and U970 (N_970,In_1983,In_608);
and U971 (N_971,In_1794,In_1433);
nand U972 (N_972,In_1384,In_865);
nor U973 (N_973,In_1317,In_264);
nor U974 (N_974,In_1056,In_1530);
and U975 (N_975,In_1458,In_1355);
nor U976 (N_976,In_1287,In_1096);
and U977 (N_977,In_1960,In_45);
and U978 (N_978,In_1329,In_1918);
or U979 (N_979,In_419,In_226);
xor U980 (N_980,In_600,In_755);
nor U981 (N_981,In_1661,In_1064);
and U982 (N_982,In_537,In_1440);
nand U983 (N_983,In_279,In_361);
xnor U984 (N_984,In_690,In_1764);
or U985 (N_985,In_980,In_942);
or U986 (N_986,In_711,In_1763);
nor U987 (N_987,In_747,In_1770);
or U988 (N_988,In_806,In_801);
nor U989 (N_989,In_1482,In_1760);
nor U990 (N_990,In_616,In_635);
or U991 (N_991,In_268,In_972);
and U992 (N_992,In_141,In_240);
or U993 (N_993,In_1685,In_1099);
or U994 (N_994,In_1808,In_1295);
nand U995 (N_995,In_1294,In_1873);
nand U996 (N_996,In_23,In_234);
nand U997 (N_997,In_559,In_1645);
or U998 (N_998,In_292,In_1393);
or U999 (N_999,In_605,In_1032);
nand U1000 (N_1000,In_1276,In_1536);
nor U1001 (N_1001,In_598,In_739);
nand U1002 (N_1002,In_1326,In_5);
nor U1003 (N_1003,In_1439,In_1624);
xnor U1004 (N_1004,In_1066,In_1087);
or U1005 (N_1005,In_443,In_1196);
or U1006 (N_1006,In_205,In_162);
xnor U1007 (N_1007,In_1250,In_851);
and U1008 (N_1008,In_119,In_679);
nand U1009 (N_1009,In_1943,In_569);
or U1010 (N_1010,In_639,In_274);
nand U1011 (N_1011,In_1472,In_1476);
xor U1012 (N_1012,In_1463,In_1553);
nor U1013 (N_1013,In_390,In_422);
nand U1014 (N_1014,In_1615,In_72);
nand U1015 (N_1015,In_112,In_385);
xor U1016 (N_1016,In_1594,In_1264);
xnor U1017 (N_1017,In_1906,In_1071);
or U1018 (N_1018,In_128,In_1653);
nand U1019 (N_1019,In_1679,In_1801);
nand U1020 (N_1020,In_598,In_563);
nand U1021 (N_1021,In_1217,In_986);
nor U1022 (N_1022,In_743,In_314);
and U1023 (N_1023,In_20,In_164);
or U1024 (N_1024,In_1175,In_579);
and U1025 (N_1025,In_119,In_1071);
and U1026 (N_1026,In_893,In_751);
nand U1027 (N_1027,In_1165,In_1099);
nor U1028 (N_1028,In_1895,In_1948);
nand U1029 (N_1029,In_1690,In_1826);
and U1030 (N_1030,In_29,In_1381);
and U1031 (N_1031,In_648,In_1277);
or U1032 (N_1032,In_823,In_1719);
and U1033 (N_1033,In_1885,In_247);
and U1034 (N_1034,In_1775,In_498);
and U1035 (N_1035,In_1661,In_1993);
nor U1036 (N_1036,In_984,In_1640);
and U1037 (N_1037,In_1017,In_392);
or U1038 (N_1038,In_996,In_1647);
nor U1039 (N_1039,In_240,In_1055);
xnor U1040 (N_1040,In_233,In_614);
nor U1041 (N_1041,In_1085,In_958);
and U1042 (N_1042,In_394,In_66);
nand U1043 (N_1043,In_1260,In_1316);
nand U1044 (N_1044,In_596,In_1384);
and U1045 (N_1045,In_603,In_1672);
nand U1046 (N_1046,In_1818,In_930);
nand U1047 (N_1047,In_894,In_1172);
nor U1048 (N_1048,In_1487,In_1750);
xor U1049 (N_1049,In_1348,In_1492);
and U1050 (N_1050,In_742,In_860);
or U1051 (N_1051,In_1367,In_729);
nor U1052 (N_1052,In_212,In_864);
or U1053 (N_1053,In_164,In_1452);
and U1054 (N_1054,In_320,In_1549);
and U1055 (N_1055,In_874,In_466);
or U1056 (N_1056,In_656,In_309);
nor U1057 (N_1057,In_526,In_774);
nor U1058 (N_1058,In_953,In_130);
nor U1059 (N_1059,In_1592,In_1574);
or U1060 (N_1060,In_981,In_273);
nand U1061 (N_1061,In_1616,In_1797);
nor U1062 (N_1062,In_918,In_1256);
xor U1063 (N_1063,In_1353,In_1879);
or U1064 (N_1064,In_1512,In_1679);
nor U1065 (N_1065,In_1962,In_817);
nor U1066 (N_1066,In_1109,In_1603);
or U1067 (N_1067,In_1659,In_1033);
or U1068 (N_1068,In_268,In_909);
or U1069 (N_1069,In_597,In_472);
or U1070 (N_1070,In_777,In_1691);
nor U1071 (N_1071,In_981,In_53);
or U1072 (N_1072,In_226,In_1339);
and U1073 (N_1073,In_1217,In_1539);
or U1074 (N_1074,In_1273,In_602);
or U1075 (N_1075,In_1196,In_478);
nand U1076 (N_1076,In_1901,In_1318);
nor U1077 (N_1077,In_1423,In_1353);
or U1078 (N_1078,In_1792,In_247);
xor U1079 (N_1079,In_50,In_339);
and U1080 (N_1080,In_672,In_1302);
and U1081 (N_1081,In_491,In_186);
nor U1082 (N_1082,In_167,In_1524);
nor U1083 (N_1083,In_785,In_1505);
nor U1084 (N_1084,In_1592,In_978);
or U1085 (N_1085,In_231,In_167);
nor U1086 (N_1086,In_145,In_855);
or U1087 (N_1087,In_1762,In_836);
nor U1088 (N_1088,In_1173,In_1371);
xor U1089 (N_1089,In_1065,In_1382);
and U1090 (N_1090,In_1106,In_15);
nand U1091 (N_1091,In_1946,In_21);
and U1092 (N_1092,In_583,In_1427);
or U1093 (N_1093,In_551,In_1328);
nand U1094 (N_1094,In_1056,In_275);
nand U1095 (N_1095,In_140,In_1199);
and U1096 (N_1096,In_1677,In_742);
and U1097 (N_1097,In_259,In_1428);
nor U1098 (N_1098,In_1472,In_319);
nand U1099 (N_1099,In_1369,In_1050);
or U1100 (N_1100,In_620,In_288);
and U1101 (N_1101,In_1131,In_1371);
nand U1102 (N_1102,In_286,In_601);
nor U1103 (N_1103,In_630,In_637);
nor U1104 (N_1104,In_97,In_852);
nand U1105 (N_1105,In_1894,In_999);
nor U1106 (N_1106,In_1375,In_640);
or U1107 (N_1107,In_1543,In_1035);
or U1108 (N_1108,In_1633,In_1161);
nor U1109 (N_1109,In_1485,In_1044);
or U1110 (N_1110,In_376,In_678);
nand U1111 (N_1111,In_1821,In_1961);
xnor U1112 (N_1112,In_1332,In_93);
or U1113 (N_1113,In_1684,In_1670);
nand U1114 (N_1114,In_708,In_1182);
or U1115 (N_1115,In_1830,In_496);
nand U1116 (N_1116,In_1938,In_1370);
nor U1117 (N_1117,In_1424,In_1423);
xnor U1118 (N_1118,In_249,In_381);
nand U1119 (N_1119,In_1049,In_202);
xor U1120 (N_1120,In_944,In_1823);
xor U1121 (N_1121,In_1590,In_549);
and U1122 (N_1122,In_433,In_948);
nand U1123 (N_1123,In_1686,In_1738);
and U1124 (N_1124,In_129,In_683);
nand U1125 (N_1125,In_1411,In_1780);
nor U1126 (N_1126,In_939,In_40);
and U1127 (N_1127,In_1931,In_1737);
nand U1128 (N_1128,In_1246,In_632);
nor U1129 (N_1129,In_1996,In_35);
nor U1130 (N_1130,In_39,In_391);
nand U1131 (N_1131,In_1669,In_657);
or U1132 (N_1132,In_1316,In_421);
and U1133 (N_1133,In_1280,In_279);
and U1134 (N_1134,In_771,In_1954);
and U1135 (N_1135,In_1734,In_435);
nor U1136 (N_1136,In_1568,In_57);
and U1137 (N_1137,In_1485,In_1173);
nand U1138 (N_1138,In_1887,In_931);
xor U1139 (N_1139,In_1990,In_1508);
xor U1140 (N_1140,In_1480,In_1859);
nor U1141 (N_1141,In_1209,In_1878);
and U1142 (N_1142,In_1979,In_492);
and U1143 (N_1143,In_430,In_1425);
nor U1144 (N_1144,In_917,In_126);
nor U1145 (N_1145,In_414,In_640);
or U1146 (N_1146,In_1204,In_1320);
and U1147 (N_1147,In_640,In_1664);
nand U1148 (N_1148,In_978,In_726);
or U1149 (N_1149,In_1378,In_635);
or U1150 (N_1150,In_547,In_540);
xor U1151 (N_1151,In_1534,In_1540);
xnor U1152 (N_1152,In_1927,In_821);
and U1153 (N_1153,In_167,In_807);
nor U1154 (N_1154,In_1667,In_1947);
or U1155 (N_1155,In_1029,In_1105);
or U1156 (N_1156,In_315,In_276);
nor U1157 (N_1157,In_1074,In_1152);
and U1158 (N_1158,In_1899,In_203);
and U1159 (N_1159,In_42,In_1384);
or U1160 (N_1160,In_1893,In_1950);
or U1161 (N_1161,In_1290,In_1114);
or U1162 (N_1162,In_129,In_202);
and U1163 (N_1163,In_1165,In_33);
nand U1164 (N_1164,In_130,In_690);
xnor U1165 (N_1165,In_267,In_1193);
or U1166 (N_1166,In_214,In_1976);
nor U1167 (N_1167,In_536,In_981);
nand U1168 (N_1168,In_608,In_514);
nor U1169 (N_1169,In_1415,In_474);
and U1170 (N_1170,In_581,In_1209);
or U1171 (N_1171,In_1240,In_388);
nor U1172 (N_1172,In_215,In_1079);
nand U1173 (N_1173,In_351,In_453);
and U1174 (N_1174,In_721,In_1934);
nor U1175 (N_1175,In_1781,In_1753);
nand U1176 (N_1176,In_150,In_1076);
or U1177 (N_1177,In_358,In_896);
nand U1178 (N_1178,In_1464,In_976);
or U1179 (N_1179,In_403,In_364);
and U1180 (N_1180,In_799,In_1248);
and U1181 (N_1181,In_1360,In_855);
or U1182 (N_1182,In_388,In_1683);
or U1183 (N_1183,In_844,In_646);
xor U1184 (N_1184,In_1925,In_1816);
and U1185 (N_1185,In_1832,In_1073);
nand U1186 (N_1186,In_1682,In_843);
nor U1187 (N_1187,In_187,In_1260);
nand U1188 (N_1188,In_1609,In_405);
or U1189 (N_1189,In_1942,In_959);
xor U1190 (N_1190,In_594,In_179);
nand U1191 (N_1191,In_158,In_1);
and U1192 (N_1192,In_154,In_1826);
xor U1193 (N_1193,In_1623,In_493);
or U1194 (N_1194,In_650,In_1558);
nor U1195 (N_1195,In_1971,In_1092);
and U1196 (N_1196,In_1526,In_735);
and U1197 (N_1197,In_1405,In_645);
nand U1198 (N_1198,In_1526,In_1242);
and U1199 (N_1199,In_891,In_1623);
nor U1200 (N_1200,In_1535,In_955);
nor U1201 (N_1201,In_1194,In_732);
nor U1202 (N_1202,In_1313,In_173);
nand U1203 (N_1203,In_397,In_430);
and U1204 (N_1204,In_719,In_1320);
nand U1205 (N_1205,In_1264,In_453);
or U1206 (N_1206,In_332,In_273);
or U1207 (N_1207,In_1910,In_153);
nor U1208 (N_1208,In_1779,In_1247);
nand U1209 (N_1209,In_101,In_1580);
xor U1210 (N_1210,In_843,In_1230);
nor U1211 (N_1211,In_1524,In_168);
nor U1212 (N_1212,In_246,In_455);
and U1213 (N_1213,In_503,In_631);
or U1214 (N_1214,In_602,In_874);
and U1215 (N_1215,In_1023,In_109);
and U1216 (N_1216,In_366,In_1861);
or U1217 (N_1217,In_501,In_373);
nand U1218 (N_1218,In_1859,In_225);
and U1219 (N_1219,In_1391,In_1163);
or U1220 (N_1220,In_1312,In_1396);
xnor U1221 (N_1221,In_1967,In_1587);
nor U1222 (N_1222,In_24,In_949);
nor U1223 (N_1223,In_1023,In_392);
or U1224 (N_1224,In_298,In_1618);
nor U1225 (N_1225,In_1699,In_1564);
or U1226 (N_1226,In_170,In_890);
or U1227 (N_1227,In_528,In_1935);
and U1228 (N_1228,In_1468,In_1029);
nor U1229 (N_1229,In_368,In_774);
xor U1230 (N_1230,In_637,In_1848);
nand U1231 (N_1231,In_1999,In_1002);
or U1232 (N_1232,In_205,In_209);
xnor U1233 (N_1233,In_523,In_1930);
nand U1234 (N_1234,In_739,In_678);
nor U1235 (N_1235,In_1817,In_1434);
or U1236 (N_1236,In_1396,In_537);
and U1237 (N_1237,In_1139,In_992);
xnor U1238 (N_1238,In_546,In_1133);
or U1239 (N_1239,In_1242,In_1079);
nor U1240 (N_1240,In_1129,In_1296);
nand U1241 (N_1241,In_751,In_781);
nor U1242 (N_1242,In_517,In_1979);
and U1243 (N_1243,In_1828,In_1267);
nor U1244 (N_1244,In_1521,In_458);
or U1245 (N_1245,In_1839,In_904);
and U1246 (N_1246,In_360,In_1463);
nor U1247 (N_1247,In_16,In_1719);
nand U1248 (N_1248,In_570,In_1524);
nor U1249 (N_1249,In_1113,In_1196);
xnor U1250 (N_1250,In_1169,In_1498);
and U1251 (N_1251,In_899,In_831);
or U1252 (N_1252,In_1147,In_1043);
nor U1253 (N_1253,In_824,In_1135);
and U1254 (N_1254,In_1925,In_121);
nand U1255 (N_1255,In_1512,In_1870);
nor U1256 (N_1256,In_19,In_1838);
nand U1257 (N_1257,In_651,In_205);
or U1258 (N_1258,In_787,In_85);
nor U1259 (N_1259,In_1454,In_921);
nor U1260 (N_1260,In_1488,In_212);
or U1261 (N_1261,In_805,In_3);
nand U1262 (N_1262,In_151,In_996);
nor U1263 (N_1263,In_739,In_1043);
xnor U1264 (N_1264,In_265,In_1415);
or U1265 (N_1265,In_1405,In_964);
nor U1266 (N_1266,In_954,In_511);
and U1267 (N_1267,In_1242,In_1662);
nand U1268 (N_1268,In_432,In_1194);
or U1269 (N_1269,In_1915,In_19);
and U1270 (N_1270,In_244,In_513);
nand U1271 (N_1271,In_1250,In_1191);
and U1272 (N_1272,In_991,In_943);
or U1273 (N_1273,In_1588,In_922);
or U1274 (N_1274,In_333,In_1955);
xor U1275 (N_1275,In_1653,In_592);
or U1276 (N_1276,In_1290,In_236);
xor U1277 (N_1277,In_1276,In_883);
nand U1278 (N_1278,In_60,In_1821);
nor U1279 (N_1279,In_1668,In_1263);
xnor U1280 (N_1280,In_407,In_788);
nor U1281 (N_1281,In_1770,In_1452);
and U1282 (N_1282,In_1222,In_381);
nor U1283 (N_1283,In_1696,In_863);
and U1284 (N_1284,In_1623,In_279);
nand U1285 (N_1285,In_1739,In_221);
nand U1286 (N_1286,In_1616,In_960);
and U1287 (N_1287,In_165,In_324);
nand U1288 (N_1288,In_194,In_843);
nand U1289 (N_1289,In_37,In_1799);
or U1290 (N_1290,In_1196,In_349);
xor U1291 (N_1291,In_1930,In_358);
and U1292 (N_1292,In_871,In_608);
nor U1293 (N_1293,In_608,In_672);
nand U1294 (N_1294,In_1648,In_935);
and U1295 (N_1295,In_1646,In_199);
xnor U1296 (N_1296,In_251,In_1961);
or U1297 (N_1297,In_1303,In_755);
or U1298 (N_1298,In_1763,In_834);
and U1299 (N_1299,In_806,In_1929);
or U1300 (N_1300,In_1314,In_400);
and U1301 (N_1301,In_327,In_657);
and U1302 (N_1302,In_617,In_1592);
nor U1303 (N_1303,In_1346,In_1222);
nand U1304 (N_1304,In_684,In_1084);
or U1305 (N_1305,In_1437,In_314);
nor U1306 (N_1306,In_44,In_389);
nand U1307 (N_1307,In_1970,In_1805);
and U1308 (N_1308,In_1060,In_1277);
or U1309 (N_1309,In_960,In_1374);
and U1310 (N_1310,In_256,In_1294);
nor U1311 (N_1311,In_1675,In_1698);
and U1312 (N_1312,In_470,In_328);
or U1313 (N_1313,In_283,In_1829);
and U1314 (N_1314,In_1121,In_14);
nor U1315 (N_1315,In_410,In_1309);
or U1316 (N_1316,In_428,In_471);
nand U1317 (N_1317,In_1627,In_723);
nor U1318 (N_1318,In_97,In_1873);
nand U1319 (N_1319,In_1557,In_434);
nor U1320 (N_1320,In_1201,In_732);
nand U1321 (N_1321,In_367,In_176);
and U1322 (N_1322,In_829,In_816);
nand U1323 (N_1323,In_1082,In_1667);
nand U1324 (N_1324,In_1977,In_278);
nor U1325 (N_1325,In_956,In_1491);
nor U1326 (N_1326,In_1404,In_250);
or U1327 (N_1327,In_186,In_1395);
nand U1328 (N_1328,In_99,In_115);
or U1329 (N_1329,In_1387,In_1328);
nor U1330 (N_1330,In_1708,In_346);
and U1331 (N_1331,In_1723,In_1242);
and U1332 (N_1332,In_623,In_1371);
or U1333 (N_1333,In_1315,In_908);
and U1334 (N_1334,In_1179,In_407);
or U1335 (N_1335,In_1598,In_1777);
and U1336 (N_1336,In_439,In_1875);
nor U1337 (N_1337,In_1133,In_887);
nor U1338 (N_1338,In_521,In_527);
xor U1339 (N_1339,In_1572,In_173);
or U1340 (N_1340,In_224,In_1365);
nor U1341 (N_1341,In_585,In_1939);
xnor U1342 (N_1342,In_1911,In_430);
and U1343 (N_1343,In_1769,In_1903);
or U1344 (N_1344,In_857,In_1030);
xor U1345 (N_1345,In_451,In_394);
nor U1346 (N_1346,In_131,In_1468);
and U1347 (N_1347,In_181,In_1373);
nand U1348 (N_1348,In_1730,In_1276);
and U1349 (N_1349,In_1999,In_109);
and U1350 (N_1350,In_1959,In_1654);
nand U1351 (N_1351,In_964,In_334);
or U1352 (N_1352,In_1128,In_607);
nand U1353 (N_1353,In_789,In_65);
or U1354 (N_1354,In_1773,In_1921);
or U1355 (N_1355,In_1201,In_108);
nor U1356 (N_1356,In_1973,In_369);
or U1357 (N_1357,In_1467,In_1640);
and U1358 (N_1358,In_1028,In_720);
and U1359 (N_1359,In_1929,In_376);
xnor U1360 (N_1360,In_1193,In_723);
or U1361 (N_1361,In_1208,In_416);
or U1362 (N_1362,In_1575,In_966);
or U1363 (N_1363,In_1359,In_1059);
nor U1364 (N_1364,In_834,In_192);
nand U1365 (N_1365,In_1795,In_1505);
or U1366 (N_1366,In_1265,In_180);
or U1367 (N_1367,In_860,In_596);
xnor U1368 (N_1368,In_1890,In_110);
or U1369 (N_1369,In_239,In_528);
nand U1370 (N_1370,In_1327,In_1895);
and U1371 (N_1371,In_1478,In_594);
and U1372 (N_1372,In_334,In_937);
nor U1373 (N_1373,In_78,In_374);
and U1374 (N_1374,In_838,In_739);
and U1375 (N_1375,In_19,In_1704);
or U1376 (N_1376,In_532,In_77);
or U1377 (N_1377,In_1091,In_1009);
nand U1378 (N_1378,In_1565,In_751);
or U1379 (N_1379,In_836,In_1364);
nor U1380 (N_1380,In_134,In_1697);
and U1381 (N_1381,In_738,In_1185);
xnor U1382 (N_1382,In_367,In_1191);
nor U1383 (N_1383,In_1278,In_1700);
or U1384 (N_1384,In_1857,In_1288);
nand U1385 (N_1385,In_570,In_1746);
nand U1386 (N_1386,In_436,In_1604);
or U1387 (N_1387,In_196,In_927);
and U1388 (N_1388,In_425,In_1033);
or U1389 (N_1389,In_1164,In_707);
nor U1390 (N_1390,In_554,In_236);
and U1391 (N_1391,In_63,In_963);
or U1392 (N_1392,In_1774,In_1614);
and U1393 (N_1393,In_1685,In_1602);
and U1394 (N_1394,In_180,In_205);
or U1395 (N_1395,In_1235,In_1788);
nor U1396 (N_1396,In_227,In_1252);
xnor U1397 (N_1397,In_523,In_1761);
or U1398 (N_1398,In_1845,In_1075);
and U1399 (N_1399,In_1892,In_103);
and U1400 (N_1400,In_821,In_1890);
and U1401 (N_1401,In_1918,In_1593);
or U1402 (N_1402,In_474,In_526);
and U1403 (N_1403,In_1370,In_397);
nand U1404 (N_1404,In_1890,In_231);
or U1405 (N_1405,In_61,In_1955);
nor U1406 (N_1406,In_1520,In_1910);
nor U1407 (N_1407,In_732,In_1407);
nor U1408 (N_1408,In_1843,In_799);
or U1409 (N_1409,In_1293,In_1627);
nor U1410 (N_1410,In_845,In_868);
nand U1411 (N_1411,In_414,In_1804);
and U1412 (N_1412,In_1185,In_1832);
or U1413 (N_1413,In_1187,In_1045);
or U1414 (N_1414,In_704,In_420);
nor U1415 (N_1415,In_712,In_1132);
or U1416 (N_1416,In_825,In_438);
nand U1417 (N_1417,In_749,In_686);
nor U1418 (N_1418,In_1355,In_825);
and U1419 (N_1419,In_654,In_1469);
nor U1420 (N_1420,In_21,In_1728);
nor U1421 (N_1421,In_1802,In_690);
or U1422 (N_1422,In_766,In_1566);
nand U1423 (N_1423,In_413,In_984);
nor U1424 (N_1424,In_1036,In_240);
nor U1425 (N_1425,In_1067,In_1843);
nor U1426 (N_1426,In_1970,In_1239);
or U1427 (N_1427,In_1898,In_1262);
nand U1428 (N_1428,In_279,In_638);
xnor U1429 (N_1429,In_892,In_1095);
nor U1430 (N_1430,In_1460,In_277);
or U1431 (N_1431,In_463,In_137);
or U1432 (N_1432,In_1682,In_478);
or U1433 (N_1433,In_1284,In_687);
or U1434 (N_1434,In_1437,In_338);
nand U1435 (N_1435,In_71,In_1896);
nand U1436 (N_1436,In_1904,In_1879);
and U1437 (N_1437,In_760,In_362);
and U1438 (N_1438,In_255,In_1598);
or U1439 (N_1439,In_1432,In_210);
nor U1440 (N_1440,In_1459,In_1044);
and U1441 (N_1441,In_1023,In_389);
or U1442 (N_1442,In_971,In_610);
and U1443 (N_1443,In_1866,In_1980);
or U1444 (N_1444,In_1839,In_606);
or U1445 (N_1445,In_1812,In_1773);
nor U1446 (N_1446,In_787,In_1271);
and U1447 (N_1447,In_1238,In_580);
and U1448 (N_1448,In_157,In_1297);
nand U1449 (N_1449,In_1354,In_1952);
nor U1450 (N_1450,In_647,In_72);
nand U1451 (N_1451,In_500,In_1494);
nor U1452 (N_1452,In_1644,In_580);
or U1453 (N_1453,In_267,In_1123);
and U1454 (N_1454,In_331,In_41);
nand U1455 (N_1455,In_103,In_210);
nand U1456 (N_1456,In_1656,In_355);
xor U1457 (N_1457,In_1351,In_528);
nand U1458 (N_1458,In_990,In_382);
xor U1459 (N_1459,In_1454,In_9);
and U1460 (N_1460,In_1663,In_297);
nand U1461 (N_1461,In_1767,In_1825);
nor U1462 (N_1462,In_1478,In_13);
nand U1463 (N_1463,In_640,In_963);
xnor U1464 (N_1464,In_596,In_1495);
or U1465 (N_1465,In_1327,In_1145);
and U1466 (N_1466,In_1849,In_339);
nand U1467 (N_1467,In_779,In_473);
or U1468 (N_1468,In_731,In_137);
nor U1469 (N_1469,In_1565,In_865);
or U1470 (N_1470,In_16,In_220);
nor U1471 (N_1471,In_64,In_371);
nor U1472 (N_1472,In_453,In_43);
nor U1473 (N_1473,In_384,In_1554);
and U1474 (N_1474,In_1356,In_1718);
and U1475 (N_1475,In_1804,In_1617);
nor U1476 (N_1476,In_1906,In_210);
or U1477 (N_1477,In_187,In_572);
and U1478 (N_1478,In_1152,In_332);
nand U1479 (N_1479,In_1784,In_1314);
nand U1480 (N_1480,In_482,In_1391);
or U1481 (N_1481,In_1298,In_5);
or U1482 (N_1482,In_342,In_1053);
or U1483 (N_1483,In_718,In_1182);
and U1484 (N_1484,In_807,In_1577);
xor U1485 (N_1485,In_954,In_390);
nor U1486 (N_1486,In_120,In_1444);
and U1487 (N_1487,In_595,In_462);
or U1488 (N_1488,In_510,In_1842);
or U1489 (N_1489,In_1356,In_1990);
and U1490 (N_1490,In_694,In_1997);
nor U1491 (N_1491,In_788,In_1808);
and U1492 (N_1492,In_113,In_1565);
nand U1493 (N_1493,In_392,In_1436);
or U1494 (N_1494,In_1066,In_313);
nand U1495 (N_1495,In_766,In_1631);
nor U1496 (N_1496,In_443,In_285);
nand U1497 (N_1497,In_1641,In_2);
and U1498 (N_1498,In_1736,In_1188);
nand U1499 (N_1499,In_212,In_990);
or U1500 (N_1500,In_772,In_1750);
nor U1501 (N_1501,In_786,In_1868);
or U1502 (N_1502,In_1442,In_1312);
and U1503 (N_1503,In_269,In_1064);
and U1504 (N_1504,In_588,In_1387);
nor U1505 (N_1505,In_936,In_225);
or U1506 (N_1506,In_1612,In_95);
or U1507 (N_1507,In_162,In_11);
nand U1508 (N_1508,In_570,In_217);
and U1509 (N_1509,In_709,In_1680);
and U1510 (N_1510,In_927,In_1886);
and U1511 (N_1511,In_1919,In_1897);
and U1512 (N_1512,In_245,In_1141);
and U1513 (N_1513,In_355,In_414);
or U1514 (N_1514,In_466,In_1824);
and U1515 (N_1515,In_1291,In_431);
nor U1516 (N_1516,In_683,In_1473);
and U1517 (N_1517,In_1818,In_842);
nor U1518 (N_1518,In_451,In_1860);
or U1519 (N_1519,In_627,In_1181);
and U1520 (N_1520,In_1518,In_1636);
and U1521 (N_1521,In_1603,In_221);
nand U1522 (N_1522,In_1336,In_106);
xor U1523 (N_1523,In_239,In_119);
xnor U1524 (N_1524,In_1950,In_616);
or U1525 (N_1525,In_1008,In_1401);
nand U1526 (N_1526,In_1891,In_575);
or U1527 (N_1527,In_1531,In_1145);
nor U1528 (N_1528,In_1812,In_1787);
and U1529 (N_1529,In_969,In_776);
and U1530 (N_1530,In_1649,In_870);
nand U1531 (N_1531,In_783,In_1589);
or U1532 (N_1532,In_317,In_11);
xnor U1533 (N_1533,In_1677,In_494);
nand U1534 (N_1534,In_173,In_883);
and U1535 (N_1535,In_252,In_34);
xor U1536 (N_1536,In_191,In_354);
xor U1537 (N_1537,In_419,In_546);
or U1538 (N_1538,In_1790,In_509);
nand U1539 (N_1539,In_1096,In_1233);
and U1540 (N_1540,In_1476,In_238);
or U1541 (N_1541,In_69,In_1837);
and U1542 (N_1542,In_133,In_1693);
or U1543 (N_1543,In_1202,In_1210);
nor U1544 (N_1544,In_1906,In_466);
nand U1545 (N_1545,In_453,In_830);
nand U1546 (N_1546,In_95,In_1984);
nor U1547 (N_1547,In_1916,In_1340);
or U1548 (N_1548,In_673,In_346);
nor U1549 (N_1549,In_1809,In_130);
and U1550 (N_1550,In_559,In_337);
or U1551 (N_1551,In_704,In_510);
or U1552 (N_1552,In_1606,In_1470);
nand U1553 (N_1553,In_1725,In_661);
or U1554 (N_1554,In_178,In_185);
or U1555 (N_1555,In_1568,In_1976);
nand U1556 (N_1556,In_796,In_197);
nand U1557 (N_1557,In_857,In_17);
and U1558 (N_1558,In_309,In_247);
nor U1559 (N_1559,In_743,In_825);
nand U1560 (N_1560,In_1299,In_398);
or U1561 (N_1561,In_986,In_1963);
nand U1562 (N_1562,In_1471,In_395);
or U1563 (N_1563,In_534,In_821);
nor U1564 (N_1564,In_1676,In_995);
nand U1565 (N_1565,In_1748,In_492);
nor U1566 (N_1566,In_1953,In_93);
nand U1567 (N_1567,In_158,In_1434);
and U1568 (N_1568,In_636,In_518);
xnor U1569 (N_1569,In_1588,In_926);
nand U1570 (N_1570,In_1917,In_384);
xnor U1571 (N_1571,In_1961,In_875);
and U1572 (N_1572,In_271,In_986);
nand U1573 (N_1573,In_1786,In_10);
and U1574 (N_1574,In_531,In_578);
or U1575 (N_1575,In_827,In_641);
nand U1576 (N_1576,In_242,In_1391);
nor U1577 (N_1577,In_84,In_1663);
or U1578 (N_1578,In_351,In_466);
or U1579 (N_1579,In_1219,In_722);
and U1580 (N_1580,In_897,In_1118);
nand U1581 (N_1581,In_1113,In_654);
nor U1582 (N_1582,In_1103,In_1015);
and U1583 (N_1583,In_549,In_1108);
and U1584 (N_1584,In_258,In_1143);
or U1585 (N_1585,In_1034,In_1980);
nand U1586 (N_1586,In_1227,In_1600);
nand U1587 (N_1587,In_624,In_568);
and U1588 (N_1588,In_1355,In_19);
nand U1589 (N_1589,In_522,In_269);
and U1590 (N_1590,In_730,In_124);
and U1591 (N_1591,In_1305,In_577);
nand U1592 (N_1592,In_1167,In_1907);
nand U1593 (N_1593,In_204,In_1011);
or U1594 (N_1594,In_1358,In_1756);
or U1595 (N_1595,In_204,In_763);
or U1596 (N_1596,In_714,In_1708);
nand U1597 (N_1597,In_102,In_1647);
nor U1598 (N_1598,In_1954,In_567);
nand U1599 (N_1599,In_1569,In_1217);
nand U1600 (N_1600,In_1074,In_147);
and U1601 (N_1601,In_483,In_750);
nand U1602 (N_1602,In_699,In_858);
nand U1603 (N_1603,In_38,In_1963);
nand U1604 (N_1604,In_1486,In_310);
nand U1605 (N_1605,In_579,In_278);
and U1606 (N_1606,In_583,In_55);
or U1607 (N_1607,In_418,In_378);
and U1608 (N_1608,In_756,In_1704);
and U1609 (N_1609,In_1427,In_363);
or U1610 (N_1610,In_1367,In_1103);
nand U1611 (N_1611,In_1169,In_776);
or U1612 (N_1612,In_1092,In_583);
and U1613 (N_1613,In_1464,In_574);
nor U1614 (N_1614,In_514,In_1845);
nor U1615 (N_1615,In_976,In_1151);
and U1616 (N_1616,In_136,In_81);
nand U1617 (N_1617,In_817,In_480);
and U1618 (N_1618,In_1581,In_1073);
and U1619 (N_1619,In_1218,In_808);
xor U1620 (N_1620,In_1781,In_887);
xor U1621 (N_1621,In_1520,In_1200);
or U1622 (N_1622,In_186,In_120);
and U1623 (N_1623,In_462,In_1524);
nand U1624 (N_1624,In_1064,In_1856);
or U1625 (N_1625,In_896,In_922);
nand U1626 (N_1626,In_1433,In_1598);
nand U1627 (N_1627,In_1415,In_1615);
or U1628 (N_1628,In_494,In_1964);
nor U1629 (N_1629,In_22,In_751);
nand U1630 (N_1630,In_765,In_1035);
or U1631 (N_1631,In_549,In_474);
and U1632 (N_1632,In_388,In_1742);
xnor U1633 (N_1633,In_1666,In_982);
nor U1634 (N_1634,In_1887,In_1738);
nand U1635 (N_1635,In_128,In_343);
or U1636 (N_1636,In_827,In_1509);
or U1637 (N_1637,In_1284,In_1881);
and U1638 (N_1638,In_1095,In_1663);
nand U1639 (N_1639,In_1547,In_173);
or U1640 (N_1640,In_776,In_344);
or U1641 (N_1641,In_1964,In_768);
nor U1642 (N_1642,In_678,In_1695);
xnor U1643 (N_1643,In_1217,In_1165);
nand U1644 (N_1644,In_362,In_598);
nand U1645 (N_1645,In_334,In_1214);
nor U1646 (N_1646,In_147,In_1563);
and U1647 (N_1647,In_1215,In_1522);
or U1648 (N_1648,In_639,In_571);
nor U1649 (N_1649,In_1043,In_1853);
or U1650 (N_1650,In_907,In_1058);
nor U1651 (N_1651,In_1221,In_1813);
nor U1652 (N_1652,In_1879,In_611);
nand U1653 (N_1653,In_1460,In_816);
nor U1654 (N_1654,In_354,In_1715);
or U1655 (N_1655,In_749,In_1541);
or U1656 (N_1656,In_1933,In_703);
nand U1657 (N_1657,In_824,In_1707);
and U1658 (N_1658,In_1725,In_551);
or U1659 (N_1659,In_389,In_56);
or U1660 (N_1660,In_1865,In_1277);
xor U1661 (N_1661,In_931,In_1906);
or U1662 (N_1662,In_715,In_1232);
nand U1663 (N_1663,In_1749,In_1552);
nand U1664 (N_1664,In_1947,In_1587);
nor U1665 (N_1665,In_1217,In_1767);
and U1666 (N_1666,In_649,In_1995);
and U1667 (N_1667,In_96,In_356);
and U1668 (N_1668,In_1121,In_886);
or U1669 (N_1669,In_284,In_1235);
nor U1670 (N_1670,In_1260,In_119);
or U1671 (N_1671,In_191,In_494);
and U1672 (N_1672,In_1934,In_545);
and U1673 (N_1673,In_1652,In_1617);
or U1674 (N_1674,In_1480,In_1330);
nand U1675 (N_1675,In_968,In_101);
xnor U1676 (N_1676,In_1800,In_475);
nor U1677 (N_1677,In_1307,In_338);
nand U1678 (N_1678,In_1848,In_703);
nor U1679 (N_1679,In_267,In_287);
and U1680 (N_1680,In_1128,In_590);
or U1681 (N_1681,In_605,In_713);
nor U1682 (N_1682,In_1082,In_381);
or U1683 (N_1683,In_1296,In_694);
nand U1684 (N_1684,In_1184,In_1310);
or U1685 (N_1685,In_359,In_1414);
nor U1686 (N_1686,In_1942,In_1099);
nor U1687 (N_1687,In_706,In_1163);
nor U1688 (N_1688,In_1819,In_224);
nor U1689 (N_1689,In_338,In_265);
and U1690 (N_1690,In_903,In_125);
or U1691 (N_1691,In_891,In_1679);
or U1692 (N_1692,In_1771,In_390);
or U1693 (N_1693,In_1321,In_1624);
and U1694 (N_1694,In_311,In_543);
nand U1695 (N_1695,In_91,In_957);
xor U1696 (N_1696,In_1604,In_1892);
nor U1697 (N_1697,In_1307,In_1627);
and U1698 (N_1698,In_540,In_1494);
and U1699 (N_1699,In_1060,In_1421);
nand U1700 (N_1700,In_1054,In_1194);
nand U1701 (N_1701,In_535,In_339);
or U1702 (N_1702,In_1806,In_1498);
xor U1703 (N_1703,In_1528,In_701);
xor U1704 (N_1704,In_1930,In_1180);
or U1705 (N_1705,In_847,In_1505);
and U1706 (N_1706,In_1902,In_1125);
nor U1707 (N_1707,In_1921,In_421);
and U1708 (N_1708,In_1202,In_1580);
or U1709 (N_1709,In_1596,In_1134);
xor U1710 (N_1710,In_1843,In_1484);
and U1711 (N_1711,In_382,In_718);
nand U1712 (N_1712,In_1300,In_129);
xnor U1713 (N_1713,In_1710,In_1485);
and U1714 (N_1714,In_1350,In_640);
and U1715 (N_1715,In_82,In_268);
or U1716 (N_1716,In_131,In_1129);
or U1717 (N_1717,In_1420,In_1220);
nand U1718 (N_1718,In_78,In_1258);
nor U1719 (N_1719,In_443,In_505);
and U1720 (N_1720,In_1398,In_1245);
and U1721 (N_1721,In_1178,In_472);
and U1722 (N_1722,In_1750,In_596);
nor U1723 (N_1723,In_247,In_1700);
or U1724 (N_1724,In_738,In_764);
xor U1725 (N_1725,In_258,In_1534);
and U1726 (N_1726,In_898,In_154);
nor U1727 (N_1727,In_1742,In_1943);
or U1728 (N_1728,In_241,In_233);
and U1729 (N_1729,In_477,In_1544);
xnor U1730 (N_1730,In_517,In_7);
nor U1731 (N_1731,In_912,In_1212);
or U1732 (N_1732,In_205,In_1255);
or U1733 (N_1733,In_421,In_1045);
xnor U1734 (N_1734,In_1074,In_1399);
or U1735 (N_1735,In_7,In_198);
and U1736 (N_1736,In_444,In_1668);
and U1737 (N_1737,In_653,In_159);
and U1738 (N_1738,In_1584,In_936);
and U1739 (N_1739,In_1662,In_1798);
nor U1740 (N_1740,In_1053,In_219);
and U1741 (N_1741,In_583,In_1483);
or U1742 (N_1742,In_1170,In_1613);
nand U1743 (N_1743,In_485,In_1071);
or U1744 (N_1744,In_404,In_1132);
or U1745 (N_1745,In_947,In_886);
nand U1746 (N_1746,In_1584,In_828);
and U1747 (N_1747,In_802,In_1367);
xnor U1748 (N_1748,In_929,In_1287);
or U1749 (N_1749,In_1189,In_904);
or U1750 (N_1750,In_335,In_1627);
nor U1751 (N_1751,In_1157,In_1071);
nand U1752 (N_1752,In_969,In_794);
and U1753 (N_1753,In_465,In_658);
and U1754 (N_1754,In_1927,In_305);
nor U1755 (N_1755,In_669,In_800);
xor U1756 (N_1756,In_626,In_628);
nand U1757 (N_1757,In_1111,In_1609);
xor U1758 (N_1758,In_1173,In_342);
nor U1759 (N_1759,In_1275,In_1651);
nor U1760 (N_1760,In_1720,In_1307);
nor U1761 (N_1761,In_537,In_809);
and U1762 (N_1762,In_728,In_498);
and U1763 (N_1763,In_1134,In_1537);
or U1764 (N_1764,In_891,In_612);
or U1765 (N_1765,In_52,In_1351);
nand U1766 (N_1766,In_1728,In_435);
or U1767 (N_1767,In_1883,In_150);
and U1768 (N_1768,In_103,In_1268);
and U1769 (N_1769,In_553,In_1314);
or U1770 (N_1770,In_1683,In_1434);
or U1771 (N_1771,In_660,In_1603);
or U1772 (N_1772,In_1044,In_258);
nor U1773 (N_1773,In_1364,In_707);
or U1774 (N_1774,In_1042,In_276);
nor U1775 (N_1775,In_1564,In_1537);
and U1776 (N_1776,In_895,In_1657);
and U1777 (N_1777,In_1766,In_1010);
nor U1778 (N_1778,In_218,In_863);
nand U1779 (N_1779,In_1141,In_1277);
and U1780 (N_1780,In_1210,In_1584);
and U1781 (N_1781,In_1095,In_392);
and U1782 (N_1782,In_1680,In_1424);
nand U1783 (N_1783,In_703,In_1251);
nand U1784 (N_1784,In_1227,In_1255);
nand U1785 (N_1785,In_1729,In_1247);
and U1786 (N_1786,In_461,In_657);
and U1787 (N_1787,In_616,In_749);
or U1788 (N_1788,In_557,In_579);
nand U1789 (N_1789,In_1593,In_624);
or U1790 (N_1790,In_522,In_342);
nand U1791 (N_1791,In_1220,In_1765);
or U1792 (N_1792,In_1609,In_804);
xor U1793 (N_1793,In_255,In_1458);
nand U1794 (N_1794,In_1290,In_287);
nor U1795 (N_1795,In_1193,In_1176);
nand U1796 (N_1796,In_253,In_52);
nor U1797 (N_1797,In_1219,In_825);
xor U1798 (N_1798,In_312,In_1706);
or U1799 (N_1799,In_1959,In_1387);
and U1800 (N_1800,In_1735,In_1452);
and U1801 (N_1801,In_1270,In_801);
and U1802 (N_1802,In_1357,In_749);
and U1803 (N_1803,In_1794,In_1029);
nand U1804 (N_1804,In_1736,In_1503);
nor U1805 (N_1805,In_845,In_1771);
or U1806 (N_1806,In_1846,In_1706);
and U1807 (N_1807,In_1523,In_1821);
and U1808 (N_1808,In_1399,In_1297);
nand U1809 (N_1809,In_1056,In_272);
and U1810 (N_1810,In_567,In_1289);
and U1811 (N_1811,In_1720,In_1259);
and U1812 (N_1812,In_1845,In_1951);
or U1813 (N_1813,In_653,In_210);
and U1814 (N_1814,In_1634,In_1124);
and U1815 (N_1815,In_744,In_1897);
nor U1816 (N_1816,In_1241,In_50);
xor U1817 (N_1817,In_10,In_1001);
and U1818 (N_1818,In_1503,In_1572);
xor U1819 (N_1819,In_679,In_120);
nor U1820 (N_1820,In_966,In_283);
nor U1821 (N_1821,In_570,In_792);
nor U1822 (N_1822,In_1687,In_1757);
and U1823 (N_1823,In_1852,In_1833);
xor U1824 (N_1824,In_189,In_720);
or U1825 (N_1825,In_1862,In_803);
nand U1826 (N_1826,In_219,In_1089);
nor U1827 (N_1827,In_1437,In_991);
or U1828 (N_1828,In_1014,In_1948);
or U1829 (N_1829,In_1935,In_1894);
or U1830 (N_1830,In_1914,In_416);
and U1831 (N_1831,In_1501,In_1800);
nand U1832 (N_1832,In_377,In_859);
xnor U1833 (N_1833,In_1734,In_781);
xor U1834 (N_1834,In_1567,In_470);
or U1835 (N_1835,In_984,In_421);
and U1836 (N_1836,In_336,In_1275);
nand U1837 (N_1837,In_620,In_246);
nor U1838 (N_1838,In_1607,In_21);
nor U1839 (N_1839,In_866,In_306);
nand U1840 (N_1840,In_868,In_1138);
xnor U1841 (N_1841,In_1645,In_1512);
nor U1842 (N_1842,In_444,In_52);
nor U1843 (N_1843,In_1415,In_147);
nand U1844 (N_1844,In_563,In_566);
nor U1845 (N_1845,In_152,In_645);
or U1846 (N_1846,In_806,In_1064);
nand U1847 (N_1847,In_1850,In_1101);
or U1848 (N_1848,In_974,In_1264);
nor U1849 (N_1849,In_399,In_631);
nor U1850 (N_1850,In_107,In_752);
nor U1851 (N_1851,In_1822,In_1993);
or U1852 (N_1852,In_319,In_612);
nor U1853 (N_1853,In_8,In_1219);
nand U1854 (N_1854,In_1781,In_838);
and U1855 (N_1855,In_1067,In_1574);
xnor U1856 (N_1856,In_329,In_609);
nor U1857 (N_1857,In_1194,In_1312);
and U1858 (N_1858,In_773,In_1412);
nor U1859 (N_1859,In_907,In_975);
and U1860 (N_1860,In_123,In_886);
nand U1861 (N_1861,In_1310,In_1983);
nand U1862 (N_1862,In_1132,In_1413);
or U1863 (N_1863,In_1422,In_1996);
nand U1864 (N_1864,In_1063,In_1870);
nand U1865 (N_1865,In_1036,In_1000);
or U1866 (N_1866,In_808,In_984);
and U1867 (N_1867,In_258,In_718);
nand U1868 (N_1868,In_1297,In_1653);
and U1869 (N_1869,In_938,In_1648);
nand U1870 (N_1870,In_1273,In_1704);
nand U1871 (N_1871,In_1902,In_1976);
and U1872 (N_1872,In_1182,In_1370);
nor U1873 (N_1873,In_1035,In_1548);
nand U1874 (N_1874,In_1626,In_1538);
nor U1875 (N_1875,In_257,In_1127);
xor U1876 (N_1876,In_746,In_1598);
or U1877 (N_1877,In_1528,In_1152);
or U1878 (N_1878,In_375,In_179);
or U1879 (N_1879,In_1350,In_1119);
and U1880 (N_1880,In_1555,In_1330);
nand U1881 (N_1881,In_1508,In_346);
nor U1882 (N_1882,In_1628,In_1339);
and U1883 (N_1883,In_917,In_43);
and U1884 (N_1884,In_462,In_195);
and U1885 (N_1885,In_249,In_1991);
or U1886 (N_1886,In_1361,In_816);
nor U1887 (N_1887,In_213,In_684);
and U1888 (N_1888,In_738,In_447);
and U1889 (N_1889,In_1788,In_487);
and U1890 (N_1890,In_1503,In_186);
and U1891 (N_1891,In_1856,In_945);
nor U1892 (N_1892,In_1146,In_415);
and U1893 (N_1893,In_993,In_1605);
or U1894 (N_1894,In_1094,In_1326);
nand U1895 (N_1895,In_313,In_21);
or U1896 (N_1896,In_483,In_1135);
nand U1897 (N_1897,In_1407,In_1890);
or U1898 (N_1898,In_1024,In_1179);
nor U1899 (N_1899,In_370,In_1548);
nor U1900 (N_1900,In_1933,In_1973);
nor U1901 (N_1901,In_662,In_476);
nand U1902 (N_1902,In_1693,In_138);
xor U1903 (N_1903,In_1139,In_1351);
and U1904 (N_1904,In_425,In_1180);
nor U1905 (N_1905,In_328,In_746);
nor U1906 (N_1906,In_308,In_52);
and U1907 (N_1907,In_1314,In_121);
nand U1908 (N_1908,In_510,In_417);
nor U1909 (N_1909,In_916,In_1815);
or U1910 (N_1910,In_554,In_1740);
nand U1911 (N_1911,In_12,In_850);
or U1912 (N_1912,In_1311,In_740);
or U1913 (N_1913,In_1453,In_1132);
nor U1914 (N_1914,In_1,In_1620);
nor U1915 (N_1915,In_1769,In_1298);
xor U1916 (N_1916,In_770,In_1537);
nand U1917 (N_1917,In_235,In_1984);
nor U1918 (N_1918,In_917,In_346);
and U1919 (N_1919,In_570,In_1348);
nand U1920 (N_1920,In_607,In_1123);
nand U1921 (N_1921,In_666,In_723);
nand U1922 (N_1922,In_548,In_172);
nor U1923 (N_1923,In_1020,In_348);
nor U1924 (N_1924,In_744,In_436);
nor U1925 (N_1925,In_769,In_110);
nand U1926 (N_1926,In_1097,In_529);
nor U1927 (N_1927,In_763,In_1217);
or U1928 (N_1928,In_1360,In_254);
and U1929 (N_1929,In_1334,In_1615);
nand U1930 (N_1930,In_1738,In_174);
nor U1931 (N_1931,In_721,In_720);
and U1932 (N_1932,In_63,In_516);
and U1933 (N_1933,In_1391,In_892);
or U1934 (N_1934,In_1764,In_1267);
and U1935 (N_1935,In_960,In_1448);
xnor U1936 (N_1936,In_1507,In_1676);
or U1937 (N_1937,In_767,In_1962);
nand U1938 (N_1938,In_1871,In_1308);
nand U1939 (N_1939,In_1107,In_1401);
or U1940 (N_1940,In_49,In_1689);
or U1941 (N_1941,In_1681,In_414);
or U1942 (N_1942,In_675,In_969);
nand U1943 (N_1943,In_1705,In_394);
nand U1944 (N_1944,In_1670,In_931);
nand U1945 (N_1945,In_1253,In_1993);
nor U1946 (N_1946,In_14,In_1032);
or U1947 (N_1947,In_1347,In_63);
nand U1948 (N_1948,In_1178,In_858);
nor U1949 (N_1949,In_208,In_1773);
and U1950 (N_1950,In_558,In_459);
and U1951 (N_1951,In_1959,In_79);
or U1952 (N_1952,In_696,In_1952);
and U1953 (N_1953,In_1128,In_221);
xor U1954 (N_1954,In_165,In_1292);
nor U1955 (N_1955,In_776,In_1608);
nor U1956 (N_1956,In_721,In_802);
xnor U1957 (N_1957,In_1419,In_1619);
xor U1958 (N_1958,In_1285,In_414);
nor U1959 (N_1959,In_11,In_1440);
nor U1960 (N_1960,In_1093,In_951);
and U1961 (N_1961,In_884,In_271);
or U1962 (N_1962,In_1409,In_923);
and U1963 (N_1963,In_1985,In_1448);
or U1964 (N_1964,In_656,In_1000);
xnor U1965 (N_1965,In_245,In_622);
nor U1966 (N_1966,In_773,In_772);
nand U1967 (N_1967,In_675,In_465);
nor U1968 (N_1968,In_1684,In_1927);
or U1969 (N_1969,In_1580,In_1052);
nor U1970 (N_1970,In_1149,In_1247);
nor U1971 (N_1971,In_872,In_1956);
nand U1972 (N_1972,In_1045,In_1192);
nor U1973 (N_1973,In_882,In_645);
or U1974 (N_1974,In_841,In_1822);
nor U1975 (N_1975,In_1202,In_1793);
nor U1976 (N_1976,In_1886,In_296);
or U1977 (N_1977,In_755,In_1639);
nor U1978 (N_1978,In_793,In_1447);
nor U1979 (N_1979,In_64,In_1182);
or U1980 (N_1980,In_1212,In_1576);
and U1981 (N_1981,In_1751,In_1833);
nand U1982 (N_1982,In_1240,In_1751);
nor U1983 (N_1983,In_1206,In_1351);
nand U1984 (N_1984,In_39,In_732);
and U1985 (N_1985,In_214,In_1563);
nor U1986 (N_1986,In_1436,In_310);
nor U1987 (N_1987,In_745,In_1043);
nor U1988 (N_1988,In_877,In_97);
nand U1989 (N_1989,In_1072,In_1430);
and U1990 (N_1990,In_1010,In_350);
nand U1991 (N_1991,In_168,In_620);
nand U1992 (N_1992,In_181,In_548);
or U1993 (N_1993,In_1225,In_1993);
xor U1994 (N_1994,In_1535,In_813);
and U1995 (N_1995,In_1478,In_773);
and U1996 (N_1996,In_1449,In_719);
nand U1997 (N_1997,In_1412,In_338);
nor U1998 (N_1998,In_357,In_1503);
or U1999 (N_1999,In_1714,In_973);
xor U2000 (N_2000,In_1310,In_912);
and U2001 (N_2001,In_1724,In_575);
nor U2002 (N_2002,In_707,In_426);
and U2003 (N_2003,In_975,In_1985);
and U2004 (N_2004,In_1026,In_65);
nand U2005 (N_2005,In_1071,In_1718);
and U2006 (N_2006,In_619,In_457);
or U2007 (N_2007,In_1306,In_1599);
and U2008 (N_2008,In_1042,In_1429);
nor U2009 (N_2009,In_912,In_793);
nand U2010 (N_2010,In_142,In_1841);
and U2011 (N_2011,In_508,In_720);
or U2012 (N_2012,In_1009,In_206);
nor U2013 (N_2013,In_1893,In_524);
nor U2014 (N_2014,In_1234,In_1889);
nor U2015 (N_2015,In_1145,In_277);
or U2016 (N_2016,In_306,In_202);
nor U2017 (N_2017,In_1568,In_330);
nor U2018 (N_2018,In_154,In_1511);
and U2019 (N_2019,In_850,In_722);
or U2020 (N_2020,In_1211,In_813);
nand U2021 (N_2021,In_1410,In_1708);
or U2022 (N_2022,In_1011,In_610);
nand U2023 (N_2023,In_845,In_1321);
or U2024 (N_2024,In_1268,In_1137);
xnor U2025 (N_2025,In_1467,In_416);
or U2026 (N_2026,In_479,In_1599);
and U2027 (N_2027,In_1416,In_1573);
or U2028 (N_2028,In_216,In_285);
or U2029 (N_2029,In_1690,In_251);
or U2030 (N_2030,In_1705,In_1577);
and U2031 (N_2031,In_740,In_1949);
nand U2032 (N_2032,In_650,In_1702);
and U2033 (N_2033,In_1770,In_359);
or U2034 (N_2034,In_1005,In_1414);
and U2035 (N_2035,In_1314,In_1720);
or U2036 (N_2036,In_1095,In_1116);
and U2037 (N_2037,In_1828,In_1897);
nor U2038 (N_2038,In_1661,In_1271);
nand U2039 (N_2039,In_323,In_1035);
or U2040 (N_2040,In_1975,In_1057);
nor U2041 (N_2041,In_1207,In_1339);
or U2042 (N_2042,In_1678,In_532);
or U2043 (N_2043,In_61,In_1655);
and U2044 (N_2044,In_1223,In_98);
or U2045 (N_2045,In_1651,In_1782);
and U2046 (N_2046,In_1690,In_483);
nand U2047 (N_2047,In_888,In_1821);
nand U2048 (N_2048,In_925,In_776);
nor U2049 (N_2049,In_1129,In_155);
or U2050 (N_2050,In_1968,In_274);
and U2051 (N_2051,In_1094,In_1594);
nor U2052 (N_2052,In_1539,In_1771);
and U2053 (N_2053,In_1570,In_1424);
and U2054 (N_2054,In_1267,In_745);
nor U2055 (N_2055,In_1885,In_38);
nor U2056 (N_2056,In_1770,In_824);
or U2057 (N_2057,In_258,In_1950);
and U2058 (N_2058,In_1693,In_1467);
nor U2059 (N_2059,In_1485,In_1904);
or U2060 (N_2060,In_470,In_1960);
xor U2061 (N_2061,In_1619,In_1350);
and U2062 (N_2062,In_1188,In_288);
and U2063 (N_2063,In_1130,In_1536);
and U2064 (N_2064,In_1587,In_1284);
nor U2065 (N_2065,In_1195,In_759);
nand U2066 (N_2066,In_18,In_286);
and U2067 (N_2067,In_1197,In_280);
and U2068 (N_2068,In_1227,In_1919);
nor U2069 (N_2069,In_324,In_115);
nand U2070 (N_2070,In_728,In_897);
nand U2071 (N_2071,In_1704,In_30);
nor U2072 (N_2072,In_1455,In_1324);
xor U2073 (N_2073,In_826,In_530);
and U2074 (N_2074,In_78,In_1377);
or U2075 (N_2075,In_927,In_16);
nor U2076 (N_2076,In_1056,In_1137);
and U2077 (N_2077,In_1952,In_1817);
and U2078 (N_2078,In_1511,In_1886);
nand U2079 (N_2079,In_832,In_158);
nor U2080 (N_2080,In_125,In_647);
or U2081 (N_2081,In_186,In_956);
nor U2082 (N_2082,In_1600,In_862);
nor U2083 (N_2083,In_659,In_1335);
nand U2084 (N_2084,In_1966,In_1845);
nor U2085 (N_2085,In_1785,In_88);
and U2086 (N_2086,In_680,In_2);
or U2087 (N_2087,In_1454,In_1510);
or U2088 (N_2088,In_1515,In_59);
or U2089 (N_2089,In_1769,In_1287);
and U2090 (N_2090,In_267,In_63);
nand U2091 (N_2091,In_1887,In_887);
nor U2092 (N_2092,In_1283,In_464);
nor U2093 (N_2093,In_1727,In_324);
nand U2094 (N_2094,In_394,In_745);
nand U2095 (N_2095,In_1950,In_427);
nor U2096 (N_2096,In_1196,In_444);
nand U2097 (N_2097,In_818,In_693);
xor U2098 (N_2098,In_889,In_452);
nor U2099 (N_2099,In_325,In_959);
nor U2100 (N_2100,In_297,In_672);
nor U2101 (N_2101,In_1379,In_1997);
nand U2102 (N_2102,In_1831,In_287);
nor U2103 (N_2103,In_1208,In_808);
xnor U2104 (N_2104,In_787,In_394);
nand U2105 (N_2105,In_1355,In_740);
nand U2106 (N_2106,In_1906,In_1854);
xnor U2107 (N_2107,In_170,In_1152);
or U2108 (N_2108,In_1489,In_1879);
and U2109 (N_2109,In_1572,In_1596);
or U2110 (N_2110,In_455,In_1473);
nand U2111 (N_2111,In_461,In_1740);
nand U2112 (N_2112,In_1712,In_118);
and U2113 (N_2113,In_1551,In_1784);
nor U2114 (N_2114,In_1096,In_1518);
and U2115 (N_2115,In_18,In_1290);
or U2116 (N_2116,In_1606,In_1124);
or U2117 (N_2117,In_1885,In_25);
nand U2118 (N_2118,In_1722,In_365);
and U2119 (N_2119,In_1113,In_1962);
nor U2120 (N_2120,In_514,In_602);
or U2121 (N_2121,In_888,In_147);
and U2122 (N_2122,In_196,In_1894);
xnor U2123 (N_2123,In_1974,In_1971);
nor U2124 (N_2124,In_975,In_1751);
nand U2125 (N_2125,In_1954,In_1643);
or U2126 (N_2126,In_108,In_896);
or U2127 (N_2127,In_1450,In_1019);
or U2128 (N_2128,In_1670,In_1501);
xnor U2129 (N_2129,In_852,In_978);
nor U2130 (N_2130,In_1048,In_1215);
xor U2131 (N_2131,In_811,In_1440);
and U2132 (N_2132,In_1512,In_1693);
and U2133 (N_2133,In_886,In_719);
and U2134 (N_2134,In_1167,In_371);
nand U2135 (N_2135,In_6,In_1023);
nor U2136 (N_2136,In_1304,In_1629);
nand U2137 (N_2137,In_1741,In_1161);
and U2138 (N_2138,In_1619,In_334);
nand U2139 (N_2139,In_247,In_876);
and U2140 (N_2140,In_659,In_1160);
nand U2141 (N_2141,In_556,In_1144);
nand U2142 (N_2142,In_716,In_125);
nand U2143 (N_2143,In_642,In_888);
nor U2144 (N_2144,In_765,In_1172);
and U2145 (N_2145,In_1931,In_1624);
nand U2146 (N_2146,In_385,In_1081);
nor U2147 (N_2147,In_1459,In_212);
nand U2148 (N_2148,In_191,In_54);
nor U2149 (N_2149,In_743,In_935);
nor U2150 (N_2150,In_1395,In_3);
and U2151 (N_2151,In_1734,In_1584);
nor U2152 (N_2152,In_1064,In_842);
nand U2153 (N_2153,In_652,In_1399);
and U2154 (N_2154,In_640,In_1246);
and U2155 (N_2155,In_812,In_1999);
nand U2156 (N_2156,In_1600,In_1490);
and U2157 (N_2157,In_938,In_440);
and U2158 (N_2158,In_1559,In_1327);
nand U2159 (N_2159,In_171,In_612);
nand U2160 (N_2160,In_1917,In_693);
or U2161 (N_2161,In_1895,In_960);
nand U2162 (N_2162,In_784,In_775);
nor U2163 (N_2163,In_1471,In_1241);
nand U2164 (N_2164,In_1247,In_1535);
or U2165 (N_2165,In_1601,In_1738);
or U2166 (N_2166,In_1922,In_573);
nor U2167 (N_2167,In_894,In_1079);
and U2168 (N_2168,In_908,In_237);
and U2169 (N_2169,In_1938,In_1797);
nor U2170 (N_2170,In_8,In_1076);
or U2171 (N_2171,In_1192,In_473);
nand U2172 (N_2172,In_251,In_1102);
nor U2173 (N_2173,In_19,In_88);
xnor U2174 (N_2174,In_156,In_1607);
nor U2175 (N_2175,In_151,In_870);
nor U2176 (N_2176,In_227,In_1248);
nor U2177 (N_2177,In_0,In_1193);
nand U2178 (N_2178,In_1345,In_1827);
and U2179 (N_2179,In_357,In_27);
xor U2180 (N_2180,In_134,In_621);
nand U2181 (N_2181,In_1333,In_147);
nand U2182 (N_2182,In_1550,In_34);
nor U2183 (N_2183,In_720,In_1359);
or U2184 (N_2184,In_406,In_219);
nor U2185 (N_2185,In_1418,In_381);
xor U2186 (N_2186,In_507,In_680);
nand U2187 (N_2187,In_1381,In_1691);
and U2188 (N_2188,In_1076,In_282);
or U2189 (N_2189,In_1494,In_417);
nand U2190 (N_2190,In_1855,In_1933);
and U2191 (N_2191,In_220,In_8);
and U2192 (N_2192,In_941,In_1412);
nand U2193 (N_2193,In_1799,In_622);
and U2194 (N_2194,In_694,In_506);
or U2195 (N_2195,In_1573,In_121);
nand U2196 (N_2196,In_1265,In_646);
nand U2197 (N_2197,In_1430,In_1544);
and U2198 (N_2198,In_1015,In_1833);
nand U2199 (N_2199,In_1823,In_1910);
nor U2200 (N_2200,In_542,In_1695);
nor U2201 (N_2201,In_1057,In_1184);
xnor U2202 (N_2202,In_259,In_1323);
nand U2203 (N_2203,In_1303,In_914);
nand U2204 (N_2204,In_1897,In_1002);
or U2205 (N_2205,In_954,In_219);
and U2206 (N_2206,In_589,In_1996);
nand U2207 (N_2207,In_93,In_1842);
nand U2208 (N_2208,In_994,In_905);
nor U2209 (N_2209,In_471,In_61);
nor U2210 (N_2210,In_1725,In_1422);
nand U2211 (N_2211,In_1225,In_1696);
xnor U2212 (N_2212,In_540,In_637);
or U2213 (N_2213,In_447,In_1151);
and U2214 (N_2214,In_1612,In_1397);
nor U2215 (N_2215,In_1244,In_1862);
or U2216 (N_2216,In_1080,In_736);
or U2217 (N_2217,In_260,In_913);
nand U2218 (N_2218,In_1297,In_20);
or U2219 (N_2219,In_1940,In_1665);
and U2220 (N_2220,In_1512,In_1240);
nand U2221 (N_2221,In_1593,In_176);
or U2222 (N_2222,In_1854,In_1614);
and U2223 (N_2223,In_1888,In_1157);
nor U2224 (N_2224,In_1916,In_1984);
nor U2225 (N_2225,In_1160,In_1418);
and U2226 (N_2226,In_549,In_1732);
nor U2227 (N_2227,In_1436,In_1732);
or U2228 (N_2228,In_1560,In_1332);
nand U2229 (N_2229,In_707,In_1187);
nor U2230 (N_2230,In_815,In_467);
nor U2231 (N_2231,In_812,In_676);
nand U2232 (N_2232,In_135,In_390);
nand U2233 (N_2233,In_1004,In_1132);
and U2234 (N_2234,In_1961,In_711);
or U2235 (N_2235,In_895,In_60);
nand U2236 (N_2236,In_731,In_172);
nor U2237 (N_2237,In_1372,In_442);
nand U2238 (N_2238,In_718,In_245);
nor U2239 (N_2239,In_641,In_1220);
xnor U2240 (N_2240,In_15,In_1622);
or U2241 (N_2241,In_512,In_1601);
and U2242 (N_2242,In_1995,In_460);
nor U2243 (N_2243,In_876,In_1757);
or U2244 (N_2244,In_77,In_1444);
nor U2245 (N_2245,In_1507,In_1336);
nand U2246 (N_2246,In_666,In_287);
nor U2247 (N_2247,In_481,In_701);
and U2248 (N_2248,In_958,In_922);
nor U2249 (N_2249,In_1149,In_1582);
and U2250 (N_2250,In_1399,In_44);
nor U2251 (N_2251,In_1880,In_986);
nand U2252 (N_2252,In_484,In_53);
nand U2253 (N_2253,In_1444,In_1207);
nand U2254 (N_2254,In_129,In_476);
nor U2255 (N_2255,In_1174,In_636);
nand U2256 (N_2256,In_263,In_1242);
or U2257 (N_2257,In_1811,In_175);
nand U2258 (N_2258,In_611,In_1929);
and U2259 (N_2259,In_8,In_347);
and U2260 (N_2260,In_709,In_1412);
and U2261 (N_2261,In_1614,In_1436);
nor U2262 (N_2262,In_227,In_545);
nand U2263 (N_2263,In_584,In_1064);
or U2264 (N_2264,In_1961,In_498);
nand U2265 (N_2265,In_990,In_1037);
nor U2266 (N_2266,In_994,In_1198);
nand U2267 (N_2267,In_458,In_448);
nor U2268 (N_2268,In_164,In_1613);
or U2269 (N_2269,In_908,In_75);
and U2270 (N_2270,In_452,In_1744);
nor U2271 (N_2271,In_1265,In_381);
and U2272 (N_2272,In_683,In_1390);
xnor U2273 (N_2273,In_684,In_1054);
nand U2274 (N_2274,In_1718,In_1101);
nor U2275 (N_2275,In_1143,In_1238);
xnor U2276 (N_2276,In_885,In_1871);
nor U2277 (N_2277,In_1430,In_1431);
xnor U2278 (N_2278,In_736,In_1470);
or U2279 (N_2279,In_1618,In_1691);
and U2280 (N_2280,In_267,In_767);
or U2281 (N_2281,In_1322,In_161);
nand U2282 (N_2282,In_969,In_1312);
or U2283 (N_2283,In_1937,In_972);
nand U2284 (N_2284,In_66,In_996);
or U2285 (N_2285,In_453,In_1559);
or U2286 (N_2286,In_172,In_1908);
and U2287 (N_2287,In_1016,In_1421);
nand U2288 (N_2288,In_1746,In_1804);
nor U2289 (N_2289,In_1035,In_1857);
nor U2290 (N_2290,In_1055,In_319);
nand U2291 (N_2291,In_784,In_1053);
or U2292 (N_2292,In_607,In_877);
nor U2293 (N_2293,In_157,In_221);
nor U2294 (N_2294,In_898,In_1508);
and U2295 (N_2295,In_1445,In_1537);
nor U2296 (N_2296,In_13,In_817);
nand U2297 (N_2297,In_1887,In_1261);
nor U2298 (N_2298,In_1243,In_1261);
and U2299 (N_2299,In_289,In_1625);
nand U2300 (N_2300,In_417,In_1236);
nor U2301 (N_2301,In_944,In_219);
and U2302 (N_2302,In_959,In_318);
nor U2303 (N_2303,In_1626,In_1962);
nor U2304 (N_2304,In_258,In_1055);
nor U2305 (N_2305,In_1295,In_607);
or U2306 (N_2306,In_823,In_1509);
nor U2307 (N_2307,In_278,In_1292);
nand U2308 (N_2308,In_1707,In_1978);
or U2309 (N_2309,In_346,In_989);
or U2310 (N_2310,In_663,In_1408);
xnor U2311 (N_2311,In_59,In_290);
nand U2312 (N_2312,In_911,In_1530);
nor U2313 (N_2313,In_1048,In_1702);
nand U2314 (N_2314,In_334,In_888);
nor U2315 (N_2315,In_1773,In_709);
nor U2316 (N_2316,In_1196,In_1928);
or U2317 (N_2317,In_123,In_1503);
and U2318 (N_2318,In_649,In_1030);
nor U2319 (N_2319,In_432,In_732);
nand U2320 (N_2320,In_74,In_393);
nand U2321 (N_2321,In_1763,In_687);
and U2322 (N_2322,In_795,In_1595);
nor U2323 (N_2323,In_249,In_1745);
xnor U2324 (N_2324,In_869,In_859);
nor U2325 (N_2325,In_685,In_466);
nand U2326 (N_2326,In_444,In_1259);
nor U2327 (N_2327,In_1129,In_911);
and U2328 (N_2328,In_1724,In_1752);
or U2329 (N_2329,In_999,In_801);
or U2330 (N_2330,In_377,In_38);
xor U2331 (N_2331,In_753,In_456);
xor U2332 (N_2332,In_926,In_249);
nor U2333 (N_2333,In_1940,In_1763);
nor U2334 (N_2334,In_1723,In_1820);
and U2335 (N_2335,In_499,In_1028);
and U2336 (N_2336,In_3,In_431);
and U2337 (N_2337,In_57,In_1689);
nand U2338 (N_2338,In_650,In_1577);
nand U2339 (N_2339,In_1198,In_1449);
and U2340 (N_2340,In_1964,In_1574);
or U2341 (N_2341,In_1194,In_1234);
nand U2342 (N_2342,In_1627,In_402);
nand U2343 (N_2343,In_524,In_1479);
and U2344 (N_2344,In_1809,In_476);
and U2345 (N_2345,In_279,In_1560);
or U2346 (N_2346,In_1996,In_1720);
nand U2347 (N_2347,In_162,In_1584);
nor U2348 (N_2348,In_1035,In_1033);
or U2349 (N_2349,In_1165,In_1242);
nor U2350 (N_2350,In_136,In_1291);
nand U2351 (N_2351,In_191,In_242);
or U2352 (N_2352,In_1212,In_1744);
nand U2353 (N_2353,In_1985,In_1855);
xor U2354 (N_2354,In_1055,In_1786);
or U2355 (N_2355,In_1872,In_6);
nand U2356 (N_2356,In_507,In_1919);
or U2357 (N_2357,In_1256,In_683);
and U2358 (N_2358,In_1524,In_1239);
and U2359 (N_2359,In_309,In_734);
and U2360 (N_2360,In_769,In_363);
or U2361 (N_2361,In_1233,In_1322);
xor U2362 (N_2362,In_1476,In_1515);
and U2363 (N_2363,In_1331,In_1757);
and U2364 (N_2364,In_1564,In_402);
xor U2365 (N_2365,In_637,In_1735);
xor U2366 (N_2366,In_454,In_770);
nor U2367 (N_2367,In_1487,In_1834);
nand U2368 (N_2368,In_1830,In_1338);
nor U2369 (N_2369,In_1541,In_126);
and U2370 (N_2370,In_497,In_116);
xnor U2371 (N_2371,In_1953,In_1035);
nor U2372 (N_2372,In_508,In_844);
nand U2373 (N_2373,In_268,In_805);
nand U2374 (N_2374,In_792,In_1236);
and U2375 (N_2375,In_490,In_1684);
and U2376 (N_2376,In_1562,In_1960);
nor U2377 (N_2377,In_606,In_1096);
nor U2378 (N_2378,In_1104,In_1478);
nor U2379 (N_2379,In_701,In_1885);
and U2380 (N_2380,In_1979,In_1661);
nor U2381 (N_2381,In_1193,In_261);
xor U2382 (N_2382,In_1115,In_478);
xnor U2383 (N_2383,In_1734,In_596);
nor U2384 (N_2384,In_65,In_1078);
xor U2385 (N_2385,In_1852,In_790);
and U2386 (N_2386,In_1283,In_168);
nor U2387 (N_2387,In_635,In_1855);
nor U2388 (N_2388,In_1458,In_500);
and U2389 (N_2389,In_31,In_500);
nor U2390 (N_2390,In_280,In_221);
or U2391 (N_2391,In_24,In_1885);
nand U2392 (N_2392,In_1557,In_1712);
nand U2393 (N_2393,In_70,In_1367);
nor U2394 (N_2394,In_820,In_408);
or U2395 (N_2395,In_1223,In_1868);
or U2396 (N_2396,In_1617,In_1996);
and U2397 (N_2397,In_1566,In_1063);
and U2398 (N_2398,In_1443,In_797);
nor U2399 (N_2399,In_725,In_919);
or U2400 (N_2400,In_1141,In_496);
xnor U2401 (N_2401,In_1728,In_857);
nor U2402 (N_2402,In_546,In_1205);
nor U2403 (N_2403,In_509,In_1454);
nor U2404 (N_2404,In_1658,In_353);
nand U2405 (N_2405,In_349,In_280);
and U2406 (N_2406,In_1085,In_379);
nor U2407 (N_2407,In_1041,In_1848);
or U2408 (N_2408,In_1366,In_779);
or U2409 (N_2409,In_408,In_402);
or U2410 (N_2410,In_458,In_734);
and U2411 (N_2411,In_1044,In_360);
nand U2412 (N_2412,In_1118,In_79);
or U2413 (N_2413,In_1288,In_1515);
nand U2414 (N_2414,In_1548,In_1840);
or U2415 (N_2415,In_87,In_1115);
or U2416 (N_2416,In_543,In_133);
and U2417 (N_2417,In_1314,In_377);
or U2418 (N_2418,In_883,In_543);
and U2419 (N_2419,In_129,In_429);
nand U2420 (N_2420,In_751,In_1756);
nor U2421 (N_2421,In_1327,In_1513);
or U2422 (N_2422,In_1096,In_7);
or U2423 (N_2423,In_331,In_316);
and U2424 (N_2424,In_1298,In_418);
nor U2425 (N_2425,In_1954,In_1847);
and U2426 (N_2426,In_1615,In_1397);
nor U2427 (N_2427,In_318,In_1936);
or U2428 (N_2428,In_12,In_195);
xor U2429 (N_2429,In_909,In_610);
or U2430 (N_2430,In_97,In_1964);
or U2431 (N_2431,In_1808,In_1803);
nand U2432 (N_2432,In_1510,In_697);
and U2433 (N_2433,In_1615,In_1178);
nand U2434 (N_2434,In_1301,In_799);
or U2435 (N_2435,In_1542,In_1599);
or U2436 (N_2436,In_1948,In_642);
and U2437 (N_2437,In_467,In_867);
nand U2438 (N_2438,In_1409,In_308);
nor U2439 (N_2439,In_310,In_142);
xnor U2440 (N_2440,In_1978,In_1240);
or U2441 (N_2441,In_1358,In_931);
nand U2442 (N_2442,In_1496,In_1420);
or U2443 (N_2443,In_828,In_1190);
and U2444 (N_2444,In_1165,In_1743);
or U2445 (N_2445,In_1487,In_19);
nand U2446 (N_2446,In_891,In_344);
xor U2447 (N_2447,In_1461,In_1867);
nor U2448 (N_2448,In_1398,In_900);
nand U2449 (N_2449,In_14,In_27);
and U2450 (N_2450,In_395,In_1230);
nor U2451 (N_2451,In_1796,In_1999);
nand U2452 (N_2452,In_1393,In_609);
xnor U2453 (N_2453,In_1167,In_825);
nand U2454 (N_2454,In_403,In_720);
xnor U2455 (N_2455,In_465,In_507);
and U2456 (N_2456,In_818,In_467);
nor U2457 (N_2457,In_1622,In_721);
or U2458 (N_2458,In_1503,In_733);
nand U2459 (N_2459,In_823,In_1123);
or U2460 (N_2460,In_1658,In_1942);
or U2461 (N_2461,In_143,In_1293);
and U2462 (N_2462,In_1157,In_1322);
nand U2463 (N_2463,In_1372,In_466);
or U2464 (N_2464,In_497,In_324);
xnor U2465 (N_2465,In_1352,In_1396);
or U2466 (N_2466,In_694,In_1696);
nand U2467 (N_2467,In_254,In_1260);
or U2468 (N_2468,In_749,In_849);
nor U2469 (N_2469,In_1224,In_597);
nand U2470 (N_2470,In_344,In_1190);
or U2471 (N_2471,In_500,In_1476);
nor U2472 (N_2472,In_1290,In_1697);
or U2473 (N_2473,In_727,In_1614);
nand U2474 (N_2474,In_1543,In_190);
nor U2475 (N_2475,In_1861,In_1122);
nand U2476 (N_2476,In_348,In_1545);
and U2477 (N_2477,In_173,In_945);
and U2478 (N_2478,In_689,In_1534);
and U2479 (N_2479,In_1880,In_1252);
nor U2480 (N_2480,In_213,In_899);
or U2481 (N_2481,In_614,In_1835);
or U2482 (N_2482,In_229,In_176);
nor U2483 (N_2483,In_664,In_871);
nor U2484 (N_2484,In_925,In_688);
xnor U2485 (N_2485,In_1498,In_1429);
or U2486 (N_2486,In_103,In_1784);
or U2487 (N_2487,In_1153,In_1548);
nor U2488 (N_2488,In_1703,In_313);
or U2489 (N_2489,In_1628,In_1887);
xnor U2490 (N_2490,In_1467,In_132);
and U2491 (N_2491,In_492,In_1133);
nand U2492 (N_2492,In_1415,In_1912);
and U2493 (N_2493,In_1708,In_1699);
or U2494 (N_2494,In_745,In_1966);
nor U2495 (N_2495,In_1706,In_447);
nand U2496 (N_2496,In_382,In_611);
or U2497 (N_2497,In_1430,In_1984);
or U2498 (N_2498,In_1634,In_1768);
or U2499 (N_2499,In_523,In_1835);
or U2500 (N_2500,In_890,In_1297);
nor U2501 (N_2501,In_1654,In_1166);
nand U2502 (N_2502,In_932,In_883);
or U2503 (N_2503,In_1052,In_1970);
nor U2504 (N_2504,In_966,In_1564);
and U2505 (N_2505,In_1017,In_1531);
nand U2506 (N_2506,In_1996,In_1439);
nand U2507 (N_2507,In_178,In_962);
nand U2508 (N_2508,In_1930,In_957);
and U2509 (N_2509,In_811,In_1121);
nand U2510 (N_2510,In_1094,In_1837);
or U2511 (N_2511,In_1380,In_951);
nor U2512 (N_2512,In_1127,In_1145);
and U2513 (N_2513,In_916,In_1469);
xnor U2514 (N_2514,In_1292,In_584);
nor U2515 (N_2515,In_1198,In_1559);
nand U2516 (N_2516,In_613,In_807);
nand U2517 (N_2517,In_594,In_54);
nand U2518 (N_2518,In_228,In_1769);
nand U2519 (N_2519,In_38,In_1014);
nor U2520 (N_2520,In_494,In_1006);
and U2521 (N_2521,In_155,In_1272);
nand U2522 (N_2522,In_1470,In_730);
nor U2523 (N_2523,In_338,In_1795);
and U2524 (N_2524,In_1682,In_383);
nor U2525 (N_2525,In_1693,In_889);
nand U2526 (N_2526,In_1566,In_546);
nand U2527 (N_2527,In_1031,In_141);
nand U2528 (N_2528,In_1102,In_599);
nor U2529 (N_2529,In_1077,In_16);
nor U2530 (N_2530,In_496,In_357);
nor U2531 (N_2531,In_96,In_1889);
xnor U2532 (N_2532,In_1183,In_1866);
or U2533 (N_2533,In_162,In_1943);
and U2534 (N_2534,In_501,In_1503);
nor U2535 (N_2535,In_1973,In_1555);
xnor U2536 (N_2536,In_1003,In_615);
or U2537 (N_2537,In_61,In_520);
and U2538 (N_2538,In_1161,In_428);
nand U2539 (N_2539,In_1983,In_267);
or U2540 (N_2540,In_70,In_1270);
xnor U2541 (N_2541,In_550,In_251);
and U2542 (N_2542,In_1759,In_1141);
xnor U2543 (N_2543,In_1496,In_935);
nand U2544 (N_2544,In_674,In_1270);
or U2545 (N_2545,In_1411,In_149);
nand U2546 (N_2546,In_380,In_1956);
or U2547 (N_2547,In_1307,In_1718);
nand U2548 (N_2548,In_1957,In_72);
and U2549 (N_2549,In_1579,In_1093);
xor U2550 (N_2550,In_1223,In_818);
nor U2551 (N_2551,In_1772,In_659);
xnor U2552 (N_2552,In_1898,In_1003);
xor U2553 (N_2553,In_593,In_1242);
xnor U2554 (N_2554,In_1115,In_570);
nor U2555 (N_2555,In_1052,In_673);
or U2556 (N_2556,In_260,In_1991);
nand U2557 (N_2557,In_1723,In_367);
or U2558 (N_2558,In_1797,In_168);
nand U2559 (N_2559,In_1608,In_1657);
nand U2560 (N_2560,In_273,In_1981);
nand U2561 (N_2561,In_779,In_409);
xnor U2562 (N_2562,In_473,In_364);
or U2563 (N_2563,In_669,In_971);
nor U2564 (N_2564,In_1055,In_150);
nand U2565 (N_2565,In_941,In_1328);
and U2566 (N_2566,In_1712,In_1724);
nand U2567 (N_2567,In_1428,In_321);
xnor U2568 (N_2568,In_1512,In_1660);
and U2569 (N_2569,In_422,In_1520);
xor U2570 (N_2570,In_405,In_276);
nor U2571 (N_2571,In_537,In_1583);
nand U2572 (N_2572,In_880,In_1775);
nand U2573 (N_2573,In_84,In_606);
nand U2574 (N_2574,In_527,In_899);
or U2575 (N_2575,In_1225,In_327);
nand U2576 (N_2576,In_378,In_544);
or U2577 (N_2577,In_637,In_1732);
or U2578 (N_2578,In_1783,In_1714);
nor U2579 (N_2579,In_1993,In_1261);
nand U2580 (N_2580,In_1070,In_611);
xnor U2581 (N_2581,In_1789,In_5);
or U2582 (N_2582,In_921,In_612);
or U2583 (N_2583,In_1982,In_210);
and U2584 (N_2584,In_743,In_810);
or U2585 (N_2585,In_702,In_1072);
nor U2586 (N_2586,In_1261,In_1743);
or U2587 (N_2587,In_1432,In_1001);
or U2588 (N_2588,In_80,In_502);
and U2589 (N_2589,In_1161,In_320);
xor U2590 (N_2590,In_1155,In_1055);
or U2591 (N_2591,In_103,In_1049);
and U2592 (N_2592,In_932,In_410);
nor U2593 (N_2593,In_987,In_75);
nor U2594 (N_2594,In_881,In_236);
nand U2595 (N_2595,In_1615,In_1859);
nand U2596 (N_2596,In_216,In_245);
nand U2597 (N_2597,In_294,In_965);
nand U2598 (N_2598,In_1578,In_1278);
and U2599 (N_2599,In_924,In_1559);
or U2600 (N_2600,In_932,In_312);
nor U2601 (N_2601,In_740,In_1739);
or U2602 (N_2602,In_1185,In_285);
and U2603 (N_2603,In_1381,In_750);
xor U2604 (N_2604,In_1196,In_1152);
nand U2605 (N_2605,In_537,In_1128);
nand U2606 (N_2606,In_1603,In_558);
or U2607 (N_2607,In_291,In_462);
and U2608 (N_2608,In_414,In_25);
and U2609 (N_2609,In_1811,In_287);
and U2610 (N_2610,In_1577,In_1447);
or U2611 (N_2611,In_811,In_582);
and U2612 (N_2612,In_1827,In_1449);
xnor U2613 (N_2613,In_1910,In_1270);
or U2614 (N_2614,In_1387,In_232);
and U2615 (N_2615,In_277,In_1284);
nor U2616 (N_2616,In_197,In_1228);
nor U2617 (N_2617,In_1108,In_1734);
and U2618 (N_2618,In_1398,In_1005);
or U2619 (N_2619,In_1847,In_1804);
nor U2620 (N_2620,In_1355,In_938);
nor U2621 (N_2621,In_1858,In_145);
xnor U2622 (N_2622,In_1138,In_235);
and U2623 (N_2623,In_1318,In_913);
nor U2624 (N_2624,In_625,In_714);
and U2625 (N_2625,In_568,In_891);
and U2626 (N_2626,In_1273,In_340);
nand U2627 (N_2627,In_1530,In_288);
or U2628 (N_2628,In_1960,In_276);
and U2629 (N_2629,In_697,In_686);
nand U2630 (N_2630,In_920,In_1041);
or U2631 (N_2631,In_1018,In_833);
nand U2632 (N_2632,In_1198,In_286);
nor U2633 (N_2633,In_1372,In_601);
or U2634 (N_2634,In_1730,In_1858);
nand U2635 (N_2635,In_1731,In_590);
xor U2636 (N_2636,In_60,In_1141);
or U2637 (N_2637,In_500,In_824);
nor U2638 (N_2638,In_1256,In_189);
nor U2639 (N_2639,In_893,In_1378);
nand U2640 (N_2640,In_1038,In_904);
and U2641 (N_2641,In_723,In_1899);
or U2642 (N_2642,In_781,In_1397);
nand U2643 (N_2643,In_908,In_255);
nor U2644 (N_2644,In_1865,In_1898);
nor U2645 (N_2645,In_1379,In_1740);
and U2646 (N_2646,In_277,In_182);
nor U2647 (N_2647,In_824,In_395);
and U2648 (N_2648,In_1441,In_1105);
xnor U2649 (N_2649,In_694,In_771);
nor U2650 (N_2650,In_1104,In_886);
nand U2651 (N_2651,In_1291,In_1217);
nor U2652 (N_2652,In_514,In_596);
nor U2653 (N_2653,In_1906,In_61);
and U2654 (N_2654,In_1780,In_1624);
nand U2655 (N_2655,In_1768,In_639);
or U2656 (N_2656,In_649,In_780);
nand U2657 (N_2657,In_1502,In_684);
nand U2658 (N_2658,In_1667,In_107);
and U2659 (N_2659,In_45,In_1165);
nor U2660 (N_2660,In_234,In_11);
nand U2661 (N_2661,In_1619,In_249);
or U2662 (N_2662,In_915,In_789);
nand U2663 (N_2663,In_1394,In_809);
or U2664 (N_2664,In_961,In_613);
or U2665 (N_2665,In_784,In_1710);
and U2666 (N_2666,In_303,In_1882);
or U2667 (N_2667,In_478,In_1104);
or U2668 (N_2668,In_1914,In_735);
nor U2669 (N_2669,In_1375,In_846);
and U2670 (N_2670,In_941,In_731);
and U2671 (N_2671,In_1921,In_49);
nor U2672 (N_2672,In_219,In_1008);
and U2673 (N_2673,In_1809,In_1845);
or U2674 (N_2674,In_339,In_1198);
nand U2675 (N_2675,In_1987,In_646);
and U2676 (N_2676,In_1007,In_1647);
nand U2677 (N_2677,In_1031,In_384);
or U2678 (N_2678,In_493,In_891);
xnor U2679 (N_2679,In_694,In_608);
xnor U2680 (N_2680,In_1152,In_644);
nand U2681 (N_2681,In_492,In_1740);
xnor U2682 (N_2682,In_687,In_1327);
nand U2683 (N_2683,In_459,In_901);
or U2684 (N_2684,In_364,In_765);
xor U2685 (N_2685,In_1422,In_1888);
nor U2686 (N_2686,In_1791,In_1089);
and U2687 (N_2687,In_839,In_161);
nand U2688 (N_2688,In_1789,In_609);
or U2689 (N_2689,In_1162,In_311);
nand U2690 (N_2690,In_306,In_1291);
or U2691 (N_2691,In_892,In_1376);
xnor U2692 (N_2692,In_1008,In_1252);
nand U2693 (N_2693,In_529,In_1373);
and U2694 (N_2694,In_1618,In_0);
or U2695 (N_2695,In_561,In_1670);
xnor U2696 (N_2696,In_1158,In_1540);
and U2697 (N_2697,In_161,In_920);
xnor U2698 (N_2698,In_783,In_1609);
nand U2699 (N_2699,In_507,In_1693);
nor U2700 (N_2700,In_1429,In_364);
nor U2701 (N_2701,In_1576,In_1110);
nor U2702 (N_2702,In_1328,In_127);
nor U2703 (N_2703,In_1605,In_1292);
or U2704 (N_2704,In_978,In_569);
or U2705 (N_2705,In_497,In_1158);
or U2706 (N_2706,In_1333,In_115);
or U2707 (N_2707,In_414,In_1898);
nor U2708 (N_2708,In_1801,In_590);
nor U2709 (N_2709,In_488,In_271);
or U2710 (N_2710,In_207,In_1957);
nand U2711 (N_2711,In_1162,In_1827);
nand U2712 (N_2712,In_1096,In_1669);
and U2713 (N_2713,In_991,In_1182);
and U2714 (N_2714,In_1716,In_485);
nor U2715 (N_2715,In_789,In_770);
or U2716 (N_2716,In_143,In_878);
and U2717 (N_2717,In_1748,In_865);
nor U2718 (N_2718,In_1744,In_543);
and U2719 (N_2719,In_743,In_681);
and U2720 (N_2720,In_1721,In_1316);
and U2721 (N_2721,In_846,In_1041);
nand U2722 (N_2722,In_1657,In_1761);
nand U2723 (N_2723,In_1915,In_1905);
nand U2724 (N_2724,In_1122,In_964);
or U2725 (N_2725,In_1733,In_695);
and U2726 (N_2726,In_118,In_952);
and U2727 (N_2727,In_1273,In_1219);
nand U2728 (N_2728,In_1449,In_1454);
nand U2729 (N_2729,In_1816,In_884);
nand U2730 (N_2730,In_1305,In_840);
or U2731 (N_2731,In_902,In_1206);
nand U2732 (N_2732,In_939,In_1468);
or U2733 (N_2733,In_1196,In_1995);
nor U2734 (N_2734,In_384,In_1945);
nor U2735 (N_2735,In_1373,In_953);
xnor U2736 (N_2736,In_1695,In_1539);
or U2737 (N_2737,In_303,In_531);
xor U2738 (N_2738,In_1601,In_1316);
xor U2739 (N_2739,In_758,In_328);
or U2740 (N_2740,In_1161,In_1511);
nor U2741 (N_2741,In_1395,In_1923);
nor U2742 (N_2742,In_1506,In_210);
and U2743 (N_2743,In_265,In_1790);
and U2744 (N_2744,In_1487,In_591);
or U2745 (N_2745,In_1887,In_1074);
nand U2746 (N_2746,In_1973,In_1393);
or U2747 (N_2747,In_1105,In_1559);
and U2748 (N_2748,In_61,In_199);
and U2749 (N_2749,In_740,In_502);
nor U2750 (N_2750,In_776,In_1009);
and U2751 (N_2751,In_808,In_717);
nor U2752 (N_2752,In_870,In_465);
and U2753 (N_2753,In_1197,In_501);
nor U2754 (N_2754,In_15,In_1471);
nor U2755 (N_2755,In_1661,In_1214);
nand U2756 (N_2756,In_679,In_1900);
or U2757 (N_2757,In_1130,In_364);
or U2758 (N_2758,In_422,In_387);
nand U2759 (N_2759,In_1312,In_1664);
and U2760 (N_2760,In_682,In_259);
or U2761 (N_2761,In_167,In_49);
and U2762 (N_2762,In_1637,In_436);
and U2763 (N_2763,In_1961,In_1899);
nand U2764 (N_2764,In_241,In_493);
or U2765 (N_2765,In_1454,In_106);
or U2766 (N_2766,In_580,In_467);
nor U2767 (N_2767,In_493,In_905);
or U2768 (N_2768,In_874,In_1079);
xor U2769 (N_2769,In_404,In_1293);
or U2770 (N_2770,In_92,In_847);
or U2771 (N_2771,In_1798,In_1385);
nand U2772 (N_2772,In_719,In_1871);
xnor U2773 (N_2773,In_375,In_78);
and U2774 (N_2774,In_1452,In_1166);
and U2775 (N_2775,In_986,In_1727);
nor U2776 (N_2776,In_1602,In_270);
or U2777 (N_2777,In_1683,In_440);
or U2778 (N_2778,In_1233,In_1367);
and U2779 (N_2779,In_969,In_1910);
xor U2780 (N_2780,In_1876,In_1446);
nand U2781 (N_2781,In_592,In_59);
nand U2782 (N_2782,In_899,In_1536);
nand U2783 (N_2783,In_922,In_334);
or U2784 (N_2784,In_828,In_1531);
nor U2785 (N_2785,In_1702,In_788);
nand U2786 (N_2786,In_1102,In_117);
nor U2787 (N_2787,In_1018,In_463);
nor U2788 (N_2788,In_1481,In_158);
and U2789 (N_2789,In_688,In_1388);
xnor U2790 (N_2790,In_775,In_467);
and U2791 (N_2791,In_321,In_231);
xor U2792 (N_2792,In_217,In_1134);
nand U2793 (N_2793,In_413,In_839);
xor U2794 (N_2794,In_195,In_1236);
nand U2795 (N_2795,In_1868,In_1646);
and U2796 (N_2796,In_558,In_832);
nand U2797 (N_2797,In_1197,In_1751);
nand U2798 (N_2798,In_1803,In_1199);
nor U2799 (N_2799,In_1722,In_242);
nor U2800 (N_2800,In_1631,In_631);
or U2801 (N_2801,In_1852,In_1899);
and U2802 (N_2802,In_179,In_1711);
nand U2803 (N_2803,In_725,In_648);
nor U2804 (N_2804,In_1733,In_1970);
nand U2805 (N_2805,In_900,In_750);
or U2806 (N_2806,In_1170,In_1581);
and U2807 (N_2807,In_407,In_349);
nor U2808 (N_2808,In_255,In_232);
nand U2809 (N_2809,In_1739,In_572);
xnor U2810 (N_2810,In_828,In_46);
or U2811 (N_2811,In_286,In_1040);
nor U2812 (N_2812,In_1258,In_858);
and U2813 (N_2813,In_313,In_987);
or U2814 (N_2814,In_548,In_1848);
nor U2815 (N_2815,In_651,In_1011);
or U2816 (N_2816,In_1128,In_1065);
or U2817 (N_2817,In_973,In_589);
nor U2818 (N_2818,In_831,In_743);
and U2819 (N_2819,In_1473,In_1424);
and U2820 (N_2820,In_1368,In_1473);
or U2821 (N_2821,In_539,In_915);
nor U2822 (N_2822,In_1740,In_1972);
nor U2823 (N_2823,In_1536,In_450);
nand U2824 (N_2824,In_20,In_441);
or U2825 (N_2825,In_1651,In_425);
nor U2826 (N_2826,In_1086,In_1508);
or U2827 (N_2827,In_63,In_1163);
or U2828 (N_2828,In_1989,In_236);
nand U2829 (N_2829,In_507,In_1400);
nor U2830 (N_2830,In_1212,In_811);
nor U2831 (N_2831,In_610,In_1440);
nor U2832 (N_2832,In_944,In_148);
xor U2833 (N_2833,In_1422,In_1401);
and U2834 (N_2834,In_455,In_1760);
nand U2835 (N_2835,In_35,In_1009);
nor U2836 (N_2836,In_272,In_108);
nand U2837 (N_2837,In_1652,In_947);
and U2838 (N_2838,In_119,In_968);
nor U2839 (N_2839,In_913,In_639);
nor U2840 (N_2840,In_430,In_853);
xnor U2841 (N_2841,In_1552,In_115);
nor U2842 (N_2842,In_234,In_732);
nand U2843 (N_2843,In_243,In_1416);
nand U2844 (N_2844,In_1085,In_63);
nor U2845 (N_2845,In_618,In_523);
or U2846 (N_2846,In_1916,In_1788);
nand U2847 (N_2847,In_1730,In_93);
xnor U2848 (N_2848,In_166,In_676);
nor U2849 (N_2849,In_1429,In_1470);
or U2850 (N_2850,In_1913,In_1893);
and U2851 (N_2851,In_1842,In_271);
nor U2852 (N_2852,In_1342,In_981);
xor U2853 (N_2853,In_618,In_520);
xnor U2854 (N_2854,In_1742,In_671);
and U2855 (N_2855,In_545,In_1659);
nor U2856 (N_2856,In_287,In_1055);
or U2857 (N_2857,In_730,In_1373);
nand U2858 (N_2858,In_1883,In_1980);
nor U2859 (N_2859,In_509,In_559);
or U2860 (N_2860,In_1733,In_394);
nor U2861 (N_2861,In_1752,In_1186);
xnor U2862 (N_2862,In_1920,In_964);
and U2863 (N_2863,In_398,In_1037);
nand U2864 (N_2864,In_1470,In_631);
nor U2865 (N_2865,In_141,In_1913);
nand U2866 (N_2866,In_1727,In_568);
and U2867 (N_2867,In_1370,In_658);
and U2868 (N_2868,In_217,In_726);
and U2869 (N_2869,In_743,In_481);
and U2870 (N_2870,In_1078,In_341);
nor U2871 (N_2871,In_1298,In_515);
nor U2872 (N_2872,In_730,In_1173);
nor U2873 (N_2873,In_1112,In_742);
nor U2874 (N_2874,In_1174,In_1948);
nor U2875 (N_2875,In_679,In_1269);
nor U2876 (N_2876,In_31,In_497);
nor U2877 (N_2877,In_1433,In_508);
or U2878 (N_2878,In_475,In_818);
nand U2879 (N_2879,In_559,In_1912);
or U2880 (N_2880,In_1408,In_1224);
or U2881 (N_2881,In_126,In_1866);
xnor U2882 (N_2882,In_1571,In_275);
nand U2883 (N_2883,In_1959,In_1113);
nand U2884 (N_2884,In_926,In_1013);
nand U2885 (N_2885,In_1306,In_1731);
or U2886 (N_2886,In_587,In_976);
nand U2887 (N_2887,In_866,In_280);
and U2888 (N_2888,In_1115,In_1279);
xor U2889 (N_2889,In_168,In_1334);
and U2890 (N_2890,In_870,In_1670);
and U2891 (N_2891,In_1630,In_661);
or U2892 (N_2892,In_528,In_312);
nor U2893 (N_2893,In_773,In_819);
and U2894 (N_2894,In_555,In_1422);
and U2895 (N_2895,In_302,In_936);
or U2896 (N_2896,In_78,In_250);
nor U2897 (N_2897,In_1215,In_536);
nand U2898 (N_2898,In_565,In_807);
nand U2899 (N_2899,In_985,In_1073);
and U2900 (N_2900,In_592,In_471);
nor U2901 (N_2901,In_1397,In_40);
nand U2902 (N_2902,In_1320,In_1215);
and U2903 (N_2903,In_1274,In_819);
and U2904 (N_2904,In_1696,In_509);
nand U2905 (N_2905,In_1062,In_563);
nand U2906 (N_2906,In_1956,In_813);
nor U2907 (N_2907,In_595,In_77);
nor U2908 (N_2908,In_216,In_1234);
and U2909 (N_2909,In_1801,In_420);
nor U2910 (N_2910,In_245,In_447);
nand U2911 (N_2911,In_130,In_1490);
xor U2912 (N_2912,In_1822,In_927);
or U2913 (N_2913,In_666,In_501);
or U2914 (N_2914,In_1320,In_981);
xor U2915 (N_2915,In_1151,In_1676);
or U2916 (N_2916,In_513,In_1165);
nor U2917 (N_2917,In_839,In_1147);
or U2918 (N_2918,In_1493,In_1500);
nand U2919 (N_2919,In_333,In_1067);
nor U2920 (N_2920,In_206,In_635);
nand U2921 (N_2921,In_718,In_112);
xnor U2922 (N_2922,In_1058,In_474);
and U2923 (N_2923,In_429,In_1297);
nand U2924 (N_2924,In_682,In_669);
nor U2925 (N_2925,In_385,In_1652);
nand U2926 (N_2926,In_1459,In_1465);
nor U2927 (N_2927,In_1490,In_655);
or U2928 (N_2928,In_38,In_1813);
xor U2929 (N_2929,In_529,In_1900);
and U2930 (N_2930,In_1608,In_305);
nor U2931 (N_2931,In_1373,In_339);
xor U2932 (N_2932,In_1624,In_1706);
xor U2933 (N_2933,In_615,In_797);
or U2934 (N_2934,In_23,In_192);
xnor U2935 (N_2935,In_616,In_1644);
nand U2936 (N_2936,In_59,In_612);
nor U2937 (N_2937,In_272,In_1268);
or U2938 (N_2938,In_1220,In_873);
or U2939 (N_2939,In_861,In_1185);
or U2940 (N_2940,In_319,In_1058);
nor U2941 (N_2941,In_173,In_1849);
and U2942 (N_2942,In_754,In_1726);
or U2943 (N_2943,In_340,In_1003);
nor U2944 (N_2944,In_1427,In_858);
and U2945 (N_2945,In_663,In_1936);
xor U2946 (N_2946,In_839,In_1033);
or U2947 (N_2947,In_1191,In_1358);
and U2948 (N_2948,In_1410,In_1127);
nand U2949 (N_2949,In_559,In_1684);
nand U2950 (N_2950,In_233,In_35);
nand U2951 (N_2951,In_225,In_1141);
nor U2952 (N_2952,In_445,In_1596);
or U2953 (N_2953,In_939,In_836);
nor U2954 (N_2954,In_1891,In_1622);
nand U2955 (N_2955,In_1426,In_1243);
nor U2956 (N_2956,In_747,In_141);
or U2957 (N_2957,In_991,In_1460);
and U2958 (N_2958,In_1321,In_1451);
or U2959 (N_2959,In_1083,In_232);
or U2960 (N_2960,In_1861,In_727);
nand U2961 (N_2961,In_1061,In_1764);
nor U2962 (N_2962,In_297,In_17);
nand U2963 (N_2963,In_286,In_1279);
xnor U2964 (N_2964,In_244,In_1832);
nor U2965 (N_2965,In_59,In_1270);
or U2966 (N_2966,In_1902,In_1077);
or U2967 (N_2967,In_468,In_1738);
or U2968 (N_2968,In_284,In_962);
nand U2969 (N_2969,In_1027,In_303);
and U2970 (N_2970,In_1956,In_1688);
and U2971 (N_2971,In_1414,In_534);
nor U2972 (N_2972,In_501,In_1697);
or U2973 (N_2973,In_1178,In_1297);
and U2974 (N_2974,In_1166,In_966);
nand U2975 (N_2975,In_168,In_1129);
nand U2976 (N_2976,In_525,In_35);
or U2977 (N_2977,In_277,In_764);
and U2978 (N_2978,In_1388,In_1407);
and U2979 (N_2979,In_1725,In_833);
or U2980 (N_2980,In_174,In_428);
and U2981 (N_2981,In_1124,In_1459);
or U2982 (N_2982,In_997,In_1431);
and U2983 (N_2983,In_468,In_774);
and U2984 (N_2984,In_1589,In_24);
xnor U2985 (N_2985,In_432,In_1802);
nor U2986 (N_2986,In_1481,In_872);
nand U2987 (N_2987,In_1466,In_352);
nand U2988 (N_2988,In_1874,In_1568);
nor U2989 (N_2989,In_649,In_1431);
xor U2990 (N_2990,In_65,In_677);
xor U2991 (N_2991,In_122,In_331);
or U2992 (N_2992,In_1500,In_1498);
nor U2993 (N_2993,In_1306,In_1929);
nor U2994 (N_2994,In_1194,In_1427);
or U2995 (N_2995,In_798,In_1748);
nor U2996 (N_2996,In_1935,In_123);
nand U2997 (N_2997,In_752,In_938);
and U2998 (N_2998,In_1252,In_473);
nor U2999 (N_2999,In_1837,In_1355);
or U3000 (N_3000,In_1720,In_667);
xor U3001 (N_3001,In_97,In_1495);
nor U3002 (N_3002,In_441,In_922);
nand U3003 (N_3003,In_1131,In_1154);
nand U3004 (N_3004,In_1278,In_1974);
and U3005 (N_3005,In_1460,In_211);
nand U3006 (N_3006,In_1368,In_763);
nor U3007 (N_3007,In_761,In_404);
and U3008 (N_3008,In_522,In_969);
nand U3009 (N_3009,In_1700,In_88);
nand U3010 (N_3010,In_422,In_9);
nor U3011 (N_3011,In_1722,In_234);
nor U3012 (N_3012,In_938,In_578);
nand U3013 (N_3013,In_494,In_1561);
nor U3014 (N_3014,In_961,In_976);
nor U3015 (N_3015,In_1727,In_1236);
nand U3016 (N_3016,In_1423,In_542);
and U3017 (N_3017,In_273,In_431);
and U3018 (N_3018,In_242,In_1529);
nand U3019 (N_3019,In_1355,In_1895);
nand U3020 (N_3020,In_1056,In_1407);
or U3021 (N_3021,In_924,In_1617);
xor U3022 (N_3022,In_789,In_461);
nand U3023 (N_3023,In_1298,In_325);
and U3024 (N_3024,In_369,In_732);
nand U3025 (N_3025,In_1220,In_1936);
nand U3026 (N_3026,In_1189,In_1732);
or U3027 (N_3027,In_224,In_1900);
and U3028 (N_3028,In_1401,In_323);
nand U3029 (N_3029,In_1737,In_1450);
nor U3030 (N_3030,In_556,In_659);
nand U3031 (N_3031,In_1819,In_1773);
nor U3032 (N_3032,In_1262,In_509);
and U3033 (N_3033,In_139,In_1187);
nor U3034 (N_3034,In_1285,In_766);
nor U3035 (N_3035,In_635,In_1680);
and U3036 (N_3036,In_889,In_471);
xor U3037 (N_3037,In_1417,In_1982);
xor U3038 (N_3038,In_557,In_1082);
nor U3039 (N_3039,In_210,In_895);
and U3040 (N_3040,In_796,In_1574);
nor U3041 (N_3041,In_1622,In_1358);
xnor U3042 (N_3042,In_49,In_1263);
nand U3043 (N_3043,In_1529,In_1624);
nand U3044 (N_3044,In_781,In_1223);
or U3045 (N_3045,In_872,In_71);
nand U3046 (N_3046,In_1943,In_241);
nor U3047 (N_3047,In_1727,In_1938);
xnor U3048 (N_3048,In_279,In_547);
and U3049 (N_3049,In_1526,In_1573);
or U3050 (N_3050,In_1102,In_1207);
xor U3051 (N_3051,In_468,In_1702);
nand U3052 (N_3052,In_1527,In_1454);
or U3053 (N_3053,In_1684,In_1223);
nor U3054 (N_3054,In_392,In_1134);
nand U3055 (N_3055,In_287,In_395);
nor U3056 (N_3056,In_372,In_1215);
or U3057 (N_3057,In_1553,In_1919);
nor U3058 (N_3058,In_1015,In_1842);
nor U3059 (N_3059,In_291,In_469);
xor U3060 (N_3060,In_347,In_1741);
nor U3061 (N_3061,In_1250,In_158);
nor U3062 (N_3062,In_917,In_521);
and U3063 (N_3063,In_474,In_92);
nand U3064 (N_3064,In_1371,In_1210);
or U3065 (N_3065,In_1698,In_1273);
nor U3066 (N_3066,In_901,In_1301);
or U3067 (N_3067,In_294,In_1989);
xnor U3068 (N_3068,In_1266,In_3);
or U3069 (N_3069,In_625,In_1430);
nand U3070 (N_3070,In_909,In_975);
or U3071 (N_3071,In_1920,In_1604);
and U3072 (N_3072,In_460,In_1732);
nand U3073 (N_3073,In_1949,In_1499);
and U3074 (N_3074,In_140,In_1553);
and U3075 (N_3075,In_1821,In_1054);
nand U3076 (N_3076,In_1250,In_753);
or U3077 (N_3077,In_1195,In_748);
and U3078 (N_3078,In_1112,In_1932);
nand U3079 (N_3079,In_662,In_1432);
and U3080 (N_3080,In_1336,In_1807);
nand U3081 (N_3081,In_1264,In_1423);
xnor U3082 (N_3082,In_651,In_937);
and U3083 (N_3083,In_1076,In_1962);
and U3084 (N_3084,In_1196,In_923);
nor U3085 (N_3085,In_452,In_1996);
or U3086 (N_3086,In_451,In_124);
and U3087 (N_3087,In_931,In_207);
nand U3088 (N_3088,In_1891,In_163);
or U3089 (N_3089,In_1870,In_1849);
nand U3090 (N_3090,In_440,In_70);
nor U3091 (N_3091,In_137,In_1964);
and U3092 (N_3092,In_1169,In_1266);
nand U3093 (N_3093,In_491,In_1898);
nor U3094 (N_3094,In_598,In_1557);
nor U3095 (N_3095,In_93,In_1265);
and U3096 (N_3096,In_1663,In_978);
nand U3097 (N_3097,In_1256,In_689);
nor U3098 (N_3098,In_1457,In_399);
or U3099 (N_3099,In_1640,In_741);
or U3100 (N_3100,In_691,In_787);
or U3101 (N_3101,In_1344,In_1508);
and U3102 (N_3102,In_289,In_1638);
or U3103 (N_3103,In_1181,In_323);
nor U3104 (N_3104,In_1773,In_3);
xnor U3105 (N_3105,In_672,In_1226);
and U3106 (N_3106,In_253,In_1301);
xnor U3107 (N_3107,In_648,In_1418);
and U3108 (N_3108,In_720,In_487);
xnor U3109 (N_3109,In_31,In_1694);
and U3110 (N_3110,In_960,In_900);
or U3111 (N_3111,In_1919,In_755);
and U3112 (N_3112,In_1618,In_372);
or U3113 (N_3113,In_1059,In_626);
or U3114 (N_3114,In_366,In_702);
nand U3115 (N_3115,In_372,In_1979);
nand U3116 (N_3116,In_56,In_1226);
xnor U3117 (N_3117,In_1842,In_153);
and U3118 (N_3118,In_1498,In_402);
nor U3119 (N_3119,In_743,In_853);
or U3120 (N_3120,In_662,In_235);
or U3121 (N_3121,In_1867,In_548);
or U3122 (N_3122,In_128,In_1452);
nor U3123 (N_3123,In_1328,In_1519);
or U3124 (N_3124,In_1222,In_1261);
xor U3125 (N_3125,In_266,In_913);
nand U3126 (N_3126,In_160,In_170);
and U3127 (N_3127,In_138,In_670);
nor U3128 (N_3128,In_1857,In_1009);
nand U3129 (N_3129,In_38,In_752);
nand U3130 (N_3130,In_686,In_679);
and U3131 (N_3131,In_1505,In_1456);
nor U3132 (N_3132,In_1490,In_1589);
and U3133 (N_3133,In_1344,In_1610);
nand U3134 (N_3134,In_1997,In_747);
nor U3135 (N_3135,In_1324,In_675);
nor U3136 (N_3136,In_1681,In_391);
and U3137 (N_3137,In_107,In_1979);
and U3138 (N_3138,In_1940,In_162);
nor U3139 (N_3139,In_1334,In_1072);
xnor U3140 (N_3140,In_262,In_1360);
and U3141 (N_3141,In_153,In_1024);
nand U3142 (N_3142,In_1681,In_647);
nand U3143 (N_3143,In_1560,In_700);
nor U3144 (N_3144,In_1044,In_1419);
or U3145 (N_3145,In_378,In_172);
and U3146 (N_3146,In_1599,In_68);
nand U3147 (N_3147,In_1684,In_1971);
and U3148 (N_3148,In_712,In_1122);
nand U3149 (N_3149,In_603,In_1490);
or U3150 (N_3150,In_1615,In_1371);
nor U3151 (N_3151,In_12,In_453);
nor U3152 (N_3152,In_1014,In_1567);
nor U3153 (N_3153,In_1213,In_1285);
and U3154 (N_3154,In_1066,In_1929);
nor U3155 (N_3155,In_1206,In_1194);
and U3156 (N_3156,In_1512,In_1990);
or U3157 (N_3157,In_289,In_552);
nor U3158 (N_3158,In_1635,In_1597);
and U3159 (N_3159,In_237,In_1751);
nor U3160 (N_3160,In_1714,In_64);
and U3161 (N_3161,In_320,In_998);
or U3162 (N_3162,In_131,In_1403);
or U3163 (N_3163,In_1823,In_499);
nand U3164 (N_3164,In_1049,In_1480);
nand U3165 (N_3165,In_1192,In_683);
nor U3166 (N_3166,In_1961,In_1419);
nand U3167 (N_3167,In_1018,In_31);
and U3168 (N_3168,In_1209,In_669);
xnor U3169 (N_3169,In_1640,In_995);
nor U3170 (N_3170,In_616,In_1062);
xnor U3171 (N_3171,In_32,In_859);
nand U3172 (N_3172,In_323,In_575);
and U3173 (N_3173,In_1728,In_1739);
and U3174 (N_3174,In_966,In_429);
nor U3175 (N_3175,In_615,In_1705);
and U3176 (N_3176,In_1159,In_908);
nand U3177 (N_3177,In_273,In_303);
nor U3178 (N_3178,In_1595,In_761);
nand U3179 (N_3179,In_1791,In_394);
nand U3180 (N_3180,In_18,In_724);
nor U3181 (N_3181,In_1513,In_976);
and U3182 (N_3182,In_1539,In_1384);
nand U3183 (N_3183,In_781,In_1053);
or U3184 (N_3184,In_183,In_1010);
nand U3185 (N_3185,In_967,In_1011);
nor U3186 (N_3186,In_1611,In_459);
or U3187 (N_3187,In_1842,In_1877);
and U3188 (N_3188,In_88,In_1643);
or U3189 (N_3189,In_31,In_1833);
or U3190 (N_3190,In_1753,In_425);
nand U3191 (N_3191,In_727,In_973);
and U3192 (N_3192,In_955,In_1714);
xor U3193 (N_3193,In_834,In_1581);
nor U3194 (N_3194,In_820,In_1216);
nand U3195 (N_3195,In_182,In_1910);
or U3196 (N_3196,In_1981,In_71);
xnor U3197 (N_3197,In_1354,In_749);
and U3198 (N_3198,In_333,In_524);
nor U3199 (N_3199,In_1337,In_1040);
nand U3200 (N_3200,In_491,In_1460);
or U3201 (N_3201,In_1773,In_1982);
nand U3202 (N_3202,In_537,In_425);
nor U3203 (N_3203,In_1573,In_416);
nand U3204 (N_3204,In_964,In_1445);
and U3205 (N_3205,In_122,In_925);
or U3206 (N_3206,In_155,In_1887);
and U3207 (N_3207,In_1824,In_714);
nand U3208 (N_3208,In_1112,In_147);
nand U3209 (N_3209,In_1471,In_1878);
nor U3210 (N_3210,In_1360,In_1651);
nand U3211 (N_3211,In_1245,In_978);
and U3212 (N_3212,In_291,In_1083);
and U3213 (N_3213,In_1871,In_1263);
and U3214 (N_3214,In_537,In_12);
and U3215 (N_3215,In_486,In_1044);
or U3216 (N_3216,In_899,In_587);
and U3217 (N_3217,In_646,In_1261);
or U3218 (N_3218,In_134,In_1156);
or U3219 (N_3219,In_1928,In_326);
xor U3220 (N_3220,In_1096,In_1606);
nand U3221 (N_3221,In_1009,In_523);
and U3222 (N_3222,In_142,In_988);
nand U3223 (N_3223,In_823,In_93);
xor U3224 (N_3224,In_1322,In_1110);
or U3225 (N_3225,In_1383,In_122);
nor U3226 (N_3226,In_487,In_473);
nor U3227 (N_3227,In_114,In_1398);
nor U3228 (N_3228,In_1876,In_718);
and U3229 (N_3229,In_98,In_1939);
or U3230 (N_3230,In_1784,In_1742);
nor U3231 (N_3231,In_1075,In_318);
nand U3232 (N_3232,In_1957,In_428);
and U3233 (N_3233,In_1673,In_1234);
nor U3234 (N_3234,In_920,In_397);
and U3235 (N_3235,In_974,In_478);
and U3236 (N_3236,In_961,In_1580);
or U3237 (N_3237,In_1883,In_492);
or U3238 (N_3238,In_1913,In_469);
or U3239 (N_3239,In_506,In_1752);
nor U3240 (N_3240,In_1122,In_118);
nor U3241 (N_3241,In_1424,In_622);
and U3242 (N_3242,In_234,In_1200);
and U3243 (N_3243,In_990,In_1936);
or U3244 (N_3244,In_1844,In_1920);
and U3245 (N_3245,In_1102,In_682);
nand U3246 (N_3246,In_33,In_1163);
nand U3247 (N_3247,In_1395,In_376);
or U3248 (N_3248,In_218,In_225);
nand U3249 (N_3249,In_1905,In_1150);
nor U3250 (N_3250,In_87,In_1190);
xnor U3251 (N_3251,In_1749,In_1520);
or U3252 (N_3252,In_526,In_1302);
xor U3253 (N_3253,In_241,In_451);
or U3254 (N_3254,In_1778,In_873);
and U3255 (N_3255,In_1072,In_1885);
or U3256 (N_3256,In_1935,In_19);
nand U3257 (N_3257,In_1162,In_1833);
xnor U3258 (N_3258,In_1753,In_1928);
and U3259 (N_3259,In_483,In_982);
nand U3260 (N_3260,In_971,In_1649);
nor U3261 (N_3261,In_818,In_642);
and U3262 (N_3262,In_256,In_522);
and U3263 (N_3263,In_224,In_1947);
xor U3264 (N_3264,In_879,In_605);
nand U3265 (N_3265,In_614,In_779);
or U3266 (N_3266,In_1807,In_181);
or U3267 (N_3267,In_382,In_8);
nand U3268 (N_3268,In_943,In_324);
xnor U3269 (N_3269,In_402,In_415);
and U3270 (N_3270,In_1134,In_716);
nor U3271 (N_3271,In_919,In_460);
or U3272 (N_3272,In_1505,In_489);
nor U3273 (N_3273,In_1563,In_179);
and U3274 (N_3274,In_1735,In_401);
and U3275 (N_3275,In_932,In_570);
xor U3276 (N_3276,In_1462,In_1832);
and U3277 (N_3277,In_1936,In_455);
and U3278 (N_3278,In_234,In_292);
and U3279 (N_3279,In_1053,In_120);
and U3280 (N_3280,In_1192,In_1489);
and U3281 (N_3281,In_1514,In_1489);
xor U3282 (N_3282,In_127,In_1670);
nor U3283 (N_3283,In_181,In_1463);
nand U3284 (N_3284,In_754,In_1809);
nand U3285 (N_3285,In_577,In_42);
and U3286 (N_3286,In_1578,In_76);
and U3287 (N_3287,In_540,In_1659);
or U3288 (N_3288,In_252,In_1847);
and U3289 (N_3289,In_1850,In_1466);
and U3290 (N_3290,In_1127,In_155);
nand U3291 (N_3291,In_103,In_264);
and U3292 (N_3292,In_1891,In_1341);
nor U3293 (N_3293,In_752,In_1962);
nand U3294 (N_3294,In_375,In_346);
nand U3295 (N_3295,In_1176,In_108);
and U3296 (N_3296,In_589,In_167);
xnor U3297 (N_3297,In_998,In_742);
and U3298 (N_3298,In_1972,In_651);
or U3299 (N_3299,In_1865,In_1974);
and U3300 (N_3300,In_1587,In_242);
or U3301 (N_3301,In_342,In_437);
nor U3302 (N_3302,In_1823,In_606);
xnor U3303 (N_3303,In_822,In_830);
and U3304 (N_3304,In_1138,In_1337);
nor U3305 (N_3305,In_1416,In_1372);
and U3306 (N_3306,In_322,In_1801);
nand U3307 (N_3307,In_1396,In_1443);
nor U3308 (N_3308,In_1477,In_1760);
or U3309 (N_3309,In_1649,In_1825);
or U3310 (N_3310,In_1318,In_1451);
or U3311 (N_3311,In_342,In_1374);
or U3312 (N_3312,In_830,In_1700);
nor U3313 (N_3313,In_371,In_713);
and U3314 (N_3314,In_1398,In_568);
and U3315 (N_3315,In_637,In_85);
nor U3316 (N_3316,In_218,In_811);
nor U3317 (N_3317,In_349,In_1511);
or U3318 (N_3318,In_23,In_1402);
nor U3319 (N_3319,In_914,In_1635);
and U3320 (N_3320,In_1860,In_1876);
nand U3321 (N_3321,In_104,In_615);
xnor U3322 (N_3322,In_1306,In_876);
nand U3323 (N_3323,In_955,In_252);
nor U3324 (N_3324,In_499,In_1557);
nand U3325 (N_3325,In_816,In_994);
nor U3326 (N_3326,In_1059,In_1069);
nand U3327 (N_3327,In_349,In_34);
nand U3328 (N_3328,In_479,In_1875);
xor U3329 (N_3329,In_1149,In_887);
nand U3330 (N_3330,In_1872,In_915);
and U3331 (N_3331,In_1115,In_1329);
nor U3332 (N_3332,In_203,In_1900);
nor U3333 (N_3333,In_824,In_1994);
and U3334 (N_3334,In_1678,In_1504);
and U3335 (N_3335,In_122,In_975);
nand U3336 (N_3336,In_14,In_522);
or U3337 (N_3337,In_1305,In_1596);
or U3338 (N_3338,In_1079,In_587);
and U3339 (N_3339,In_1594,In_1373);
and U3340 (N_3340,In_1498,In_1174);
nor U3341 (N_3341,In_1318,In_527);
nor U3342 (N_3342,In_1885,In_250);
nand U3343 (N_3343,In_1964,In_1069);
or U3344 (N_3344,In_1556,In_1852);
nand U3345 (N_3345,In_1135,In_429);
and U3346 (N_3346,In_87,In_1038);
or U3347 (N_3347,In_1518,In_471);
nor U3348 (N_3348,In_457,In_1977);
or U3349 (N_3349,In_236,In_218);
nand U3350 (N_3350,In_242,In_1043);
and U3351 (N_3351,In_1549,In_740);
or U3352 (N_3352,In_1294,In_637);
nand U3353 (N_3353,In_918,In_359);
xor U3354 (N_3354,In_477,In_1712);
or U3355 (N_3355,In_217,In_124);
nor U3356 (N_3356,In_1685,In_51);
nor U3357 (N_3357,In_1139,In_728);
and U3358 (N_3358,In_29,In_18);
nand U3359 (N_3359,In_162,In_836);
nor U3360 (N_3360,In_1087,In_1879);
and U3361 (N_3361,In_2,In_1790);
nor U3362 (N_3362,In_1480,In_888);
and U3363 (N_3363,In_474,In_1134);
and U3364 (N_3364,In_847,In_360);
xnor U3365 (N_3365,In_840,In_1822);
nand U3366 (N_3366,In_325,In_564);
nor U3367 (N_3367,In_154,In_20);
or U3368 (N_3368,In_1990,In_742);
nand U3369 (N_3369,In_373,In_4);
or U3370 (N_3370,In_1322,In_1679);
and U3371 (N_3371,In_198,In_221);
nand U3372 (N_3372,In_1963,In_1988);
or U3373 (N_3373,In_1230,In_1287);
and U3374 (N_3374,In_1340,In_1871);
nor U3375 (N_3375,In_1171,In_505);
or U3376 (N_3376,In_1114,In_367);
or U3377 (N_3377,In_132,In_1300);
nand U3378 (N_3378,In_473,In_1343);
xnor U3379 (N_3379,In_1257,In_653);
or U3380 (N_3380,In_1010,In_1007);
and U3381 (N_3381,In_1732,In_1932);
or U3382 (N_3382,In_229,In_914);
or U3383 (N_3383,In_1972,In_755);
nor U3384 (N_3384,In_1910,In_1834);
and U3385 (N_3385,In_8,In_563);
xor U3386 (N_3386,In_1624,In_84);
xnor U3387 (N_3387,In_188,In_730);
nor U3388 (N_3388,In_1961,In_1150);
nand U3389 (N_3389,In_778,In_1449);
nor U3390 (N_3390,In_1913,In_1452);
nand U3391 (N_3391,In_1583,In_970);
and U3392 (N_3392,In_1693,In_1061);
and U3393 (N_3393,In_1299,In_91);
and U3394 (N_3394,In_706,In_1368);
and U3395 (N_3395,In_998,In_937);
nor U3396 (N_3396,In_1420,In_90);
and U3397 (N_3397,In_783,In_964);
nand U3398 (N_3398,In_598,In_1827);
or U3399 (N_3399,In_398,In_1878);
nand U3400 (N_3400,In_488,In_1042);
xor U3401 (N_3401,In_1090,In_323);
nor U3402 (N_3402,In_892,In_799);
and U3403 (N_3403,In_1162,In_1691);
or U3404 (N_3404,In_1652,In_103);
and U3405 (N_3405,In_1574,In_113);
xor U3406 (N_3406,In_648,In_795);
or U3407 (N_3407,In_1324,In_1710);
nand U3408 (N_3408,In_1772,In_969);
or U3409 (N_3409,In_761,In_888);
and U3410 (N_3410,In_749,In_1542);
nand U3411 (N_3411,In_355,In_564);
nand U3412 (N_3412,In_28,In_47);
or U3413 (N_3413,In_599,In_1461);
nor U3414 (N_3414,In_478,In_1342);
xor U3415 (N_3415,In_1837,In_323);
or U3416 (N_3416,In_1142,In_742);
and U3417 (N_3417,In_588,In_838);
or U3418 (N_3418,In_1761,In_1048);
xnor U3419 (N_3419,In_725,In_96);
nand U3420 (N_3420,In_1259,In_22);
or U3421 (N_3421,In_1211,In_450);
or U3422 (N_3422,In_1717,In_1562);
and U3423 (N_3423,In_606,In_1244);
xnor U3424 (N_3424,In_1019,In_749);
nand U3425 (N_3425,In_704,In_1973);
and U3426 (N_3426,In_1199,In_889);
or U3427 (N_3427,In_1275,In_377);
nand U3428 (N_3428,In_725,In_494);
nor U3429 (N_3429,In_147,In_1830);
xnor U3430 (N_3430,In_1207,In_338);
xor U3431 (N_3431,In_1797,In_1819);
nor U3432 (N_3432,In_17,In_655);
and U3433 (N_3433,In_1110,In_830);
nor U3434 (N_3434,In_1658,In_778);
and U3435 (N_3435,In_378,In_841);
nor U3436 (N_3436,In_1792,In_188);
and U3437 (N_3437,In_574,In_188);
nor U3438 (N_3438,In_151,In_835);
or U3439 (N_3439,In_1773,In_1542);
nor U3440 (N_3440,In_1339,In_601);
nand U3441 (N_3441,In_1623,In_1421);
nor U3442 (N_3442,In_1616,In_956);
and U3443 (N_3443,In_661,In_792);
and U3444 (N_3444,In_1237,In_1963);
nor U3445 (N_3445,In_548,In_913);
nand U3446 (N_3446,In_155,In_403);
xnor U3447 (N_3447,In_1933,In_1555);
nand U3448 (N_3448,In_407,In_404);
nand U3449 (N_3449,In_1112,In_1321);
nand U3450 (N_3450,In_655,In_1967);
nand U3451 (N_3451,In_276,In_39);
nor U3452 (N_3452,In_557,In_1721);
and U3453 (N_3453,In_1464,In_1186);
nor U3454 (N_3454,In_876,In_254);
and U3455 (N_3455,In_1238,In_1992);
and U3456 (N_3456,In_1229,In_551);
and U3457 (N_3457,In_1902,In_435);
and U3458 (N_3458,In_1711,In_1145);
nand U3459 (N_3459,In_1284,In_1319);
xnor U3460 (N_3460,In_904,In_1385);
or U3461 (N_3461,In_215,In_2);
or U3462 (N_3462,In_230,In_1673);
xnor U3463 (N_3463,In_1923,In_1132);
and U3464 (N_3464,In_103,In_1916);
nor U3465 (N_3465,In_1114,In_1229);
or U3466 (N_3466,In_1558,In_1492);
or U3467 (N_3467,In_815,In_1140);
nor U3468 (N_3468,In_807,In_68);
and U3469 (N_3469,In_263,In_226);
xnor U3470 (N_3470,In_1510,In_305);
and U3471 (N_3471,In_1093,In_433);
nor U3472 (N_3472,In_47,In_1968);
and U3473 (N_3473,In_1036,In_1650);
or U3474 (N_3474,In_1921,In_431);
nand U3475 (N_3475,In_309,In_1138);
nor U3476 (N_3476,In_591,In_1823);
or U3477 (N_3477,In_333,In_155);
nor U3478 (N_3478,In_112,In_713);
xnor U3479 (N_3479,In_234,In_833);
nor U3480 (N_3480,In_1523,In_1548);
and U3481 (N_3481,In_1860,In_46);
and U3482 (N_3482,In_1696,In_150);
xor U3483 (N_3483,In_486,In_1508);
nand U3484 (N_3484,In_1962,In_352);
nand U3485 (N_3485,In_148,In_1791);
or U3486 (N_3486,In_1225,In_1530);
nor U3487 (N_3487,In_905,In_869);
nor U3488 (N_3488,In_1045,In_843);
nand U3489 (N_3489,In_465,In_1548);
nor U3490 (N_3490,In_1769,In_214);
or U3491 (N_3491,In_916,In_1156);
nor U3492 (N_3492,In_1725,In_162);
nand U3493 (N_3493,In_636,In_1384);
nor U3494 (N_3494,In_1706,In_1009);
nand U3495 (N_3495,In_1037,In_890);
and U3496 (N_3496,In_975,In_1526);
or U3497 (N_3497,In_1226,In_1974);
and U3498 (N_3498,In_1598,In_1727);
xnor U3499 (N_3499,In_164,In_434);
and U3500 (N_3500,In_577,In_743);
or U3501 (N_3501,In_742,In_1510);
nand U3502 (N_3502,In_579,In_1767);
nand U3503 (N_3503,In_1463,In_1077);
nor U3504 (N_3504,In_667,In_1562);
or U3505 (N_3505,In_1295,In_614);
and U3506 (N_3506,In_1803,In_192);
nor U3507 (N_3507,In_1433,In_1435);
nand U3508 (N_3508,In_1981,In_97);
nand U3509 (N_3509,In_1122,In_479);
and U3510 (N_3510,In_323,In_1993);
nor U3511 (N_3511,In_1491,In_7);
or U3512 (N_3512,In_1422,In_972);
nor U3513 (N_3513,In_1753,In_907);
and U3514 (N_3514,In_1311,In_1927);
nand U3515 (N_3515,In_1425,In_1748);
nor U3516 (N_3516,In_1838,In_766);
or U3517 (N_3517,In_725,In_1712);
xnor U3518 (N_3518,In_1467,In_108);
nor U3519 (N_3519,In_443,In_1120);
xnor U3520 (N_3520,In_108,In_1387);
nor U3521 (N_3521,In_1963,In_1320);
nand U3522 (N_3522,In_186,In_1436);
or U3523 (N_3523,In_181,In_682);
or U3524 (N_3524,In_1288,In_1702);
nand U3525 (N_3525,In_609,In_1335);
nor U3526 (N_3526,In_235,In_1821);
xnor U3527 (N_3527,In_1969,In_1489);
nor U3528 (N_3528,In_1060,In_1838);
and U3529 (N_3529,In_619,In_305);
nand U3530 (N_3530,In_885,In_1006);
nor U3531 (N_3531,In_1286,In_1627);
or U3532 (N_3532,In_632,In_658);
and U3533 (N_3533,In_1153,In_1613);
nand U3534 (N_3534,In_732,In_25);
or U3535 (N_3535,In_1761,In_1930);
or U3536 (N_3536,In_1057,In_1718);
or U3537 (N_3537,In_338,In_1039);
or U3538 (N_3538,In_1974,In_808);
xnor U3539 (N_3539,In_1477,In_987);
or U3540 (N_3540,In_1767,In_1944);
nand U3541 (N_3541,In_69,In_1543);
nand U3542 (N_3542,In_1080,In_1948);
nor U3543 (N_3543,In_177,In_403);
nand U3544 (N_3544,In_1354,In_1582);
nor U3545 (N_3545,In_1444,In_89);
nand U3546 (N_3546,In_1460,In_1240);
and U3547 (N_3547,In_960,In_1012);
or U3548 (N_3548,In_1655,In_406);
or U3549 (N_3549,In_1710,In_1550);
and U3550 (N_3550,In_735,In_817);
nor U3551 (N_3551,In_1272,In_1768);
and U3552 (N_3552,In_1506,In_1686);
or U3553 (N_3553,In_909,In_1094);
or U3554 (N_3554,In_308,In_437);
nand U3555 (N_3555,In_1686,In_1570);
nand U3556 (N_3556,In_601,In_110);
and U3557 (N_3557,In_1056,In_1813);
nor U3558 (N_3558,In_184,In_355);
nand U3559 (N_3559,In_986,In_528);
nand U3560 (N_3560,In_1497,In_1127);
nand U3561 (N_3561,In_1098,In_1710);
or U3562 (N_3562,In_1529,In_1934);
nor U3563 (N_3563,In_1728,In_1455);
and U3564 (N_3564,In_881,In_762);
xor U3565 (N_3565,In_1608,In_1341);
nand U3566 (N_3566,In_905,In_1895);
nor U3567 (N_3567,In_959,In_1836);
or U3568 (N_3568,In_991,In_440);
and U3569 (N_3569,In_1161,In_327);
nor U3570 (N_3570,In_1664,In_225);
nor U3571 (N_3571,In_341,In_1222);
and U3572 (N_3572,In_18,In_353);
nand U3573 (N_3573,In_812,In_1406);
nor U3574 (N_3574,In_646,In_1742);
nand U3575 (N_3575,In_592,In_863);
nor U3576 (N_3576,In_938,In_817);
or U3577 (N_3577,In_485,In_668);
nand U3578 (N_3578,In_215,In_1991);
and U3579 (N_3579,In_1613,In_673);
nand U3580 (N_3580,In_1618,In_1881);
nor U3581 (N_3581,In_1019,In_1736);
or U3582 (N_3582,In_16,In_1355);
or U3583 (N_3583,In_1361,In_1400);
nand U3584 (N_3584,In_1579,In_556);
nand U3585 (N_3585,In_1661,In_1505);
xor U3586 (N_3586,In_1720,In_674);
and U3587 (N_3587,In_1970,In_542);
and U3588 (N_3588,In_1307,In_1615);
nand U3589 (N_3589,In_1043,In_1888);
nand U3590 (N_3590,In_947,In_651);
or U3591 (N_3591,In_668,In_62);
nand U3592 (N_3592,In_760,In_1433);
or U3593 (N_3593,In_0,In_661);
nor U3594 (N_3594,In_377,In_657);
nor U3595 (N_3595,In_1711,In_410);
nand U3596 (N_3596,In_151,In_528);
and U3597 (N_3597,In_1031,In_1869);
xnor U3598 (N_3598,In_410,In_1251);
nor U3599 (N_3599,In_85,In_228);
nand U3600 (N_3600,In_1610,In_925);
or U3601 (N_3601,In_834,In_240);
and U3602 (N_3602,In_940,In_158);
xnor U3603 (N_3603,In_1086,In_1293);
nand U3604 (N_3604,In_1932,In_1681);
xor U3605 (N_3605,In_1765,In_1725);
nand U3606 (N_3606,In_1815,In_1216);
and U3607 (N_3607,In_737,In_541);
and U3608 (N_3608,In_919,In_591);
nand U3609 (N_3609,In_1435,In_1824);
and U3610 (N_3610,In_1846,In_1955);
nand U3611 (N_3611,In_517,In_605);
nand U3612 (N_3612,In_86,In_1443);
and U3613 (N_3613,In_1721,In_1691);
or U3614 (N_3614,In_1084,In_747);
and U3615 (N_3615,In_408,In_933);
nand U3616 (N_3616,In_1157,In_1421);
nand U3617 (N_3617,In_363,In_1213);
or U3618 (N_3618,In_1201,In_368);
nand U3619 (N_3619,In_1002,In_1667);
nand U3620 (N_3620,In_1580,In_1451);
nor U3621 (N_3621,In_1371,In_1710);
nand U3622 (N_3622,In_553,In_753);
or U3623 (N_3623,In_1335,In_1267);
nand U3624 (N_3624,In_1984,In_1951);
nand U3625 (N_3625,In_828,In_334);
nand U3626 (N_3626,In_1459,In_1364);
nor U3627 (N_3627,In_1689,In_1718);
or U3628 (N_3628,In_350,In_1546);
or U3629 (N_3629,In_1999,In_965);
and U3630 (N_3630,In_12,In_1548);
nor U3631 (N_3631,In_641,In_51);
nand U3632 (N_3632,In_1071,In_1095);
or U3633 (N_3633,In_1660,In_1610);
xnor U3634 (N_3634,In_412,In_1963);
xor U3635 (N_3635,In_1538,In_450);
nor U3636 (N_3636,In_1769,In_902);
nor U3637 (N_3637,In_1129,In_410);
or U3638 (N_3638,In_1561,In_1562);
nor U3639 (N_3639,In_1330,In_1420);
and U3640 (N_3640,In_864,In_1449);
or U3641 (N_3641,In_1002,In_1341);
or U3642 (N_3642,In_744,In_1487);
nand U3643 (N_3643,In_971,In_961);
nor U3644 (N_3644,In_853,In_785);
or U3645 (N_3645,In_697,In_971);
nand U3646 (N_3646,In_1238,In_379);
nand U3647 (N_3647,In_1681,In_1916);
nand U3648 (N_3648,In_1146,In_408);
or U3649 (N_3649,In_784,In_1298);
and U3650 (N_3650,In_240,In_835);
nand U3651 (N_3651,In_1736,In_816);
nor U3652 (N_3652,In_1115,In_1109);
and U3653 (N_3653,In_1457,In_834);
nand U3654 (N_3654,In_905,In_1704);
or U3655 (N_3655,In_250,In_1320);
nor U3656 (N_3656,In_198,In_429);
and U3657 (N_3657,In_1671,In_597);
and U3658 (N_3658,In_1595,In_514);
and U3659 (N_3659,In_1488,In_1623);
nor U3660 (N_3660,In_130,In_1765);
nor U3661 (N_3661,In_1664,In_1295);
nor U3662 (N_3662,In_1632,In_692);
nand U3663 (N_3663,In_1468,In_1387);
nor U3664 (N_3664,In_1772,In_1660);
nand U3665 (N_3665,In_1824,In_437);
or U3666 (N_3666,In_1423,In_389);
nor U3667 (N_3667,In_473,In_1836);
and U3668 (N_3668,In_897,In_1853);
or U3669 (N_3669,In_242,In_1680);
nand U3670 (N_3670,In_1703,In_316);
nand U3671 (N_3671,In_125,In_824);
and U3672 (N_3672,In_1505,In_1433);
nand U3673 (N_3673,In_1866,In_354);
or U3674 (N_3674,In_476,In_1182);
and U3675 (N_3675,In_805,In_1208);
nor U3676 (N_3676,In_1651,In_1049);
and U3677 (N_3677,In_756,In_1406);
nand U3678 (N_3678,In_1327,In_109);
nor U3679 (N_3679,In_223,In_1688);
xnor U3680 (N_3680,In_1513,In_59);
nor U3681 (N_3681,In_926,In_1358);
nand U3682 (N_3682,In_1823,In_1906);
xor U3683 (N_3683,In_1636,In_71);
nor U3684 (N_3684,In_1757,In_465);
and U3685 (N_3685,In_296,In_14);
and U3686 (N_3686,In_466,In_360);
and U3687 (N_3687,In_1221,In_1091);
nand U3688 (N_3688,In_992,In_361);
nor U3689 (N_3689,In_1337,In_1960);
nand U3690 (N_3690,In_795,In_1191);
or U3691 (N_3691,In_1697,In_551);
or U3692 (N_3692,In_1414,In_527);
xnor U3693 (N_3693,In_420,In_1288);
or U3694 (N_3694,In_316,In_842);
or U3695 (N_3695,In_730,In_1375);
nand U3696 (N_3696,In_454,In_83);
nand U3697 (N_3697,In_483,In_44);
and U3698 (N_3698,In_230,In_814);
nor U3699 (N_3699,In_972,In_1889);
and U3700 (N_3700,In_1168,In_1961);
or U3701 (N_3701,In_168,In_445);
nand U3702 (N_3702,In_1867,In_26);
and U3703 (N_3703,In_1531,In_1285);
nand U3704 (N_3704,In_1671,In_1726);
or U3705 (N_3705,In_1884,In_685);
nor U3706 (N_3706,In_33,In_509);
or U3707 (N_3707,In_851,In_1755);
nand U3708 (N_3708,In_1915,In_1537);
and U3709 (N_3709,In_657,In_1718);
and U3710 (N_3710,In_439,In_1460);
or U3711 (N_3711,In_1685,In_701);
or U3712 (N_3712,In_331,In_1387);
and U3713 (N_3713,In_300,In_83);
nand U3714 (N_3714,In_61,In_1692);
nor U3715 (N_3715,In_707,In_1663);
or U3716 (N_3716,In_1537,In_742);
nor U3717 (N_3717,In_288,In_300);
and U3718 (N_3718,In_1075,In_131);
and U3719 (N_3719,In_1748,In_74);
nand U3720 (N_3720,In_85,In_1122);
nand U3721 (N_3721,In_429,In_59);
and U3722 (N_3722,In_1094,In_696);
nor U3723 (N_3723,In_351,In_1728);
and U3724 (N_3724,In_635,In_690);
nor U3725 (N_3725,In_99,In_395);
and U3726 (N_3726,In_1344,In_1564);
nor U3727 (N_3727,In_432,In_419);
and U3728 (N_3728,In_1829,In_1231);
or U3729 (N_3729,In_1892,In_763);
nand U3730 (N_3730,In_1944,In_928);
nor U3731 (N_3731,In_1560,In_829);
and U3732 (N_3732,In_1319,In_585);
nand U3733 (N_3733,In_1195,In_211);
nor U3734 (N_3734,In_127,In_1439);
and U3735 (N_3735,In_476,In_1351);
and U3736 (N_3736,In_537,In_80);
nand U3737 (N_3737,In_1249,In_1997);
and U3738 (N_3738,In_649,In_1282);
nor U3739 (N_3739,In_1465,In_1352);
nand U3740 (N_3740,In_945,In_1165);
xor U3741 (N_3741,In_834,In_32);
or U3742 (N_3742,In_1113,In_90);
xor U3743 (N_3743,In_1450,In_389);
xnor U3744 (N_3744,In_1070,In_827);
or U3745 (N_3745,In_1328,In_1240);
nand U3746 (N_3746,In_343,In_1275);
nand U3747 (N_3747,In_369,In_1515);
nand U3748 (N_3748,In_1793,In_69);
nor U3749 (N_3749,In_1780,In_1771);
or U3750 (N_3750,In_1550,In_221);
nor U3751 (N_3751,In_1457,In_1516);
xnor U3752 (N_3752,In_1892,In_1594);
nor U3753 (N_3753,In_1718,In_933);
or U3754 (N_3754,In_1640,In_145);
nor U3755 (N_3755,In_671,In_1886);
xnor U3756 (N_3756,In_1432,In_1807);
nor U3757 (N_3757,In_1865,In_1091);
or U3758 (N_3758,In_1088,In_1725);
nand U3759 (N_3759,In_98,In_1648);
nand U3760 (N_3760,In_385,In_851);
nor U3761 (N_3761,In_695,In_863);
nand U3762 (N_3762,In_544,In_896);
or U3763 (N_3763,In_1271,In_856);
nand U3764 (N_3764,In_1406,In_1766);
nor U3765 (N_3765,In_38,In_1536);
nand U3766 (N_3766,In_1959,In_460);
or U3767 (N_3767,In_1406,In_690);
and U3768 (N_3768,In_1850,In_403);
nor U3769 (N_3769,In_241,In_490);
nand U3770 (N_3770,In_1697,In_1335);
nand U3771 (N_3771,In_1452,In_205);
nor U3772 (N_3772,In_1615,In_1001);
and U3773 (N_3773,In_1257,In_1326);
or U3774 (N_3774,In_1107,In_1976);
xnor U3775 (N_3775,In_1138,In_675);
nand U3776 (N_3776,In_497,In_1218);
nor U3777 (N_3777,In_667,In_1741);
xnor U3778 (N_3778,In_1760,In_778);
xnor U3779 (N_3779,In_1417,In_864);
or U3780 (N_3780,In_1234,In_88);
nand U3781 (N_3781,In_355,In_296);
nand U3782 (N_3782,In_649,In_1810);
or U3783 (N_3783,In_34,In_835);
or U3784 (N_3784,In_678,In_849);
nor U3785 (N_3785,In_394,In_559);
and U3786 (N_3786,In_1736,In_1344);
or U3787 (N_3787,In_625,In_486);
or U3788 (N_3788,In_246,In_1093);
nor U3789 (N_3789,In_306,In_1048);
nand U3790 (N_3790,In_1174,In_348);
or U3791 (N_3791,In_1666,In_1027);
xnor U3792 (N_3792,In_100,In_121);
and U3793 (N_3793,In_634,In_1927);
nand U3794 (N_3794,In_1577,In_54);
or U3795 (N_3795,In_1260,In_706);
and U3796 (N_3796,In_1989,In_1928);
or U3797 (N_3797,In_1241,In_1535);
nand U3798 (N_3798,In_174,In_724);
nor U3799 (N_3799,In_1296,In_437);
nand U3800 (N_3800,In_1048,In_1750);
or U3801 (N_3801,In_734,In_985);
nand U3802 (N_3802,In_428,In_1524);
xnor U3803 (N_3803,In_859,In_1617);
and U3804 (N_3804,In_1088,In_819);
nand U3805 (N_3805,In_115,In_1710);
nand U3806 (N_3806,In_1529,In_646);
nand U3807 (N_3807,In_69,In_1403);
nand U3808 (N_3808,In_1094,In_99);
and U3809 (N_3809,In_1307,In_493);
xor U3810 (N_3810,In_460,In_1958);
or U3811 (N_3811,In_966,In_1073);
nand U3812 (N_3812,In_661,In_1515);
and U3813 (N_3813,In_1647,In_1558);
or U3814 (N_3814,In_1102,In_422);
nor U3815 (N_3815,In_1726,In_137);
nand U3816 (N_3816,In_1777,In_811);
and U3817 (N_3817,In_60,In_479);
and U3818 (N_3818,In_465,In_788);
and U3819 (N_3819,In_305,In_953);
and U3820 (N_3820,In_1551,In_1373);
nand U3821 (N_3821,In_1130,In_1501);
or U3822 (N_3822,In_1131,In_1544);
xnor U3823 (N_3823,In_1129,In_1108);
nand U3824 (N_3824,In_671,In_180);
xnor U3825 (N_3825,In_466,In_666);
nand U3826 (N_3826,In_1964,In_1610);
nor U3827 (N_3827,In_468,In_836);
nand U3828 (N_3828,In_1437,In_256);
nand U3829 (N_3829,In_1641,In_716);
or U3830 (N_3830,In_1221,In_1722);
nor U3831 (N_3831,In_1162,In_284);
and U3832 (N_3832,In_294,In_303);
nor U3833 (N_3833,In_322,In_273);
nor U3834 (N_3834,In_1582,In_173);
nand U3835 (N_3835,In_1454,In_1271);
and U3836 (N_3836,In_402,In_1890);
and U3837 (N_3837,In_1768,In_1073);
nand U3838 (N_3838,In_1849,In_1253);
nand U3839 (N_3839,In_454,In_1170);
and U3840 (N_3840,In_1785,In_1153);
nor U3841 (N_3841,In_1864,In_1682);
nand U3842 (N_3842,In_1529,In_382);
nor U3843 (N_3843,In_220,In_1924);
and U3844 (N_3844,In_1523,In_1476);
and U3845 (N_3845,In_622,In_333);
or U3846 (N_3846,In_12,In_284);
nor U3847 (N_3847,In_1427,In_53);
and U3848 (N_3848,In_525,In_947);
or U3849 (N_3849,In_19,In_82);
or U3850 (N_3850,In_1867,In_296);
nand U3851 (N_3851,In_53,In_255);
nor U3852 (N_3852,In_1682,In_1099);
and U3853 (N_3853,In_792,In_1549);
xnor U3854 (N_3854,In_1725,In_440);
nand U3855 (N_3855,In_577,In_1527);
xnor U3856 (N_3856,In_735,In_1235);
nand U3857 (N_3857,In_1641,In_1250);
and U3858 (N_3858,In_1873,In_618);
and U3859 (N_3859,In_1499,In_1135);
and U3860 (N_3860,In_774,In_1366);
nand U3861 (N_3861,In_45,In_1875);
or U3862 (N_3862,In_1169,In_1286);
nand U3863 (N_3863,In_43,In_437);
nand U3864 (N_3864,In_1145,In_596);
xnor U3865 (N_3865,In_1577,In_1147);
nor U3866 (N_3866,In_1767,In_364);
nor U3867 (N_3867,In_1146,In_516);
and U3868 (N_3868,In_907,In_1060);
nand U3869 (N_3869,In_709,In_1559);
or U3870 (N_3870,In_232,In_553);
and U3871 (N_3871,In_756,In_485);
and U3872 (N_3872,In_1556,In_410);
nor U3873 (N_3873,In_1473,In_1639);
nand U3874 (N_3874,In_518,In_446);
or U3875 (N_3875,In_1254,In_603);
nor U3876 (N_3876,In_540,In_1023);
or U3877 (N_3877,In_1038,In_231);
or U3878 (N_3878,In_1849,In_431);
nand U3879 (N_3879,In_98,In_1406);
nor U3880 (N_3880,In_1866,In_534);
nand U3881 (N_3881,In_318,In_934);
nor U3882 (N_3882,In_1358,In_349);
nor U3883 (N_3883,In_1001,In_1962);
and U3884 (N_3884,In_75,In_101);
nor U3885 (N_3885,In_861,In_1448);
and U3886 (N_3886,In_171,In_876);
and U3887 (N_3887,In_1248,In_1168);
or U3888 (N_3888,In_82,In_1057);
nor U3889 (N_3889,In_1998,In_588);
nand U3890 (N_3890,In_1795,In_825);
nand U3891 (N_3891,In_1809,In_1617);
nor U3892 (N_3892,In_185,In_1203);
nor U3893 (N_3893,In_1742,In_1345);
xnor U3894 (N_3894,In_1979,In_1985);
nand U3895 (N_3895,In_1815,In_1412);
nor U3896 (N_3896,In_446,In_1273);
nand U3897 (N_3897,In_1387,In_1837);
or U3898 (N_3898,In_1418,In_281);
and U3899 (N_3899,In_98,In_948);
or U3900 (N_3900,In_1742,In_230);
xnor U3901 (N_3901,In_1595,In_1103);
nand U3902 (N_3902,In_1259,In_440);
nor U3903 (N_3903,In_511,In_631);
or U3904 (N_3904,In_1520,In_1411);
nor U3905 (N_3905,In_870,In_1387);
and U3906 (N_3906,In_434,In_1814);
nand U3907 (N_3907,In_1658,In_308);
or U3908 (N_3908,In_1840,In_1489);
and U3909 (N_3909,In_916,In_1101);
or U3910 (N_3910,In_678,In_217);
nand U3911 (N_3911,In_251,In_838);
or U3912 (N_3912,In_1093,In_1853);
nor U3913 (N_3913,In_1365,In_590);
or U3914 (N_3914,In_1716,In_1567);
nor U3915 (N_3915,In_938,In_1358);
or U3916 (N_3916,In_1035,In_1115);
nor U3917 (N_3917,In_114,In_1944);
or U3918 (N_3918,In_1888,In_1738);
nor U3919 (N_3919,In_1191,In_1787);
xnor U3920 (N_3920,In_365,In_752);
and U3921 (N_3921,In_688,In_845);
nand U3922 (N_3922,In_641,In_1107);
nand U3923 (N_3923,In_1733,In_1568);
or U3924 (N_3924,In_1200,In_241);
and U3925 (N_3925,In_857,In_926);
nor U3926 (N_3926,In_859,In_1406);
nand U3927 (N_3927,In_401,In_310);
xor U3928 (N_3928,In_138,In_1593);
nand U3929 (N_3929,In_699,In_1102);
nand U3930 (N_3930,In_1901,In_1053);
nand U3931 (N_3931,In_1178,In_1900);
or U3932 (N_3932,In_1914,In_99);
or U3933 (N_3933,In_1440,In_505);
and U3934 (N_3934,In_1948,In_1952);
nand U3935 (N_3935,In_1399,In_1028);
or U3936 (N_3936,In_1606,In_513);
xor U3937 (N_3937,In_1214,In_1);
nor U3938 (N_3938,In_1725,In_1682);
and U3939 (N_3939,In_1995,In_454);
and U3940 (N_3940,In_1427,In_215);
nand U3941 (N_3941,In_530,In_836);
or U3942 (N_3942,In_123,In_451);
or U3943 (N_3943,In_1398,In_387);
and U3944 (N_3944,In_1669,In_183);
or U3945 (N_3945,In_601,In_1592);
nand U3946 (N_3946,In_734,In_1617);
nor U3947 (N_3947,In_197,In_1058);
nand U3948 (N_3948,In_706,In_1113);
nor U3949 (N_3949,In_274,In_1197);
and U3950 (N_3950,In_1987,In_1528);
nand U3951 (N_3951,In_175,In_38);
nor U3952 (N_3952,In_226,In_1079);
and U3953 (N_3953,In_1281,In_1753);
and U3954 (N_3954,In_1663,In_1754);
and U3955 (N_3955,In_1463,In_325);
and U3956 (N_3956,In_158,In_840);
and U3957 (N_3957,In_519,In_599);
and U3958 (N_3958,In_363,In_73);
and U3959 (N_3959,In_797,In_1717);
nand U3960 (N_3960,In_747,In_377);
and U3961 (N_3961,In_881,In_1936);
xor U3962 (N_3962,In_1856,In_967);
nand U3963 (N_3963,In_1199,In_1648);
nand U3964 (N_3964,In_1441,In_492);
nor U3965 (N_3965,In_1123,In_245);
nor U3966 (N_3966,In_1289,In_295);
nand U3967 (N_3967,In_1718,In_833);
nor U3968 (N_3968,In_1560,In_150);
nand U3969 (N_3969,In_331,In_792);
xnor U3970 (N_3970,In_578,In_415);
or U3971 (N_3971,In_1722,In_1296);
nand U3972 (N_3972,In_900,In_1804);
nor U3973 (N_3973,In_1807,In_1107);
nor U3974 (N_3974,In_616,In_507);
and U3975 (N_3975,In_1835,In_1628);
xor U3976 (N_3976,In_183,In_693);
nor U3977 (N_3977,In_203,In_1865);
or U3978 (N_3978,In_350,In_909);
nor U3979 (N_3979,In_1089,In_524);
and U3980 (N_3980,In_1238,In_124);
or U3981 (N_3981,In_47,In_256);
nand U3982 (N_3982,In_1813,In_1907);
nand U3983 (N_3983,In_786,In_1945);
nor U3984 (N_3984,In_1553,In_1157);
and U3985 (N_3985,In_936,In_548);
or U3986 (N_3986,In_402,In_1153);
nor U3987 (N_3987,In_1261,In_340);
or U3988 (N_3988,In_1839,In_212);
xnor U3989 (N_3989,In_1182,In_968);
and U3990 (N_3990,In_1997,In_1134);
or U3991 (N_3991,In_1667,In_1174);
nand U3992 (N_3992,In_490,In_843);
nand U3993 (N_3993,In_1193,In_809);
nand U3994 (N_3994,In_1396,In_1351);
xor U3995 (N_3995,In_1712,In_797);
nand U3996 (N_3996,In_1776,In_1923);
and U3997 (N_3997,In_1044,In_334);
and U3998 (N_3998,In_739,In_1127);
nor U3999 (N_3999,In_1576,In_1287);
or U4000 (N_4000,N_418,N_1924);
xnor U4001 (N_4001,N_3644,N_985);
and U4002 (N_4002,N_3404,N_3512);
nand U4003 (N_4003,N_3005,N_18);
xor U4004 (N_4004,N_1658,N_521);
or U4005 (N_4005,N_3344,N_3618);
or U4006 (N_4006,N_1294,N_2926);
or U4007 (N_4007,N_1961,N_882);
xnor U4008 (N_4008,N_2460,N_2719);
nor U4009 (N_4009,N_718,N_2676);
nor U4010 (N_4010,N_2645,N_590);
nand U4011 (N_4011,N_3761,N_268);
or U4012 (N_4012,N_105,N_3995);
xor U4013 (N_4013,N_3985,N_2907);
or U4014 (N_4014,N_63,N_1111);
or U4015 (N_4015,N_3540,N_1552);
or U4016 (N_4016,N_2277,N_1041);
xor U4017 (N_4017,N_523,N_2289);
and U4018 (N_4018,N_993,N_3851);
nand U4019 (N_4019,N_1689,N_2048);
or U4020 (N_4020,N_1458,N_371);
or U4021 (N_4021,N_433,N_561);
or U4022 (N_4022,N_1340,N_2989);
or U4023 (N_4023,N_747,N_857);
nand U4024 (N_4024,N_1663,N_3613);
and U4025 (N_4025,N_1138,N_3658);
or U4026 (N_4026,N_3726,N_711);
or U4027 (N_4027,N_3201,N_2133);
nor U4028 (N_4028,N_692,N_139);
or U4029 (N_4029,N_2835,N_3155);
nand U4030 (N_4030,N_859,N_2107);
and U4031 (N_4031,N_1272,N_2468);
nor U4032 (N_4032,N_3522,N_1886);
and U4033 (N_4033,N_94,N_3146);
or U4034 (N_4034,N_2484,N_121);
nand U4035 (N_4035,N_3162,N_1889);
and U4036 (N_4036,N_3511,N_228);
or U4037 (N_4037,N_1185,N_2440);
nand U4038 (N_4038,N_3434,N_1387);
nand U4039 (N_4039,N_1003,N_1516);
and U4040 (N_4040,N_2503,N_3941);
nor U4041 (N_4041,N_2581,N_3854);
or U4042 (N_4042,N_1607,N_1585);
nor U4043 (N_4043,N_1519,N_1157);
and U4044 (N_4044,N_680,N_357);
or U4045 (N_4045,N_2909,N_3362);
nor U4046 (N_4046,N_2718,N_45);
and U4047 (N_4047,N_2112,N_2208);
or U4048 (N_4048,N_1888,N_3841);
or U4049 (N_4049,N_380,N_3961);
and U4050 (N_4050,N_2128,N_3315);
or U4051 (N_4051,N_2281,N_3364);
and U4052 (N_4052,N_2722,N_3248);
or U4053 (N_4053,N_569,N_1567);
nor U4054 (N_4054,N_272,N_3786);
and U4055 (N_4055,N_2955,N_1483);
nor U4056 (N_4056,N_2652,N_2780);
nand U4057 (N_4057,N_1861,N_1600);
xnor U4058 (N_4058,N_3017,N_366);
and U4059 (N_4059,N_1477,N_1357);
nor U4060 (N_4060,N_3552,N_2459);
nand U4061 (N_4061,N_3097,N_1947);
nand U4062 (N_4062,N_748,N_1301);
nor U4063 (N_4063,N_1964,N_2467);
and U4064 (N_4064,N_2579,N_2479);
xnor U4065 (N_4065,N_1619,N_731);
and U4066 (N_4066,N_741,N_3307);
or U4067 (N_4067,N_1838,N_1461);
nand U4068 (N_4068,N_3982,N_3935);
nor U4069 (N_4069,N_3326,N_2951);
or U4070 (N_4070,N_1803,N_492);
nand U4071 (N_4071,N_738,N_1827);
and U4072 (N_4072,N_3564,N_740);
nand U4073 (N_4073,N_2414,N_3044);
nor U4074 (N_4074,N_2219,N_1900);
nor U4075 (N_4075,N_3389,N_354);
nand U4076 (N_4076,N_1231,N_239);
nand U4077 (N_4077,N_504,N_2760);
and U4078 (N_4078,N_2721,N_3451);
nor U4079 (N_4079,N_3497,N_1877);
or U4080 (N_4080,N_2668,N_2711);
nand U4081 (N_4081,N_2313,N_2191);
or U4082 (N_4082,N_799,N_1783);
nand U4083 (N_4083,N_1314,N_2055);
or U4084 (N_4084,N_3733,N_2160);
nor U4085 (N_4085,N_1471,N_1089);
and U4086 (N_4086,N_53,N_3177);
xnor U4087 (N_4087,N_1278,N_1743);
xnor U4088 (N_4088,N_2103,N_1184);
nand U4089 (N_4089,N_3927,N_1640);
xor U4090 (N_4090,N_2229,N_1636);
nor U4091 (N_4091,N_2430,N_2605);
nor U4092 (N_4092,N_888,N_3126);
nand U4093 (N_4093,N_1160,N_1595);
nor U4094 (N_4094,N_2084,N_2895);
or U4095 (N_4095,N_3690,N_1922);
nor U4096 (N_4096,N_3021,N_294);
and U4097 (N_4097,N_2373,N_557);
or U4098 (N_4098,N_3244,N_1059);
nor U4099 (N_4099,N_3744,N_3372);
nand U4100 (N_4100,N_3758,N_2236);
xnor U4101 (N_4101,N_3458,N_256);
nor U4102 (N_4102,N_1329,N_2530);
and U4103 (N_4103,N_2940,N_3719);
nand U4104 (N_4104,N_1420,N_2728);
or U4105 (N_4105,N_2851,N_3);
and U4106 (N_4106,N_3352,N_2022);
and U4107 (N_4107,N_2456,N_3297);
or U4108 (N_4108,N_1153,N_3863);
nand U4109 (N_4109,N_2777,N_328);
and U4110 (N_4110,N_3308,N_1047);
and U4111 (N_4111,N_714,N_1255);
or U4112 (N_4112,N_562,N_2498);
or U4113 (N_4113,N_1647,N_2746);
xor U4114 (N_4114,N_3240,N_1851);
and U4115 (N_4115,N_2602,N_568);
nand U4116 (N_4116,N_3101,N_1050);
nand U4117 (N_4117,N_2045,N_930);
or U4118 (N_4118,N_3489,N_949);
nand U4119 (N_4119,N_2221,N_1418);
or U4120 (N_4120,N_2376,N_2170);
nor U4121 (N_4121,N_1751,N_1234);
or U4122 (N_4122,N_2608,N_1762);
or U4123 (N_4123,N_323,N_5);
nor U4124 (N_4124,N_3537,N_906);
and U4125 (N_4125,N_3908,N_3846);
or U4126 (N_4126,N_242,N_2611);
or U4127 (N_4127,N_2988,N_2238);
xor U4128 (N_4128,N_1805,N_2408);
and U4129 (N_4129,N_3238,N_321);
or U4130 (N_4130,N_1912,N_2395);
or U4131 (N_4131,N_2396,N_3526);
nor U4132 (N_4132,N_1662,N_3460);
nor U4133 (N_4133,N_1131,N_1685);
and U4134 (N_4134,N_451,N_1722);
nand U4135 (N_4135,N_1645,N_752);
and U4136 (N_4136,N_3514,N_2454);
or U4137 (N_4137,N_2059,N_291);
nand U4138 (N_4138,N_3650,N_1732);
xor U4139 (N_4139,N_3797,N_1507);
or U4140 (N_4140,N_1996,N_2300);
and U4141 (N_4141,N_1885,N_2528);
or U4142 (N_4142,N_825,N_3600);
or U4143 (N_4143,N_2756,N_3082);
or U4144 (N_4144,N_3598,N_1720);
or U4145 (N_4145,N_3066,N_484);
and U4146 (N_4146,N_3542,N_2572);
or U4147 (N_4147,N_3322,N_315);
nor U4148 (N_4148,N_783,N_3055);
and U4149 (N_4149,N_1593,N_3815);
and U4150 (N_4150,N_3243,N_2158);
and U4151 (N_4151,N_3734,N_3158);
nand U4152 (N_4152,N_1150,N_3621);
nor U4153 (N_4153,N_2399,N_905);
and U4154 (N_4154,N_737,N_2670);
or U4155 (N_4155,N_858,N_1528);
nor U4156 (N_4156,N_3033,N_635);
and U4157 (N_4157,N_1313,N_1578);
or U4158 (N_4158,N_3046,N_1938);
and U4159 (N_4159,N_2570,N_3309);
nand U4160 (N_4160,N_1752,N_2069);
or U4161 (N_4161,N_3790,N_1355);
nor U4162 (N_4162,N_2730,N_10);
or U4163 (N_4163,N_1123,N_1086);
nor U4164 (N_4164,N_3675,N_3350);
and U4165 (N_4165,N_2280,N_2681);
or U4166 (N_4166,N_917,N_1857);
or U4167 (N_4167,N_1206,N_410);
nor U4168 (N_4168,N_2561,N_3090);
nand U4169 (N_4169,N_277,N_3902);
xor U4170 (N_4170,N_2911,N_2098);
nand U4171 (N_4171,N_1328,N_1773);
nand U4172 (N_4172,N_476,N_576);
nand U4173 (N_4173,N_1068,N_174);
and U4174 (N_4174,N_3660,N_2063);
and U4175 (N_4175,N_3229,N_2379);
and U4176 (N_4176,N_2637,N_1262);
or U4177 (N_4177,N_2862,N_97);
nor U4178 (N_4178,N_3380,N_1438);
nor U4179 (N_4179,N_2083,N_3314);
or U4180 (N_4180,N_3121,N_2000);
and U4181 (N_4181,N_2997,N_3933);
nand U4182 (N_4182,N_1077,N_3812);
or U4183 (N_4183,N_3356,N_96);
or U4184 (N_4184,N_2117,N_3197);
and U4185 (N_4185,N_643,N_3704);
or U4186 (N_4186,N_3345,N_2322);
and U4187 (N_4187,N_2812,N_2419);
or U4188 (N_4188,N_2226,N_3709);
or U4189 (N_4189,N_206,N_1425);
nor U4190 (N_4190,N_3979,N_219);
nor U4191 (N_4191,N_2639,N_1141);
nor U4192 (N_4192,N_2402,N_787);
nand U4193 (N_4193,N_2148,N_1655);
and U4194 (N_4194,N_2129,N_3396);
nor U4195 (N_4195,N_273,N_37);
and U4196 (N_4196,N_2825,N_3864);
xor U4197 (N_4197,N_3614,N_1914);
nor U4198 (N_4198,N_3518,N_3169);
nand U4199 (N_4199,N_325,N_2123);
or U4200 (N_4200,N_3701,N_2687);
or U4201 (N_4201,N_3775,N_1460);
or U4202 (N_4202,N_2305,N_1470);
and U4203 (N_4203,N_1181,N_707);
nand U4204 (N_4204,N_3479,N_962);
nand U4205 (N_4205,N_3640,N_773);
nor U4206 (N_4206,N_664,N_2776);
nand U4207 (N_4207,N_3508,N_3042);
and U4208 (N_4208,N_1613,N_1033);
nand U4209 (N_4209,N_1983,N_3799);
or U4210 (N_4210,N_275,N_2493);
nor U4211 (N_4211,N_1687,N_3471);
nor U4212 (N_4212,N_3305,N_1998);
nand U4213 (N_4213,N_3020,N_520);
nand U4214 (N_4214,N_3871,N_2883);
or U4215 (N_4215,N_3228,N_522);
nand U4216 (N_4216,N_2377,N_436);
xnor U4217 (N_4217,N_3943,N_1538);
nand U4218 (N_4218,N_3837,N_326);
nand U4219 (N_4219,N_1285,N_3065);
nor U4220 (N_4220,N_1739,N_3847);
and U4221 (N_4221,N_1412,N_113);
or U4222 (N_4222,N_1368,N_1383);
nor U4223 (N_4223,N_866,N_3431);
and U4224 (N_4224,N_3279,N_959);
or U4225 (N_4225,N_404,N_1030);
nor U4226 (N_4226,N_3610,N_2400);
and U4227 (N_4227,N_964,N_2380);
or U4228 (N_4228,N_3707,N_3679);
nand U4229 (N_4229,N_1795,N_1002);
nor U4230 (N_4230,N_2844,N_3168);
and U4231 (N_4231,N_2319,N_2032);
nand U4232 (N_4232,N_2949,N_1537);
nor U4233 (N_4233,N_3139,N_2630);
and U4234 (N_4234,N_1779,N_610);
nor U4235 (N_4235,N_2632,N_3688);
nand U4236 (N_4236,N_1839,N_3772);
nand U4237 (N_4237,N_2976,N_3413);
xnor U4238 (N_4238,N_1445,N_827);
or U4239 (N_4239,N_3237,N_1994);
nor U4240 (N_4240,N_2869,N_2854);
or U4241 (N_4241,N_2905,N_2049);
xor U4242 (N_4242,N_3195,N_1616);
or U4243 (N_4243,N_2209,N_1800);
nor U4244 (N_4244,N_3768,N_140);
nor U4245 (N_4245,N_1081,N_3608);
nand U4246 (N_4246,N_6,N_1563);
and U4247 (N_4247,N_1289,N_1604);
or U4248 (N_4248,N_148,N_2180);
nand U4249 (N_4249,N_182,N_593);
nand U4250 (N_4250,N_2551,N_2842);
xnor U4251 (N_4251,N_1865,N_2324);
nor U4252 (N_4252,N_2496,N_3009);
nand U4253 (N_4253,N_1032,N_1060);
xnor U4254 (N_4254,N_3683,N_1550);
or U4255 (N_4255,N_2397,N_1660);
and U4256 (N_4256,N_1337,N_1824);
xnor U4257 (N_4257,N_3999,N_911);
or U4258 (N_4258,N_3691,N_2432);
and U4259 (N_4259,N_1706,N_2426);
xnor U4260 (N_4260,N_1592,N_3298);
xor U4261 (N_4261,N_1807,N_3032);
nor U4262 (N_4262,N_3232,N_3106);
and U4263 (N_4263,N_1351,N_3947);
nand U4264 (N_4264,N_599,N_2071);
and U4265 (N_4265,N_3390,N_1723);
or U4266 (N_4266,N_1457,N_1837);
nand U4267 (N_4267,N_518,N_2298);
or U4268 (N_4268,N_419,N_64);
and U4269 (N_4269,N_570,N_3502);
nand U4270 (N_4270,N_2183,N_751);
nand U4271 (N_4271,N_1750,N_1731);
and U4272 (N_4272,N_2470,N_588);
nand U4273 (N_4273,N_1629,N_2125);
nor U4274 (N_4274,N_2534,N_1214);
and U4275 (N_4275,N_151,N_1200);
nor U4276 (N_4276,N_1918,N_3885);
or U4277 (N_4277,N_3070,N_2688);
nor U4278 (N_4278,N_112,N_2709);
nand U4279 (N_4279,N_2434,N_611);
nor U4280 (N_4280,N_943,N_3213);
or U4281 (N_4281,N_3482,N_2700);
nor U4282 (N_4282,N_1695,N_2953);
or U4283 (N_4283,N_2575,N_3071);
and U4284 (N_4284,N_1499,N_2783);
nor U4285 (N_4285,N_721,N_2030);
xnor U4286 (N_4286,N_3879,N_2110);
nand U4287 (N_4287,N_2891,N_3246);
nor U4288 (N_4288,N_3891,N_813);
nor U4289 (N_4289,N_2995,N_877);
nand U4290 (N_4290,N_1623,N_1866);
or U4291 (N_4291,N_1701,N_403);
nand U4292 (N_4292,N_3874,N_870);
xnor U4293 (N_4293,N_289,N_3636);
and U4294 (N_4294,N_3186,N_2809);
or U4295 (N_4295,N_3716,N_3111);
nor U4296 (N_4296,N_2475,N_3385);
or U4297 (N_4297,N_3260,N_2539);
nand U4298 (N_4298,N_2950,N_3109);
and U4299 (N_4299,N_938,N_3154);
and U4300 (N_4300,N_744,N_1842);
xnor U4301 (N_4301,N_2985,N_2513);
xor U4302 (N_4302,N_812,N_2114);
nor U4303 (N_4303,N_636,N_2983);
nor U4304 (N_4304,N_3916,N_1187);
and U4305 (N_4305,N_178,N_68);
or U4306 (N_4306,N_500,N_1652);
nor U4307 (N_4307,N_2308,N_1844);
nand U4308 (N_4308,N_2478,N_743);
or U4309 (N_4309,N_895,N_2175);
or U4310 (N_4310,N_3446,N_3634);
nor U4311 (N_4311,N_560,N_3409);
and U4312 (N_4312,N_1835,N_1905);
nor U4313 (N_4313,N_1121,N_3727);
and U4314 (N_4314,N_3140,N_3157);
nor U4315 (N_4315,N_3964,N_1758);
nand U4316 (N_4316,N_3967,N_591);
nor U4317 (N_4317,N_3737,N_1071);
nor U4318 (N_4318,N_1572,N_3004);
nand U4319 (N_4319,N_392,N_1946);
nand U4320 (N_4320,N_1674,N_3736);
nand U4321 (N_4321,N_1223,N_2364);
xor U4322 (N_4322,N_3207,N_379);
nand U4323 (N_4323,N_1566,N_1118);
nor U4324 (N_4324,N_2531,N_1063);
or U4325 (N_4325,N_578,N_1444);
and U4326 (N_4326,N_3003,N_699);
and U4327 (N_4327,N_1919,N_1478);
or U4328 (N_4328,N_59,N_3043);
xor U4329 (N_4329,N_3507,N_2898);
and U4330 (N_4330,N_2177,N_192);
and U4331 (N_4331,N_972,N_1980);
and U4332 (N_4332,N_57,N_1710);
and U4333 (N_4333,N_2301,N_2713);
nor U4334 (N_4334,N_55,N_2011);
nor U4335 (N_4335,N_3193,N_3304);
or U4336 (N_4336,N_2800,N_3699);
or U4337 (N_4337,N_3960,N_2421);
nor U4338 (N_4338,N_2269,N_1283);
or U4339 (N_4339,N_66,N_2973);
nand U4340 (N_4340,N_3234,N_815);
or U4341 (N_4341,N_848,N_3519);
or U4342 (N_4342,N_3755,N_211);
or U4343 (N_4343,N_903,N_3665);
nor U4344 (N_4344,N_2628,N_261);
nand U4345 (N_4345,N_627,N_545);
or U4346 (N_4346,N_909,N_2715);
or U4347 (N_4347,N_1811,N_2494);
or U4348 (N_4348,N_1381,N_579);
nor U4349 (N_4349,N_3324,N_123);
nor U4350 (N_4350,N_2559,N_3682);
or U4351 (N_4351,N_67,N_1801);
nand U4352 (N_4352,N_655,N_1057);
nor U4353 (N_4353,N_2734,N_3406);
and U4354 (N_4354,N_2387,N_3853);
or U4355 (N_4355,N_1279,N_3420);
and U4356 (N_4356,N_1416,N_3627);
nand U4357 (N_4357,N_1053,N_755);
and U4358 (N_4358,N_1523,N_1920);
nor U4359 (N_4359,N_873,N_1261);
and U4360 (N_4360,N_1869,N_1364);
nor U4361 (N_4361,N_1943,N_3814);
nand U4362 (N_4362,N_1124,N_1394);
and U4363 (N_4363,N_2463,N_3052);
or U4364 (N_4364,N_785,N_1429);
nor U4365 (N_4365,N_2742,N_1659);
nor U4366 (N_4366,N_9,N_1814);
and U4367 (N_4367,N_1197,N_1522);
nand U4368 (N_4368,N_2540,N_3029);
or U4369 (N_4369,N_3398,N_2127);
or U4370 (N_4370,N_2025,N_661);
nand U4371 (N_4371,N_806,N_1763);
nor U4372 (N_4372,N_805,N_2879);
nor U4373 (N_4373,N_2014,N_1910);
and U4374 (N_4374,N_1067,N_1316);
or U4375 (N_4375,N_1870,N_853);
nand U4376 (N_4376,N_493,N_2872);
nand U4377 (N_4377,N_1892,N_1873);
nor U4378 (N_4378,N_937,N_3646);
nand U4379 (N_4379,N_986,N_2873);
xor U4380 (N_4380,N_954,N_1854);
nand U4381 (N_4381,N_1448,N_2714);
and U4382 (N_4382,N_1242,N_1986);
and U4383 (N_4383,N_3647,N_2613);
nor U4384 (N_4384,N_1005,N_2710);
xor U4385 (N_4385,N_136,N_3194);
and U4386 (N_4386,N_1106,N_128);
or U4387 (N_4387,N_1426,N_372);
nand U4388 (N_4388,N_169,N_2369);
nand U4389 (N_4389,N_2607,N_2403);
or U4390 (N_4390,N_2801,N_698);
nor U4391 (N_4391,N_2405,N_1492);
xor U4392 (N_4392,N_3366,N_102);
and U4393 (N_4393,N_3118,N_958);
nand U4394 (N_4394,N_3787,N_1828);
nand U4395 (N_4395,N_3637,N_1711);
or U4396 (N_4396,N_2230,N_1271);
xor U4397 (N_4397,N_3373,N_3784);
nand U4398 (N_4398,N_2355,N_526);
and U4399 (N_4399,N_715,N_2027);
and U4400 (N_4400,N_2187,N_199);
and U4401 (N_4401,N_330,N_2625);
xor U4402 (N_4402,N_2987,N_1450);
or U4403 (N_4403,N_46,N_512);
nand U4404 (N_4404,N_965,N_1681);
or U4405 (N_4405,N_2947,N_2145);
nand U4406 (N_4406,N_2193,N_704);
or U4407 (N_4407,N_2488,N_3723);
xnor U4408 (N_4408,N_3831,N_3597);
nand U4409 (N_4409,N_3354,N_1440);
or U4410 (N_4410,N_2051,N_2136);
or U4411 (N_4411,N_975,N_686);
or U4412 (N_4412,N_3412,N_2860);
and U4413 (N_4413,N_1926,N_3554);
nor U4414 (N_4414,N_3441,N_449);
or U4415 (N_4415,N_2109,N_1560);
nor U4416 (N_4416,N_444,N_1353);
and U4417 (N_4417,N_2624,N_1867);
nand U4418 (N_4418,N_2699,N_1598);
xnor U4419 (N_4419,N_2684,N_2597);
and U4420 (N_4420,N_1698,N_2392);
nand U4421 (N_4421,N_193,N_150);
xor U4422 (N_4422,N_1001,N_1901);
or U4423 (N_4423,N_142,N_1709);
and U4424 (N_4424,N_2338,N_823);
xnor U4425 (N_4425,N_3265,N_2388);
nor U4426 (N_4426,N_235,N_2139);
xnor U4427 (N_4427,N_1302,N_1992);
nand U4428 (N_4428,N_957,N_682);
and U4429 (N_4429,N_229,N_999);
nand U4430 (N_4430,N_940,N_3226);
and U4431 (N_4431,N_2847,N_3942);
nor U4432 (N_4432,N_3416,N_1456);
nor U4433 (N_4433,N_2569,N_577);
nand U4434 (N_4434,N_1630,N_233);
nand U4435 (N_4435,N_3762,N_3687);
nor U4436 (N_4436,N_1721,N_2694);
and U4437 (N_4437,N_426,N_3068);
xnor U4438 (N_4438,N_2930,N_2691);
and U4439 (N_4439,N_2260,N_1384);
nor U4440 (N_4440,N_3190,N_1576);
and U4441 (N_4441,N_2075,N_3645);
and U4442 (N_4442,N_362,N_3069);
or U4443 (N_4443,N_2435,N_1699);
nand U4444 (N_4444,N_1392,N_1096);
and U4445 (N_4445,N_3612,N_149);
xnor U4446 (N_4446,N_2986,N_3206);
nand U4447 (N_4447,N_3290,N_3865);
or U4448 (N_4448,N_154,N_1973);
nor U4449 (N_4449,N_1291,N_1095);
or U4450 (N_4450,N_3287,N_2198);
and U4451 (N_4451,N_2696,N_879);
nor U4452 (N_4452,N_543,N_3463);
and U4453 (N_4453,N_2339,N_1974);
xnor U4454 (N_4454,N_622,N_423);
and U4455 (N_4455,N_989,N_318);
or U4456 (N_4456,N_2431,N_3253);
nor U4457 (N_4457,N_420,N_2367);
and U4458 (N_4458,N_3435,N_728);
and U4459 (N_4459,N_1476,N_1250);
or U4460 (N_4460,N_1380,N_2272);
nand U4461 (N_4461,N_1288,N_771);
and U4462 (N_4462,N_1939,N_3873);
nor U4463 (N_4463,N_3376,N_646);
nor U4464 (N_4464,N_1517,N_152);
and U4465 (N_4465,N_2267,N_3866);
or U4466 (N_4466,N_458,N_3250);
and U4467 (N_4467,N_1883,N_2088);
or U4468 (N_4468,N_3459,N_2775);
or U4469 (N_4469,N_2622,N_880);
and U4470 (N_4470,N_3303,N_1407);
nand U4471 (N_4471,N_3670,N_892);
nand U4472 (N_4472,N_2233,N_1521);
and U4473 (N_4473,N_1052,N_2254);
and U4474 (N_4474,N_1791,N_2795);
nand U4475 (N_4475,N_145,N_3249);
nor U4476 (N_4476,N_3087,N_2261);
nand U4477 (N_4477,N_2293,N_1836);
nand U4478 (N_4478,N_3590,N_1588);
nand U4479 (N_4479,N_3653,N_1682);
nand U4480 (N_4480,N_1562,N_2085);
xnor U4481 (N_4481,N_1748,N_2781);
nor U4482 (N_4482,N_2237,N_1804);
nor U4483 (N_4483,N_2287,N_2867);
or U4484 (N_4484,N_3785,N_1960);
nor U4485 (N_4485,N_2641,N_1236);
nor U4486 (N_4486,N_2234,N_3649);
or U4487 (N_4487,N_1847,N_2707);
nor U4488 (N_4488,N_2124,N_2271);
and U4489 (N_4489,N_3414,N_3132);
xnor U4490 (N_4490,N_131,N_990);
and U4491 (N_4491,N_3745,N_2766);
nand U4492 (N_4492,N_3626,N_2677);
and U4493 (N_4493,N_3342,N_3906);
nand U4494 (N_4494,N_2195,N_393);
and U4495 (N_4495,N_3657,N_3977);
or U4496 (N_4496,N_1495,N_2525);
xor U4497 (N_4497,N_1561,N_2303);
nand U4498 (N_4498,N_3513,N_2453);
and U4499 (N_4499,N_2,N_2247);
and U4500 (N_4500,N_2156,N_2587);
or U4501 (N_4501,N_1639,N_1789);
nand U4502 (N_4502,N_1670,N_2176);
or U4503 (N_4503,N_3583,N_1534);
and U4504 (N_4504,N_2481,N_1239);
and U4505 (N_4505,N_974,N_1366);
or U4506 (N_4506,N_2972,N_970);
and U4507 (N_4507,N_3832,N_1755);
nor U4508 (N_4508,N_1266,N_1072);
and U4509 (N_4509,N_257,N_3408);
nor U4510 (N_4510,N_2471,N_2061);
nor U4511 (N_4511,N_122,N_666);
nand U4512 (N_4512,N_378,N_1896);
nor U4513 (N_4513,N_2813,N_2593);
or U4514 (N_4514,N_78,N_1863);
nor U4515 (N_4515,N_2040,N_563);
or U4516 (N_4516,N_246,N_89);
nor U4517 (N_4517,N_3291,N_1580);
and U4518 (N_4518,N_2753,N_1044);
and U4519 (N_4519,N_1265,N_1858);
nor U4520 (N_4520,N_1207,N_2934);
nand U4521 (N_4521,N_2603,N_777);
or U4522 (N_4522,N_2329,N_963);
and U4523 (N_4523,N_3478,N_3926);
or U4524 (N_4524,N_2487,N_3769);
nor U4525 (N_4525,N_2465,N_3254);
nor U4526 (N_4526,N_3351,N_333);
and U4527 (N_4527,N_2994,N_3487);
and U4528 (N_4528,N_1376,N_2827);
xor U4529 (N_4529,N_416,N_2650);
nand U4530 (N_4530,N_447,N_1342);
xnor U4531 (N_4531,N_1930,N_3302);
nand U4532 (N_4532,N_1775,N_3115);
and U4533 (N_4533,N_1818,N_3818);
xnor U4534 (N_4534,N_1140,N_3081);
and U4535 (N_4535,N_3886,N_1671);
or U4536 (N_4536,N_3652,N_2149);
and U4537 (N_4537,N_3181,N_3602);
and U4538 (N_4538,N_2634,N_535);
nor U4539 (N_4539,N_1903,N_2619);
and U4540 (N_4540,N_689,N_373);
nor U4541 (N_4541,N_2469,N_2919);
and U4542 (N_4542,N_3607,N_1423);
or U4543 (N_4543,N_3661,N_1152);
and U4544 (N_4544,N_674,N_3599);
or U4545 (N_4545,N_1054,N_2331);
nor U4546 (N_4546,N_3993,N_1601);
or U4547 (N_4547,N_3363,N_1729);
or U4548 (N_4548,N_3387,N_3083);
nor U4549 (N_4549,N_2604,N_2921);
nand U4550 (N_4550,N_133,N_428);
or U4551 (N_4551,N_3791,N_3897);
or U4552 (N_4552,N_2076,N_933);
nand U4553 (N_4553,N_1802,N_3485);
or U4554 (N_4554,N_2595,N_2653);
or U4555 (N_4555,N_3631,N_3718);
or U4556 (N_4556,N_3317,N_2660);
nand U4557 (N_4557,N_2012,N_2394);
xnor U4558 (N_4558,N_3123,N_2480);
nand U4559 (N_4559,N_370,N_670);
and U4560 (N_4560,N_2119,N_3896);
nor U4561 (N_4561,N_3427,N_0);
nand U4562 (N_4562,N_1042,N_1897);
and U4563 (N_4563,N_3107,N_1841);
nor U4564 (N_4564,N_1718,N_3129);
or U4565 (N_4565,N_2999,N_168);
and U4566 (N_4566,N_2667,N_3208);
nor U4567 (N_4567,N_1904,N_30);
nor U4568 (N_4568,N_1617,N_2344);
nand U4569 (N_4569,N_546,N_1794);
xnor U4570 (N_4570,N_2749,N_3203);
nand U4571 (N_4571,N_934,N_3022);
or U4572 (N_4572,N_1916,N_3860);
nand U4573 (N_4573,N_3681,N_1415);
or U4574 (N_4574,N_1252,N_1275);
or U4575 (N_4575,N_1345,N_1307);
nand U4576 (N_4576,N_2391,N_3731);
and U4577 (N_4577,N_3088,N_1646);
nor U4578 (N_4578,N_177,N_2213);
and U4579 (N_4579,N_609,N_3383);
and U4580 (N_4580,N_1104,N_3062);
nand U4581 (N_4581,N_730,N_3375);
and U4582 (N_4582,N_1948,N_195);
nand U4583 (N_4583,N_2859,N_3209);
xnor U4584 (N_4584,N_1568,N_534);
and U4585 (N_4585,N_928,N_3689);
nand U4586 (N_4586,N_343,N_2981);
nand U4587 (N_4587,N_3040,N_1108);
xor U4588 (N_4588,N_1,N_1171);
nand U4589 (N_4589,N_3403,N_2818);
xnor U4590 (N_4590,N_2938,N_158);
nor U4591 (N_4591,N_2937,N_2946);
xnor U4592 (N_4592,N_2422,N_1066);
nand U4593 (N_4593,N_691,N_1962);
or U4594 (N_4594,N_1019,N_2965);
and U4595 (N_4595,N_2082,N_1970);
nand U4596 (N_4596,N_3076,N_2258);
and U4597 (N_4597,N_1875,N_1917);
and U4598 (N_4598,N_1642,N_3078);
xnor U4599 (N_4599,N_916,N_2351);
and U4600 (N_4600,N_3861,N_808);
and U4601 (N_4601,N_1968,N_29);
nand U4602 (N_4602,N_3929,N_2880);
nor U4603 (N_4603,N_1006,N_3759);
nand U4604 (N_4604,N_240,N_778);
or U4605 (N_4605,N_833,N_1178);
or U4606 (N_4606,N_3953,N_2356);
nand U4607 (N_4607,N_411,N_2621);
or U4608 (N_4608,N_1090,N_1332);
xor U4609 (N_4609,N_450,N_1374);
or U4610 (N_4610,N_1277,N_109);
and U4611 (N_4611,N_301,N_1690);
or U4612 (N_4612,N_948,N_1921);
or U4613 (N_4613,N_1324,N_467);
or U4614 (N_4614,N_3561,N_1350);
nor U4615 (N_4615,N_894,N_1254);
and U4616 (N_4616,N_2697,N_3161);
and U4617 (N_4617,N_1439,N_1764);
or U4618 (N_4618,N_596,N_2189);
nand U4619 (N_4619,N_555,N_2831);
or U4620 (N_4620,N_3028,N_3300);
and U4621 (N_4621,N_31,N_2325);
and U4622 (N_4622,N_460,N_2897);
xnor U4623 (N_4623,N_3750,N_2294);
nor U4624 (N_4624,N_1245,N_1008);
nor U4625 (N_4625,N_3368,N_1000);
or U4626 (N_4626,N_2428,N_795);
or U4627 (N_4627,N_1648,N_337);
nand U4628 (N_4628,N_2359,N_2924);
or U4629 (N_4629,N_471,N_3267);
nand U4630 (N_4630,N_2121,N_1369);
nand U4631 (N_4631,N_1370,N_3185);
and U4632 (N_4632,N_310,N_360);
and U4633 (N_4633,N_3242,N_1009);
or U4634 (N_4634,N_678,N_2750);
nor U4635 (N_4635,N_1031,N_3536);
or U4636 (N_4636,N_792,N_3781);
or U4637 (N_4637,N_2784,N_3027);
and U4638 (N_4638,N_2887,N_630);
nand U4639 (N_4639,N_2548,N_602);
and U4640 (N_4640,N_127,N_601);
nand U4641 (N_4641,N_375,N_3923);
and U4642 (N_4642,N_2599,N_597);
nand U4643 (N_4643,N_82,N_3360);
nor U4644 (N_4644,N_3259,N_2218);
or U4645 (N_4645,N_3705,N_2629);
and U4646 (N_4646,N_2635,N_3018);
nand U4647 (N_4647,N_683,N_791);
nor U4648 (N_4648,N_935,N_248);
or U4649 (N_4649,N_1098,N_559);
nor U4650 (N_4650,N_1693,N_3576);
and U4651 (N_4651,N_1631,N_3411);
and U4652 (N_4652,N_1297,N_696);
or U4653 (N_4653,N_3778,N_2410);
or U4654 (N_4654,N_2858,N_2120);
xor U4655 (N_4655,N_3934,N_1767);
nand U4656 (N_4656,N_2612,N_1115);
or U4657 (N_4657,N_3227,N_516);
nor U4658 (N_4658,N_1813,N_2565);
or U4659 (N_4659,N_1727,N_453);
nand U4660 (N_4660,N_3579,N_135);
nor U4661 (N_4661,N_3400,N_679);
and U4662 (N_4662,N_3819,N_1216);
or U4663 (N_4663,N_1982,N_2288);
nor U4664 (N_4664,N_3603,N_734);
xnor U4665 (N_4665,N_781,N_2816);
nor U4666 (N_4666,N_3456,N_782);
and U4667 (N_4667,N_3543,N_260);
and U4668 (N_4668,N_3549,N_1954);
xnor U4669 (N_4669,N_346,N_1437);
nand U4670 (N_4670,N_2497,N_1466);
nand U4671 (N_4671,N_759,N_3520);
and U4672 (N_4672,N_776,N_860);
xnor U4673 (N_4673,N_2249,N_3664);
nor U4674 (N_4674,N_3138,N_207);
nand U4675 (N_4675,N_1343,N_547);
nand U4676 (N_4676,N_1577,N_3437);
and U4677 (N_4677,N_1692,N_3025);
and U4678 (N_4678,N_3903,N_2547);
nor U4679 (N_4679,N_251,N_656);
nor U4680 (N_4680,N_2505,N_878);
xnor U4681 (N_4681,N_2520,N_24);
xor U4682 (N_4682,N_3525,N_114);
and U4683 (N_4683,N_2805,N_2015);
xor U4684 (N_4684,N_3720,N_2223);
nand U4685 (N_4685,N_3674,N_835);
nand U4686 (N_4686,N_3280,N_3810);
nor U4687 (N_4687,N_2115,N_1868);
nor U4688 (N_4688,N_3179,N_3320);
and U4689 (N_4689,N_1130,N_3095);
and U4690 (N_4690,N_3870,N_3651);
and U4691 (N_4691,N_549,N_2792);
and U4692 (N_4692,N_1621,N_2600);
or U4693 (N_4693,N_2659,N_1975);
and U4694 (N_4694,N_1367,N_384);
nand U4695 (N_4695,N_4,N_1608);
and U4696 (N_4696,N_1548,N_2970);
and U4697 (N_4697,N_2906,N_2332);
nand U4698 (N_4698,N_3659,N_27);
and U4699 (N_4699,N_1292,N_1719);
nor U4700 (N_4700,N_3706,N_2996);
nor U4701 (N_4701,N_3059,N_584);
and U4702 (N_4702,N_2253,N_2457);
xor U4703 (N_4703,N_1240,N_3261);
nand U4704 (N_4704,N_608,N_753);
or U4705 (N_4705,N_1190,N_1226);
nor U4706 (N_4706,N_3930,N_847);
xnor U4707 (N_4707,N_2929,N_2518);
nor U4708 (N_4708,N_3568,N_3211);
and U4709 (N_4709,N_984,N_1846);
nor U4710 (N_4710,N_829,N_1188);
nor U4711 (N_4711,N_1408,N_2449);
nor U4712 (N_4712,N_119,N_1880);
nor U4713 (N_4713,N_942,N_2004);
nand U4714 (N_4714,N_960,N_3036);
and U4715 (N_4715,N_3060,N_2056);
nor U4716 (N_4716,N_1990,N_1320);
or U4717 (N_4717,N_264,N_1389);
nor U4718 (N_4718,N_912,N_1399);
nor U4719 (N_4719,N_1787,N_1945);
nor U4720 (N_4720,N_837,N_1584);
nor U4721 (N_4721,N_129,N_1991);
nand U4722 (N_4722,N_455,N_1853);
nand U4723 (N_4723,N_2007,N_695);
or U4724 (N_4724,N_432,N_3676);
and U4725 (N_4725,N_2510,N_3306);
xnor U4726 (N_4726,N_565,N_160);
or U4727 (N_4727,N_3795,N_279);
or U4728 (N_4728,N_464,N_941);
or U4729 (N_4729,N_3822,N_2002);
nand U4730 (N_4730,N_2633,N_987);
or U4731 (N_4731,N_914,N_3767);
or U4732 (N_4732,N_1087,N_3149);
xnor U4733 (N_4733,N_3798,N_1318);
xor U4734 (N_4734,N_3937,N_3012);
nor U4735 (N_4735,N_3980,N_313);
xor U4736 (N_4736,N_1023,N_2594);
nor U4737 (N_4737,N_3624,N_2378);
nand U4738 (N_4738,N_1257,N_430);
nand U4739 (N_4739,N_1997,N_2340);
nand U4740 (N_4740,N_1045,N_2217);
or U4741 (N_4741,N_3394,N_377);
or U4742 (N_4742,N_100,N_209);
nor U4743 (N_4743,N_1469,N_98);
or U4744 (N_4744,N_869,N_1599);
nand U4745 (N_4745,N_1323,N_475);
or U4746 (N_4746,N_3183,N_2638);
and U4747 (N_4747,N_2242,N_3804);
nor U4748 (N_4748,N_2578,N_3285);
nand U4749 (N_4749,N_3475,N_2491);
nor U4750 (N_4750,N_1501,N_1944);
xnor U4751 (N_4751,N_2220,N_1191);
nand U4752 (N_4752,N_3473,N_3100);
nor U4753 (N_4753,N_3754,N_342);
nand U4754 (N_4754,N_3992,N_3278);
xnor U4755 (N_4755,N_2644,N_3057);
nand U4756 (N_4756,N_12,N_3780);
nor U4757 (N_4757,N_1872,N_2935);
and U4758 (N_4758,N_258,N_3551);
nor U4759 (N_4759,N_1541,N_2008);
and U4760 (N_4760,N_159,N_2678);
and U4761 (N_4761,N_3273,N_1128);
and U4762 (N_4762,N_3725,N_2462);
or U4763 (N_4763,N_2507,N_1170);
and U4764 (N_4764,N_3830,N_3465);
or U4765 (N_4765,N_3739,N_3048);
nor U4766 (N_4766,N_2057,N_3877);
nor U4767 (N_4767,N_831,N_750);
nand U4768 (N_4768,N_3135,N_2102);
and U4769 (N_4769,N_1144,N_3919);
nor U4770 (N_4770,N_69,N_2444);
or U4771 (N_4771,N_77,N_185);
nand U4772 (N_4772,N_2024,N_3742);
or U4773 (N_4773,N_3231,N_2211);
and U4774 (N_4774,N_3189,N_290);
nor U4775 (N_4775,N_196,N_2876);
and U4776 (N_4776,N_1386,N_657);
and U4777 (N_4777,N_3578,N_992);
and U4778 (N_4778,N_1549,N_3802);
or U4779 (N_4779,N_3876,N_3779);
or U4780 (N_4780,N_3843,N_2153);
nand U4781 (N_4781,N_1251,N_1155);
or U4782 (N_4782,N_70,N_2990);
nand U4783 (N_4783,N_2782,N_3058);
nor U4784 (N_4784,N_1734,N_241);
or U4785 (N_4785,N_2932,N_3756);
or U4786 (N_4786,N_1015,N_1558);
or U4787 (N_4787,N_3439,N_2314);
or U4788 (N_4788,N_1235,N_95);
and U4789 (N_4789,N_1116,N_3288);
or U4790 (N_4790,N_2093,N_687);
xnor U4791 (N_4791,N_2358,N_1753);
or U4792 (N_4792,N_1204,N_3589);
or U4793 (N_4793,N_1966,N_709);
xnor U4794 (N_4794,N_3887,N_3697);
and U4795 (N_4795,N_789,N_2197);
xor U4796 (N_4796,N_344,N_7);
nand U4797 (N_4797,N_1158,N_3581);
and U4798 (N_4798,N_702,N_308);
xor U4799 (N_4799,N_3274,N_3419);
or U4800 (N_4800,N_2517,N_3760);
or U4801 (N_4801,N_1653,N_1702);
and U4802 (N_4802,N_3823,N_1097);
or U4803 (N_4803,N_3272,N_3997);
nand U4804 (N_4804,N_3921,N_191);
or U4805 (N_4805,N_1075,N_595);
nor U4806 (N_4806,N_126,N_3480);
nand U4807 (N_4807,N_2586,N_1061);
nand U4808 (N_4808,N_3293,N_175);
and U4809 (N_4809,N_3477,N_3091);
or U4810 (N_4810,N_2618,N_1817);
nor U4811 (N_4811,N_1536,N_3880);
nor U4812 (N_4812,N_3604,N_1940);
nor U4813 (N_4813,N_3685,N_3532);
nand U4814 (N_4814,N_1151,N_162);
and U4815 (N_4815,N_1487,N_973);
nor U4816 (N_4816,N_265,N_1480);
or U4817 (N_4817,N_3067,N_573);
nand U4818 (N_4818,N_2870,N_437);
nand U4819 (N_4819,N_2370,N_1627);
or U4820 (N_4820,N_1286,N_2104);
xnor U4821 (N_4821,N_2347,N_1678);
or U4822 (N_4822,N_2589,N_1142);
or U4823 (N_4823,N_3539,N_3959);
nor U4824 (N_4824,N_2648,N_1082);
or U4825 (N_4825,N_3321,N_1784);
xnor U4826 (N_4826,N_409,N_3523);
and U4827 (N_4827,N_2447,N_498);
or U4828 (N_4828,N_3295,N_1428);
or U4829 (N_4829,N_3378,N_1179);
nor U4830 (N_4830,N_587,N_1213);
nand U4831 (N_4831,N_1571,N_2778);
or U4832 (N_4832,N_1183,N_2979);
or U4833 (N_4833,N_994,N_3538);
xor U4834 (N_4834,N_3517,N_3562);
nand U4835 (N_4835,N_1122,N_645);
nor U4836 (N_4836,N_1656,N_927);
xnor U4837 (N_4837,N_3774,N_14);
and U4838 (N_4838,N_334,N_3130);
and U4839 (N_4839,N_1531,N_3998);
and U4840 (N_4840,N_3041,N_2524);
xor U4841 (N_4841,N_3715,N_217);
and U4842 (N_4842,N_3116,N_3192);
and U4843 (N_4843,N_479,N_439);
xnor U4844 (N_4844,N_3686,N_3156);
xnor U4845 (N_4845,N_944,N_270);
or U4846 (N_4846,N_2461,N_921);
nor U4847 (N_4847,N_1893,N_2250);
nand U4848 (N_4848,N_3103,N_2923);
and U4849 (N_4849,N_2819,N_1378);
nor U4850 (N_4850,N_3367,N_224);
or U4851 (N_4851,N_3900,N_3711);
and U4852 (N_4852,N_1166,N_574);
nor U4853 (N_4853,N_2284,N_2884);
xnor U4854 (N_4854,N_44,N_34);
nand U4855 (N_4855,N_1198,N_2441);
and U4856 (N_4856,N_844,N_19);
nor U4857 (N_4857,N_1512,N_3013);
or U4858 (N_4858,N_1589,N_1891);
or U4859 (N_4859,N_115,N_49);
nor U4860 (N_4860,N_1344,N_1371);
nor U4861 (N_4861,N_2748,N_1154);
nor U4862 (N_4862,N_1246,N_3011);
and U4863 (N_4863,N_1159,N_3628);
nand U4864 (N_4864,N_3401,N_3438);
nand U4865 (N_4865,N_1309,N_3341);
nor U4866 (N_4866,N_1125,N_1569);
and U4867 (N_4867,N_3550,N_1430);
nor U4868 (N_4868,N_3630,N_1635);
and U4869 (N_4869,N_1410,N_3198);
or U4870 (N_4870,N_374,N_3230);
or U4871 (N_4871,N_2826,N_2159);
and U4872 (N_4872,N_1447,N_505);
nand U4873 (N_4873,N_710,N_288);
or U4874 (N_4874,N_572,N_1941);
xor U4875 (N_4875,N_2512,N_3617);
and U4876 (N_4876,N_99,N_463);
nor U4877 (N_4877,N_991,N_2747);
or U4878 (N_4878,N_1906,N_1282);
and U4879 (N_4879,N_1339,N_249);
or U4880 (N_4880,N_1756,N_2759);
nor U4881 (N_4881,N_339,N_1338);
and U4882 (N_4882,N_200,N_2323);
xnor U4883 (N_4883,N_1913,N_1049);
or U4884 (N_4884,N_640,N_3703);
and U4885 (N_4885,N_2669,N_745);
xnor U4886 (N_4886,N_582,N_603);
or U4887 (N_4887,N_1745,N_3488);
and U4888 (N_4888,N_1304,N_3811);
nand U4889 (N_4889,N_1145,N_3662);
xor U4890 (N_4890,N_3826,N_2786);
nor U4891 (N_4891,N_669,N_2966);
nand U4892 (N_4892,N_1280,N_788);
nor U4893 (N_4893,N_1276,N_3808);
and U4894 (N_4894,N_2150,N_3984);
nand U4895 (N_4895,N_2902,N_106);
and U4896 (N_4896,N_3467,N_2843);
or U4897 (N_4897,N_3708,N_3611);
nand U4898 (N_4898,N_606,N_1110);
and U4899 (N_4899,N_1675,N_3813);
and U4900 (N_4900,N_383,N_3642);
xnor U4901 (N_4901,N_915,N_3105);
nand U4902 (N_4902,N_2203,N_1064);
xor U4903 (N_4903,N_1615,N_23);
or U4904 (N_4904,N_3771,N_1212);
nand U4905 (N_4905,N_2886,N_2099);
nand U4906 (N_4906,N_2712,N_2553);
nand U4907 (N_4907,N_1219,N_1583);
xnor U4908 (N_4908,N_3049,N_2466);
and U4909 (N_4909,N_2855,N_717);
nand U4910 (N_4910,N_3370,N_890);
or U4911 (N_4911,N_1210,N_2758);
nor U4912 (N_4912,N_2875,N_564);
and U4913 (N_4913,N_2169,N_3379);
and U4914 (N_4914,N_1402,N_519);
nand U4915 (N_4915,N_3931,N_2841);
nand U4916 (N_4916,N_2166,N_604);
xor U4917 (N_4917,N_865,N_1076);
or U4918 (N_4918,N_722,N_3331);
or U4919 (N_4919,N_3257,N_2474);
nor U4920 (N_4920,N_3019,N_2200);
nand U4921 (N_4921,N_3428,N_624);
or U4922 (N_4922,N_1696,N_465);
and U4923 (N_4923,N_3638,N_3145);
or U4924 (N_4924,N_407,N_3484);
nor U4925 (N_4925,N_2346,N_3741);
nor U4926 (N_4926,N_3503,N_1707);
or U4927 (N_4927,N_2785,N_1134);
xor U4928 (N_4928,N_3494,N_2060);
and U4929 (N_4929,N_3800,N_2366);
nor U4930 (N_4930,N_1315,N_3498);
xor U4931 (N_4931,N_1065,N_3553);
nand U4932 (N_4932,N_1594,N_924);
or U4933 (N_4933,N_2890,N_925);
and U4934 (N_4934,N_1786,N_41);
nor U4935 (N_4935,N_936,N_468);
and U4936 (N_4936,N_1186,N_2372);
nand U4937 (N_4937,N_1391,N_3560);
or U4938 (N_4938,N_3178,N_2857);
and U4939 (N_4939,N_2222,N_1117);
or U4940 (N_4940,N_2146,N_3845);
and U4941 (N_4941,N_641,N_2140);
or U4942 (N_4942,N_1668,N_3382);
or U4943 (N_4943,N_1691,N_3848);
nor U4944 (N_4944,N_1493,N_202);
nand U4945 (N_4945,N_1273,N_2960);
xor U4946 (N_4946,N_3079,N_3968);
and U4947 (N_4947,N_74,N_2942);
nor U4948 (N_4948,N_1247,N_2874);
and U4949 (N_4949,N_3890,N_852);
nor U4950 (N_4950,N_2087,N_2773);
nand U4951 (N_4951,N_138,N_1884);
and U4952 (N_4952,N_1677,N_2941);
and U4953 (N_4953,N_1004,N_2583);
or U4954 (N_4954,N_809,N_1777);
and U4955 (N_4955,N_3884,N_1925);
and U4956 (N_4956,N_3667,N_1705);
and U4957 (N_4957,N_1942,N_861);
or U4958 (N_4958,N_2389,N_3641);
nor U4959 (N_4959,N_62,N_2577);
and U4960 (N_4960,N_1505,N_2216);
nor U4961 (N_4961,N_2446,N_532);
nand U4962 (N_4962,N_259,N_1573);
nor U4963 (N_4963,N_2010,N_3580);
nand U4964 (N_4964,N_502,N_881);
xnor U4965 (N_4965,N_652,N_2656);
or U4966 (N_4966,N_3978,N_1733);
nand U4967 (N_4967,N_3971,N_1361);
and U4968 (N_4968,N_1395,N_351);
nor U4969 (N_4969,N_1203,N_1632);
nor U4970 (N_4970,N_807,N_1356);
or U4971 (N_4971,N_2173,N_770);
nor U4972 (N_4972,N_335,N_278);
and U4973 (N_4973,N_2179,N_749);
nor U4974 (N_4974,N_651,N_3418);
nand U4975 (N_4975,N_3593,N_90);
nand U4976 (N_4976,N_1174,N_3974);
or U4977 (N_4977,N_3166,N_134);
and U4978 (N_4978,N_1700,N_3654);
nor U4979 (N_4979,N_3125,N_531);
and U4980 (N_4980,N_1774,N_3575);
xnor U4981 (N_4981,N_1358,N_3462);
nor U4982 (N_4982,N_225,N_236);
nand U4983 (N_4983,N_2536,N_2174);
xnor U4984 (N_4984,N_1027,N_1661);
and U4985 (N_4985,N_2967,N_2799);
nand U4986 (N_4986,N_1017,N_1379);
nor U4987 (N_4987,N_1874,N_3577);
or U4988 (N_4988,N_1020,N_1643);
nor U4989 (N_4989,N_2273,N_1797);
nand U4990 (N_4990,N_2817,N_1331);
nor U4991 (N_4991,N_2916,N_1069);
nor U4992 (N_4992,N_385,N_1781);
nand U4993 (N_4993,N_2144,N_843);
nand U4994 (N_4994,N_822,N_644);
xnor U4995 (N_4995,N_1555,N_2672);
nor U4996 (N_4996,N_398,N_3114);
nor U4997 (N_4997,N_1169,N_2404);
nand U4998 (N_4998,N_2840,N_1498);
and U4999 (N_4999,N_2535,N_667);
nor U5000 (N_5000,N_2090,N_1634);
nor U5001 (N_5001,N_1535,N_1793);
nor U5002 (N_5002,N_1127,N_446);
nand U5003 (N_5003,N_1895,N_1333);
xnor U5004 (N_5004,N_1024,N_2215);
nor U5005 (N_5005,N_726,N_3965);
nor U5006 (N_5006,N_312,N_3722);
or U5007 (N_5007,N_1951,N_2908);
and U5008 (N_5008,N_2849,N_2732);
nand U5009 (N_5009,N_425,N_3486);
and U5010 (N_5010,N_234,N_2590);
nor U5011 (N_5011,N_3160,N_266);
nor U5012 (N_5012,N_2567,N_2543);
nor U5013 (N_5013,N_1382,N_3239);
nor U5014 (N_5014,N_2142,N_3696);
nor U5015 (N_5015,N_2382,N_760);
nand U5016 (N_5016,N_1390,N_2917);
and U5017 (N_5017,N_3515,N_3147);
and U5018 (N_5018,N_1354,N_2674);
or U5019 (N_5019,N_3084,N_3858);
nand U5020 (N_5020,N_3159,N_761);
and U5021 (N_5021,N_2519,N_2546);
xnor U5022 (N_5022,N_1666,N_2499);
xor U5023 (N_5023,N_88,N_2936);
xnor U5024 (N_5024,N_167,N_3753);
or U5025 (N_5025,N_144,N_2134);
nor U5026 (N_5026,N_2852,N_1467);
or U5027 (N_5027,N_2365,N_3735);
nor U5028 (N_5028,N_1590,N_480);
or U5029 (N_5029,N_2155,N_2549);
nand U5030 (N_5030,N_2393,N_632);
and U5031 (N_5031,N_2167,N_2803);
nor U5032 (N_5032,N_3371,N_3442);
nand U5033 (N_5033,N_429,N_797);
nand U5034 (N_5034,N_2162,N_1375);
and U5035 (N_5035,N_3918,N_2054);
xnor U5036 (N_5036,N_2521,N_3895);
xor U5037 (N_5037,N_25,N_677);
and U5038 (N_5038,N_1497,N_887);
and U5039 (N_5039,N_2768,N_2477);
nor U5040 (N_5040,N_3310,N_2689);
nand U5041 (N_5041,N_253,N_1937);
and U5042 (N_5042,N_884,N_2885);
nor U5043 (N_5043,N_754,N_1205);
nor U5044 (N_5044,N_1021,N_2845);
or U5045 (N_5045,N_3165,N_571);
or U5046 (N_5046,N_2651,N_1274);
and U5047 (N_5047,N_929,N_3803);
and U5048 (N_5048,N_1167,N_359);
or U5049 (N_5049,N_2035,N_3991);
and U5050 (N_5050,N_3962,N_3085);
nor U5051 (N_5051,N_1602,N_1574);
nor U5052 (N_5052,N_2815,N_2508);
xnor U5053 (N_5053,N_1268,N_3595);
nor U5054 (N_5054,N_832,N_284);
and U5055 (N_5055,N_605,N_697);
nor U5056 (N_5056,N_483,N_1101);
and U5057 (N_5057,N_387,N_981);
nand U5058 (N_5058,N_402,N_390);
or U5059 (N_5059,N_314,N_388);
or U5060 (N_5060,N_600,N_3924);
xnor U5061 (N_5061,N_32,N_901);
and U5062 (N_5062,N_1760,N_3782);
nand U5063 (N_5063,N_1806,N_845);
and U5064 (N_5064,N_2643,N_311);
xnor U5065 (N_5065,N_486,N_2787);
nand U5066 (N_5066,N_198,N_1308);
or U5067 (N_5067,N_15,N_3566);
or U5068 (N_5068,N_1464,N_2232);
xor U5069 (N_5069,N_3531,N_1224);
and U5070 (N_5070,N_811,N_188);
and U5071 (N_5071,N_1051,N_2154);
or U5072 (N_5072,N_2956,N_871);
xor U5073 (N_5073,N_13,N_1139);
nand U5074 (N_5074,N_3233,N_638);
nor U5075 (N_5075,N_988,N_2894);
and U5076 (N_5076,N_1093,N_2761);
or U5077 (N_5077,N_1119,N_3357);
and U5078 (N_5078,N_1241,N_80);
xor U5079 (N_5079,N_2108,N_3766);
or U5080 (N_5080,N_769,N_1725);
nand U5081 (N_5081,N_3563,N_1928);
or U5082 (N_5082,N_1143,N_1890);
and U5083 (N_5083,N_700,N_1073);
and U5084 (N_5084,N_889,N_2239);
and U5085 (N_5085,N_1349,N_1649);
or U5086 (N_5086,N_3346,N_369);
or U5087 (N_5087,N_2945,N_2336);
nand U5088 (N_5088,N_1398,N_65);
and U5089 (N_5089,N_3051,N_1812);
nor U5090 (N_5090,N_269,N_978);
nor U5091 (N_5091,N_1688,N_1728);
and U5092 (N_5092,N_389,N_2771);
and U5093 (N_5093,N_2122,N_3330);
or U5094 (N_5094,N_1832,N_201);
nand U5095 (N_5095,N_1201,N_3910);
and U5096 (N_5096,N_1243,N_2720);
nand U5097 (N_5097,N_1253,N_2736);
and U5098 (N_5098,N_1401,N_2472);
nor U5099 (N_5099,N_1963,N_155);
and U5100 (N_5100,N_2627,N_541);
or U5101 (N_5101,N_3476,N_2727);
or U5102 (N_5102,N_2703,N_1433);
nor U5103 (N_5103,N_1526,N_3615);
nor U5104 (N_5104,N_1596,N_3432);
nor U5105 (N_5105,N_618,N_172);
or U5106 (N_5106,N_503,N_2527);
nand U5107 (N_5107,N_2762,N_1035);
and U5108 (N_5108,N_2243,N_230);
or U5109 (N_5109,N_101,N_497);
nand U5110 (N_5110,N_3976,N_2251);
nand U5111 (N_5111,N_3633,N_2779);
or U5112 (N_5112,N_3421,N_2334);
or U5113 (N_5113,N_904,N_1299);
and U5114 (N_5114,N_3151,N_8);
xor U5115 (N_5115,N_469,N_2172);
and U5116 (N_5116,N_1978,N_3415);
or U5117 (N_5117,N_2664,N_1776);
nand U5118 (N_5118,N_132,N_3572);
or U5119 (N_5119,N_979,N_1641);
or U5120 (N_5120,N_3868,N_2171);
nand U5121 (N_5121,N_2371,N_1849);
xor U5122 (N_5122,N_2974,N_305);
nor U5123 (N_5123,N_3588,N_2751);
xor U5124 (N_5124,N_3449,N_40);
and U5125 (N_5125,N_3948,N_705);
nor U5126 (N_5126,N_2086,N_2111);
and U5127 (N_5127,N_3796,N_161);
nor U5128 (N_5128,N_694,N_1591);
and U5129 (N_5129,N_117,N_2092);
nand U5130 (N_5130,N_1965,N_3541);
nor U5131 (N_5131,N_3505,N_802);
and U5132 (N_5132,N_1511,N_720);
and U5133 (N_5133,N_2566,N_2537);
and U5134 (N_5134,N_1409,N_2246);
nand U5135 (N_5135,N_967,N_1833);
and U5136 (N_5136,N_2839,N_3928);
xnor U5137 (N_5137,N_775,N_3289);
nand U5138 (N_5138,N_1221,N_1959);
or U5139 (N_5139,N_3878,N_2598);
nand U5140 (N_5140,N_2384,N_1432);
nor U5141 (N_5141,N_2285,N_3410);
or U5142 (N_5142,N_2882,N_955);
and U5143 (N_5143,N_2969,N_855);
xnor U5144 (N_5144,N_2295,N_2693);
or U5145 (N_5145,N_1672,N_3236);
nand U5146 (N_5146,N_79,N_3141);
xor U5147 (N_5147,N_690,N_3496);
nand U5148 (N_5148,N_668,N_765);
or U5149 (N_5149,N_316,N_3672);
nand U5150 (N_5150,N_237,N_2135);
nor U5151 (N_5151,N_1778,N_3256);
or U5152 (N_5152,N_840,N_189);
nand U5153 (N_5153,N_3089,N_3182);
and U5154 (N_5154,N_3872,N_1971);
and U5155 (N_5155,N_163,N_2482);
nor U5156 (N_5156,N_2584,N_1396);
nand U5157 (N_5157,N_61,N_1993);
nand U5158 (N_5158,N_1845,N_1113);
nand U5159 (N_5159,N_1650,N_1468);
or U5160 (N_5160,N_2838,N_3263);
nor U5161 (N_5161,N_293,N_3807);
nand U5162 (N_5162,N_3283,N_1303);
xor U5163 (N_5163,N_2913,N_3557);
or U5164 (N_5164,N_2126,N_47);
or U5165 (N_5165,N_1740,N_821);
or U5166 (N_5166,N_3712,N_2235);
and U5167 (N_5167,N_3889,N_2327);
xor U5168 (N_5168,N_2361,N_3472);
and U5169 (N_5169,N_3915,N_2094);
nor U5170 (N_5170,N_2201,N_1256);
nand U5171 (N_5171,N_2912,N_488);
nor U5172 (N_5172,N_1296,N_1435);
nor U5173 (N_5173,N_719,N_3037);
nand U5174 (N_5174,N_285,N_2206);
nor U5175 (N_5175,N_3509,N_1427);
nor U5176 (N_5176,N_215,N_3987);
nor U5177 (N_5177,N_3258,N_1133);
and U5178 (N_5178,N_262,N_804);
nand U5179 (N_5179,N_553,N_800);
nor U5180 (N_5180,N_617,N_2797);
and U5181 (N_5181,N_1673,N_3424);
nor U5182 (N_5182,N_474,N_2349);
or U5183 (N_5183,N_3296,N_2501);
and U5184 (N_5184,N_226,N_3695);
or U5185 (N_5185,N_1654,N_3187);
nor U5186 (N_5186,N_81,N_2157);
or U5187 (N_5187,N_1326,N_2515);
or U5188 (N_5188,N_2302,N_461);
xor U5189 (N_5189,N_1708,N_2888);
and U5190 (N_5190,N_3205,N_2291);
xor U5191 (N_5191,N_633,N_899);
nor U5192 (N_5192,N_36,N_659);
nand U5193 (N_5193,N_2182,N_3348);
xnor U5194 (N_5194,N_2614,N_1738);
nand U5195 (N_5195,N_3241,N_650);
nor U5196 (N_5196,N_1742,N_3825);
or U5197 (N_5197,N_2863,N_299);
nand U5198 (N_5198,N_1025,N_3565);
nand U5199 (N_5199,N_2436,N_634);
nor U5200 (N_5200,N_2601,N_3920);
or U5201 (N_5201,N_3524,N_3738);
nor U5202 (N_5202,N_1237,N_3112);
nand U5203 (N_5203,N_1735,N_197);
and U5204 (N_5204,N_3086,N_3990);
nand U5205 (N_5205,N_1074,N_1683);
nand U5206 (N_5206,N_3217,N_317);
nand U5207 (N_5207,N_897,N_2018);
and U5208 (N_5208,N_1132,N_3529);
or U5209 (N_5209,N_1199,N_1485);
nand U5210 (N_5210,N_1923,N_348);
and U5211 (N_5211,N_1244,N_2743);
or U5212 (N_5212,N_996,N_386);
nand U5213 (N_5213,N_1088,N_2933);
nor U5214 (N_5214,N_396,N_2096);
nor U5215 (N_5215,N_1744,N_626);
or U5216 (N_5216,N_623,N_456);
nand U5217 (N_5217,N_3469,N_2079);
or U5218 (N_5218,N_3124,N_1714);
xnor U5219 (N_5219,N_898,N_1581);
and U5220 (N_5220,N_250,N_2341);
nor U5221 (N_5221,N_1258,N_2592);
nor U5222 (N_5222,N_3835,N_544);
and U5223 (N_5223,N_3824,N_1644);
nor U5224 (N_5224,N_3006,N_153);
and U5225 (N_5225,N_3752,N_445);
nand U5226 (N_5226,N_2606,N_349);
nand U5227 (N_5227,N_16,N_1192);
and U5228 (N_5228,N_2975,N_3639);
or U5229 (N_5229,N_2409,N_22);
nor U5230 (N_5230,N_414,N_3635);
nor U5231 (N_5231,N_3461,N_2489);
nand U5232 (N_5232,N_3875,N_1300);
nand U5233 (N_5233,N_3443,N_2473);
nor U5234 (N_5234,N_1372,N_327);
nand U5235 (N_5235,N_1385,N_3061);
nor U5236 (N_5236,N_896,N_2490);
xor U5237 (N_5237,N_1749,N_2270);
nand U5238 (N_5238,N_11,N_187);
or U5239 (N_5239,N_3801,N_3457);
nor U5240 (N_5240,N_621,N_3144);
and U5241 (N_5241,N_3150,N_1957);
nand U5242 (N_5242,N_2978,N_3901);
or U5243 (N_5243,N_3235,N_3955);
and U5244 (N_5244,N_3007,N_130);
nand U5245 (N_5245,N_405,N_1759);
nand U5246 (N_5246,N_2977,N_2864);
nand U5247 (N_5247,N_2701,N_3113);
nor U5248 (N_5248,N_3972,N_648);
nand U5249 (N_5249,N_1182,N_17);
nand U5250 (N_5250,N_361,N_966);
nor U5251 (N_5251,N_345,N_1754);
nor U5252 (N_5252,N_442,N_3163);
nand U5253 (N_5253,N_2026,N_2914);
nor U5254 (N_5254,N_440,N_3904);
or U5255 (N_5255,N_2244,N_2675);
nand U5256 (N_5256,N_358,N_3102);
nor U5257 (N_5257,N_3134,N_397);
nor U5258 (N_5258,N_2959,N_3892);
and U5259 (N_5259,N_3063,N_2558);
and U5260 (N_5260,N_3817,N_1503);
nor U5261 (N_5261,N_3204,N_2192);
nor U5262 (N_5262,N_72,N_2058);
or U5263 (N_5263,N_3429,N_2296);
or U5264 (N_5264,N_1070,N_1149);
and U5265 (N_5265,N_1882,N_1424);
or U5266 (N_5266,N_2958,N_1414);
nor U5267 (N_5267,N_2716,N_1287);
or U5268 (N_5268,N_452,N_3355);
and U5269 (N_5269,N_1156,N_660);
and U5270 (N_5270,N_350,N_3417);
nand U5271 (N_5271,N_3064,N_2039);
nand U5272 (N_5272,N_1393,N_1229);
nor U5273 (N_5273,N_907,N_1684);
nor U5274 (N_5274,N_3867,N_1010);
xor U5275 (N_5275,N_3592,N_1525);
xor U5276 (N_5276,N_3423,N_3184);
xor U5277 (N_5277,N_2188,N_1988);
or U5278 (N_5278,N_1726,N_2706);
and U5279 (N_5279,N_1809,N_3313);
nand U5280 (N_5280,N_818,N_850);
nor U5281 (N_5281,N_764,N_1712);
nand U5282 (N_5282,N_3594,N_3840);
nor U5283 (N_5283,N_1894,N_3833);
nand U5284 (N_5284,N_922,N_2695);
and U5285 (N_5285,N_424,N_2665);
nor U5286 (N_5286,N_2588,N_868);
nand U5287 (N_5287,N_2770,N_3773);
xnor U5288 (N_5288,N_2509,N_509);
and U5289 (N_5289,N_181,N_2574);
and U5290 (N_5290,N_2647,N_2455);
and U5291 (N_5291,N_2964,N_2767);
xnor U5292 (N_5292,N_856,N_1228);
nor U5293 (N_5293,N_3905,N_676);
nand U5294 (N_5294,N_1189,N_3327);
xor U5295 (N_5295,N_296,N_413);
nand U5296 (N_5296,N_1411,N_1995);
and U5297 (N_5297,N_2089,N_2623);
or U5298 (N_5298,N_1079,N_2212);
xnor U5299 (N_5299,N_1757,N_111);
and U5300 (N_5300,N_2077,N_947);
nand U5301 (N_5301,N_2763,N_2661);
or U5302 (N_5302,N_3619,N_2041);
or U5303 (N_5303,N_1834,N_1730);
nor U5304 (N_5304,N_3499,N_2448);
and U5305 (N_5305,N_1488,N_2925);
nor U5306 (N_5306,N_3000,N_3023);
or U5307 (N_5307,N_3325,N_2091);
nor U5308 (N_5308,N_3605,N_3333);
nand U5309 (N_5309,N_368,N_2343);
nor U5310 (N_5310,N_2892,N_2342);
nor U5311 (N_5311,N_2013,N_51);
and U5312 (N_5312,N_3757,N_3131);
and U5313 (N_5313,N_619,N_1902);
xor U5314 (N_5314,N_300,N_3392);
and U5315 (N_5315,N_2881,N_2214);
xor U5316 (N_5316,N_324,N_3777);
nor U5317 (N_5317,N_472,N_3073);
nand U5318 (N_5318,N_2231,N_462);
and U5319 (N_5319,N_1542,N_3510);
nand U5320 (N_5320,N_920,N_2735);
and U5321 (N_5321,N_1579,N_3016);
nand U5322 (N_5322,N_716,N_3911);
or U5323 (N_5323,N_2846,N_1856);
nor U5324 (N_5324,N_819,N_891);
and U5325 (N_5325,N_254,N_2464);
nor U5326 (N_5326,N_103,N_3582);
and U5327 (N_5327,N_84,N_2196);
and U5328 (N_5328,N_2116,N_1509);
xor U5329 (N_5329,N_2225,N_2830);
xor U5330 (N_5330,N_2962,N_1442);
nor U5331 (N_5331,N_1091,N_3946);
nand U5332 (N_5332,N_1506,N_3792);
and U5333 (N_5333,N_3120,N_2292);
and U5334 (N_5334,N_2451,N_1105);
nand U5335 (N_5335,N_3913,N_21);
and U5336 (N_5336,N_3002,N_2557);
or U5337 (N_5337,N_629,N_2143);
or U5338 (N_5338,N_3788,N_1058);
or U5339 (N_5339,N_883,N_3839);
xor U5340 (N_5340,N_2576,N_1018);
or U5341 (N_5341,N_1825,N_3010);
nand U5342 (N_5342,N_1667,N_3031);
or U5343 (N_5343,N_1148,N_3764);
and U5344 (N_5344,N_2636,N_1881);
and U5345 (N_5345,N_2034,N_1999);
nor U5346 (N_5346,N_2374,N_2037);
nand U5347 (N_5347,N_1860,N_1554);
nor U5348 (N_5348,N_2755,N_2429);
and U5349 (N_5349,N_3128,N_3334);
or U5350 (N_5350,N_1766,N_35);
nand U5351 (N_5351,N_271,N_3196);
or U5352 (N_5352,N_3136,N_732);
and U5353 (N_5353,N_1195,N_2545);
or U5354 (N_5354,N_1360,N_3548);
xnor U5355 (N_5355,N_329,N_530);
and U5356 (N_5356,N_3223,N_3620);
xor U5357 (N_5357,N_708,N_2019);
nand U5358 (N_5358,N_614,N_1958);
nor U5359 (N_5359,N_3395,N_3655);
nor U5360 (N_5360,N_1611,N_1056);
nor U5361 (N_5361,N_3749,N_3648);
xor U5362 (N_5362,N_2275,N_231);
nand U5363 (N_5363,N_220,N_3692);
or U5364 (N_5364,N_1908,N_1909);
or U5365 (N_5365,N_427,N_3504);
and U5366 (N_5366,N_499,N_2297);
xor U5367 (N_5367,N_3047,N_3713);
nor U5368 (N_5368,N_3821,N_347);
nand U5369 (N_5369,N_1330,N_2416);
nor U5370 (N_5370,N_1290,N_685);
nand U5371 (N_5371,N_281,N_836);
xor U5372 (N_5372,N_1481,N_540);
and U5373 (N_5373,N_2984,N_3983);
nor U5374 (N_5374,N_1193,N_550);
nand U5375 (N_5375,N_3783,N_179);
and U5376 (N_5376,N_631,N_1486);
and U5377 (N_5377,N_1765,N_902);
and U5378 (N_5378,N_2915,N_303);
or U5379 (N_5379,N_3275,N_2033);
or U5380 (N_5380,N_2132,N_3585);
nor U5381 (N_5381,N_2686,N_533);
nor U5382 (N_5382,N_2582,N_218);
and U5383 (N_5383,N_2807,N_238);
or U5384 (N_5384,N_3133,N_2486);
or U5385 (N_5385,N_567,N_525);
and U5386 (N_5386,N_2304,N_2036);
nor U5387 (N_5387,N_3202,N_1474);
or U5388 (N_5388,N_3220,N_1967);
or U5389 (N_5389,N_1267,N_3883);
or U5390 (N_5390,N_1007,N_1352);
nor U5391 (N_5391,N_1614,N_2357);
or U5392 (N_5392,N_2005,N_2274);
xnor U5393 (N_5393,N_3836,N_2207);
nor U5394 (N_5394,N_1527,N_2381);
and U5395 (N_5395,N_3386,N_2824);
or U5396 (N_5396,N_1625,N_1036);
or U5397 (N_5397,N_1336,N_2789);
or U5398 (N_5398,N_2550,N_3717);
xnor U5399 (N_5399,N_1215,N_2205);
nor U5400 (N_5400,N_826,N_2811);
nand U5401 (N_5401,N_1515,N_2450);
nor U5402 (N_5402,N_2425,N_3152);
or U5403 (N_5403,N_1348,N_2317);
xor U5404 (N_5404,N_976,N_298);
or U5405 (N_5405,N_1887,N_3347);
nand U5406 (N_5406,N_1100,N_263);
nor U5407 (N_5407,N_244,N_3199);
nand U5408 (N_5408,N_3917,N_552);
nor U5409 (N_5409,N_2516,N_3174);
xnor U5410 (N_5410,N_1099,N_2310);
nand U5411 (N_5411,N_1936,N_1768);
xor U5412 (N_5412,N_932,N_3215);
nand U5413 (N_5413,N_1233,N_2417);
and U5414 (N_5414,N_507,N_575);
and U5415 (N_5415,N_3039,N_3949);
nand U5416 (N_5416,N_3958,N_3728);
or U5417 (N_5417,N_2282,N_2256);
or U5418 (N_5418,N_1147,N_1606);
nand U5419 (N_5419,N_2692,N_969);
nand U5420 (N_5420,N_75,N_2526);
and U5421 (N_5421,N_854,N_2963);
nor U5422 (N_5422,N_3216,N_1441);
nor U5423 (N_5423,N_3393,N_365);
nor U5424 (N_5424,N_2998,N_1788);
nor U5425 (N_5425,N_3632,N_1451);
or U5426 (N_5426,N_3732,N_867);
and U5427 (N_5427,N_3893,N_816);
nor U5428 (N_5428,N_1094,N_1500);
or U5429 (N_5429,N_3527,N_2662);
nand U5430 (N_5430,N_515,N_583);
or U5431 (N_5431,N_2837,N_104);
and U5432 (N_5432,N_1112,N_1180);
nor U5433 (N_5433,N_406,N_267);
nor U5434 (N_5434,N_2739,N_586);
or U5435 (N_5435,N_83,N_2368);
or U5436 (N_5436,N_60,N_1848);
and U5437 (N_5437,N_42,N_998);
and U5438 (N_5438,N_2311,N_1137);
nand U5439 (N_5439,N_1543,N_529);
nor U5440 (N_5440,N_340,N_1792);
nor U5441 (N_5441,N_1855,N_214);
nand U5442 (N_5442,N_3436,N_3212);
nor U5443 (N_5443,N_243,N_2903);
or U5444 (N_5444,N_3481,N_3859);
and U5445 (N_5445,N_820,N_2348);
and U5446 (N_5446,N_1084,N_3038);
nand U5447 (N_5447,N_766,N_2560);
or U5448 (N_5448,N_1587,N_1208);
nand U5449 (N_5449,N_3377,N_2649);
and U5450 (N_5450,N_2290,N_3493);
nand U5451 (N_5451,N_2406,N_1624);
and U5452 (N_5452,N_3533,N_1164);
and U5453 (N_5453,N_3951,N_1092);
nand U5454 (N_5454,N_3622,N_3492);
and U5455 (N_5455,N_322,N_3789);
or U5456 (N_5456,N_3671,N_2796);
nor U5457 (N_5457,N_2564,N_3932);
or U5458 (N_5458,N_3724,N_2445);
or U5459 (N_5459,N_2562,N_401);
or U5460 (N_5460,N_491,N_2413);
and U5461 (N_5461,N_2834,N_2823);
xor U5462 (N_5462,N_3751,N_2717);
nor U5463 (N_5463,N_356,N_58);
nor U5464 (N_5464,N_3255,N_3957);
nor U5465 (N_5465,N_1933,N_1502);
or U5466 (N_5466,N_931,N_513);
nand U5467 (N_5467,N_2554,N_3569);
nor U5468 (N_5468,N_1417,N_2407);
and U5469 (N_5469,N_839,N_286);
nand U5470 (N_5470,N_810,N_2016);
nand U5471 (N_5471,N_3391,N_1612);
xnor U5472 (N_5472,N_786,N_1981);
and U5473 (N_5473,N_585,N_2047);
or U5474 (N_5474,N_2105,N_1637);
or U5475 (N_5475,N_3669,N_3264);
or U5476 (N_5476,N_3381,N_834);
nor U5477 (N_5477,N_556,N_1799);
or U5478 (N_5478,N_3053,N_3829);
nor U5479 (N_5479,N_3015,N_1259);
nand U5480 (N_5480,N_3464,N_2227);
xnor U5481 (N_5481,N_2657,N_1724);
or U5482 (N_5482,N_2663,N_222);
xor U5483 (N_5483,N_1341,N_971);
nand U5484 (N_5484,N_3663,N_295);
nor U5485 (N_5485,N_2307,N_1175);
or U5486 (N_5486,N_3956,N_983);
nor U5487 (N_5487,N_2001,N_208);
nor U5488 (N_5488,N_862,N_3374);
nor U5489 (N_5489,N_1039,N_1546);
nand U5490 (N_5490,N_3173,N_1114);
nand U5491 (N_5491,N_3606,N_3008);
or U5492 (N_5492,N_1609,N_3444);
or U5493 (N_5493,N_2532,N_1984);
nor U5494 (N_5494,N_3573,N_1716);
nor U5495 (N_5495,N_2021,N_3730);
nor U5496 (N_5496,N_3328,N_2957);
or U5497 (N_5497,N_1346,N_1305);
nand U5498 (N_5498,N_3765,N_1772);
or U5499 (N_5499,N_3849,N_3301);
xor U5500 (N_5500,N_3700,N_364);
or U5501 (N_5501,N_2424,N_1168);
nor U5502 (N_5502,N_1494,N_2066);
nor U5503 (N_5503,N_2744,N_511);
nor U5504 (N_5504,N_496,N_2184);
and U5505 (N_5505,N_2330,N_2853);
or U5506 (N_5506,N_2420,N_2017);
and U5507 (N_5507,N_3122,N_1618);
or U5508 (N_5508,N_1222,N_2992);
nand U5509 (N_5509,N_3268,N_2968);
nand U5510 (N_5510,N_1551,N_2822);
or U5511 (N_5511,N_3556,N_2335);
and U5512 (N_5512,N_367,N_2118);
nand U5513 (N_5513,N_2680,N_1898);
xor U5514 (N_5514,N_1513,N_1109);
nand U5515 (N_5515,N_2878,N_477);
or U5516 (N_5516,N_1524,N_796);
nor U5517 (N_5517,N_1404,N_2993);
nand U5518 (N_5518,N_2555,N_3219);
nand U5519 (N_5519,N_280,N_2053);
nand U5520 (N_5520,N_2262,N_1202);
nor U5521 (N_5521,N_919,N_2257);
nand U5522 (N_5522,N_1405,N_1741);
nor U5523 (N_5523,N_1559,N_615);
nor U5524 (N_5524,N_3148,N_1327);
nand U5525 (N_5525,N_2255,N_165);
and U5526 (N_5526,N_56,N_1048);
nand U5527 (N_5527,N_968,N_3746);
nor U5528 (N_5528,N_886,N_2029);
or U5529 (N_5529,N_1406,N_341);
or U5530 (N_5530,N_276,N_2788);
or U5531 (N_5531,N_2020,N_2889);
nand U5532 (N_5532,N_2866,N_2326);
nand U5533 (N_5533,N_2168,N_73);
and U5534 (N_5534,N_3245,N_2194);
and U5535 (N_5535,N_1878,N_1540);
nor U5536 (N_5536,N_1782,N_3407);
or U5537 (N_5537,N_2401,N_3748);
and U5538 (N_5538,N_817,N_3643);
and U5539 (N_5539,N_1796,N_828);
nor U5540 (N_5540,N_1769,N_706);
and U5541 (N_5541,N_2097,N_1633);
xnor U5542 (N_5542,N_2806,N_3340);
or U5543 (N_5543,N_3994,N_252);
nand U5544 (N_5544,N_2658,N_658);
or U5545 (N_5545,N_110,N_1013);
or U5546 (N_5546,N_2299,N_1932);
or U5547 (N_5547,N_2939,N_2671);
nand U5548 (N_5548,N_654,N_616);
nor U5549 (N_5549,N_146,N_3856);
and U5550 (N_5550,N_441,N_514);
nor U5551 (N_5551,N_1260,N_2138);
nor U5552 (N_5552,N_412,N_3358);
nor U5553 (N_5553,N_363,N_71);
and U5554 (N_5554,N_1311,N_772);
or U5555 (N_5555,N_3842,N_86);
and U5556 (N_5556,N_1679,N_282);
nand U5557 (N_5557,N_443,N_1533);
nor U5558 (N_5558,N_3335,N_1575);
nor U5559 (N_5559,N_141,N_801);
or U5560 (N_5560,N_2829,N_408);
nor U5561 (N_5561,N_3050,N_1107);
nor U5562 (N_5562,N_2542,N_1704);
xor U5563 (N_5563,N_1703,N_125);
nand U5564 (N_5564,N_2263,N_3170);
or U5565 (N_5565,N_203,N_2802);
nor U5566 (N_5566,N_758,N_3721);
nor U5567 (N_5567,N_1570,N_1985);
or U5568 (N_5568,N_3099,N_3311);
nand U5569 (N_5569,N_331,N_2279);
or U5570 (N_5570,N_3282,N_307);
nand U5571 (N_5571,N_703,N_1102);
nand U5572 (N_5572,N_1934,N_536);
xor U5573 (N_5573,N_3072,N_194);
or U5574 (N_5574,N_2765,N_872);
nand U5575 (N_5575,N_3567,N_594);
or U5576 (N_5576,N_589,N_1230);
or U5577 (N_5577,N_2729,N_1694);
and U5578 (N_5578,N_2003,N_662);
nor U5579 (N_5579,N_1717,N_3452);
xnor U5580 (N_5580,N_2165,N_2820);
xnor U5581 (N_5581,N_3214,N_3276);
or U5582 (N_5582,N_2023,N_3077);
and U5583 (N_5583,N_2178,N_566);
nor U5584 (N_5584,N_2268,N_3143);
nand U5585 (N_5585,N_1664,N_2306);
and U5586 (N_5586,N_3056,N_2724);
nand U5587 (N_5587,N_746,N_3898);
nor U5588 (N_5588,N_1582,N_245);
and U5589 (N_5589,N_2360,N_3117);
and U5590 (N_5590,N_1269,N_2609);
nand U5591 (N_5591,N_2585,N_2333);
nor U5592 (N_5592,N_2130,N_1976);
nand U5593 (N_5593,N_2241,N_3093);
nand U5594 (N_5594,N_779,N_3266);
xnor U5595 (N_5595,N_2072,N_170);
nor U5596 (N_5596,N_2522,N_3422);
and U5597 (N_5597,N_3225,N_1915);
or U5598 (N_5598,N_2856,N_1989);
and U5599 (N_5599,N_2943,N_3361);
nand U5600 (N_5600,N_482,N_3433);
nand U5601 (N_5601,N_3677,N_1556);
nand U5602 (N_5602,N_3850,N_1931);
nand U5603 (N_5603,N_1085,N_147);
nand U5604 (N_5604,N_673,N_1949);
nand U5605 (N_5605,N_1565,N_3026);
nand U5606 (N_5606,N_2286,N_43);
nand U5607 (N_5607,N_1843,N_3680);
nor U5608 (N_5608,N_3176,N_2070);
nor U5609 (N_5609,N_3702,N_3545);
and U5610 (N_5610,N_1173,N_639);
nand U5611 (N_5611,N_1530,N_3402);
or U5612 (N_5612,N_1747,N_1586);
nor U5613 (N_5613,N_2533,N_3909);
nor U5614 (N_5614,N_1638,N_1373);
and U5615 (N_5615,N_2095,N_2141);
and U5616 (N_5616,N_1306,N_2354);
or U5617 (N_5617,N_3448,N_793);
and U5618 (N_5618,N_2848,N_183);
nor U5619 (N_5619,N_3966,N_2804);
and U5620 (N_5620,N_137,N_1979);
and U5621 (N_5621,N_2928,N_918);
or U5622 (N_5622,N_2224,N_2620);
or U5623 (N_5623,N_995,N_473);
xor U5624 (N_5624,N_2901,N_1270);
nor U5625 (N_5625,N_180,N_2511);
nor U5626 (N_5626,N_3470,N_733);
nand U5627 (N_5627,N_1831,N_2774);
nand U5628 (N_5628,N_2240,N_400);
and U5629 (N_5629,N_2485,N_2147);
nor U5630 (N_5630,N_3323,N_489);
and U5631 (N_5631,N_415,N_2278);
and U5632 (N_5632,N_3881,N_665);
nor U5633 (N_5633,N_422,N_309);
and U5634 (N_5634,N_1686,N_2363);
or U5635 (N_5635,N_3668,N_2685);
nor U5636 (N_5636,N_2199,N_581);
or U5637 (N_5637,N_459,N_3353);
nor U5638 (N_5638,N_3986,N_2861);
or U5639 (N_5639,N_1443,N_3714);
nor U5640 (N_5640,N_3834,N_1434);
nand U5641 (N_5641,N_1852,N_3944);
and U5642 (N_5642,N_2900,N_2046);
or U5643 (N_5643,N_2492,N_2458);
and U5644 (N_5644,N_1798,N_688);
and U5645 (N_5645,N_2131,N_213);
nor U5646 (N_5646,N_3337,N_297);
nor U5647 (N_5647,N_457,N_2113);
nor U5648 (N_5648,N_2794,N_2439);
nand U5649 (N_5649,N_2740,N_3936);
and U5650 (N_5650,N_2626,N_625);
nor U5651 (N_5651,N_1120,N_184);
and U5652 (N_5652,N_3950,N_2031);
xnor U5653 (N_5653,N_977,N_2769);
or U5654 (N_5654,N_1161,N_2443);
nor U5655 (N_5655,N_1136,N_28);
nor U5656 (N_5656,N_923,N_118);
or U5657 (N_5657,N_54,N_3430);
or U5658 (N_5658,N_255,N_1907);
nand U5659 (N_5659,N_3996,N_1489);
xor U5660 (N_5660,N_1298,N_1539);
or U5661 (N_5661,N_1626,N_3252);
nand U5662 (N_5662,N_2798,N_524);
or U5663 (N_5663,N_2640,N_945);
or U5664 (N_5664,N_798,N_3912);
xor U5665 (N_5665,N_2952,N_2164);
or U5666 (N_5666,N_1176,N_3809);
nor U5667 (N_5667,N_3001,N_3528);
nand U5668 (N_5668,N_2252,N_2375);
nand U5669 (N_5669,N_2573,N_1037);
or U5670 (N_5670,N_3740,N_3210);
xor U5671 (N_5671,N_3827,N_2318);
nand U5672 (N_5672,N_3332,N_87);
nor U5673 (N_5673,N_1810,N_736);
nand U5674 (N_5674,N_2064,N_2006);
nor U5675 (N_5675,N_3075,N_952);
xor U5676 (N_5676,N_2309,N_1310);
nand U5677 (N_5677,N_2836,N_319);
or U5678 (N_5678,N_3973,N_33);
or U5679 (N_5679,N_1227,N_3104);
nor U5680 (N_5680,N_2312,N_1547);
nor U5681 (N_5681,N_116,N_1815);
nand U5682 (N_5682,N_774,N_1544);
or U5683 (N_5683,N_50,N_1103);
or U5684 (N_5684,N_3609,N_3110);
and U5685 (N_5685,N_3535,N_3838);
nand U5686 (N_5686,N_863,N_1771);
nor U5687 (N_5687,N_2538,N_1826);
and U5688 (N_5688,N_1790,N_2495);
nand U5689 (N_5689,N_558,N_2723);
xnor U5690 (N_5690,N_1977,N_3534);
and U5691 (N_5691,N_3629,N_3558);
nand U5692 (N_5692,N_926,N_2666);
or U5693 (N_5693,N_3218,N_713);
xor U5694 (N_5694,N_3495,N_3440);
xnor U5695 (N_5695,N_2186,N_501);
or U5696 (N_5696,N_2733,N_592);
nor U5697 (N_5697,N_2137,N_3318);
and U5698 (N_5698,N_1564,N_824);
xor U5699 (N_5699,N_1325,N_1165);
nand U5700 (N_5700,N_1211,N_76);
nand U5701 (N_5701,N_3521,N_3656);
and U5702 (N_5702,N_1046,N_2910);
xor U5703 (N_5703,N_675,N_434);
nor U5704 (N_5704,N_3729,N_2427);
and U5705 (N_5705,N_1840,N_739);
nand U5706 (N_5706,N_431,N_2264);
and U5707 (N_5707,N_653,N_1557);
and U5708 (N_5708,N_2698,N_52);
nand U5709 (N_5709,N_3338,N_1012);
and U5710 (N_5710,N_3405,N_1490);
and U5711 (N_5711,N_527,N_763);
nor U5712 (N_5712,N_1377,N_448);
nand U5713 (N_5713,N_2276,N_2616);
nand U5714 (N_5714,N_1597,N_1862);
nor U5715 (N_5715,N_803,N_2044);
and U5716 (N_5716,N_1028,N_908);
or U5717 (N_5717,N_1449,N_2568);
and U5718 (N_5718,N_1676,N_2745);
xnor U5719 (N_5719,N_2893,N_3491);
or U5720 (N_5720,N_2764,N_3981);
or U5721 (N_5721,N_2954,N_3862);
nor U5722 (N_5722,N_1040,N_537);
and U5723 (N_5723,N_950,N_1334);
nand U5724 (N_5724,N_287,N_913);
nand U5725 (N_5725,N_780,N_1935);
and U5726 (N_5726,N_3559,N_164);
xor U5727 (N_5727,N_3952,N_186);
nand U5728 (N_5728,N_466,N_864);
nor U5729 (N_5729,N_2043,N_1473);
nand U5730 (N_5730,N_1238,N_1829);
or U5731 (N_5731,N_306,N_2248);
nand U5732 (N_5732,N_2904,N_1514);
or U5733 (N_5733,N_1532,N_1317);
xor U5734 (N_5734,N_3080,N_663);
or U5735 (N_5735,N_1780,N_3281);
nand U5736 (N_5736,N_3474,N_3343);
xor U5737 (N_5737,N_980,N_1436);
nand U5738 (N_5738,N_2411,N_1504);
nand U5739 (N_5739,N_2808,N_1078);
nand U5740 (N_5740,N_3172,N_1465);
nor U5741 (N_5741,N_3188,N_2814);
nand U5742 (N_5742,N_2028,N_910);
nor U5743 (N_5743,N_283,N_2362);
xor U5744 (N_5744,N_3591,N_1785);
nor U5745 (N_5745,N_3570,N_3500);
or U5746 (N_5746,N_2738,N_1713);
or U5747 (N_5747,N_2204,N_3445);
or U5748 (N_5748,N_3571,N_506);
xnor U5749 (N_5749,N_3625,N_85);
nand U5750 (N_5750,N_2552,N_3175);
or U5751 (N_5751,N_1146,N_838);
or U5752 (N_5752,N_2080,N_1479);
nor U5753 (N_5753,N_693,N_227);
nand U5754 (N_5754,N_3888,N_3693);
nor U5755 (N_5755,N_1455,N_3096);
xor U5756 (N_5756,N_1194,N_1879);
xnor U5757 (N_5757,N_3806,N_2931);
or U5758 (N_5758,N_3108,N_2106);
xnor U5759 (N_5759,N_2556,N_3349);
nand U5760 (N_5760,N_2352,N_320);
and U5761 (N_5761,N_223,N_1736);
xnor U5762 (N_5762,N_3925,N_2828);
nand U5763 (N_5763,N_173,N_3098);
nor U5764 (N_5764,N_580,N_1080);
xor U5765 (N_5765,N_2245,N_2433);
or U5766 (N_5766,N_3501,N_3271);
or U5767 (N_5767,N_956,N_2259);
nor U5768 (N_5768,N_3794,N_2922);
or U5769 (N_5769,N_1955,N_1620);
nor U5770 (N_5770,N_1062,N_1972);
nand U5771 (N_5771,N_3137,N_3277);
nor U5772 (N_5772,N_3970,N_742);
or U5773 (N_5773,N_2283,N_1322);
nand U5774 (N_5774,N_2832,N_628);
or U5775 (N_5775,N_3544,N_3466);
or U5776 (N_5776,N_3596,N_3171);
or U5777 (N_5777,N_2705,N_2673);
or U5778 (N_5778,N_26,N_551);
and U5779 (N_5779,N_1819,N_613);
nor U5780 (N_5780,N_830,N_3678);
and U5781 (N_5781,N_1055,N_3450);
nor U5782 (N_5782,N_2821,N_982);
and U5783 (N_5783,N_1876,N_2655);
nand U5784 (N_5784,N_1715,N_1697);
and U5785 (N_5785,N_2514,N_3384);
nand U5786 (N_5786,N_124,N_701);
or U5787 (N_5787,N_1026,N_3770);
xor U5788 (N_5788,N_1952,N_1510);
nor U5789 (N_5789,N_3447,N_3262);
nor U5790 (N_5790,N_1680,N_1603);
nor U5791 (N_5791,N_355,N_2702);
nand U5792 (N_5792,N_1929,N_612);
and U5793 (N_5793,N_712,N_3453);
nand U5794 (N_5794,N_2065,N_2181);
nor U5795 (N_5795,N_1911,N_2265);
nor U5796 (N_5796,N_2642,N_1129);
or U5797 (N_5797,N_684,N_2927);
or U5798 (N_5798,N_382,N_1746);
or U5799 (N_5799,N_3142,N_1518);
nand U5800 (N_5800,N_1126,N_794);
nand U5801 (N_5801,N_338,N_1987);
nand U5802 (N_5802,N_3828,N_2202);
xor U5803 (N_5803,N_2646,N_3035);
and U5804 (N_5804,N_2328,N_767);
nand U5805 (N_5805,N_671,N_2791);
nor U5806 (N_5806,N_1665,N_647);
xor U5807 (N_5807,N_3963,N_1293);
xor U5808 (N_5808,N_176,N_539);
xnor U5809 (N_5809,N_3221,N_1622);
nand U5810 (N_5810,N_1319,N_3425);
and U5811 (N_5811,N_2865,N_2737);
and U5812 (N_5812,N_2081,N_961);
or U5813 (N_5813,N_421,N_642);
nor U5814 (N_5814,N_1761,N_2591);
nand U5815 (N_5815,N_93,N_3694);
or U5816 (N_5816,N_790,N_1218);
or U5817 (N_5817,N_399,N_3855);
or U5818 (N_5818,N_435,N_120);
nand U5819 (N_5819,N_1335,N_3426);
or U5820 (N_5820,N_1196,N_494);
and U5821 (N_5821,N_391,N_1431);
and U5822 (N_5822,N_3747,N_1899);
nor U5823 (N_5823,N_1669,N_3024);
nor U5824 (N_5824,N_3490,N_3988);
and U5825 (N_5825,N_3365,N_997);
nand U5826 (N_5826,N_3894,N_2320);
or U5827 (N_5827,N_3584,N_2731);
nand U5828 (N_5828,N_2315,N_1083);
or U5829 (N_5829,N_2185,N_2228);
nor U5830 (N_5830,N_1022,N_735);
nand U5831 (N_5831,N_3336,N_381);
nor U5832 (N_5832,N_2790,N_1463);
or U5833 (N_5833,N_3616,N_2752);
nand U5834 (N_5834,N_2772,N_2982);
and U5835 (N_5835,N_542,N_672);
and U5836 (N_5836,N_3247,N_1264);
nor U5837 (N_5837,N_1529,N_1217);
nand U5838 (N_5838,N_3516,N_1459);
nor U5839 (N_5839,N_485,N_2679);
nor U5840 (N_5840,N_1397,N_2610);
or U5841 (N_5841,N_3776,N_495);
and U5842 (N_5842,N_2596,N_3388);
and U5843 (N_5843,N_3547,N_3153);
nand U5844 (N_5844,N_3483,N_3270);
nor U5845 (N_5845,N_171,N_3299);
nor U5846 (N_5846,N_1248,N_2321);
nor U5847 (N_5847,N_3922,N_1969);
or U5848 (N_5848,N_2415,N_1496);
or U5849 (N_5849,N_1553,N_3805);
nand U5850 (N_5850,N_1808,N_2654);
nor U5851 (N_5851,N_2423,N_454);
nor U5852 (N_5852,N_39,N_3034);
xor U5853 (N_5853,N_1820,N_723);
or U5854 (N_5854,N_1312,N_1816);
nand U5855 (N_5855,N_939,N_2529);
xnor U5856 (N_5856,N_607,N_3359);
nor U5857 (N_5857,N_1135,N_304);
nor U5858 (N_5858,N_874,N_487);
nand U5859 (N_5859,N_247,N_1823);
nand U5860 (N_5860,N_1491,N_1610);
nor U5861 (N_5861,N_3312,N_2971);
xnor U5862 (N_5862,N_3763,N_3939);
nor U5863 (N_5863,N_2704,N_2754);
nand U5864 (N_5864,N_2390,N_2100);
and U5865 (N_5865,N_3286,N_841);
or U5866 (N_5866,N_3397,N_1162);
or U5867 (N_5867,N_727,N_1520);
nand U5868 (N_5868,N_1830,N_3319);
and U5869 (N_5869,N_1482,N_2151);
or U5870 (N_5870,N_2353,N_353);
or U5871 (N_5871,N_352,N_1403);
nand U5872 (N_5872,N_2948,N_757);
nor U5873 (N_5873,N_1413,N_3710);
nor U5874 (N_5874,N_2877,N_2483);
and U5875 (N_5875,N_2210,N_1472);
or U5876 (N_5876,N_3743,N_3251);
or U5877 (N_5877,N_143,N_1484);
or U5878 (N_5878,N_417,N_2050);
or U5879 (N_5879,N_1454,N_91);
nand U5880 (N_5880,N_842,N_3269);
or U5881 (N_5881,N_2708,N_2437);
nand U5882 (N_5882,N_3945,N_2682);
nand U5883 (N_5883,N_2810,N_3454);
and U5884 (N_5884,N_2944,N_814);
and U5885 (N_5885,N_292,N_875);
nand U5886 (N_5886,N_212,N_3666);
nor U5887 (N_5887,N_3191,N_1038);
nor U5888 (N_5888,N_2920,N_190);
nand U5889 (N_5889,N_3546,N_3200);
nor U5890 (N_5890,N_724,N_510);
and U5891 (N_5891,N_3907,N_2161);
nand U5892 (N_5892,N_2741,N_1220);
and U5893 (N_5893,N_2961,N_637);
xor U5894 (N_5894,N_2580,N_649);
nand U5895 (N_5895,N_893,N_232);
or U5896 (N_5896,N_2523,N_1446);
nor U5897 (N_5897,N_48,N_3989);
xor U5898 (N_5898,N_953,N_3455);
nand U5899 (N_5899,N_210,N_2899);
and U5900 (N_5900,N_1651,N_2385);
and U5901 (N_5901,N_846,N_3092);
and U5902 (N_5902,N_1284,N_1347);
and U5903 (N_5903,N_3940,N_2101);
or U5904 (N_5904,N_1232,N_3816);
nor U5905 (N_5905,N_2563,N_1850);
or U5906 (N_5906,N_1956,N_395);
nand U5907 (N_5907,N_1363,N_1462);
nor U5908 (N_5908,N_1281,N_1605);
and U5909 (N_5909,N_478,N_3857);
or U5910 (N_5910,N_538,N_946);
and U5911 (N_5911,N_1225,N_2383);
or U5912 (N_5912,N_332,N_681);
and U5913 (N_5913,N_1657,N_885);
nor U5914 (N_5914,N_3292,N_166);
and U5915 (N_5915,N_108,N_3294);
and U5916 (N_5916,N_2980,N_2052);
nand U5917 (N_5917,N_1209,N_2038);
nor U5918 (N_5918,N_1822,N_1014);
xor U5919 (N_5919,N_1737,N_2571);
or U5920 (N_5920,N_204,N_1388);
nor U5921 (N_5921,N_3468,N_1927);
nand U5922 (N_5922,N_3167,N_1422);
or U5923 (N_5923,N_1871,N_2345);
nand U5924 (N_5924,N_3127,N_1950);
and U5925 (N_5925,N_3684,N_1172);
nand U5926 (N_5926,N_1770,N_3914);
and U5927 (N_5927,N_3586,N_3601);
and U5928 (N_5928,N_1163,N_3119);
and U5929 (N_5929,N_2452,N_3054);
and U5930 (N_5930,N_481,N_2871);
nand U5931 (N_5931,N_3316,N_1864);
and U5932 (N_5932,N_1362,N_3969);
and U5933 (N_5933,N_756,N_1029);
nand U5934 (N_5934,N_548,N_3882);
or U5935 (N_5935,N_3224,N_1628);
or U5936 (N_5936,N_2833,N_336);
nand U5937 (N_5937,N_1177,N_2073);
and U5938 (N_5938,N_876,N_394);
nor U5939 (N_5939,N_3844,N_2398);
and U5940 (N_5940,N_3284,N_768);
nor U5941 (N_5941,N_1453,N_725);
nand U5942 (N_5942,N_2190,N_2617);
and U5943 (N_5943,N_3045,N_3623);
and U5944 (N_5944,N_2793,N_2502);
xnor U5945 (N_5945,N_92,N_2850);
nand U5946 (N_5946,N_1953,N_156);
nor U5947 (N_5947,N_221,N_107);
or U5948 (N_5948,N_1263,N_2152);
nand U5949 (N_5949,N_2062,N_2386);
nand U5950 (N_5950,N_3869,N_598);
nand U5951 (N_5951,N_851,N_3954);
xor U5952 (N_5952,N_2504,N_2918);
nand U5953 (N_5953,N_470,N_2506);
and U5954 (N_5954,N_2541,N_1421);
nand U5955 (N_5955,N_2544,N_1043);
or U5956 (N_5956,N_3030,N_1859);
nor U5957 (N_5957,N_2418,N_274);
nor U5958 (N_5958,N_2074,N_157);
nand U5959 (N_5959,N_2337,N_3339);
and U5960 (N_5960,N_1016,N_3222);
nor U5961 (N_5961,N_1400,N_3587);
nor U5962 (N_5962,N_2725,N_3014);
and U5963 (N_5963,N_3074,N_3506);
nor U5964 (N_5964,N_517,N_762);
xor U5965 (N_5965,N_784,N_2631);
and U5966 (N_5966,N_216,N_2442);
nand U5967 (N_5967,N_2266,N_2009);
or U5968 (N_5968,N_1365,N_3530);
nand U5969 (N_5969,N_1359,N_2615);
and U5970 (N_5970,N_2163,N_302);
xnor U5971 (N_5971,N_1295,N_3399);
xor U5972 (N_5972,N_3938,N_3852);
nor U5973 (N_5973,N_1475,N_951);
and U5974 (N_5974,N_1545,N_20);
nand U5975 (N_5975,N_2078,N_3369);
xnor U5976 (N_5976,N_508,N_38);
or U5977 (N_5977,N_490,N_2690);
and U5978 (N_5978,N_2068,N_1011);
nor U5979 (N_5979,N_2067,N_1452);
nand U5980 (N_5980,N_620,N_3698);
nand U5981 (N_5981,N_2991,N_2042);
nand U5982 (N_5982,N_205,N_1821);
nor U5983 (N_5983,N_2896,N_849);
and U5984 (N_5984,N_1508,N_1419);
and U5985 (N_5985,N_3793,N_2412);
or U5986 (N_5986,N_3975,N_2757);
nor U5987 (N_5987,N_2683,N_3164);
and U5988 (N_5988,N_3673,N_3094);
nand U5989 (N_5989,N_2316,N_2476);
or U5990 (N_5990,N_3574,N_376);
and U5991 (N_5991,N_3555,N_438);
nor U5992 (N_5992,N_1034,N_2350);
or U5993 (N_5993,N_3180,N_528);
and U5994 (N_5994,N_900,N_1249);
or U5995 (N_5995,N_2868,N_729);
nor U5996 (N_5996,N_2726,N_2500);
or U5997 (N_5997,N_554,N_1321);
nand U5998 (N_5998,N_2438,N_3329);
and U5999 (N_5999,N_3899,N_3820);
xor U6000 (N_6000,N_332,N_550);
or U6001 (N_6001,N_3355,N_537);
or U6002 (N_6002,N_729,N_741);
nor U6003 (N_6003,N_3969,N_823);
nor U6004 (N_6004,N_735,N_1046);
and U6005 (N_6005,N_1353,N_3221);
nand U6006 (N_6006,N_713,N_467);
nand U6007 (N_6007,N_2190,N_1529);
nor U6008 (N_6008,N_161,N_3586);
nor U6009 (N_6009,N_2928,N_153);
xnor U6010 (N_6010,N_3686,N_2509);
and U6011 (N_6011,N_2144,N_831);
or U6012 (N_6012,N_751,N_2983);
and U6013 (N_6013,N_3641,N_3510);
xor U6014 (N_6014,N_3230,N_1024);
nor U6015 (N_6015,N_1521,N_1142);
nand U6016 (N_6016,N_263,N_3001);
nor U6017 (N_6017,N_2115,N_755);
nor U6018 (N_6018,N_3760,N_1891);
xnor U6019 (N_6019,N_1404,N_651);
and U6020 (N_6020,N_1944,N_3239);
nand U6021 (N_6021,N_472,N_1842);
and U6022 (N_6022,N_3559,N_3530);
nor U6023 (N_6023,N_3284,N_55);
nor U6024 (N_6024,N_2598,N_3451);
xor U6025 (N_6025,N_2383,N_2678);
or U6026 (N_6026,N_2757,N_425);
or U6027 (N_6027,N_2819,N_3113);
or U6028 (N_6028,N_2415,N_687);
and U6029 (N_6029,N_769,N_403);
or U6030 (N_6030,N_1603,N_3154);
and U6031 (N_6031,N_1635,N_564);
nand U6032 (N_6032,N_2843,N_2604);
nor U6033 (N_6033,N_2147,N_3952);
xor U6034 (N_6034,N_2590,N_2328);
nor U6035 (N_6035,N_3806,N_535);
nand U6036 (N_6036,N_215,N_3127);
and U6037 (N_6037,N_3887,N_740);
xor U6038 (N_6038,N_89,N_727);
nor U6039 (N_6039,N_1405,N_2291);
or U6040 (N_6040,N_2035,N_2716);
nand U6041 (N_6041,N_2363,N_150);
or U6042 (N_6042,N_2858,N_878);
or U6043 (N_6043,N_3005,N_3830);
nand U6044 (N_6044,N_2056,N_3544);
nand U6045 (N_6045,N_2302,N_2192);
xor U6046 (N_6046,N_1170,N_3659);
nor U6047 (N_6047,N_2105,N_3398);
nand U6048 (N_6048,N_369,N_873);
and U6049 (N_6049,N_667,N_2659);
xor U6050 (N_6050,N_1726,N_3574);
nand U6051 (N_6051,N_2061,N_3106);
xor U6052 (N_6052,N_3965,N_974);
or U6053 (N_6053,N_451,N_3361);
nor U6054 (N_6054,N_1539,N_3168);
or U6055 (N_6055,N_2201,N_2758);
and U6056 (N_6056,N_2293,N_2377);
nor U6057 (N_6057,N_250,N_2776);
or U6058 (N_6058,N_3852,N_3624);
nand U6059 (N_6059,N_3815,N_1144);
or U6060 (N_6060,N_687,N_1388);
xnor U6061 (N_6061,N_982,N_3415);
nor U6062 (N_6062,N_1993,N_1789);
or U6063 (N_6063,N_3574,N_2230);
and U6064 (N_6064,N_1618,N_1554);
xor U6065 (N_6065,N_1874,N_1098);
nand U6066 (N_6066,N_2420,N_3457);
or U6067 (N_6067,N_221,N_3532);
and U6068 (N_6068,N_1577,N_3584);
nand U6069 (N_6069,N_169,N_3639);
or U6070 (N_6070,N_592,N_1247);
nand U6071 (N_6071,N_1180,N_2284);
or U6072 (N_6072,N_753,N_3907);
nand U6073 (N_6073,N_3058,N_1960);
xor U6074 (N_6074,N_1399,N_2027);
nand U6075 (N_6075,N_2315,N_1967);
nor U6076 (N_6076,N_1211,N_2022);
or U6077 (N_6077,N_456,N_1769);
or U6078 (N_6078,N_1647,N_3446);
or U6079 (N_6079,N_3064,N_625);
or U6080 (N_6080,N_267,N_1646);
nor U6081 (N_6081,N_1992,N_446);
and U6082 (N_6082,N_838,N_2660);
nor U6083 (N_6083,N_2836,N_3652);
or U6084 (N_6084,N_2105,N_2485);
xor U6085 (N_6085,N_1717,N_1343);
xnor U6086 (N_6086,N_3770,N_3445);
and U6087 (N_6087,N_3497,N_3282);
and U6088 (N_6088,N_2565,N_441);
nand U6089 (N_6089,N_2547,N_1471);
and U6090 (N_6090,N_600,N_2388);
nand U6091 (N_6091,N_856,N_2153);
or U6092 (N_6092,N_1003,N_2621);
and U6093 (N_6093,N_575,N_1049);
and U6094 (N_6094,N_939,N_2548);
nor U6095 (N_6095,N_2163,N_1176);
and U6096 (N_6096,N_2904,N_1874);
nand U6097 (N_6097,N_1167,N_2405);
xor U6098 (N_6098,N_3415,N_3287);
nand U6099 (N_6099,N_907,N_193);
nor U6100 (N_6100,N_2349,N_1691);
nand U6101 (N_6101,N_3071,N_870);
and U6102 (N_6102,N_2211,N_3227);
and U6103 (N_6103,N_1159,N_1271);
and U6104 (N_6104,N_1253,N_3524);
xnor U6105 (N_6105,N_1065,N_3374);
and U6106 (N_6106,N_1276,N_2353);
nand U6107 (N_6107,N_1837,N_754);
nand U6108 (N_6108,N_3067,N_3886);
nand U6109 (N_6109,N_1531,N_3306);
nand U6110 (N_6110,N_1752,N_2722);
and U6111 (N_6111,N_24,N_917);
xnor U6112 (N_6112,N_2900,N_2908);
and U6113 (N_6113,N_2386,N_2846);
or U6114 (N_6114,N_1408,N_2397);
and U6115 (N_6115,N_2122,N_1317);
nand U6116 (N_6116,N_3386,N_1716);
or U6117 (N_6117,N_1283,N_42);
xnor U6118 (N_6118,N_3561,N_3512);
xnor U6119 (N_6119,N_130,N_3301);
or U6120 (N_6120,N_2423,N_2071);
and U6121 (N_6121,N_3022,N_1694);
and U6122 (N_6122,N_3708,N_2930);
nand U6123 (N_6123,N_650,N_397);
nand U6124 (N_6124,N_2924,N_840);
or U6125 (N_6125,N_2716,N_1139);
and U6126 (N_6126,N_387,N_2734);
and U6127 (N_6127,N_1822,N_2131);
nor U6128 (N_6128,N_1622,N_3691);
nor U6129 (N_6129,N_2920,N_3128);
nor U6130 (N_6130,N_2965,N_1021);
nor U6131 (N_6131,N_1794,N_2690);
or U6132 (N_6132,N_3289,N_3790);
or U6133 (N_6133,N_1232,N_159);
and U6134 (N_6134,N_514,N_2806);
nor U6135 (N_6135,N_769,N_107);
nor U6136 (N_6136,N_3772,N_58);
or U6137 (N_6137,N_3623,N_3977);
and U6138 (N_6138,N_3702,N_2645);
xnor U6139 (N_6139,N_1810,N_1282);
or U6140 (N_6140,N_843,N_2710);
or U6141 (N_6141,N_2845,N_124);
and U6142 (N_6142,N_410,N_2377);
xnor U6143 (N_6143,N_3420,N_261);
nand U6144 (N_6144,N_2740,N_1706);
nor U6145 (N_6145,N_3360,N_3277);
xor U6146 (N_6146,N_2505,N_988);
xnor U6147 (N_6147,N_776,N_3517);
and U6148 (N_6148,N_3156,N_3757);
nor U6149 (N_6149,N_3152,N_2751);
or U6150 (N_6150,N_3723,N_2985);
nor U6151 (N_6151,N_2845,N_2650);
or U6152 (N_6152,N_2394,N_1699);
xor U6153 (N_6153,N_2605,N_497);
or U6154 (N_6154,N_21,N_2358);
and U6155 (N_6155,N_0,N_820);
or U6156 (N_6156,N_524,N_3157);
and U6157 (N_6157,N_598,N_1425);
or U6158 (N_6158,N_3843,N_2996);
nand U6159 (N_6159,N_1742,N_3489);
xnor U6160 (N_6160,N_2920,N_2925);
or U6161 (N_6161,N_405,N_3225);
nor U6162 (N_6162,N_3032,N_2064);
or U6163 (N_6163,N_2420,N_2736);
nand U6164 (N_6164,N_633,N_3542);
and U6165 (N_6165,N_1209,N_61);
and U6166 (N_6166,N_155,N_3587);
nand U6167 (N_6167,N_1151,N_925);
or U6168 (N_6168,N_2362,N_2759);
or U6169 (N_6169,N_1280,N_2793);
nor U6170 (N_6170,N_2758,N_1695);
and U6171 (N_6171,N_3676,N_651);
or U6172 (N_6172,N_802,N_168);
or U6173 (N_6173,N_2494,N_2929);
nor U6174 (N_6174,N_3065,N_2935);
nand U6175 (N_6175,N_1559,N_3932);
nand U6176 (N_6176,N_2732,N_3821);
nor U6177 (N_6177,N_784,N_1194);
nand U6178 (N_6178,N_1065,N_76);
nor U6179 (N_6179,N_2017,N_3721);
nand U6180 (N_6180,N_2601,N_3563);
nand U6181 (N_6181,N_428,N_2464);
and U6182 (N_6182,N_354,N_1692);
and U6183 (N_6183,N_1562,N_3864);
and U6184 (N_6184,N_3504,N_1429);
and U6185 (N_6185,N_2876,N_2593);
nand U6186 (N_6186,N_1478,N_1747);
and U6187 (N_6187,N_1820,N_3570);
nor U6188 (N_6188,N_2773,N_997);
or U6189 (N_6189,N_3043,N_1750);
nand U6190 (N_6190,N_2828,N_2781);
nor U6191 (N_6191,N_776,N_1824);
nand U6192 (N_6192,N_1651,N_2646);
nand U6193 (N_6193,N_419,N_1471);
and U6194 (N_6194,N_1017,N_3057);
nand U6195 (N_6195,N_3728,N_1878);
nor U6196 (N_6196,N_1655,N_916);
and U6197 (N_6197,N_1433,N_3233);
or U6198 (N_6198,N_987,N_3586);
nor U6199 (N_6199,N_1809,N_245);
and U6200 (N_6200,N_1212,N_2265);
and U6201 (N_6201,N_2621,N_1489);
and U6202 (N_6202,N_257,N_1730);
nor U6203 (N_6203,N_1624,N_2832);
nor U6204 (N_6204,N_1193,N_52);
nand U6205 (N_6205,N_780,N_2996);
and U6206 (N_6206,N_193,N_2950);
nand U6207 (N_6207,N_3282,N_50);
or U6208 (N_6208,N_3212,N_3749);
or U6209 (N_6209,N_1429,N_7);
nor U6210 (N_6210,N_371,N_2931);
nor U6211 (N_6211,N_123,N_2374);
or U6212 (N_6212,N_3843,N_3012);
and U6213 (N_6213,N_372,N_2083);
or U6214 (N_6214,N_840,N_2782);
xor U6215 (N_6215,N_2612,N_3263);
nand U6216 (N_6216,N_3116,N_1574);
nand U6217 (N_6217,N_679,N_1786);
nand U6218 (N_6218,N_1209,N_3712);
and U6219 (N_6219,N_2767,N_1667);
and U6220 (N_6220,N_478,N_794);
nand U6221 (N_6221,N_1669,N_1635);
nor U6222 (N_6222,N_2568,N_3691);
and U6223 (N_6223,N_1408,N_2133);
and U6224 (N_6224,N_2010,N_2131);
or U6225 (N_6225,N_802,N_2607);
nor U6226 (N_6226,N_2290,N_1515);
and U6227 (N_6227,N_525,N_2875);
nor U6228 (N_6228,N_114,N_2377);
nand U6229 (N_6229,N_3294,N_3789);
and U6230 (N_6230,N_3749,N_2712);
nor U6231 (N_6231,N_2312,N_2612);
or U6232 (N_6232,N_2561,N_534);
or U6233 (N_6233,N_627,N_3458);
or U6234 (N_6234,N_959,N_1118);
and U6235 (N_6235,N_3356,N_3528);
nor U6236 (N_6236,N_1818,N_878);
and U6237 (N_6237,N_1606,N_461);
or U6238 (N_6238,N_3663,N_2418);
or U6239 (N_6239,N_3356,N_2552);
xor U6240 (N_6240,N_1768,N_638);
nor U6241 (N_6241,N_490,N_720);
or U6242 (N_6242,N_2101,N_3090);
nor U6243 (N_6243,N_1121,N_1126);
and U6244 (N_6244,N_3426,N_1040);
xor U6245 (N_6245,N_1441,N_603);
and U6246 (N_6246,N_936,N_2658);
nand U6247 (N_6247,N_3633,N_1732);
nor U6248 (N_6248,N_78,N_2982);
xnor U6249 (N_6249,N_435,N_1134);
nor U6250 (N_6250,N_2020,N_0);
nand U6251 (N_6251,N_3948,N_340);
nand U6252 (N_6252,N_765,N_1869);
nor U6253 (N_6253,N_3109,N_1806);
nor U6254 (N_6254,N_690,N_1380);
or U6255 (N_6255,N_2453,N_1268);
or U6256 (N_6256,N_1452,N_3289);
nor U6257 (N_6257,N_2860,N_2977);
xnor U6258 (N_6258,N_3588,N_2110);
and U6259 (N_6259,N_3202,N_1984);
or U6260 (N_6260,N_2086,N_1096);
nand U6261 (N_6261,N_3217,N_746);
nor U6262 (N_6262,N_3198,N_3480);
nand U6263 (N_6263,N_316,N_539);
nor U6264 (N_6264,N_2892,N_1104);
nor U6265 (N_6265,N_1946,N_1816);
or U6266 (N_6266,N_1469,N_276);
nand U6267 (N_6267,N_2523,N_3255);
nand U6268 (N_6268,N_672,N_1946);
and U6269 (N_6269,N_2619,N_2137);
nand U6270 (N_6270,N_2032,N_511);
and U6271 (N_6271,N_3812,N_1613);
and U6272 (N_6272,N_212,N_1224);
or U6273 (N_6273,N_2959,N_3208);
and U6274 (N_6274,N_1723,N_3885);
nor U6275 (N_6275,N_3568,N_2972);
and U6276 (N_6276,N_2777,N_1336);
nand U6277 (N_6277,N_2569,N_2750);
xor U6278 (N_6278,N_3128,N_1153);
nand U6279 (N_6279,N_2057,N_1788);
or U6280 (N_6280,N_3672,N_529);
and U6281 (N_6281,N_2165,N_2101);
nor U6282 (N_6282,N_2117,N_2503);
nand U6283 (N_6283,N_862,N_1750);
and U6284 (N_6284,N_2525,N_1486);
or U6285 (N_6285,N_675,N_1020);
nand U6286 (N_6286,N_2074,N_2042);
nand U6287 (N_6287,N_1,N_3358);
or U6288 (N_6288,N_2633,N_2421);
or U6289 (N_6289,N_571,N_2446);
and U6290 (N_6290,N_435,N_3925);
or U6291 (N_6291,N_1519,N_3185);
or U6292 (N_6292,N_590,N_783);
nand U6293 (N_6293,N_3421,N_1160);
nand U6294 (N_6294,N_1572,N_1125);
nor U6295 (N_6295,N_2951,N_17);
nor U6296 (N_6296,N_2600,N_833);
nand U6297 (N_6297,N_2776,N_3871);
nand U6298 (N_6298,N_2480,N_343);
nand U6299 (N_6299,N_2183,N_52);
or U6300 (N_6300,N_889,N_3881);
nor U6301 (N_6301,N_2590,N_513);
or U6302 (N_6302,N_3646,N_1523);
nand U6303 (N_6303,N_818,N_2123);
or U6304 (N_6304,N_3371,N_3237);
nor U6305 (N_6305,N_884,N_3556);
nor U6306 (N_6306,N_3249,N_2182);
or U6307 (N_6307,N_3485,N_571);
xor U6308 (N_6308,N_3974,N_338);
and U6309 (N_6309,N_3105,N_548);
or U6310 (N_6310,N_3269,N_2116);
xor U6311 (N_6311,N_2552,N_2684);
nor U6312 (N_6312,N_3156,N_2055);
nand U6313 (N_6313,N_65,N_363);
and U6314 (N_6314,N_3779,N_3418);
xor U6315 (N_6315,N_3858,N_3182);
nand U6316 (N_6316,N_2695,N_2546);
or U6317 (N_6317,N_3480,N_3745);
or U6318 (N_6318,N_3399,N_1628);
xor U6319 (N_6319,N_268,N_1939);
or U6320 (N_6320,N_3506,N_2887);
or U6321 (N_6321,N_1374,N_1587);
and U6322 (N_6322,N_3027,N_1714);
or U6323 (N_6323,N_1216,N_3018);
nor U6324 (N_6324,N_1167,N_337);
xnor U6325 (N_6325,N_2747,N_1498);
xor U6326 (N_6326,N_3170,N_1811);
nor U6327 (N_6327,N_1534,N_2566);
xor U6328 (N_6328,N_573,N_255);
nor U6329 (N_6329,N_314,N_943);
nor U6330 (N_6330,N_1652,N_392);
or U6331 (N_6331,N_2189,N_1123);
or U6332 (N_6332,N_2354,N_3602);
xor U6333 (N_6333,N_2339,N_3700);
and U6334 (N_6334,N_2157,N_2519);
and U6335 (N_6335,N_505,N_3632);
and U6336 (N_6336,N_3912,N_79);
and U6337 (N_6337,N_3572,N_2715);
nor U6338 (N_6338,N_3153,N_852);
nand U6339 (N_6339,N_2087,N_3131);
nor U6340 (N_6340,N_240,N_2375);
or U6341 (N_6341,N_44,N_1663);
and U6342 (N_6342,N_1571,N_492);
and U6343 (N_6343,N_941,N_2709);
or U6344 (N_6344,N_751,N_1967);
and U6345 (N_6345,N_885,N_684);
nand U6346 (N_6346,N_3620,N_546);
nand U6347 (N_6347,N_1646,N_3883);
or U6348 (N_6348,N_346,N_967);
xor U6349 (N_6349,N_153,N_1107);
nor U6350 (N_6350,N_2319,N_464);
nand U6351 (N_6351,N_450,N_16);
or U6352 (N_6352,N_822,N_2085);
nor U6353 (N_6353,N_3091,N_2569);
and U6354 (N_6354,N_2337,N_2620);
nor U6355 (N_6355,N_1805,N_1749);
nand U6356 (N_6356,N_3291,N_1031);
and U6357 (N_6357,N_3932,N_155);
nand U6358 (N_6358,N_1151,N_2064);
nand U6359 (N_6359,N_2613,N_3467);
nand U6360 (N_6360,N_565,N_915);
and U6361 (N_6361,N_1454,N_660);
nor U6362 (N_6362,N_303,N_3422);
nand U6363 (N_6363,N_3607,N_80);
or U6364 (N_6364,N_1800,N_3600);
nand U6365 (N_6365,N_3873,N_587);
or U6366 (N_6366,N_1121,N_3690);
nor U6367 (N_6367,N_1967,N_802);
nor U6368 (N_6368,N_3225,N_207);
nand U6369 (N_6369,N_2797,N_1414);
and U6370 (N_6370,N_3617,N_85);
nor U6371 (N_6371,N_757,N_1409);
nand U6372 (N_6372,N_3573,N_3262);
or U6373 (N_6373,N_3518,N_1719);
nand U6374 (N_6374,N_538,N_2774);
or U6375 (N_6375,N_2751,N_2335);
nor U6376 (N_6376,N_602,N_1931);
or U6377 (N_6377,N_2901,N_3293);
and U6378 (N_6378,N_2201,N_3344);
or U6379 (N_6379,N_3100,N_2464);
and U6380 (N_6380,N_1818,N_3092);
or U6381 (N_6381,N_898,N_3085);
xnor U6382 (N_6382,N_2709,N_3923);
nor U6383 (N_6383,N_568,N_3130);
or U6384 (N_6384,N_482,N_1274);
or U6385 (N_6385,N_1711,N_1404);
and U6386 (N_6386,N_957,N_3317);
nand U6387 (N_6387,N_2705,N_384);
nor U6388 (N_6388,N_3672,N_1145);
and U6389 (N_6389,N_543,N_3378);
and U6390 (N_6390,N_3541,N_241);
nor U6391 (N_6391,N_1103,N_3304);
nand U6392 (N_6392,N_3139,N_2300);
nand U6393 (N_6393,N_189,N_7);
xnor U6394 (N_6394,N_2680,N_380);
or U6395 (N_6395,N_2710,N_2061);
nor U6396 (N_6396,N_304,N_2470);
and U6397 (N_6397,N_3066,N_3035);
or U6398 (N_6398,N_3419,N_1245);
nand U6399 (N_6399,N_3513,N_2227);
and U6400 (N_6400,N_1697,N_419);
or U6401 (N_6401,N_1457,N_2500);
nor U6402 (N_6402,N_2352,N_3126);
nand U6403 (N_6403,N_3487,N_2045);
and U6404 (N_6404,N_2171,N_3960);
nor U6405 (N_6405,N_2735,N_1230);
or U6406 (N_6406,N_550,N_493);
or U6407 (N_6407,N_1152,N_666);
and U6408 (N_6408,N_1660,N_1063);
nor U6409 (N_6409,N_3585,N_1422);
nand U6410 (N_6410,N_1546,N_2775);
nand U6411 (N_6411,N_1287,N_1665);
nand U6412 (N_6412,N_476,N_1000);
nor U6413 (N_6413,N_1657,N_2007);
or U6414 (N_6414,N_3310,N_912);
xnor U6415 (N_6415,N_2131,N_851);
or U6416 (N_6416,N_1942,N_684);
and U6417 (N_6417,N_3525,N_1962);
nor U6418 (N_6418,N_2739,N_3079);
nand U6419 (N_6419,N_324,N_674);
nor U6420 (N_6420,N_121,N_3003);
and U6421 (N_6421,N_329,N_2291);
and U6422 (N_6422,N_3546,N_1703);
nor U6423 (N_6423,N_2309,N_1774);
and U6424 (N_6424,N_35,N_1572);
xnor U6425 (N_6425,N_863,N_2727);
nand U6426 (N_6426,N_2098,N_1352);
and U6427 (N_6427,N_2794,N_43);
or U6428 (N_6428,N_2811,N_156);
or U6429 (N_6429,N_3760,N_1189);
or U6430 (N_6430,N_869,N_1029);
or U6431 (N_6431,N_508,N_3169);
nor U6432 (N_6432,N_3777,N_2334);
and U6433 (N_6433,N_1780,N_1534);
xor U6434 (N_6434,N_2929,N_1104);
or U6435 (N_6435,N_2402,N_1299);
or U6436 (N_6436,N_1044,N_3055);
or U6437 (N_6437,N_3375,N_2487);
nor U6438 (N_6438,N_851,N_726);
nand U6439 (N_6439,N_3207,N_1824);
nor U6440 (N_6440,N_2555,N_1993);
nand U6441 (N_6441,N_720,N_3239);
or U6442 (N_6442,N_3118,N_886);
or U6443 (N_6443,N_1494,N_2439);
nand U6444 (N_6444,N_2428,N_1006);
and U6445 (N_6445,N_150,N_2735);
and U6446 (N_6446,N_3122,N_3722);
and U6447 (N_6447,N_2425,N_2901);
nor U6448 (N_6448,N_1887,N_2080);
or U6449 (N_6449,N_683,N_1891);
nor U6450 (N_6450,N_748,N_3602);
nand U6451 (N_6451,N_2545,N_2272);
nor U6452 (N_6452,N_3445,N_1968);
or U6453 (N_6453,N_2083,N_455);
nor U6454 (N_6454,N_2744,N_3727);
nand U6455 (N_6455,N_2425,N_834);
nor U6456 (N_6456,N_1170,N_2486);
xnor U6457 (N_6457,N_1131,N_1985);
xor U6458 (N_6458,N_807,N_3155);
nand U6459 (N_6459,N_1330,N_1771);
and U6460 (N_6460,N_2108,N_3747);
nand U6461 (N_6461,N_2993,N_921);
and U6462 (N_6462,N_2814,N_3097);
xor U6463 (N_6463,N_724,N_3071);
nand U6464 (N_6464,N_434,N_2899);
nor U6465 (N_6465,N_1445,N_3405);
or U6466 (N_6466,N_1781,N_2662);
nor U6467 (N_6467,N_3931,N_1310);
xnor U6468 (N_6468,N_744,N_3407);
nand U6469 (N_6469,N_2606,N_1120);
nor U6470 (N_6470,N_1655,N_3458);
and U6471 (N_6471,N_967,N_3311);
or U6472 (N_6472,N_529,N_1379);
nand U6473 (N_6473,N_313,N_2676);
nor U6474 (N_6474,N_824,N_1551);
nor U6475 (N_6475,N_2285,N_666);
or U6476 (N_6476,N_2910,N_188);
or U6477 (N_6477,N_665,N_2310);
xor U6478 (N_6478,N_1025,N_2058);
or U6479 (N_6479,N_1527,N_2067);
or U6480 (N_6480,N_3545,N_3695);
and U6481 (N_6481,N_3506,N_1078);
and U6482 (N_6482,N_777,N_2766);
or U6483 (N_6483,N_3659,N_1111);
or U6484 (N_6484,N_3463,N_769);
nand U6485 (N_6485,N_1222,N_1418);
nor U6486 (N_6486,N_3458,N_726);
or U6487 (N_6487,N_2866,N_1176);
nand U6488 (N_6488,N_3089,N_626);
nor U6489 (N_6489,N_1959,N_2647);
nand U6490 (N_6490,N_2131,N_790);
nand U6491 (N_6491,N_1571,N_2610);
nor U6492 (N_6492,N_1656,N_718);
nand U6493 (N_6493,N_3886,N_2223);
nor U6494 (N_6494,N_746,N_3788);
nor U6495 (N_6495,N_2612,N_2559);
or U6496 (N_6496,N_114,N_3116);
nor U6497 (N_6497,N_2288,N_3233);
and U6498 (N_6498,N_2804,N_3511);
nand U6499 (N_6499,N_1779,N_1175);
xnor U6500 (N_6500,N_3384,N_562);
and U6501 (N_6501,N_2470,N_1427);
or U6502 (N_6502,N_285,N_1063);
nand U6503 (N_6503,N_3548,N_323);
nor U6504 (N_6504,N_381,N_124);
and U6505 (N_6505,N_925,N_3683);
xor U6506 (N_6506,N_2461,N_2127);
nor U6507 (N_6507,N_3102,N_2080);
nand U6508 (N_6508,N_1289,N_2735);
and U6509 (N_6509,N_3140,N_3259);
or U6510 (N_6510,N_461,N_1018);
and U6511 (N_6511,N_3601,N_2593);
nor U6512 (N_6512,N_1370,N_2332);
and U6513 (N_6513,N_2681,N_3443);
nand U6514 (N_6514,N_1405,N_1413);
or U6515 (N_6515,N_3496,N_1283);
nor U6516 (N_6516,N_762,N_143);
nand U6517 (N_6517,N_1435,N_985);
nor U6518 (N_6518,N_1414,N_3382);
nor U6519 (N_6519,N_3337,N_1812);
nor U6520 (N_6520,N_1018,N_1964);
or U6521 (N_6521,N_1347,N_2433);
nand U6522 (N_6522,N_1984,N_3180);
xor U6523 (N_6523,N_1404,N_2995);
or U6524 (N_6524,N_2477,N_1770);
and U6525 (N_6525,N_3264,N_202);
and U6526 (N_6526,N_2662,N_90);
nand U6527 (N_6527,N_1159,N_1187);
and U6528 (N_6528,N_2840,N_1140);
xor U6529 (N_6529,N_3018,N_3568);
or U6530 (N_6530,N_251,N_668);
nor U6531 (N_6531,N_1255,N_745);
nand U6532 (N_6532,N_1573,N_998);
nand U6533 (N_6533,N_2544,N_1772);
and U6534 (N_6534,N_932,N_1730);
nand U6535 (N_6535,N_1346,N_3622);
or U6536 (N_6536,N_3178,N_2253);
and U6537 (N_6537,N_3392,N_3718);
nor U6538 (N_6538,N_3168,N_2699);
or U6539 (N_6539,N_2903,N_547);
nor U6540 (N_6540,N_2545,N_1040);
or U6541 (N_6541,N_1410,N_859);
nor U6542 (N_6542,N_2886,N_968);
and U6543 (N_6543,N_3354,N_2852);
nand U6544 (N_6544,N_2346,N_3975);
or U6545 (N_6545,N_3044,N_2481);
xor U6546 (N_6546,N_3086,N_2102);
or U6547 (N_6547,N_1838,N_355);
or U6548 (N_6548,N_1011,N_3487);
nand U6549 (N_6549,N_2710,N_984);
nand U6550 (N_6550,N_2270,N_50);
or U6551 (N_6551,N_2447,N_3377);
nor U6552 (N_6552,N_384,N_3315);
nand U6553 (N_6553,N_2563,N_2918);
nand U6554 (N_6554,N_1820,N_261);
or U6555 (N_6555,N_691,N_153);
or U6556 (N_6556,N_2833,N_3466);
nand U6557 (N_6557,N_3558,N_3863);
and U6558 (N_6558,N_989,N_1325);
or U6559 (N_6559,N_3241,N_1567);
nor U6560 (N_6560,N_3477,N_676);
and U6561 (N_6561,N_1068,N_2035);
and U6562 (N_6562,N_1752,N_1445);
nor U6563 (N_6563,N_3442,N_1201);
or U6564 (N_6564,N_1432,N_374);
nand U6565 (N_6565,N_2308,N_1051);
or U6566 (N_6566,N_518,N_3197);
nand U6567 (N_6567,N_2453,N_1428);
and U6568 (N_6568,N_2639,N_3861);
xnor U6569 (N_6569,N_381,N_2456);
and U6570 (N_6570,N_2422,N_3329);
nor U6571 (N_6571,N_3405,N_3279);
or U6572 (N_6572,N_2395,N_1665);
nand U6573 (N_6573,N_2167,N_1307);
xor U6574 (N_6574,N_3785,N_1460);
or U6575 (N_6575,N_3693,N_3811);
xor U6576 (N_6576,N_1824,N_1130);
nand U6577 (N_6577,N_3827,N_3166);
nor U6578 (N_6578,N_3545,N_530);
nand U6579 (N_6579,N_3563,N_3161);
or U6580 (N_6580,N_1002,N_1933);
and U6581 (N_6581,N_2879,N_810);
nor U6582 (N_6582,N_3953,N_2571);
and U6583 (N_6583,N_3656,N_2548);
and U6584 (N_6584,N_3458,N_2207);
or U6585 (N_6585,N_40,N_3637);
nand U6586 (N_6586,N_2210,N_2381);
and U6587 (N_6587,N_1021,N_2306);
nor U6588 (N_6588,N_1852,N_2955);
nor U6589 (N_6589,N_3750,N_2680);
nor U6590 (N_6590,N_1082,N_791);
and U6591 (N_6591,N_2692,N_848);
and U6592 (N_6592,N_2823,N_3885);
or U6593 (N_6593,N_2779,N_520);
or U6594 (N_6594,N_1267,N_2930);
nor U6595 (N_6595,N_1550,N_3064);
and U6596 (N_6596,N_1404,N_568);
nor U6597 (N_6597,N_456,N_965);
nand U6598 (N_6598,N_2699,N_1013);
nand U6599 (N_6599,N_2130,N_2740);
nand U6600 (N_6600,N_1207,N_987);
nand U6601 (N_6601,N_287,N_2146);
and U6602 (N_6602,N_3124,N_3279);
nor U6603 (N_6603,N_1090,N_2514);
or U6604 (N_6604,N_2436,N_914);
nand U6605 (N_6605,N_3058,N_2700);
and U6606 (N_6606,N_2421,N_1725);
nor U6607 (N_6607,N_3241,N_2958);
and U6608 (N_6608,N_3936,N_881);
xor U6609 (N_6609,N_1870,N_3249);
and U6610 (N_6610,N_1133,N_1490);
and U6611 (N_6611,N_3572,N_1314);
and U6612 (N_6612,N_399,N_1202);
and U6613 (N_6613,N_183,N_1970);
and U6614 (N_6614,N_3982,N_2686);
nor U6615 (N_6615,N_1880,N_3040);
nor U6616 (N_6616,N_583,N_2297);
nand U6617 (N_6617,N_3159,N_939);
and U6618 (N_6618,N_3203,N_346);
nor U6619 (N_6619,N_2045,N_1565);
or U6620 (N_6620,N_2429,N_3512);
xor U6621 (N_6621,N_3731,N_1600);
nor U6622 (N_6622,N_2549,N_67);
or U6623 (N_6623,N_1381,N_2007);
nand U6624 (N_6624,N_1943,N_299);
or U6625 (N_6625,N_1756,N_3820);
nand U6626 (N_6626,N_1204,N_246);
and U6627 (N_6627,N_806,N_407);
or U6628 (N_6628,N_1463,N_833);
nand U6629 (N_6629,N_106,N_1327);
nand U6630 (N_6630,N_1779,N_1492);
nand U6631 (N_6631,N_298,N_1961);
and U6632 (N_6632,N_2317,N_2521);
nand U6633 (N_6633,N_3708,N_1278);
or U6634 (N_6634,N_3007,N_2101);
xnor U6635 (N_6635,N_487,N_950);
nor U6636 (N_6636,N_251,N_3613);
xor U6637 (N_6637,N_2074,N_3195);
or U6638 (N_6638,N_2684,N_2282);
nand U6639 (N_6639,N_55,N_2317);
or U6640 (N_6640,N_832,N_3429);
or U6641 (N_6641,N_2413,N_3528);
nor U6642 (N_6642,N_808,N_1655);
nand U6643 (N_6643,N_3989,N_556);
nor U6644 (N_6644,N_1745,N_722);
or U6645 (N_6645,N_255,N_3323);
or U6646 (N_6646,N_3665,N_3432);
or U6647 (N_6647,N_3807,N_298);
or U6648 (N_6648,N_37,N_3060);
nor U6649 (N_6649,N_3863,N_1070);
or U6650 (N_6650,N_956,N_754);
and U6651 (N_6651,N_834,N_1723);
or U6652 (N_6652,N_2219,N_2848);
and U6653 (N_6653,N_3707,N_1047);
or U6654 (N_6654,N_1099,N_1997);
or U6655 (N_6655,N_2030,N_2647);
or U6656 (N_6656,N_507,N_2084);
or U6657 (N_6657,N_437,N_991);
and U6658 (N_6658,N_2380,N_1343);
nand U6659 (N_6659,N_1990,N_1342);
or U6660 (N_6660,N_1311,N_2562);
and U6661 (N_6661,N_1225,N_1530);
nand U6662 (N_6662,N_2297,N_1260);
nor U6663 (N_6663,N_913,N_3939);
or U6664 (N_6664,N_3829,N_1904);
or U6665 (N_6665,N_2348,N_2976);
nand U6666 (N_6666,N_2681,N_2213);
nor U6667 (N_6667,N_2811,N_2543);
and U6668 (N_6668,N_3113,N_50);
and U6669 (N_6669,N_656,N_40);
or U6670 (N_6670,N_3462,N_640);
and U6671 (N_6671,N_2665,N_3869);
or U6672 (N_6672,N_504,N_3954);
or U6673 (N_6673,N_3212,N_1257);
nor U6674 (N_6674,N_2042,N_3729);
or U6675 (N_6675,N_919,N_2171);
and U6676 (N_6676,N_3341,N_2971);
xnor U6677 (N_6677,N_1169,N_742);
xnor U6678 (N_6678,N_1165,N_1461);
nand U6679 (N_6679,N_3773,N_535);
nor U6680 (N_6680,N_485,N_2938);
nor U6681 (N_6681,N_1608,N_2848);
nor U6682 (N_6682,N_3978,N_320);
nor U6683 (N_6683,N_1010,N_3615);
and U6684 (N_6684,N_1403,N_2495);
nand U6685 (N_6685,N_864,N_2146);
and U6686 (N_6686,N_798,N_1228);
or U6687 (N_6687,N_981,N_1621);
and U6688 (N_6688,N_1552,N_76);
nand U6689 (N_6689,N_1874,N_415);
and U6690 (N_6690,N_228,N_2754);
or U6691 (N_6691,N_1761,N_1463);
or U6692 (N_6692,N_1771,N_2664);
or U6693 (N_6693,N_3086,N_201);
or U6694 (N_6694,N_1303,N_170);
nor U6695 (N_6695,N_49,N_1149);
xnor U6696 (N_6696,N_1841,N_835);
nor U6697 (N_6697,N_3751,N_3816);
nand U6698 (N_6698,N_1142,N_1208);
nand U6699 (N_6699,N_3435,N_3207);
nand U6700 (N_6700,N_3184,N_717);
or U6701 (N_6701,N_2538,N_189);
nor U6702 (N_6702,N_2769,N_100);
or U6703 (N_6703,N_2260,N_313);
or U6704 (N_6704,N_956,N_3082);
xnor U6705 (N_6705,N_3196,N_1944);
xnor U6706 (N_6706,N_1381,N_3717);
and U6707 (N_6707,N_598,N_1147);
nand U6708 (N_6708,N_1736,N_444);
nor U6709 (N_6709,N_1374,N_566);
nand U6710 (N_6710,N_3969,N_2204);
xor U6711 (N_6711,N_1639,N_1975);
nand U6712 (N_6712,N_1293,N_3003);
or U6713 (N_6713,N_3098,N_815);
or U6714 (N_6714,N_2098,N_2013);
and U6715 (N_6715,N_1075,N_353);
or U6716 (N_6716,N_2416,N_3620);
or U6717 (N_6717,N_969,N_3633);
nand U6718 (N_6718,N_3261,N_3997);
and U6719 (N_6719,N_3428,N_2602);
nand U6720 (N_6720,N_585,N_610);
and U6721 (N_6721,N_155,N_3087);
nand U6722 (N_6722,N_2886,N_2777);
and U6723 (N_6723,N_2573,N_348);
or U6724 (N_6724,N_1896,N_2475);
nor U6725 (N_6725,N_1708,N_2863);
or U6726 (N_6726,N_865,N_1656);
and U6727 (N_6727,N_1785,N_303);
nand U6728 (N_6728,N_1727,N_2459);
xor U6729 (N_6729,N_1659,N_2002);
nand U6730 (N_6730,N_442,N_1937);
nand U6731 (N_6731,N_1856,N_2182);
nor U6732 (N_6732,N_1834,N_3657);
and U6733 (N_6733,N_1923,N_1443);
or U6734 (N_6734,N_2767,N_2386);
nor U6735 (N_6735,N_1317,N_3919);
and U6736 (N_6736,N_1617,N_201);
or U6737 (N_6737,N_3126,N_2993);
nor U6738 (N_6738,N_3514,N_2989);
xnor U6739 (N_6739,N_1830,N_1703);
and U6740 (N_6740,N_680,N_3076);
and U6741 (N_6741,N_1591,N_3846);
nand U6742 (N_6742,N_1893,N_983);
or U6743 (N_6743,N_304,N_2902);
nor U6744 (N_6744,N_1856,N_1466);
and U6745 (N_6745,N_3261,N_2809);
nand U6746 (N_6746,N_151,N_86);
and U6747 (N_6747,N_2449,N_1001);
and U6748 (N_6748,N_52,N_2799);
nand U6749 (N_6749,N_2139,N_776);
and U6750 (N_6750,N_2395,N_427);
or U6751 (N_6751,N_2978,N_3752);
nor U6752 (N_6752,N_193,N_1973);
nor U6753 (N_6753,N_1975,N_1822);
nor U6754 (N_6754,N_45,N_1766);
nor U6755 (N_6755,N_2427,N_3980);
and U6756 (N_6756,N_3339,N_2409);
and U6757 (N_6757,N_1196,N_2283);
or U6758 (N_6758,N_3438,N_156);
nand U6759 (N_6759,N_3965,N_1001);
and U6760 (N_6760,N_2802,N_3329);
or U6761 (N_6761,N_3611,N_2078);
xnor U6762 (N_6762,N_927,N_2320);
nand U6763 (N_6763,N_486,N_3234);
nand U6764 (N_6764,N_3530,N_764);
and U6765 (N_6765,N_3906,N_3063);
and U6766 (N_6766,N_1023,N_711);
nand U6767 (N_6767,N_1606,N_1687);
xnor U6768 (N_6768,N_2049,N_2584);
nor U6769 (N_6769,N_1382,N_3254);
and U6770 (N_6770,N_2002,N_181);
nand U6771 (N_6771,N_1786,N_2332);
or U6772 (N_6772,N_3592,N_608);
nand U6773 (N_6773,N_977,N_69);
nand U6774 (N_6774,N_2235,N_2046);
or U6775 (N_6775,N_2975,N_1167);
and U6776 (N_6776,N_1236,N_3726);
xor U6777 (N_6777,N_3593,N_2596);
or U6778 (N_6778,N_49,N_1226);
nor U6779 (N_6779,N_2681,N_522);
or U6780 (N_6780,N_2411,N_3079);
and U6781 (N_6781,N_2766,N_3874);
xor U6782 (N_6782,N_1276,N_1035);
and U6783 (N_6783,N_2644,N_2942);
and U6784 (N_6784,N_3746,N_2781);
or U6785 (N_6785,N_1684,N_3275);
nand U6786 (N_6786,N_2774,N_2043);
and U6787 (N_6787,N_2033,N_66);
nand U6788 (N_6788,N_2497,N_887);
or U6789 (N_6789,N_388,N_1919);
or U6790 (N_6790,N_572,N_3788);
nand U6791 (N_6791,N_1710,N_751);
nor U6792 (N_6792,N_1635,N_1856);
or U6793 (N_6793,N_1115,N_2628);
nor U6794 (N_6794,N_1695,N_3621);
nand U6795 (N_6795,N_3531,N_1494);
and U6796 (N_6796,N_2257,N_842);
nand U6797 (N_6797,N_2295,N_2559);
and U6798 (N_6798,N_1591,N_2820);
and U6799 (N_6799,N_2719,N_889);
nor U6800 (N_6800,N_980,N_3197);
nand U6801 (N_6801,N_3300,N_2402);
or U6802 (N_6802,N_2898,N_1321);
and U6803 (N_6803,N_1983,N_2393);
xnor U6804 (N_6804,N_3161,N_1110);
nand U6805 (N_6805,N_3823,N_1918);
nand U6806 (N_6806,N_883,N_38);
nand U6807 (N_6807,N_3334,N_3388);
or U6808 (N_6808,N_1622,N_2174);
nand U6809 (N_6809,N_3788,N_696);
nor U6810 (N_6810,N_560,N_691);
nor U6811 (N_6811,N_2086,N_3542);
and U6812 (N_6812,N_3824,N_3432);
nand U6813 (N_6813,N_3772,N_984);
nand U6814 (N_6814,N_2547,N_537);
nand U6815 (N_6815,N_1143,N_866);
or U6816 (N_6816,N_2055,N_3006);
and U6817 (N_6817,N_2845,N_1572);
and U6818 (N_6818,N_2934,N_3590);
nor U6819 (N_6819,N_1276,N_2240);
xor U6820 (N_6820,N_2497,N_1458);
nor U6821 (N_6821,N_1676,N_3679);
nor U6822 (N_6822,N_2615,N_3516);
nand U6823 (N_6823,N_944,N_1906);
nand U6824 (N_6824,N_3072,N_1229);
or U6825 (N_6825,N_356,N_2378);
nor U6826 (N_6826,N_951,N_1924);
and U6827 (N_6827,N_1616,N_986);
xnor U6828 (N_6828,N_1239,N_3266);
nand U6829 (N_6829,N_2578,N_1232);
xnor U6830 (N_6830,N_726,N_1723);
nand U6831 (N_6831,N_456,N_1192);
xor U6832 (N_6832,N_2664,N_1341);
and U6833 (N_6833,N_1902,N_438);
nor U6834 (N_6834,N_1026,N_2110);
nor U6835 (N_6835,N_330,N_680);
nor U6836 (N_6836,N_1181,N_1253);
and U6837 (N_6837,N_3017,N_2041);
nand U6838 (N_6838,N_2618,N_1161);
nor U6839 (N_6839,N_151,N_1655);
nor U6840 (N_6840,N_1060,N_1021);
nor U6841 (N_6841,N_727,N_1416);
and U6842 (N_6842,N_3779,N_1148);
and U6843 (N_6843,N_1803,N_1394);
nor U6844 (N_6844,N_346,N_2096);
or U6845 (N_6845,N_1836,N_323);
nand U6846 (N_6846,N_2455,N_2322);
nor U6847 (N_6847,N_60,N_3829);
nand U6848 (N_6848,N_2077,N_430);
and U6849 (N_6849,N_273,N_2687);
nand U6850 (N_6850,N_1743,N_3612);
and U6851 (N_6851,N_519,N_299);
nand U6852 (N_6852,N_3201,N_2558);
or U6853 (N_6853,N_2659,N_956);
or U6854 (N_6854,N_2693,N_2355);
nor U6855 (N_6855,N_3290,N_1609);
and U6856 (N_6856,N_3498,N_1474);
or U6857 (N_6857,N_1053,N_174);
xnor U6858 (N_6858,N_2738,N_277);
xor U6859 (N_6859,N_3214,N_1666);
nand U6860 (N_6860,N_371,N_1371);
xor U6861 (N_6861,N_3917,N_2488);
xor U6862 (N_6862,N_2834,N_3923);
or U6863 (N_6863,N_423,N_558);
or U6864 (N_6864,N_2814,N_2048);
or U6865 (N_6865,N_1081,N_1778);
xnor U6866 (N_6866,N_2963,N_1488);
and U6867 (N_6867,N_3440,N_631);
nand U6868 (N_6868,N_1523,N_3126);
nor U6869 (N_6869,N_2855,N_1360);
and U6870 (N_6870,N_2287,N_2576);
nand U6871 (N_6871,N_1486,N_1628);
nor U6872 (N_6872,N_3767,N_2439);
or U6873 (N_6873,N_1461,N_1905);
or U6874 (N_6874,N_2106,N_1254);
and U6875 (N_6875,N_2425,N_614);
nand U6876 (N_6876,N_3920,N_1038);
xnor U6877 (N_6877,N_2063,N_3389);
and U6878 (N_6878,N_3512,N_2180);
or U6879 (N_6879,N_516,N_1004);
xor U6880 (N_6880,N_2752,N_2957);
xnor U6881 (N_6881,N_2339,N_1582);
and U6882 (N_6882,N_575,N_1667);
nor U6883 (N_6883,N_2497,N_295);
nor U6884 (N_6884,N_3694,N_1680);
and U6885 (N_6885,N_3982,N_2571);
nand U6886 (N_6886,N_174,N_2385);
nor U6887 (N_6887,N_1944,N_3426);
or U6888 (N_6888,N_1095,N_1167);
or U6889 (N_6889,N_1529,N_1382);
nand U6890 (N_6890,N_3822,N_3288);
and U6891 (N_6891,N_3295,N_689);
xor U6892 (N_6892,N_66,N_2963);
and U6893 (N_6893,N_1555,N_1081);
nand U6894 (N_6894,N_615,N_2630);
or U6895 (N_6895,N_927,N_1717);
and U6896 (N_6896,N_1915,N_59);
xnor U6897 (N_6897,N_1166,N_109);
nand U6898 (N_6898,N_519,N_973);
and U6899 (N_6899,N_1385,N_2241);
and U6900 (N_6900,N_3870,N_3926);
or U6901 (N_6901,N_3015,N_2221);
xnor U6902 (N_6902,N_3417,N_3478);
nand U6903 (N_6903,N_3019,N_3236);
or U6904 (N_6904,N_725,N_3070);
nor U6905 (N_6905,N_1472,N_2641);
and U6906 (N_6906,N_2430,N_1361);
nor U6907 (N_6907,N_1224,N_3808);
xnor U6908 (N_6908,N_2099,N_1535);
or U6909 (N_6909,N_1758,N_732);
or U6910 (N_6910,N_2179,N_2700);
nor U6911 (N_6911,N_450,N_122);
and U6912 (N_6912,N_1633,N_217);
nand U6913 (N_6913,N_594,N_1307);
nor U6914 (N_6914,N_2386,N_993);
or U6915 (N_6915,N_1615,N_2782);
nand U6916 (N_6916,N_2842,N_572);
nor U6917 (N_6917,N_2450,N_705);
xnor U6918 (N_6918,N_1856,N_1507);
or U6919 (N_6919,N_1590,N_959);
or U6920 (N_6920,N_2781,N_3201);
nand U6921 (N_6921,N_1300,N_1050);
and U6922 (N_6922,N_3110,N_630);
or U6923 (N_6923,N_978,N_111);
nand U6924 (N_6924,N_1315,N_65);
nand U6925 (N_6925,N_1388,N_3702);
and U6926 (N_6926,N_1980,N_525);
or U6927 (N_6927,N_1234,N_3364);
or U6928 (N_6928,N_2293,N_977);
nand U6929 (N_6929,N_1925,N_349);
nand U6930 (N_6930,N_1362,N_1580);
and U6931 (N_6931,N_727,N_29);
nand U6932 (N_6932,N_759,N_3823);
and U6933 (N_6933,N_1981,N_486);
or U6934 (N_6934,N_2134,N_592);
nor U6935 (N_6935,N_1025,N_397);
xnor U6936 (N_6936,N_3033,N_861);
and U6937 (N_6937,N_1313,N_1654);
nor U6938 (N_6938,N_2747,N_3885);
nand U6939 (N_6939,N_323,N_3232);
nand U6940 (N_6940,N_243,N_1552);
nor U6941 (N_6941,N_2691,N_1577);
nor U6942 (N_6942,N_3451,N_3610);
nand U6943 (N_6943,N_419,N_2251);
or U6944 (N_6944,N_1933,N_3670);
or U6945 (N_6945,N_3301,N_3984);
nor U6946 (N_6946,N_1843,N_3640);
or U6947 (N_6947,N_434,N_1875);
or U6948 (N_6948,N_2961,N_1470);
and U6949 (N_6949,N_2654,N_1231);
nor U6950 (N_6950,N_3916,N_204);
and U6951 (N_6951,N_2682,N_3861);
xnor U6952 (N_6952,N_1767,N_2909);
nor U6953 (N_6953,N_2397,N_3970);
or U6954 (N_6954,N_1847,N_3775);
xor U6955 (N_6955,N_832,N_1757);
xnor U6956 (N_6956,N_3383,N_227);
nand U6957 (N_6957,N_3194,N_106);
nor U6958 (N_6958,N_3232,N_3271);
xor U6959 (N_6959,N_2311,N_1633);
nand U6960 (N_6960,N_2634,N_2269);
or U6961 (N_6961,N_268,N_397);
xor U6962 (N_6962,N_3214,N_1247);
and U6963 (N_6963,N_140,N_1830);
or U6964 (N_6964,N_1708,N_2810);
nor U6965 (N_6965,N_673,N_300);
nand U6966 (N_6966,N_13,N_1470);
nor U6967 (N_6967,N_3589,N_293);
or U6968 (N_6968,N_2896,N_3192);
and U6969 (N_6969,N_3171,N_1199);
and U6970 (N_6970,N_3264,N_3263);
and U6971 (N_6971,N_1602,N_1697);
nor U6972 (N_6972,N_2959,N_2592);
or U6973 (N_6973,N_3458,N_1819);
and U6974 (N_6974,N_2941,N_1790);
xor U6975 (N_6975,N_2485,N_567);
or U6976 (N_6976,N_3901,N_801);
and U6977 (N_6977,N_2566,N_2666);
nor U6978 (N_6978,N_1213,N_499);
xor U6979 (N_6979,N_3783,N_2525);
nor U6980 (N_6980,N_2819,N_1327);
nor U6981 (N_6981,N_271,N_2159);
nand U6982 (N_6982,N_1353,N_1984);
nand U6983 (N_6983,N_686,N_180);
nor U6984 (N_6984,N_3398,N_2360);
nor U6985 (N_6985,N_683,N_1195);
nand U6986 (N_6986,N_2427,N_3185);
xnor U6987 (N_6987,N_1245,N_1156);
and U6988 (N_6988,N_3296,N_247);
nand U6989 (N_6989,N_3375,N_1);
or U6990 (N_6990,N_3773,N_498);
or U6991 (N_6991,N_3391,N_243);
nor U6992 (N_6992,N_1485,N_2454);
xnor U6993 (N_6993,N_1689,N_1734);
or U6994 (N_6994,N_3536,N_2509);
and U6995 (N_6995,N_3988,N_2765);
and U6996 (N_6996,N_299,N_1908);
nor U6997 (N_6997,N_1079,N_1628);
or U6998 (N_6998,N_2777,N_3271);
xor U6999 (N_6999,N_2266,N_784);
or U7000 (N_7000,N_948,N_3032);
nor U7001 (N_7001,N_3049,N_2009);
or U7002 (N_7002,N_2892,N_668);
and U7003 (N_7003,N_3952,N_2766);
xor U7004 (N_7004,N_1575,N_2269);
or U7005 (N_7005,N_361,N_2431);
and U7006 (N_7006,N_3182,N_1523);
nor U7007 (N_7007,N_761,N_3034);
and U7008 (N_7008,N_3525,N_718);
or U7009 (N_7009,N_2141,N_2795);
nand U7010 (N_7010,N_2170,N_1765);
and U7011 (N_7011,N_520,N_1078);
and U7012 (N_7012,N_2917,N_1174);
or U7013 (N_7013,N_1206,N_358);
or U7014 (N_7014,N_48,N_1437);
or U7015 (N_7015,N_137,N_646);
and U7016 (N_7016,N_3086,N_3046);
and U7017 (N_7017,N_2029,N_2303);
nor U7018 (N_7018,N_396,N_3032);
and U7019 (N_7019,N_1316,N_2024);
nor U7020 (N_7020,N_701,N_3643);
or U7021 (N_7021,N_3012,N_2314);
nor U7022 (N_7022,N_902,N_2396);
or U7023 (N_7023,N_351,N_1514);
nand U7024 (N_7024,N_2396,N_685);
nand U7025 (N_7025,N_1903,N_2114);
and U7026 (N_7026,N_941,N_3234);
and U7027 (N_7027,N_141,N_52);
nand U7028 (N_7028,N_3201,N_591);
and U7029 (N_7029,N_153,N_12);
and U7030 (N_7030,N_3871,N_1769);
nand U7031 (N_7031,N_3853,N_3415);
nor U7032 (N_7032,N_2646,N_185);
nand U7033 (N_7033,N_2507,N_2961);
or U7034 (N_7034,N_3869,N_1534);
and U7035 (N_7035,N_3823,N_3893);
and U7036 (N_7036,N_3887,N_1662);
nor U7037 (N_7037,N_209,N_2662);
nor U7038 (N_7038,N_1722,N_166);
nand U7039 (N_7039,N_3370,N_2236);
and U7040 (N_7040,N_3999,N_3004);
or U7041 (N_7041,N_443,N_1068);
nand U7042 (N_7042,N_2865,N_3676);
or U7043 (N_7043,N_2640,N_2804);
or U7044 (N_7044,N_619,N_638);
or U7045 (N_7045,N_1098,N_3295);
nor U7046 (N_7046,N_405,N_55);
nor U7047 (N_7047,N_3214,N_3719);
nor U7048 (N_7048,N_2212,N_1489);
xor U7049 (N_7049,N_2002,N_1288);
xnor U7050 (N_7050,N_1171,N_40);
nor U7051 (N_7051,N_3997,N_137);
or U7052 (N_7052,N_95,N_1232);
or U7053 (N_7053,N_2534,N_3525);
nor U7054 (N_7054,N_2832,N_7);
nand U7055 (N_7055,N_2029,N_1704);
nand U7056 (N_7056,N_785,N_1500);
and U7057 (N_7057,N_1088,N_2437);
nor U7058 (N_7058,N_1849,N_1341);
or U7059 (N_7059,N_3110,N_1875);
xor U7060 (N_7060,N_3857,N_953);
nor U7061 (N_7061,N_1791,N_3513);
nor U7062 (N_7062,N_527,N_3574);
and U7063 (N_7063,N_2155,N_2205);
nor U7064 (N_7064,N_1533,N_1337);
and U7065 (N_7065,N_1255,N_1205);
or U7066 (N_7066,N_501,N_3321);
and U7067 (N_7067,N_2874,N_3016);
nand U7068 (N_7068,N_2904,N_745);
nor U7069 (N_7069,N_3713,N_2605);
nor U7070 (N_7070,N_359,N_1371);
xor U7071 (N_7071,N_2004,N_2897);
nor U7072 (N_7072,N_3347,N_923);
and U7073 (N_7073,N_3918,N_2122);
nor U7074 (N_7074,N_3660,N_2144);
and U7075 (N_7075,N_2820,N_2422);
nand U7076 (N_7076,N_1455,N_119);
nor U7077 (N_7077,N_2076,N_617);
and U7078 (N_7078,N_929,N_3370);
or U7079 (N_7079,N_3696,N_753);
or U7080 (N_7080,N_1108,N_3125);
nor U7081 (N_7081,N_1181,N_3656);
or U7082 (N_7082,N_3270,N_1848);
nor U7083 (N_7083,N_3980,N_3967);
nor U7084 (N_7084,N_19,N_1475);
and U7085 (N_7085,N_77,N_2526);
nand U7086 (N_7086,N_4,N_1715);
nand U7087 (N_7087,N_1574,N_1846);
or U7088 (N_7088,N_1997,N_2402);
and U7089 (N_7089,N_1489,N_3154);
and U7090 (N_7090,N_2450,N_3526);
or U7091 (N_7091,N_1490,N_1837);
or U7092 (N_7092,N_1565,N_1073);
or U7093 (N_7093,N_1824,N_3112);
nand U7094 (N_7094,N_2924,N_3924);
and U7095 (N_7095,N_1849,N_2165);
or U7096 (N_7096,N_3215,N_3030);
and U7097 (N_7097,N_2547,N_1865);
xor U7098 (N_7098,N_2998,N_467);
and U7099 (N_7099,N_285,N_956);
or U7100 (N_7100,N_465,N_2635);
and U7101 (N_7101,N_3324,N_1481);
or U7102 (N_7102,N_2263,N_2179);
or U7103 (N_7103,N_3171,N_152);
nand U7104 (N_7104,N_993,N_1262);
nor U7105 (N_7105,N_723,N_2607);
xor U7106 (N_7106,N_3775,N_1458);
nand U7107 (N_7107,N_64,N_1869);
or U7108 (N_7108,N_2373,N_664);
nand U7109 (N_7109,N_1705,N_207);
nor U7110 (N_7110,N_636,N_1236);
nor U7111 (N_7111,N_1293,N_2243);
nor U7112 (N_7112,N_1255,N_3947);
or U7113 (N_7113,N_1168,N_2346);
and U7114 (N_7114,N_3825,N_2362);
nor U7115 (N_7115,N_2634,N_3622);
xor U7116 (N_7116,N_2481,N_3296);
nor U7117 (N_7117,N_1705,N_2198);
and U7118 (N_7118,N_2080,N_3642);
nor U7119 (N_7119,N_3915,N_1309);
and U7120 (N_7120,N_754,N_3952);
nor U7121 (N_7121,N_3671,N_874);
or U7122 (N_7122,N_1027,N_342);
xor U7123 (N_7123,N_3261,N_266);
and U7124 (N_7124,N_2432,N_138);
nand U7125 (N_7125,N_2364,N_2480);
and U7126 (N_7126,N_3969,N_1812);
or U7127 (N_7127,N_1294,N_410);
nor U7128 (N_7128,N_3181,N_1020);
and U7129 (N_7129,N_2621,N_3356);
nor U7130 (N_7130,N_3015,N_3114);
xnor U7131 (N_7131,N_2247,N_2472);
nand U7132 (N_7132,N_1005,N_3907);
and U7133 (N_7133,N_656,N_2972);
nor U7134 (N_7134,N_3599,N_3368);
or U7135 (N_7135,N_2496,N_2039);
nor U7136 (N_7136,N_2296,N_1595);
nor U7137 (N_7137,N_3293,N_694);
and U7138 (N_7138,N_2593,N_1563);
or U7139 (N_7139,N_126,N_1311);
nor U7140 (N_7140,N_3451,N_1068);
or U7141 (N_7141,N_2165,N_304);
or U7142 (N_7142,N_2192,N_3958);
nor U7143 (N_7143,N_358,N_1276);
nor U7144 (N_7144,N_1850,N_889);
nor U7145 (N_7145,N_2338,N_1596);
or U7146 (N_7146,N_2302,N_1162);
or U7147 (N_7147,N_350,N_327);
and U7148 (N_7148,N_381,N_3501);
nor U7149 (N_7149,N_923,N_766);
or U7150 (N_7150,N_217,N_2420);
xnor U7151 (N_7151,N_2749,N_2467);
or U7152 (N_7152,N_1654,N_2617);
nand U7153 (N_7153,N_36,N_2796);
and U7154 (N_7154,N_712,N_3902);
xor U7155 (N_7155,N_3521,N_3869);
nand U7156 (N_7156,N_532,N_889);
or U7157 (N_7157,N_289,N_617);
and U7158 (N_7158,N_1595,N_281);
nand U7159 (N_7159,N_592,N_2800);
nand U7160 (N_7160,N_2909,N_2401);
xor U7161 (N_7161,N_3225,N_2198);
or U7162 (N_7162,N_1901,N_2609);
or U7163 (N_7163,N_1313,N_3527);
nand U7164 (N_7164,N_485,N_1449);
or U7165 (N_7165,N_69,N_293);
nand U7166 (N_7166,N_1013,N_1807);
or U7167 (N_7167,N_2124,N_2141);
nand U7168 (N_7168,N_2309,N_1070);
or U7169 (N_7169,N_2626,N_711);
and U7170 (N_7170,N_2661,N_634);
nor U7171 (N_7171,N_157,N_22);
nand U7172 (N_7172,N_2233,N_1310);
or U7173 (N_7173,N_2583,N_3947);
nand U7174 (N_7174,N_3098,N_49);
and U7175 (N_7175,N_438,N_1038);
nor U7176 (N_7176,N_106,N_2128);
or U7177 (N_7177,N_3358,N_2120);
or U7178 (N_7178,N_3278,N_2015);
and U7179 (N_7179,N_2356,N_3409);
nand U7180 (N_7180,N_2028,N_1328);
and U7181 (N_7181,N_3979,N_358);
nor U7182 (N_7182,N_3391,N_2313);
nand U7183 (N_7183,N_2820,N_653);
or U7184 (N_7184,N_101,N_2256);
or U7185 (N_7185,N_652,N_1800);
or U7186 (N_7186,N_800,N_3563);
xnor U7187 (N_7187,N_2410,N_3681);
or U7188 (N_7188,N_567,N_1554);
nand U7189 (N_7189,N_1884,N_2235);
or U7190 (N_7190,N_1983,N_16);
nor U7191 (N_7191,N_1817,N_1440);
nor U7192 (N_7192,N_3403,N_1946);
nand U7193 (N_7193,N_580,N_3208);
and U7194 (N_7194,N_219,N_1134);
and U7195 (N_7195,N_2186,N_52);
nor U7196 (N_7196,N_338,N_2606);
nand U7197 (N_7197,N_365,N_2881);
nand U7198 (N_7198,N_958,N_2755);
nand U7199 (N_7199,N_2912,N_2297);
nor U7200 (N_7200,N_2914,N_788);
and U7201 (N_7201,N_2991,N_1003);
nor U7202 (N_7202,N_2217,N_328);
nor U7203 (N_7203,N_436,N_167);
nand U7204 (N_7204,N_1275,N_797);
nand U7205 (N_7205,N_2556,N_788);
and U7206 (N_7206,N_2588,N_3655);
and U7207 (N_7207,N_1564,N_2334);
and U7208 (N_7208,N_373,N_1765);
nor U7209 (N_7209,N_3289,N_3753);
nor U7210 (N_7210,N_2952,N_3969);
nor U7211 (N_7211,N_1241,N_3795);
nand U7212 (N_7212,N_1950,N_2159);
xnor U7213 (N_7213,N_1983,N_2920);
nand U7214 (N_7214,N_707,N_2768);
nor U7215 (N_7215,N_1553,N_3958);
nor U7216 (N_7216,N_378,N_1015);
nand U7217 (N_7217,N_934,N_3729);
nor U7218 (N_7218,N_1546,N_3957);
or U7219 (N_7219,N_948,N_8);
and U7220 (N_7220,N_3627,N_330);
and U7221 (N_7221,N_3873,N_2253);
and U7222 (N_7222,N_1242,N_1922);
nor U7223 (N_7223,N_1546,N_2362);
nor U7224 (N_7224,N_2439,N_1021);
nand U7225 (N_7225,N_3197,N_3592);
nand U7226 (N_7226,N_362,N_1797);
nand U7227 (N_7227,N_2149,N_2933);
or U7228 (N_7228,N_641,N_3481);
nand U7229 (N_7229,N_3295,N_3653);
or U7230 (N_7230,N_1115,N_3608);
nand U7231 (N_7231,N_2824,N_2765);
nor U7232 (N_7232,N_1268,N_1567);
or U7233 (N_7233,N_3502,N_1756);
nand U7234 (N_7234,N_1725,N_2905);
and U7235 (N_7235,N_3081,N_433);
nor U7236 (N_7236,N_2187,N_1445);
or U7237 (N_7237,N_1171,N_3332);
xor U7238 (N_7238,N_3352,N_1295);
and U7239 (N_7239,N_554,N_1922);
or U7240 (N_7240,N_2032,N_1293);
nor U7241 (N_7241,N_2616,N_2631);
and U7242 (N_7242,N_3700,N_3283);
xnor U7243 (N_7243,N_1195,N_3213);
or U7244 (N_7244,N_2349,N_1174);
or U7245 (N_7245,N_1745,N_1861);
and U7246 (N_7246,N_2233,N_42);
or U7247 (N_7247,N_1012,N_3585);
or U7248 (N_7248,N_3883,N_1325);
and U7249 (N_7249,N_1205,N_3869);
nand U7250 (N_7250,N_3680,N_2539);
and U7251 (N_7251,N_3038,N_2686);
nand U7252 (N_7252,N_1279,N_1744);
and U7253 (N_7253,N_3434,N_3949);
nor U7254 (N_7254,N_2497,N_1013);
nor U7255 (N_7255,N_879,N_2530);
or U7256 (N_7256,N_476,N_1319);
nand U7257 (N_7257,N_2927,N_507);
and U7258 (N_7258,N_1121,N_3783);
nor U7259 (N_7259,N_3938,N_680);
or U7260 (N_7260,N_2273,N_3488);
and U7261 (N_7261,N_1923,N_422);
xor U7262 (N_7262,N_1052,N_1228);
or U7263 (N_7263,N_2360,N_3861);
and U7264 (N_7264,N_1433,N_972);
nor U7265 (N_7265,N_3821,N_2395);
nand U7266 (N_7266,N_3159,N_1675);
nor U7267 (N_7267,N_667,N_1273);
and U7268 (N_7268,N_2814,N_138);
nand U7269 (N_7269,N_3752,N_2217);
xnor U7270 (N_7270,N_2508,N_492);
or U7271 (N_7271,N_2944,N_455);
nor U7272 (N_7272,N_2785,N_3181);
nor U7273 (N_7273,N_2898,N_3029);
or U7274 (N_7274,N_680,N_559);
or U7275 (N_7275,N_2529,N_356);
or U7276 (N_7276,N_1933,N_1793);
and U7277 (N_7277,N_3317,N_1506);
nand U7278 (N_7278,N_38,N_3290);
xor U7279 (N_7279,N_3941,N_1543);
or U7280 (N_7280,N_23,N_2065);
or U7281 (N_7281,N_3267,N_1938);
or U7282 (N_7282,N_1439,N_124);
nor U7283 (N_7283,N_506,N_2730);
xor U7284 (N_7284,N_506,N_1330);
nand U7285 (N_7285,N_793,N_1681);
or U7286 (N_7286,N_1259,N_943);
or U7287 (N_7287,N_690,N_973);
or U7288 (N_7288,N_801,N_996);
nor U7289 (N_7289,N_2749,N_1227);
or U7290 (N_7290,N_1645,N_1477);
or U7291 (N_7291,N_291,N_795);
or U7292 (N_7292,N_1530,N_682);
or U7293 (N_7293,N_454,N_2955);
and U7294 (N_7294,N_2436,N_2632);
nand U7295 (N_7295,N_1507,N_663);
xnor U7296 (N_7296,N_148,N_377);
nand U7297 (N_7297,N_855,N_3115);
nand U7298 (N_7298,N_136,N_22);
nor U7299 (N_7299,N_2246,N_3466);
nand U7300 (N_7300,N_1957,N_2029);
nor U7301 (N_7301,N_2931,N_1204);
or U7302 (N_7302,N_1837,N_3160);
nor U7303 (N_7303,N_1358,N_718);
nor U7304 (N_7304,N_528,N_3091);
and U7305 (N_7305,N_1177,N_1705);
nor U7306 (N_7306,N_1885,N_2847);
or U7307 (N_7307,N_1525,N_16);
xor U7308 (N_7308,N_1577,N_2702);
and U7309 (N_7309,N_651,N_2432);
xor U7310 (N_7310,N_1066,N_803);
and U7311 (N_7311,N_2809,N_30);
nand U7312 (N_7312,N_2545,N_1315);
xor U7313 (N_7313,N_154,N_3518);
nand U7314 (N_7314,N_611,N_2177);
nand U7315 (N_7315,N_1447,N_2886);
and U7316 (N_7316,N_438,N_1351);
nor U7317 (N_7317,N_850,N_3623);
and U7318 (N_7318,N_3811,N_1601);
nand U7319 (N_7319,N_2035,N_343);
and U7320 (N_7320,N_3476,N_450);
or U7321 (N_7321,N_2164,N_303);
xnor U7322 (N_7322,N_2569,N_3699);
or U7323 (N_7323,N_1810,N_1671);
nand U7324 (N_7324,N_3620,N_3547);
xor U7325 (N_7325,N_3510,N_2810);
or U7326 (N_7326,N_1710,N_2995);
nand U7327 (N_7327,N_1603,N_3601);
xnor U7328 (N_7328,N_2090,N_1128);
xor U7329 (N_7329,N_1268,N_452);
xnor U7330 (N_7330,N_3563,N_3662);
and U7331 (N_7331,N_2397,N_1226);
xnor U7332 (N_7332,N_3977,N_549);
nand U7333 (N_7333,N_1429,N_1857);
or U7334 (N_7334,N_3935,N_1683);
and U7335 (N_7335,N_2672,N_1920);
nor U7336 (N_7336,N_911,N_576);
nor U7337 (N_7337,N_2339,N_3588);
nor U7338 (N_7338,N_344,N_3235);
nand U7339 (N_7339,N_1998,N_1902);
nor U7340 (N_7340,N_514,N_3431);
nor U7341 (N_7341,N_2222,N_1191);
nand U7342 (N_7342,N_1128,N_1075);
nand U7343 (N_7343,N_2302,N_918);
and U7344 (N_7344,N_345,N_3562);
or U7345 (N_7345,N_2051,N_1801);
nand U7346 (N_7346,N_3533,N_3696);
and U7347 (N_7347,N_1370,N_3667);
or U7348 (N_7348,N_2383,N_928);
or U7349 (N_7349,N_1892,N_3942);
or U7350 (N_7350,N_292,N_3575);
and U7351 (N_7351,N_953,N_413);
xnor U7352 (N_7352,N_38,N_1943);
or U7353 (N_7353,N_1154,N_3204);
xnor U7354 (N_7354,N_232,N_1779);
nor U7355 (N_7355,N_853,N_1491);
or U7356 (N_7356,N_1023,N_1858);
and U7357 (N_7357,N_2115,N_2613);
nor U7358 (N_7358,N_1201,N_1315);
or U7359 (N_7359,N_1952,N_808);
nor U7360 (N_7360,N_1774,N_2884);
xor U7361 (N_7361,N_973,N_2113);
nor U7362 (N_7362,N_619,N_2328);
nor U7363 (N_7363,N_1565,N_492);
nor U7364 (N_7364,N_2155,N_965);
nor U7365 (N_7365,N_3651,N_2561);
nand U7366 (N_7366,N_3574,N_1285);
or U7367 (N_7367,N_155,N_3599);
or U7368 (N_7368,N_856,N_2494);
nor U7369 (N_7369,N_3525,N_837);
xor U7370 (N_7370,N_479,N_524);
and U7371 (N_7371,N_2698,N_857);
nand U7372 (N_7372,N_1931,N_2867);
nor U7373 (N_7373,N_369,N_3029);
nand U7374 (N_7374,N_3929,N_3251);
xnor U7375 (N_7375,N_2086,N_3944);
or U7376 (N_7376,N_3731,N_2497);
or U7377 (N_7377,N_3142,N_183);
nand U7378 (N_7378,N_968,N_1427);
nor U7379 (N_7379,N_2727,N_729);
xnor U7380 (N_7380,N_3288,N_3275);
nand U7381 (N_7381,N_1949,N_2029);
or U7382 (N_7382,N_3097,N_2346);
and U7383 (N_7383,N_16,N_3651);
and U7384 (N_7384,N_3055,N_2702);
nor U7385 (N_7385,N_2387,N_2910);
and U7386 (N_7386,N_2879,N_1694);
or U7387 (N_7387,N_37,N_2621);
nor U7388 (N_7388,N_3569,N_3216);
nand U7389 (N_7389,N_3830,N_2385);
and U7390 (N_7390,N_3254,N_3160);
and U7391 (N_7391,N_125,N_333);
and U7392 (N_7392,N_3122,N_2856);
nor U7393 (N_7393,N_3893,N_3313);
nand U7394 (N_7394,N_972,N_1374);
or U7395 (N_7395,N_3926,N_2371);
and U7396 (N_7396,N_3551,N_14);
xnor U7397 (N_7397,N_3980,N_2404);
nor U7398 (N_7398,N_3589,N_1207);
nand U7399 (N_7399,N_3825,N_3621);
nand U7400 (N_7400,N_3641,N_1623);
nand U7401 (N_7401,N_1064,N_2538);
and U7402 (N_7402,N_1041,N_557);
nand U7403 (N_7403,N_622,N_1183);
or U7404 (N_7404,N_3219,N_154);
nand U7405 (N_7405,N_84,N_1488);
nand U7406 (N_7406,N_1177,N_1203);
nand U7407 (N_7407,N_1548,N_288);
and U7408 (N_7408,N_3291,N_3096);
nand U7409 (N_7409,N_430,N_3760);
and U7410 (N_7410,N_22,N_2880);
or U7411 (N_7411,N_1931,N_1000);
nor U7412 (N_7412,N_2787,N_816);
and U7413 (N_7413,N_2468,N_526);
nor U7414 (N_7414,N_2873,N_1252);
or U7415 (N_7415,N_1651,N_1473);
or U7416 (N_7416,N_182,N_2998);
or U7417 (N_7417,N_3701,N_1578);
nand U7418 (N_7418,N_1343,N_3735);
and U7419 (N_7419,N_2661,N_2222);
nand U7420 (N_7420,N_3169,N_3322);
or U7421 (N_7421,N_2371,N_3396);
and U7422 (N_7422,N_1735,N_2407);
nand U7423 (N_7423,N_3368,N_3639);
nand U7424 (N_7424,N_786,N_1018);
nor U7425 (N_7425,N_577,N_3452);
nand U7426 (N_7426,N_968,N_156);
or U7427 (N_7427,N_2137,N_2840);
nor U7428 (N_7428,N_2160,N_3488);
or U7429 (N_7429,N_1754,N_3076);
xor U7430 (N_7430,N_3375,N_3284);
nor U7431 (N_7431,N_2245,N_1823);
nor U7432 (N_7432,N_277,N_2712);
and U7433 (N_7433,N_1644,N_1673);
xor U7434 (N_7434,N_1979,N_2315);
nand U7435 (N_7435,N_2260,N_527);
or U7436 (N_7436,N_934,N_1225);
and U7437 (N_7437,N_949,N_1254);
or U7438 (N_7438,N_1353,N_2404);
or U7439 (N_7439,N_701,N_2061);
or U7440 (N_7440,N_3491,N_2219);
nand U7441 (N_7441,N_3523,N_1645);
nand U7442 (N_7442,N_1359,N_3724);
xor U7443 (N_7443,N_394,N_669);
and U7444 (N_7444,N_470,N_2018);
and U7445 (N_7445,N_2228,N_857);
nand U7446 (N_7446,N_121,N_2802);
nand U7447 (N_7447,N_3012,N_1465);
nand U7448 (N_7448,N_1349,N_3511);
and U7449 (N_7449,N_3933,N_1393);
xnor U7450 (N_7450,N_2902,N_104);
or U7451 (N_7451,N_1608,N_1623);
or U7452 (N_7452,N_2448,N_3032);
or U7453 (N_7453,N_1194,N_3571);
nor U7454 (N_7454,N_1601,N_2121);
or U7455 (N_7455,N_2609,N_2385);
nand U7456 (N_7456,N_1789,N_2310);
nor U7457 (N_7457,N_1752,N_3783);
and U7458 (N_7458,N_2459,N_1485);
and U7459 (N_7459,N_3774,N_1381);
and U7460 (N_7460,N_336,N_478);
nor U7461 (N_7461,N_418,N_109);
or U7462 (N_7462,N_3187,N_2887);
nand U7463 (N_7463,N_3722,N_3673);
nand U7464 (N_7464,N_1438,N_3468);
and U7465 (N_7465,N_1908,N_2923);
or U7466 (N_7466,N_2808,N_1516);
nor U7467 (N_7467,N_1822,N_1619);
nor U7468 (N_7468,N_3395,N_1022);
nand U7469 (N_7469,N_378,N_2971);
nand U7470 (N_7470,N_764,N_1932);
or U7471 (N_7471,N_428,N_838);
nand U7472 (N_7472,N_3430,N_1568);
and U7473 (N_7473,N_3709,N_2425);
and U7474 (N_7474,N_306,N_1688);
nor U7475 (N_7475,N_3994,N_3947);
nor U7476 (N_7476,N_1636,N_3733);
and U7477 (N_7477,N_3978,N_1171);
or U7478 (N_7478,N_354,N_1982);
or U7479 (N_7479,N_2143,N_3148);
nor U7480 (N_7480,N_1123,N_790);
xnor U7481 (N_7481,N_3976,N_1192);
nor U7482 (N_7482,N_1646,N_782);
or U7483 (N_7483,N_2504,N_1128);
or U7484 (N_7484,N_3097,N_2274);
or U7485 (N_7485,N_3330,N_3823);
and U7486 (N_7486,N_1499,N_3260);
and U7487 (N_7487,N_2051,N_2060);
nand U7488 (N_7488,N_96,N_2832);
or U7489 (N_7489,N_1690,N_276);
nand U7490 (N_7490,N_671,N_3326);
and U7491 (N_7491,N_1848,N_2322);
nand U7492 (N_7492,N_3052,N_1937);
and U7493 (N_7493,N_2477,N_3676);
nand U7494 (N_7494,N_968,N_724);
nand U7495 (N_7495,N_605,N_1859);
nand U7496 (N_7496,N_828,N_2532);
nor U7497 (N_7497,N_3931,N_3327);
or U7498 (N_7498,N_3681,N_2057);
nor U7499 (N_7499,N_2909,N_3871);
xor U7500 (N_7500,N_1114,N_199);
nand U7501 (N_7501,N_1342,N_1489);
or U7502 (N_7502,N_1815,N_2406);
and U7503 (N_7503,N_607,N_3384);
and U7504 (N_7504,N_853,N_3948);
or U7505 (N_7505,N_2835,N_1740);
nand U7506 (N_7506,N_1646,N_3164);
nor U7507 (N_7507,N_2557,N_2617);
xor U7508 (N_7508,N_993,N_1662);
nand U7509 (N_7509,N_2223,N_201);
xor U7510 (N_7510,N_511,N_344);
nand U7511 (N_7511,N_864,N_1313);
nand U7512 (N_7512,N_718,N_3741);
nand U7513 (N_7513,N_3456,N_3575);
nand U7514 (N_7514,N_3332,N_3396);
nand U7515 (N_7515,N_1203,N_1749);
nand U7516 (N_7516,N_2835,N_149);
or U7517 (N_7517,N_1006,N_2027);
nand U7518 (N_7518,N_3078,N_3928);
or U7519 (N_7519,N_3973,N_1921);
and U7520 (N_7520,N_1812,N_748);
nand U7521 (N_7521,N_231,N_2099);
nor U7522 (N_7522,N_2231,N_2803);
or U7523 (N_7523,N_1360,N_322);
nand U7524 (N_7524,N_2250,N_3293);
and U7525 (N_7525,N_2009,N_3924);
xor U7526 (N_7526,N_2636,N_648);
xnor U7527 (N_7527,N_382,N_2317);
nand U7528 (N_7528,N_970,N_3186);
and U7529 (N_7529,N_1283,N_3076);
nor U7530 (N_7530,N_3310,N_1389);
or U7531 (N_7531,N_508,N_264);
nand U7532 (N_7532,N_781,N_316);
xor U7533 (N_7533,N_3501,N_2145);
and U7534 (N_7534,N_3627,N_2893);
nand U7535 (N_7535,N_220,N_2020);
nor U7536 (N_7536,N_2010,N_354);
xor U7537 (N_7537,N_272,N_2361);
nand U7538 (N_7538,N_1942,N_1199);
xor U7539 (N_7539,N_3372,N_2243);
and U7540 (N_7540,N_2104,N_1358);
nor U7541 (N_7541,N_3951,N_3879);
or U7542 (N_7542,N_945,N_2711);
nand U7543 (N_7543,N_2183,N_1402);
and U7544 (N_7544,N_464,N_1660);
and U7545 (N_7545,N_700,N_1220);
and U7546 (N_7546,N_3498,N_316);
nand U7547 (N_7547,N_386,N_933);
nor U7548 (N_7548,N_3110,N_1151);
and U7549 (N_7549,N_1749,N_3455);
and U7550 (N_7550,N_987,N_667);
xor U7551 (N_7551,N_1539,N_3686);
nand U7552 (N_7552,N_3256,N_1968);
and U7553 (N_7553,N_2112,N_233);
or U7554 (N_7554,N_3025,N_1544);
nand U7555 (N_7555,N_3043,N_3051);
nand U7556 (N_7556,N_1578,N_2645);
nor U7557 (N_7557,N_1796,N_1778);
nor U7558 (N_7558,N_2284,N_746);
nor U7559 (N_7559,N_3053,N_372);
xor U7560 (N_7560,N_409,N_2720);
and U7561 (N_7561,N_531,N_2477);
nand U7562 (N_7562,N_1630,N_1847);
nand U7563 (N_7563,N_1409,N_634);
nand U7564 (N_7564,N_1367,N_1636);
and U7565 (N_7565,N_1364,N_3023);
and U7566 (N_7566,N_3526,N_2722);
and U7567 (N_7567,N_901,N_2296);
xnor U7568 (N_7568,N_828,N_390);
nor U7569 (N_7569,N_118,N_3063);
or U7570 (N_7570,N_2748,N_3646);
or U7571 (N_7571,N_1488,N_3424);
nand U7572 (N_7572,N_2472,N_2029);
nand U7573 (N_7573,N_3213,N_1319);
and U7574 (N_7574,N_2236,N_812);
nand U7575 (N_7575,N_2277,N_3540);
nor U7576 (N_7576,N_960,N_3899);
xor U7577 (N_7577,N_3777,N_2878);
nand U7578 (N_7578,N_3895,N_3783);
or U7579 (N_7579,N_1283,N_3260);
nor U7580 (N_7580,N_2392,N_2231);
xor U7581 (N_7581,N_2049,N_1153);
and U7582 (N_7582,N_3421,N_3093);
and U7583 (N_7583,N_471,N_3104);
nor U7584 (N_7584,N_554,N_725);
nor U7585 (N_7585,N_1285,N_1100);
or U7586 (N_7586,N_2085,N_3710);
nand U7587 (N_7587,N_3147,N_3818);
nor U7588 (N_7588,N_2090,N_54);
or U7589 (N_7589,N_149,N_45);
nand U7590 (N_7590,N_3669,N_2666);
nand U7591 (N_7591,N_2154,N_2219);
nand U7592 (N_7592,N_1616,N_3727);
and U7593 (N_7593,N_403,N_2142);
nand U7594 (N_7594,N_3490,N_36);
nand U7595 (N_7595,N_3759,N_1435);
or U7596 (N_7596,N_227,N_3300);
or U7597 (N_7597,N_1958,N_2876);
and U7598 (N_7598,N_3249,N_2959);
xnor U7599 (N_7599,N_871,N_1029);
nor U7600 (N_7600,N_748,N_277);
nand U7601 (N_7601,N_2047,N_3339);
and U7602 (N_7602,N_3415,N_2560);
nand U7603 (N_7603,N_2632,N_1802);
and U7604 (N_7604,N_1624,N_692);
or U7605 (N_7605,N_3469,N_3967);
and U7606 (N_7606,N_3592,N_2151);
and U7607 (N_7607,N_2976,N_104);
nand U7608 (N_7608,N_3100,N_668);
or U7609 (N_7609,N_3000,N_3716);
or U7610 (N_7610,N_1164,N_628);
xnor U7611 (N_7611,N_3375,N_611);
nor U7612 (N_7612,N_1800,N_1104);
or U7613 (N_7613,N_3576,N_493);
nand U7614 (N_7614,N_2127,N_2818);
xor U7615 (N_7615,N_3026,N_2682);
and U7616 (N_7616,N_2404,N_3770);
nor U7617 (N_7617,N_188,N_3634);
nand U7618 (N_7618,N_526,N_1893);
or U7619 (N_7619,N_1759,N_3654);
nor U7620 (N_7620,N_1842,N_1773);
and U7621 (N_7621,N_3559,N_1101);
or U7622 (N_7622,N_2470,N_2272);
nor U7623 (N_7623,N_407,N_3987);
and U7624 (N_7624,N_2305,N_3953);
or U7625 (N_7625,N_729,N_1567);
or U7626 (N_7626,N_28,N_3980);
nand U7627 (N_7627,N_470,N_3570);
nor U7628 (N_7628,N_922,N_2230);
or U7629 (N_7629,N_2284,N_3033);
nand U7630 (N_7630,N_2400,N_828);
nor U7631 (N_7631,N_3712,N_1681);
and U7632 (N_7632,N_479,N_1212);
nand U7633 (N_7633,N_1126,N_2422);
and U7634 (N_7634,N_429,N_648);
nand U7635 (N_7635,N_991,N_623);
or U7636 (N_7636,N_1234,N_3169);
xnor U7637 (N_7637,N_1431,N_3892);
nand U7638 (N_7638,N_691,N_2635);
or U7639 (N_7639,N_1710,N_3715);
and U7640 (N_7640,N_2641,N_2252);
nand U7641 (N_7641,N_1539,N_2759);
and U7642 (N_7642,N_1523,N_977);
or U7643 (N_7643,N_1254,N_1815);
nand U7644 (N_7644,N_323,N_3521);
and U7645 (N_7645,N_517,N_2010);
or U7646 (N_7646,N_553,N_1704);
and U7647 (N_7647,N_1324,N_3468);
nor U7648 (N_7648,N_2062,N_1458);
nand U7649 (N_7649,N_2160,N_1981);
nand U7650 (N_7650,N_3481,N_1801);
or U7651 (N_7651,N_1447,N_3440);
or U7652 (N_7652,N_3831,N_63);
nor U7653 (N_7653,N_730,N_3368);
and U7654 (N_7654,N_2127,N_1455);
or U7655 (N_7655,N_3936,N_2185);
or U7656 (N_7656,N_407,N_1465);
xnor U7657 (N_7657,N_2740,N_2244);
nor U7658 (N_7658,N_2922,N_3704);
nand U7659 (N_7659,N_2730,N_2183);
and U7660 (N_7660,N_3698,N_295);
and U7661 (N_7661,N_846,N_721);
nand U7662 (N_7662,N_274,N_3561);
nor U7663 (N_7663,N_3808,N_1379);
nor U7664 (N_7664,N_3734,N_1825);
nand U7665 (N_7665,N_176,N_458);
and U7666 (N_7666,N_2122,N_1799);
and U7667 (N_7667,N_3678,N_2780);
xnor U7668 (N_7668,N_3276,N_1279);
xor U7669 (N_7669,N_1377,N_1991);
nor U7670 (N_7670,N_1587,N_2621);
xnor U7671 (N_7671,N_83,N_3789);
xnor U7672 (N_7672,N_1574,N_3358);
or U7673 (N_7673,N_3,N_125);
and U7674 (N_7674,N_3884,N_98);
xnor U7675 (N_7675,N_2992,N_1328);
nand U7676 (N_7676,N_852,N_1089);
xor U7677 (N_7677,N_1183,N_3542);
xnor U7678 (N_7678,N_413,N_3390);
xnor U7679 (N_7679,N_1404,N_3884);
xor U7680 (N_7680,N_1983,N_509);
nand U7681 (N_7681,N_3962,N_2606);
nor U7682 (N_7682,N_1067,N_3137);
nor U7683 (N_7683,N_2463,N_3045);
nand U7684 (N_7684,N_3390,N_991);
nand U7685 (N_7685,N_436,N_3625);
nor U7686 (N_7686,N_3082,N_2217);
nand U7687 (N_7687,N_620,N_144);
or U7688 (N_7688,N_794,N_3872);
nor U7689 (N_7689,N_1379,N_1008);
nand U7690 (N_7690,N_301,N_3347);
nor U7691 (N_7691,N_3924,N_542);
nand U7692 (N_7692,N_2237,N_755);
nand U7693 (N_7693,N_3655,N_3621);
nor U7694 (N_7694,N_2688,N_1819);
nand U7695 (N_7695,N_2567,N_3858);
and U7696 (N_7696,N_2944,N_1135);
or U7697 (N_7697,N_485,N_240);
and U7698 (N_7698,N_3863,N_2968);
or U7699 (N_7699,N_2051,N_2289);
or U7700 (N_7700,N_3310,N_1872);
or U7701 (N_7701,N_2175,N_688);
or U7702 (N_7702,N_2319,N_1695);
or U7703 (N_7703,N_1020,N_2700);
nand U7704 (N_7704,N_488,N_548);
xor U7705 (N_7705,N_2627,N_924);
nand U7706 (N_7706,N_2391,N_2096);
or U7707 (N_7707,N_445,N_2604);
nand U7708 (N_7708,N_2194,N_2921);
or U7709 (N_7709,N_3787,N_1706);
or U7710 (N_7710,N_412,N_2998);
and U7711 (N_7711,N_89,N_1168);
nand U7712 (N_7712,N_936,N_1915);
and U7713 (N_7713,N_1259,N_3575);
nand U7714 (N_7714,N_78,N_3339);
nor U7715 (N_7715,N_3774,N_3739);
and U7716 (N_7716,N_698,N_2521);
xnor U7717 (N_7717,N_363,N_1076);
and U7718 (N_7718,N_435,N_3968);
and U7719 (N_7719,N_1293,N_1069);
nor U7720 (N_7720,N_3175,N_1367);
or U7721 (N_7721,N_2805,N_3367);
or U7722 (N_7722,N_326,N_3233);
or U7723 (N_7723,N_2468,N_3347);
or U7724 (N_7724,N_3230,N_2715);
or U7725 (N_7725,N_2484,N_747);
and U7726 (N_7726,N_3054,N_1054);
xor U7727 (N_7727,N_3793,N_2936);
nand U7728 (N_7728,N_3202,N_1352);
and U7729 (N_7729,N_226,N_1158);
nand U7730 (N_7730,N_3555,N_2642);
nand U7731 (N_7731,N_1146,N_3296);
nand U7732 (N_7732,N_2558,N_2645);
or U7733 (N_7733,N_1391,N_1466);
nand U7734 (N_7734,N_1239,N_1508);
nor U7735 (N_7735,N_3605,N_2182);
nand U7736 (N_7736,N_225,N_368);
nand U7737 (N_7737,N_3173,N_1171);
nand U7738 (N_7738,N_1276,N_2546);
and U7739 (N_7739,N_1037,N_2219);
xor U7740 (N_7740,N_3618,N_906);
and U7741 (N_7741,N_68,N_1767);
or U7742 (N_7742,N_2860,N_496);
xnor U7743 (N_7743,N_2815,N_46);
or U7744 (N_7744,N_2215,N_2967);
or U7745 (N_7745,N_1478,N_2714);
nor U7746 (N_7746,N_1710,N_1865);
xor U7747 (N_7747,N_3478,N_396);
nand U7748 (N_7748,N_2798,N_1511);
nand U7749 (N_7749,N_97,N_963);
xor U7750 (N_7750,N_3570,N_1795);
nand U7751 (N_7751,N_1962,N_1850);
nor U7752 (N_7752,N_3049,N_3461);
nand U7753 (N_7753,N_3176,N_839);
xnor U7754 (N_7754,N_3209,N_2671);
or U7755 (N_7755,N_824,N_1491);
nand U7756 (N_7756,N_3884,N_2724);
or U7757 (N_7757,N_2090,N_3678);
and U7758 (N_7758,N_1156,N_2651);
nand U7759 (N_7759,N_1408,N_1508);
xnor U7760 (N_7760,N_895,N_1694);
nor U7761 (N_7761,N_2649,N_758);
nand U7762 (N_7762,N_811,N_3725);
xor U7763 (N_7763,N_669,N_3058);
xor U7764 (N_7764,N_415,N_2452);
and U7765 (N_7765,N_1234,N_551);
and U7766 (N_7766,N_2267,N_3455);
xnor U7767 (N_7767,N_1630,N_165);
or U7768 (N_7768,N_2426,N_3441);
nand U7769 (N_7769,N_3904,N_549);
nor U7770 (N_7770,N_2134,N_3227);
nor U7771 (N_7771,N_263,N_3026);
and U7772 (N_7772,N_1799,N_401);
and U7773 (N_7773,N_3252,N_3802);
and U7774 (N_7774,N_151,N_3637);
xnor U7775 (N_7775,N_388,N_3530);
nand U7776 (N_7776,N_109,N_1657);
nor U7777 (N_7777,N_2045,N_2675);
nand U7778 (N_7778,N_2857,N_768);
nor U7779 (N_7779,N_3988,N_3127);
nor U7780 (N_7780,N_820,N_1953);
nand U7781 (N_7781,N_36,N_1946);
or U7782 (N_7782,N_3120,N_3224);
nand U7783 (N_7783,N_2228,N_3953);
or U7784 (N_7784,N_346,N_179);
nor U7785 (N_7785,N_1183,N_838);
or U7786 (N_7786,N_1774,N_388);
and U7787 (N_7787,N_3472,N_3936);
nor U7788 (N_7788,N_2719,N_3697);
nor U7789 (N_7789,N_991,N_3700);
and U7790 (N_7790,N_3731,N_819);
nand U7791 (N_7791,N_1574,N_3507);
or U7792 (N_7792,N_2586,N_694);
and U7793 (N_7793,N_657,N_3436);
nand U7794 (N_7794,N_3214,N_3569);
nor U7795 (N_7795,N_2483,N_2580);
or U7796 (N_7796,N_2240,N_3265);
and U7797 (N_7797,N_1713,N_2051);
nand U7798 (N_7798,N_1635,N_3062);
or U7799 (N_7799,N_2924,N_3287);
or U7800 (N_7800,N_1971,N_524);
or U7801 (N_7801,N_3028,N_2441);
or U7802 (N_7802,N_3689,N_824);
and U7803 (N_7803,N_2734,N_27);
xnor U7804 (N_7804,N_380,N_3730);
nand U7805 (N_7805,N_2394,N_1888);
or U7806 (N_7806,N_1608,N_2205);
xnor U7807 (N_7807,N_2027,N_1311);
nor U7808 (N_7808,N_3887,N_558);
nand U7809 (N_7809,N_3672,N_3530);
nand U7810 (N_7810,N_555,N_3745);
nor U7811 (N_7811,N_655,N_772);
xor U7812 (N_7812,N_3752,N_1033);
and U7813 (N_7813,N_2964,N_2222);
and U7814 (N_7814,N_1158,N_2963);
nor U7815 (N_7815,N_3151,N_3749);
nor U7816 (N_7816,N_2755,N_2113);
nor U7817 (N_7817,N_3257,N_3792);
xnor U7818 (N_7818,N_915,N_2607);
nor U7819 (N_7819,N_836,N_2033);
nand U7820 (N_7820,N_289,N_348);
nor U7821 (N_7821,N_2667,N_523);
nor U7822 (N_7822,N_484,N_961);
nand U7823 (N_7823,N_992,N_505);
and U7824 (N_7824,N_3487,N_2164);
or U7825 (N_7825,N_3192,N_3247);
nor U7826 (N_7826,N_1741,N_361);
nand U7827 (N_7827,N_1076,N_2203);
nor U7828 (N_7828,N_3790,N_348);
and U7829 (N_7829,N_1673,N_1549);
xnor U7830 (N_7830,N_300,N_2047);
xor U7831 (N_7831,N_1946,N_436);
or U7832 (N_7832,N_3644,N_1886);
and U7833 (N_7833,N_1216,N_890);
nand U7834 (N_7834,N_887,N_1260);
and U7835 (N_7835,N_3667,N_1339);
or U7836 (N_7836,N_2451,N_3108);
nor U7837 (N_7837,N_774,N_2943);
or U7838 (N_7838,N_3677,N_1030);
and U7839 (N_7839,N_526,N_2061);
nand U7840 (N_7840,N_253,N_838);
nor U7841 (N_7841,N_300,N_2748);
nand U7842 (N_7842,N_2491,N_2201);
and U7843 (N_7843,N_2678,N_2765);
and U7844 (N_7844,N_735,N_3741);
nand U7845 (N_7845,N_2323,N_516);
xnor U7846 (N_7846,N_37,N_3857);
nand U7847 (N_7847,N_520,N_3554);
or U7848 (N_7848,N_37,N_1906);
nand U7849 (N_7849,N_3839,N_1137);
nand U7850 (N_7850,N_2942,N_1797);
or U7851 (N_7851,N_214,N_298);
xnor U7852 (N_7852,N_3071,N_852);
nor U7853 (N_7853,N_56,N_889);
and U7854 (N_7854,N_2638,N_2142);
or U7855 (N_7855,N_2994,N_3563);
nor U7856 (N_7856,N_1137,N_2789);
or U7857 (N_7857,N_751,N_2827);
or U7858 (N_7858,N_428,N_3518);
or U7859 (N_7859,N_1848,N_3615);
and U7860 (N_7860,N_742,N_2236);
or U7861 (N_7861,N_3193,N_1890);
nor U7862 (N_7862,N_1354,N_3664);
and U7863 (N_7863,N_3735,N_1578);
nor U7864 (N_7864,N_998,N_1196);
or U7865 (N_7865,N_3988,N_1814);
nand U7866 (N_7866,N_511,N_3622);
nand U7867 (N_7867,N_3048,N_2858);
nand U7868 (N_7868,N_1439,N_1046);
and U7869 (N_7869,N_1563,N_3867);
xnor U7870 (N_7870,N_1184,N_2030);
nor U7871 (N_7871,N_254,N_2022);
or U7872 (N_7872,N_3282,N_3293);
and U7873 (N_7873,N_450,N_2458);
nand U7874 (N_7874,N_2040,N_1826);
or U7875 (N_7875,N_2039,N_799);
and U7876 (N_7876,N_1859,N_1019);
and U7877 (N_7877,N_1359,N_3522);
nor U7878 (N_7878,N_507,N_1642);
nor U7879 (N_7879,N_84,N_880);
and U7880 (N_7880,N_2349,N_3526);
nand U7881 (N_7881,N_225,N_141);
nor U7882 (N_7882,N_1533,N_2705);
nor U7883 (N_7883,N_111,N_1788);
xor U7884 (N_7884,N_3860,N_2089);
nand U7885 (N_7885,N_1762,N_2937);
nor U7886 (N_7886,N_1421,N_1269);
nor U7887 (N_7887,N_1768,N_2406);
or U7888 (N_7888,N_1451,N_3162);
nor U7889 (N_7889,N_3090,N_1838);
nor U7890 (N_7890,N_1066,N_1685);
nand U7891 (N_7891,N_543,N_1500);
and U7892 (N_7892,N_986,N_2485);
xor U7893 (N_7893,N_2150,N_2216);
nor U7894 (N_7894,N_1757,N_1737);
nand U7895 (N_7895,N_3509,N_1720);
and U7896 (N_7896,N_588,N_807);
nand U7897 (N_7897,N_840,N_1607);
nor U7898 (N_7898,N_1713,N_1559);
nor U7899 (N_7899,N_13,N_2935);
nor U7900 (N_7900,N_3973,N_1732);
nand U7901 (N_7901,N_2911,N_3685);
nand U7902 (N_7902,N_285,N_2399);
or U7903 (N_7903,N_2667,N_1081);
and U7904 (N_7904,N_2695,N_3391);
nor U7905 (N_7905,N_1525,N_3615);
or U7906 (N_7906,N_574,N_3571);
or U7907 (N_7907,N_1565,N_2138);
or U7908 (N_7908,N_397,N_2242);
or U7909 (N_7909,N_2176,N_1666);
nand U7910 (N_7910,N_2596,N_74);
nor U7911 (N_7911,N_182,N_2977);
nor U7912 (N_7912,N_1919,N_2633);
xnor U7913 (N_7913,N_562,N_1394);
nor U7914 (N_7914,N_3581,N_1330);
nand U7915 (N_7915,N_2050,N_2408);
and U7916 (N_7916,N_3914,N_2808);
or U7917 (N_7917,N_2463,N_3377);
or U7918 (N_7918,N_2215,N_3886);
or U7919 (N_7919,N_3812,N_3781);
nand U7920 (N_7920,N_1618,N_2428);
xor U7921 (N_7921,N_3932,N_1837);
nor U7922 (N_7922,N_1331,N_621);
and U7923 (N_7923,N_3295,N_2857);
nor U7924 (N_7924,N_2245,N_1034);
or U7925 (N_7925,N_1976,N_3651);
nand U7926 (N_7926,N_978,N_3522);
nor U7927 (N_7927,N_1138,N_2227);
nor U7928 (N_7928,N_1849,N_2037);
or U7929 (N_7929,N_2688,N_1254);
nand U7930 (N_7930,N_683,N_1795);
nor U7931 (N_7931,N_365,N_1782);
xor U7932 (N_7932,N_282,N_1215);
xnor U7933 (N_7933,N_1340,N_2276);
nand U7934 (N_7934,N_1898,N_3493);
xor U7935 (N_7935,N_2683,N_380);
nand U7936 (N_7936,N_1112,N_2804);
or U7937 (N_7937,N_1804,N_671);
and U7938 (N_7938,N_3329,N_911);
or U7939 (N_7939,N_900,N_2761);
and U7940 (N_7940,N_2249,N_3465);
nand U7941 (N_7941,N_129,N_1922);
and U7942 (N_7942,N_3186,N_511);
nor U7943 (N_7943,N_3949,N_2518);
nor U7944 (N_7944,N_2884,N_2832);
nand U7945 (N_7945,N_1714,N_1440);
nand U7946 (N_7946,N_1959,N_766);
nand U7947 (N_7947,N_18,N_2907);
or U7948 (N_7948,N_1231,N_984);
nor U7949 (N_7949,N_3886,N_3252);
and U7950 (N_7950,N_3825,N_3130);
nand U7951 (N_7951,N_2129,N_1296);
and U7952 (N_7952,N_1587,N_1593);
nand U7953 (N_7953,N_996,N_3935);
nor U7954 (N_7954,N_3384,N_3887);
nor U7955 (N_7955,N_397,N_1748);
and U7956 (N_7956,N_258,N_3193);
and U7957 (N_7957,N_628,N_2762);
or U7958 (N_7958,N_2897,N_3372);
nand U7959 (N_7959,N_2729,N_1357);
or U7960 (N_7960,N_322,N_227);
or U7961 (N_7961,N_1605,N_1475);
or U7962 (N_7962,N_3319,N_2573);
and U7963 (N_7963,N_1503,N_3266);
or U7964 (N_7964,N_832,N_895);
nand U7965 (N_7965,N_2457,N_1608);
nand U7966 (N_7966,N_1819,N_1031);
and U7967 (N_7967,N_957,N_3132);
nor U7968 (N_7968,N_2880,N_3524);
and U7969 (N_7969,N_1225,N_1963);
or U7970 (N_7970,N_2211,N_2431);
and U7971 (N_7971,N_2612,N_200);
and U7972 (N_7972,N_490,N_2982);
nor U7973 (N_7973,N_3883,N_3743);
nand U7974 (N_7974,N_3816,N_987);
or U7975 (N_7975,N_3152,N_1973);
and U7976 (N_7976,N_1842,N_588);
or U7977 (N_7977,N_1419,N_1901);
nand U7978 (N_7978,N_3429,N_3144);
or U7979 (N_7979,N_988,N_696);
or U7980 (N_7980,N_1798,N_3709);
nor U7981 (N_7981,N_1221,N_529);
nor U7982 (N_7982,N_2210,N_3645);
nand U7983 (N_7983,N_1464,N_3968);
nor U7984 (N_7984,N_3623,N_2934);
nor U7985 (N_7985,N_1049,N_3998);
or U7986 (N_7986,N_820,N_1441);
or U7987 (N_7987,N_2392,N_882);
nor U7988 (N_7988,N_2871,N_3687);
nand U7989 (N_7989,N_65,N_2476);
or U7990 (N_7990,N_2635,N_3439);
or U7991 (N_7991,N_1630,N_1526);
nor U7992 (N_7992,N_469,N_1133);
nand U7993 (N_7993,N_839,N_1618);
or U7994 (N_7994,N_3329,N_1817);
and U7995 (N_7995,N_1033,N_3371);
nand U7996 (N_7996,N_1380,N_1535);
nor U7997 (N_7997,N_3363,N_2831);
nand U7998 (N_7998,N_674,N_3408);
nor U7999 (N_7999,N_1541,N_681);
or U8000 (N_8000,N_7077,N_5856);
nand U8001 (N_8001,N_5649,N_5661);
nand U8002 (N_8002,N_7973,N_4808);
nand U8003 (N_8003,N_4716,N_7733);
nor U8004 (N_8004,N_4103,N_6898);
nor U8005 (N_8005,N_5434,N_6103);
nand U8006 (N_8006,N_7683,N_6236);
nand U8007 (N_8007,N_4405,N_7576);
nand U8008 (N_8008,N_6663,N_7656);
or U8009 (N_8009,N_7991,N_7422);
xnor U8010 (N_8010,N_4752,N_5672);
or U8011 (N_8011,N_7200,N_7857);
nor U8012 (N_8012,N_6509,N_4574);
nand U8013 (N_8013,N_4925,N_7229);
nor U8014 (N_8014,N_4313,N_6413);
or U8015 (N_8015,N_5113,N_5387);
xnor U8016 (N_8016,N_7541,N_5280);
nand U8017 (N_8017,N_6015,N_5605);
nand U8018 (N_8018,N_6642,N_4408);
or U8019 (N_8019,N_5878,N_4144);
nand U8020 (N_8020,N_5376,N_7043);
nand U8021 (N_8021,N_7842,N_6360);
nor U8022 (N_8022,N_6829,N_7676);
xnor U8023 (N_8023,N_4460,N_5256);
nand U8024 (N_8024,N_5989,N_7421);
nand U8025 (N_8025,N_6448,N_5528);
or U8026 (N_8026,N_4109,N_5178);
and U8027 (N_8027,N_5821,N_6925);
nand U8028 (N_8028,N_5899,N_5704);
or U8029 (N_8029,N_6504,N_6011);
nand U8030 (N_8030,N_4899,N_4528);
or U8031 (N_8031,N_6200,N_5272);
or U8032 (N_8032,N_5552,N_7803);
or U8033 (N_8033,N_7906,N_7603);
nor U8034 (N_8034,N_5205,N_7832);
and U8035 (N_8035,N_4805,N_7053);
and U8036 (N_8036,N_5334,N_5909);
and U8037 (N_8037,N_7258,N_4216);
or U8038 (N_8038,N_4960,N_6049);
or U8039 (N_8039,N_5812,N_7032);
and U8040 (N_8040,N_5053,N_6094);
or U8041 (N_8041,N_6393,N_4613);
and U8042 (N_8042,N_5163,N_4484);
and U8043 (N_8043,N_7849,N_7372);
xor U8044 (N_8044,N_7402,N_5841);
and U8045 (N_8045,N_7256,N_5832);
nor U8046 (N_8046,N_7942,N_7390);
xnor U8047 (N_8047,N_7764,N_6538);
and U8048 (N_8048,N_6331,N_6432);
and U8049 (N_8049,N_6778,N_6842);
nor U8050 (N_8050,N_4547,N_7648);
and U8051 (N_8051,N_5910,N_5515);
and U8052 (N_8052,N_7954,N_5249);
or U8053 (N_8053,N_4247,N_7412);
nand U8054 (N_8054,N_4041,N_6499);
nor U8055 (N_8055,N_6831,N_7451);
and U8056 (N_8056,N_4929,N_6548);
nor U8057 (N_8057,N_6553,N_5602);
nand U8058 (N_8058,N_4178,N_5212);
nor U8059 (N_8059,N_7356,N_7270);
nor U8060 (N_8060,N_4994,N_4243);
nand U8061 (N_8061,N_4399,N_6173);
nor U8062 (N_8062,N_6300,N_7584);
or U8063 (N_8063,N_7978,N_7135);
nor U8064 (N_8064,N_6027,N_6709);
or U8065 (N_8065,N_4560,N_7086);
or U8066 (N_8066,N_6157,N_7345);
and U8067 (N_8067,N_4757,N_6068);
and U8068 (N_8068,N_6557,N_6617);
and U8069 (N_8069,N_4162,N_5202);
or U8070 (N_8070,N_4636,N_4588);
and U8071 (N_8071,N_4219,N_4827);
or U8072 (N_8072,N_4346,N_5028);
or U8073 (N_8073,N_5019,N_5677);
nand U8074 (N_8074,N_5965,N_7953);
xor U8075 (N_8075,N_5669,N_6927);
nor U8076 (N_8076,N_6612,N_6799);
or U8077 (N_8077,N_4421,N_5009);
nand U8078 (N_8078,N_5162,N_7686);
and U8079 (N_8079,N_6710,N_5988);
nand U8080 (N_8080,N_6256,N_7429);
nor U8081 (N_8081,N_6754,N_6694);
nand U8082 (N_8082,N_6138,N_7231);
or U8083 (N_8083,N_6420,N_7493);
nand U8084 (N_8084,N_7209,N_4812);
and U8085 (N_8085,N_7932,N_7678);
nor U8086 (N_8086,N_6823,N_4485);
or U8087 (N_8087,N_7638,N_5340);
xnor U8088 (N_8088,N_6184,N_5996);
and U8089 (N_8089,N_6127,N_6382);
nand U8090 (N_8090,N_6240,N_7650);
or U8091 (N_8091,N_6116,N_7715);
nor U8092 (N_8092,N_5597,N_4428);
and U8093 (N_8093,N_5355,N_6916);
nand U8094 (N_8094,N_4133,N_4034);
and U8095 (N_8095,N_4623,N_4285);
or U8096 (N_8096,N_7261,N_5460);
or U8097 (N_8097,N_4909,N_5186);
nor U8098 (N_8098,N_7623,N_7639);
xnor U8099 (N_8099,N_4089,N_4815);
nand U8100 (N_8100,N_7708,N_6903);
or U8101 (N_8101,N_5763,N_4958);
and U8102 (N_8102,N_4748,N_5466);
nor U8103 (N_8103,N_7195,N_7950);
nor U8104 (N_8104,N_7166,N_4085);
or U8105 (N_8105,N_6503,N_7250);
and U8106 (N_8106,N_5201,N_5080);
and U8107 (N_8107,N_6700,N_6628);
or U8108 (N_8108,N_6301,N_4440);
nand U8109 (N_8109,N_6813,N_4657);
and U8110 (N_8110,N_4728,N_5316);
xor U8111 (N_8111,N_4214,N_4493);
xnor U8112 (N_8112,N_4443,N_7401);
or U8113 (N_8113,N_5916,N_5550);
nor U8114 (N_8114,N_5521,N_5500);
and U8115 (N_8115,N_7113,N_5033);
and U8116 (N_8116,N_4300,N_6544);
nand U8117 (N_8117,N_5265,N_5148);
nor U8118 (N_8118,N_6645,N_7843);
nor U8119 (N_8119,N_6653,N_6691);
nor U8120 (N_8120,N_6262,N_4101);
or U8121 (N_8121,N_4818,N_6824);
nand U8122 (N_8122,N_7546,N_6471);
nor U8123 (N_8123,N_5433,N_7613);
and U8124 (N_8124,N_5772,N_7153);
and U8125 (N_8125,N_4856,N_7004);
or U8126 (N_8126,N_5694,N_7123);
and U8127 (N_8127,N_5285,N_7500);
and U8128 (N_8128,N_5585,N_5819);
and U8129 (N_8129,N_5182,N_6789);
xor U8130 (N_8130,N_7288,N_6220);
and U8131 (N_8131,N_5332,N_5850);
nor U8132 (N_8132,N_6580,N_4385);
xor U8133 (N_8133,N_5563,N_6947);
and U8134 (N_8134,N_5302,N_7727);
and U8135 (N_8135,N_5663,N_5258);
nor U8136 (N_8136,N_7736,N_5138);
nor U8137 (N_8137,N_5818,N_5096);
nor U8138 (N_8138,N_4212,N_4531);
nand U8139 (N_8139,N_5099,N_4306);
nand U8140 (N_8140,N_4668,N_4427);
xnor U8141 (N_8141,N_6266,N_6041);
xor U8142 (N_8142,N_4038,N_4833);
nor U8143 (N_8143,N_4609,N_4107);
nor U8144 (N_8144,N_6915,N_6878);
nand U8145 (N_8145,N_4483,N_6441);
nand U8146 (N_8146,N_6456,N_4849);
and U8147 (N_8147,N_5975,N_5496);
and U8148 (N_8148,N_6371,N_4165);
and U8149 (N_8149,N_4556,N_5396);
nand U8150 (N_8150,N_4284,N_7640);
and U8151 (N_8151,N_4314,N_7001);
and U8152 (N_8152,N_7168,N_6464);
and U8153 (N_8153,N_7621,N_5351);
and U8154 (N_8154,N_5510,N_5278);
nand U8155 (N_8155,N_7267,N_4937);
and U8156 (N_8156,N_6000,N_7349);
xnor U8157 (N_8157,N_6550,N_6746);
nand U8158 (N_8158,N_6110,N_5685);
nand U8159 (N_8159,N_5705,N_6846);
xor U8160 (N_8160,N_5871,N_5638);
nand U8161 (N_8161,N_4648,N_6232);
nor U8162 (N_8162,N_5259,N_7711);
nor U8163 (N_8163,N_4110,N_4763);
xor U8164 (N_8164,N_6678,N_7306);
and U8165 (N_8165,N_4244,N_4148);
nor U8166 (N_8166,N_7337,N_7347);
nand U8167 (N_8167,N_4396,N_4775);
or U8168 (N_8168,N_6610,N_4772);
and U8169 (N_8169,N_4131,N_5077);
or U8170 (N_8170,N_6293,N_5948);
and U8171 (N_8171,N_6951,N_5224);
xnor U8172 (N_8172,N_4802,N_4690);
and U8173 (N_8173,N_4468,N_7757);
and U8174 (N_8174,N_7431,N_5015);
nor U8175 (N_8175,N_6261,N_6163);
nor U8176 (N_8176,N_4942,N_6463);
nor U8177 (N_8177,N_7798,N_6198);
xnor U8178 (N_8178,N_5063,N_4544);
or U8179 (N_8179,N_5740,N_6031);
nand U8180 (N_8180,N_5655,N_6359);
and U8181 (N_8181,N_4024,N_6913);
nand U8182 (N_8182,N_7911,N_5027);
nor U8183 (N_8183,N_6687,N_5848);
nor U8184 (N_8184,N_5294,N_4670);
nand U8185 (N_8185,N_4414,N_5445);
or U8186 (N_8186,N_5397,N_6943);
nand U8187 (N_8187,N_5583,N_5102);
nand U8188 (N_8188,N_6906,N_5365);
nand U8189 (N_8189,N_7693,N_6938);
nand U8190 (N_8190,N_5925,N_4832);
and U8191 (N_8191,N_6931,N_4477);
or U8192 (N_8192,N_4218,N_6762);
and U8193 (N_8193,N_7377,N_7398);
nor U8194 (N_8194,N_5643,N_5727);
or U8195 (N_8195,N_6102,N_4451);
nor U8196 (N_8196,N_5309,N_5745);
and U8197 (N_8197,N_5974,N_5554);
xor U8198 (N_8198,N_6433,N_6206);
nand U8199 (N_8199,N_5110,N_4316);
nor U8200 (N_8200,N_6564,N_7805);
and U8201 (N_8201,N_6322,N_5593);
nand U8202 (N_8202,N_7877,N_6954);
and U8203 (N_8203,N_5516,N_5230);
nand U8204 (N_8204,N_6790,N_4237);
or U8205 (N_8205,N_5065,N_7327);
xor U8206 (N_8206,N_5070,N_5736);
xnor U8207 (N_8207,N_7382,N_5068);
nand U8208 (N_8208,N_5407,N_6034);
nand U8209 (N_8209,N_6641,N_7188);
nand U8210 (N_8210,N_5699,N_7794);
nand U8211 (N_8211,N_7517,N_7015);
nand U8212 (N_8212,N_6987,N_4712);
or U8213 (N_8213,N_7698,N_4866);
and U8214 (N_8214,N_7782,N_7170);
and U8215 (N_8215,N_6204,N_4630);
or U8216 (N_8216,N_6469,N_4683);
and U8217 (N_8217,N_6515,N_4324);
nand U8218 (N_8218,N_7552,N_5125);
or U8219 (N_8219,N_4208,N_7420);
xor U8220 (N_8220,N_7065,N_4055);
nand U8221 (N_8221,N_5250,N_7643);
and U8222 (N_8222,N_6844,N_7821);
nand U8223 (N_8223,N_4173,N_4126);
xnor U8224 (N_8224,N_4215,N_7918);
or U8225 (N_8225,N_6984,N_4020);
nor U8226 (N_8226,N_7467,N_4241);
or U8227 (N_8227,N_4660,N_7284);
nand U8228 (N_8228,N_5357,N_6271);
nand U8229 (N_8229,N_7082,N_6277);
nor U8230 (N_8230,N_7454,N_5236);
and U8231 (N_8231,N_6111,N_4418);
or U8232 (N_8232,N_6107,N_4721);
nand U8233 (N_8233,N_7442,N_6815);
or U8234 (N_8234,N_7155,N_4074);
nor U8235 (N_8235,N_5847,N_6238);
and U8236 (N_8236,N_7407,N_4159);
or U8237 (N_8237,N_5419,N_4600);
and U8238 (N_8238,N_6583,N_6424);
nand U8239 (N_8239,N_5518,N_6028);
and U8240 (N_8240,N_6542,N_6358);
and U8241 (N_8241,N_4249,N_6519);
and U8242 (N_8242,N_5431,N_6969);
nand U8243 (N_8243,N_6730,N_4844);
and U8244 (N_8244,N_6212,N_4652);
nand U8245 (N_8245,N_4417,N_7182);
xor U8246 (N_8246,N_5846,N_6452);
nor U8247 (N_8247,N_5632,N_5668);
and U8248 (N_8248,N_5568,N_4449);
nand U8249 (N_8249,N_5582,N_6618);
nor U8250 (N_8250,N_4662,N_5043);
and U8251 (N_8251,N_6263,N_6723);
nor U8252 (N_8252,N_5895,N_4202);
nor U8253 (N_8253,N_6890,N_4745);
or U8254 (N_8254,N_7901,N_5581);
nor U8255 (N_8255,N_6769,N_6834);
and U8256 (N_8256,N_4147,N_6311);
and U8257 (N_8257,N_5007,N_5385);
xnor U8258 (N_8258,N_7974,N_7120);
and U8259 (N_8259,N_6404,N_4064);
and U8260 (N_8260,N_7192,N_6197);
and U8261 (N_8261,N_4529,N_7202);
and U8262 (N_8262,N_4321,N_5945);
xnor U8263 (N_8263,N_4480,N_6662);
nor U8264 (N_8264,N_4262,N_4222);
nand U8265 (N_8265,N_7259,N_4186);
and U8266 (N_8266,N_5831,N_6837);
nand U8267 (N_8267,N_6123,N_7759);
nor U8268 (N_8268,N_5891,N_4627);
or U8269 (N_8269,N_4582,N_4319);
or U8270 (N_8270,N_5506,N_4658);
or U8271 (N_8271,N_7941,N_4629);
xor U8272 (N_8272,N_4393,N_4277);
and U8273 (N_8273,N_6155,N_7561);
nand U8274 (N_8274,N_4195,N_4703);
nor U8275 (N_8275,N_5322,N_6633);
or U8276 (N_8276,N_4674,N_5588);
and U8277 (N_8277,N_4590,N_6217);
or U8278 (N_8278,N_4268,N_5416);
nand U8279 (N_8279,N_7511,N_7062);
nor U8280 (N_8280,N_5479,N_6254);
and U8281 (N_8281,N_6039,N_7020);
nor U8282 (N_8282,N_6250,N_4568);
nand U8283 (N_8283,N_5135,N_5900);
nand U8284 (N_8284,N_7283,N_6899);
xor U8285 (N_8285,N_7361,N_6934);
nand U8286 (N_8286,N_7406,N_7784);
or U8287 (N_8287,N_6506,N_4564);
or U8288 (N_8288,N_7738,N_5219);
nand U8289 (N_8289,N_7900,N_4895);
or U8290 (N_8290,N_5780,N_6387);
nand U8291 (N_8291,N_6342,N_7884);
xor U8292 (N_8292,N_4618,N_4365);
nor U8293 (N_8293,N_5088,N_6026);
or U8294 (N_8294,N_7460,N_5543);
and U8295 (N_8295,N_5696,N_5362);
or U8296 (N_8296,N_6679,N_7714);
nor U8297 (N_8297,N_4117,N_7479);
and U8298 (N_8298,N_6479,N_7786);
nor U8299 (N_8299,N_5714,N_7988);
or U8300 (N_8300,N_4552,N_4998);
and U8301 (N_8301,N_4153,N_7801);
nand U8302 (N_8302,N_6063,N_6482);
and U8303 (N_8303,N_7658,N_5659);
nand U8304 (N_8304,N_6446,N_4213);
nor U8305 (N_8305,N_5888,N_4146);
nand U8306 (N_8306,N_6447,N_5599);
xor U8307 (N_8307,N_4143,N_4593);
nand U8308 (N_8308,N_5901,N_6900);
nand U8309 (N_8309,N_4021,N_5321);
and U8310 (N_8310,N_7140,N_4388);
nand U8311 (N_8311,N_7626,N_5475);
nor U8312 (N_8312,N_5657,N_7958);
nor U8313 (N_8313,N_7161,N_6229);
or U8314 (N_8314,N_4869,N_6600);
nor U8315 (N_8315,N_7824,N_6705);
nand U8316 (N_8316,N_7696,N_6351);
and U8317 (N_8317,N_7934,N_6333);
nor U8318 (N_8318,N_5003,N_6370);
or U8319 (N_8319,N_5555,N_7052);
nor U8320 (N_8320,N_6502,N_4035);
and U8321 (N_8321,N_6388,N_4707);
nor U8322 (N_8322,N_7569,N_4134);
or U8323 (N_8323,N_7755,N_6779);
or U8324 (N_8324,N_7927,N_7047);
or U8325 (N_8325,N_7718,N_7018);
or U8326 (N_8326,N_4139,N_5048);
and U8327 (N_8327,N_6821,N_4053);
and U8328 (N_8328,N_6367,N_7960);
xnor U8329 (N_8329,N_6081,N_5379);
nand U8330 (N_8330,N_5912,N_4723);
and U8331 (N_8331,N_4447,N_5432);
and U8332 (N_8332,N_6952,N_5562);
or U8333 (N_8333,N_6245,N_6873);
nand U8334 (N_8334,N_4982,N_7854);
xnor U8335 (N_8335,N_6632,N_7326);
xor U8336 (N_8336,N_4934,N_5625);
nor U8337 (N_8337,N_7304,N_4647);
nor U8338 (N_8338,N_5284,N_7596);
nand U8339 (N_8339,N_5546,N_5786);
or U8340 (N_8340,N_7516,N_7712);
nor U8341 (N_8341,N_7299,N_7870);
or U8342 (N_8342,N_5534,N_7444);
nand U8343 (N_8343,N_5060,N_6084);
xor U8344 (N_8344,N_4442,N_6398);
nor U8345 (N_8345,N_6828,N_5777);
nand U8346 (N_8346,N_6429,N_4458);
nand U8347 (N_8347,N_5412,N_6272);
nand U8348 (N_8348,N_7427,N_5544);
xor U8349 (N_8349,N_5042,N_7970);
or U8350 (N_8350,N_6978,N_4160);
nor U8351 (N_8351,N_4913,N_6325);
and U8352 (N_8352,N_6819,N_5670);
and U8353 (N_8353,N_5606,N_5074);
nor U8354 (N_8354,N_7699,N_4836);
and U8355 (N_8355,N_7629,N_7474);
nor U8356 (N_8356,N_6534,N_7318);
or U8357 (N_8357,N_5629,N_7088);
nand U8358 (N_8358,N_7308,N_5111);
and U8359 (N_8359,N_7920,N_7743);
nor U8360 (N_8360,N_5799,N_5938);
and U8361 (N_8361,N_7277,N_6869);
and U8362 (N_8362,N_5306,N_5020);
and U8363 (N_8363,N_5741,N_5454);
nand U8364 (N_8364,N_4010,N_4888);
nor U8365 (N_8365,N_6714,N_7346);
nor U8366 (N_8366,N_4611,N_6753);
or U8367 (N_8367,N_5724,N_4307);
nor U8368 (N_8368,N_6183,N_5002);
nand U8369 (N_8369,N_5811,N_6314);
or U8370 (N_8370,N_5540,N_5990);
or U8371 (N_8371,N_5398,N_7239);
and U8372 (N_8372,N_5737,N_7606);
nor U8373 (N_8373,N_6231,N_4364);
and U8374 (N_8374,N_6814,N_4309);
nand U8375 (N_8375,N_5530,N_5173);
and U8376 (N_8376,N_4387,N_6919);
nand U8377 (N_8377,N_6914,N_4691);
nor U8378 (N_8378,N_4872,N_4586);
nor U8379 (N_8379,N_6029,N_4149);
or U8380 (N_8380,N_7614,N_5854);
xor U8381 (N_8381,N_6248,N_4584);
and U8382 (N_8382,N_4696,N_6121);
xor U8383 (N_8383,N_6785,N_5804);
and U8384 (N_8384,N_7694,N_7531);
nor U8385 (N_8385,N_5373,N_4949);
nor U8386 (N_8386,N_4308,N_7137);
nor U8387 (N_8387,N_4536,N_4766);
nand U8388 (N_8388,N_7682,N_6402);
or U8389 (N_8389,N_7199,N_4372);
and U8390 (N_8390,N_5660,N_7430);
xnor U8391 (N_8391,N_4492,N_4006);
nor U8392 (N_8392,N_6010,N_6167);
nand U8393 (N_8393,N_6721,N_5464);
nor U8394 (N_8394,N_5650,N_6803);
and U8395 (N_8395,N_5766,N_7985);
and U8396 (N_8396,N_4445,N_4979);
xor U8397 (N_8397,N_6287,N_7588);
or U8398 (N_8398,N_4181,N_7502);
xnor U8399 (N_8399,N_7031,N_6381);
nand U8400 (N_8400,N_4508,N_4233);
nor U8401 (N_8401,N_4090,N_5414);
or U8402 (N_8402,N_7859,N_6948);
nand U8403 (N_8403,N_6562,N_7262);
nand U8404 (N_8404,N_5803,N_6451);
nand U8405 (N_8405,N_5381,N_6520);
or U8406 (N_8406,N_7989,N_6988);
and U8407 (N_8407,N_6939,N_4514);
nor U8408 (N_8408,N_4826,N_4358);
nand U8409 (N_8409,N_5116,N_4127);
nand U8410 (N_8410,N_7050,N_6945);
and U8411 (N_8411,N_4831,N_6363);
or U8412 (N_8412,N_6323,N_5031);
or U8413 (N_8413,N_5611,N_7280);
xor U8414 (N_8414,N_7296,N_4635);
nor U8415 (N_8415,N_7765,N_6624);
nand U8416 (N_8416,N_6764,N_6604);
nor U8417 (N_8417,N_6349,N_7242);
and U8418 (N_8418,N_5641,N_4654);
or U8419 (N_8419,N_6809,N_7840);
nand U8420 (N_8420,N_4473,N_6894);
nor U8421 (N_8421,N_7815,N_5782);
xnor U8422 (N_8422,N_4550,N_5281);
nand U8423 (N_8423,N_6445,N_4290);
or U8424 (N_8424,N_4028,N_7829);
or U8425 (N_8425,N_7882,N_5769);
nor U8426 (N_8426,N_5000,N_4059);
xnor U8427 (N_8427,N_6082,N_5188);
nor U8428 (N_8428,N_6996,N_7172);
nand U8429 (N_8429,N_7286,N_5275);
and U8430 (N_8430,N_6505,N_6805);
or U8431 (N_8431,N_7009,N_6165);
and U8432 (N_8432,N_7036,N_5171);
or U8433 (N_8433,N_6794,N_7331);
and U8434 (N_8434,N_4397,N_5478);
nand U8435 (N_8435,N_4932,N_7788);
nand U8436 (N_8436,N_7847,N_7084);
nor U8437 (N_8437,N_4410,N_5817);
or U8438 (N_8438,N_6926,N_7373);
nor U8439 (N_8439,N_5152,N_6876);
nor U8440 (N_8440,N_4376,N_6995);
xnor U8441 (N_8441,N_7013,N_5961);
and U8442 (N_8442,N_7706,N_7732);
or U8443 (N_8443,N_6575,N_4490);
xor U8444 (N_8444,N_6715,N_5487);
nand U8445 (N_8445,N_7813,N_7826);
and U8446 (N_8446,N_5404,N_7498);
or U8447 (N_8447,N_7679,N_5503);
and U8448 (N_8448,N_5232,N_7367);
xnor U8449 (N_8449,N_6991,N_6462);
nor U8450 (N_8450,N_4179,N_5688);
and U8451 (N_8451,N_6535,N_6098);
xnor U8452 (N_8452,N_7837,N_5548);
nor U8453 (N_8453,N_7435,N_7750);
or U8454 (N_8454,N_4163,N_6185);
nand U8455 (N_8455,N_4196,N_6064);
nor U8456 (N_8456,N_7831,N_4641);
or U8457 (N_8457,N_6343,N_4779);
nor U8458 (N_8458,N_6755,N_6494);
nand U8459 (N_8459,N_7823,N_4742);
nor U8460 (N_8460,N_5126,N_6702);
nand U8461 (N_8461,N_6552,N_5119);
xor U8462 (N_8462,N_7181,N_7769);
and U8463 (N_8463,N_7856,N_6338);
nand U8464 (N_8464,N_6724,N_5880);
nand U8465 (N_8465,N_4205,N_7665);
or U8466 (N_8466,N_5656,N_6781);
or U8467 (N_8467,N_6410,N_4709);
and U8468 (N_8468,N_4964,N_7994);
nand U8469 (N_8469,N_7524,N_6362);
nor U8470 (N_8470,N_4140,N_4811);
or U8471 (N_8471,N_7287,N_7152);
and U8472 (N_8472,N_5814,N_6457);
nor U8473 (N_8473,N_6982,N_5350);
or U8474 (N_8474,N_4494,N_7581);
xor U8475 (N_8475,N_5810,N_6350);
nor U8476 (N_8476,N_4572,N_7107);
xnor U8477 (N_8477,N_5915,N_4169);
and U8478 (N_8478,N_6792,N_6734);
or U8479 (N_8479,N_5537,N_7409);
and U8480 (N_8480,N_7159,N_6239);
or U8481 (N_8481,N_5998,N_5318);
or U8482 (N_8482,N_7993,N_5353);
nand U8483 (N_8483,N_4429,N_4435);
or U8484 (N_8484,N_7707,N_5160);
nor U8485 (N_8485,N_4279,N_5755);
nor U8486 (N_8486,N_7103,N_6832);
nand U8487 (N_8487,N_5082,N_4197);
nor U8488 (N_8488,N_6292,N_4706);
and U8489 (N_8489,N_5865,N_4482);
nor U8490 (N_8490,N_6141,N_4803);
nor U8491 (N_8491,N_6378,N_4031);
nor U8492 (N_8492,N_7146,N_6001);
nand U8493 (N_8493,N_5637,N_7587);
nand U8494 (N_8494,N_4295,N_6704);
and U8495 (N_8495,N_5295,N_6008);
or U8496 (N_8496,N_5098,N_5017);
and U8497 (N_8497,N_5145,N_6806);
nor U8498 (N_8498,N_7624,N_4232);
nor U8499 (N_8499,N_6330,N_6346);
and U8500 (N_8500,N_4332,N_7664);
and U8501 (N_8501,N_6380,N_4953);
and U8502 (N_8502,N_4955,N_6521);
nand U8503 (N_8503,N_5150,N_6093);
nor U8504 (N_8504,N_5842,N_7768);
nor U8505 (N_8505,N_7909,N_4130);
and U8506 (N_8506,N_5750,N_6983);
nor U8507 (N_8507,N_5209,N_4765);
and U8508 (N_8508,N_7616,N_7321);
xnor U8509 (N_8509,N_4680,N_7893);
or U8510 (N_8510,N_6025,N_7074);
or U8511 (N_8511,N_7709,N_5687);
and U8512 (N_8512,N_6537,N_4180);
nand U8513 (N_8513,N_7205,N_5525);
nand U8514 (N_8514,N_6602,N_7449);
nand U8515 (N_8515,N_5337,N_4667);
nand U8516 (N_8516,N_7341,N_6924);
nand U8517 (N_8517,N_6332,N_4082);
nor U8518 (N_8518,N_7128,N_5083);
nand U8519 (N_8519,N_5231,N_5700);
xor U8520 (N_8520,N_6863,N_5873);
xor U8521 (N_8521,N_6046,N_4591);
xnor U8522 (N_8522,N_5245,N_6215);
nor U8523 (N_8523,N_5469,N_6765);
nand U8524 (N_8524,N_4653,N_6897);
nor U8525 (N_8525,N_6522,N_7029);
or U8526 (N_8526,N_4094,N_7314);
or U8527 (N_8527,N_5855,N_4322);
nand U8528 (N_8528,N_4644,N_5078);
and U8529 (N_8529,N_6970,N_4362);
and U8530 (N_8530,N_4991,N_6032);
or U8531 (N_8531,N_5726,N_7923);
and U8532 (N_8532,N_6836,N_7796);
nor U8533 (N_8533,N_7636,N_6054);
nor U8534 (N_8534,N_7542,N_7812);
nand U8535 (N_8535,N_5545,N_4054);
or U8536 (N_8536,N_5718,N_4527);
or U8537 (N_8537,N_7539,N_4708);
and U8538 (N_8538,N_4320,N_4915);
or U8539 (N_8539,N_7212,N_4669);
nand U8540 (N_8540,N_6357,N_4500);
or U8541 (N_8541,N_4768,N_6965);
nor U8542 (N_8542,N_5197,N_6851);
and U8543 (N_8543,N_7867,N_4154);
xnor U8544 (N_8544,N_6541,N_5049);
nor U8545 (N_8545,N_6591,N_4338);
xnor U8546 (N_8546,N_6475,N_7207);
nor U8547 (N_8547,N_7563,N_4814);
and U8548 (N_8548,N_6902,N_4495);
nand U8549 (N_8549,N_4538,N_7144);
nand U8550 (N_8550,N_5992,N_7834);
nand U8551 (N_8551,N_5613,N_6406);
nand U8552 (N_8552,N_5738,N_5367);
nand U8553 (N_8553,N_4347,N_7688);
xor U8554 (N_8554,N_6887,N_7221);
or U8555 (N_8555,N_7963,N_7169);
or U8556 (N_8556,N_6072,N_4481);
or U8557 (N_8557,N_6336,N_7265);
or U8558 (N_8558,N_5929,N_4446);
nand U8559 (N_8559,N_5137,N_6646);
and U8560 (N_8560,N_6929,N_6156);
nand U8561 (N_8561,N_7487,N_5519);
nand U8562 (N_8562,N_6568,N_7058);
and U8563 (N_8563,N_7293,N_6202);
nor U8564 (N_8564,N_4759,N_6288);
nor U8565 (N_8565,N_7090,N_5954);
or U8566 (N_8566,N_6253,N_6129);
and U8567 (N_8567,N_5131,N_6090);
or U8568 (N_8568,N_7889,N_4753);
and U8569 (N_8569,N_7654,N_6423);
or U8570 (N_8570,N_7203,N_7853);
or U8571 (N_8571,N_7023,N_4351);
nand U8572 (N_8572,N_7167,N_7206);
xor U8573 (N_8573,N_4463,N_7608);
or U8574 (N_8574,N_6316,N_6385);
nand U8575 (N_8575,N_4957,N_5221);
and U8576 (N_8576,N_7040,N_6567);
and U8577 (N_8577,N_4227,N_5893);
and U8578 (N_8578,N_7440,N_7381);
or U8579 (N_8579,N_5170,N_4734);
or U8580 (N_8580,N_5439,N_5867);
nand U8581 (N_8581,N_5767,N_5147);
and U8582 (N_8582,N_7556,N_7630);
nand U8583 (N_8583,N_4079,N_6595);
and U8584 (N_8584,N_4398,N_6334);
or U8585 (N_8585,N_7907,N_5403);
nor U8586 (N_8586,N_5913,N_4839);
and U8587 (N_8587,N_4060,N_7548);
or U8588 (N_8588,N_5936,N_5430);
xor U8589 (N_8589,N_5305,N_5361);
or U8590 (N_8590,N_6209,N_5935);
nand U8591 (N_8591,N_4311,N_7855);
or U8592 (N_8592,N_5117,N_4796);
nor U8593 (N_8593,N_5520,N_6979);
and U8594 (N_8594,N_6112,N_7661);
and U8595 (N_8595,N_6719,N_6295);
nor U8596 (N_8596,N_6324,N_5813);
or U8597 (N_8597,N_5959,N_7282);
nand U8598 (N_8598,N_6545,N_6117);
and U8599 (N_8599,N_5237,N_4904);
nand U8600 (N_8600,N_6576,N_7424);
or U8601 (N_8601,N_4870,N_5723);
nand U8602 (N_8602,N_6327,N_6153);
and U8603 (N_8603,N_7224,N_6175);
nand U8604 (N_8604,N_4631,N_4897);
nor U8605 (N_8605,N_6820,N_4158);
nand U8606 (N_8606,N_5577,N_6695);
and U8607 (N_8607,N_6546,N_7568);
xnor U8608 (N_8608,N_6666,N_5809);
nand U8609 (N_8609,N_5759,N_4749);
or U8610 (N_8610,N_7737,N_5222);
and U8611 (N_8611,N_6422,N_4235);
nor U8612 (N_8612,N_5616,N_5999);
nor U8613 (N_8613,N_4050,N_6585);
and U8614 (N_8614,N_4892,N_6891);
or U8615 (N_8615,N_4945,N_5370);
nor U8616 (N_8616,N_4225,N_7641);
and U8617 (N_8617,N_7564,N_4341);
or U8618 (N_8618,N_5986,N_7245);
or U8619 (N_8619,N_4136,N_7513);
nor U8620 (N_8620,N_7957,N_5485);
nor U8621 (N_8621,N_6396,N_6717);
nand U8622 (N_8622,N_5462,N_6470);
or U8623 (N_8623,N_7218,N_6106);
xor U8624 (N_8624,N_7374,N_4077);
nand U8625 (N_8625,N_7995,N_4066);
and U8626 (N_8626,N_4113,N_6905);
and U8627 (N_8627,N_5504,N_5183);
nor U8628 (N_8628,N_4640,N_7285);
nand U8629 (N_8629,N_5507,N_7671);
or U8630 (N_8630,N_7562,N_7836);
or U8631 (N_8631,N_4185,N_6500);
and U8632 (N_8632,N_4935,N_4520);
and U8633 (N_8633,N_7266,N_7895);
or U8634 (N_8634,N_4735,N_5829);
or U8635 (N_8635,N_4969,N_7173);
and U8636 (N_8636,N_4104,N_4874);
and U8637 (N_8637,N_4822,N_4947);
and U8638 (N_8638,N_6812,N_6203);
or U8639 (N_8639,N_4203,N_4392);
or U8640 (N_8640,N_7617,N_5626);
nor U8641 (N_8641,N_6614,N_5363);
nor U8642 (N_8642,N_7045,N_4533);
or U8643 (N_8643,N_5177,N_7247);
and U8644 (N_8644,N_4686,N_5141);
or U8645 (N_8645,N_7360,N_6921);
and U8646 (N_8646,N_5601,N_6871);
nand U8647 (N_8647,N_5692,N_6196);
or U8648 (N_8648,N_5776,N_4923);
nand U8649 (N_8649,N_5529,N_6021);
nor U8650 (N_8650,N_6967,N_6593);
or U8651 (N_8651,N_6088,N_7446);
nor U8652 (N_8652,N_7662,N_4333);
nor U8653 (N_8653,N_4095,N_4702);
nor U8654 (N_8654,N_7225,N_4737);
or U8655 (N_8655,N_6852,N_4069);
and U8656 (N_8656,N_7359,N_7721);
nor U8657 (N_8657,N_5269,N_4961);
and U8658 (N_8658,N_4521,N_4210);
nor U8659 (N_8659,N_6549,N_5238);
and U8660 (N_8660,N_4304,N_6784);
or U8661 (N_8661,N_4794,N_5791);
and U8662 (N_8662,N_5524,N_6609);
xor U8663 (N_8663,N_7760,N_6881);
nor U8664 (N_8664,N_4330,N_7607);
or U8665 (N_8665,N_4784,N_6772);
nor U8666 (N_8666,N_5438,N_6193);
or U8667 (N_8667,N_6606,N_6150);
and U8668 (N_8668,N_6810,N_7992);
and U8669 (N_8669,N_4859,N_7919);
nand U8670 (N_8670,N_7291,N_7928);
nand U8671 (N_8671,N_5674,N_7408);
or U8672 (N_8672,N_4956,N_7543);
nor U8673 (N_8673,N_6514,N_6884);
nand U8674 (N_8674,N_5934,N_6397);
and U8675 (N_8675,N_5869,N_7273);
and U8676 (N_8676,N_4426,N_7844);
xor U8677 (N_8677,N_7729,N_4264);
nand U8678 (N_8678,N_4357,N_6860);
nand U8679 (N_8679,N_5095,N_4246);
or U8680 (N_8680,N_7687,N_4367);
nand U8681 (N_8681,N_4067,N_7996);
nor U8682 (N_8682,N_6569,N_7201);
nor U8683 (N_8683,N_5598,N_6187);
and U8684 (N_8684,N_6230,N_7028);
nor U8685 (N_8685,N_7292,N_4543);
and U8686 (N_8686,N_5270,N_6172);
or U8687 (N_8687,N_4340,N_5488);
and U8688 (N_8688,N_5081,N_7366);
or U8689 (N_8689,N_7486,N_7891);
and U8690 (N_8690,N_4088,N_7819);
or U8691 (N_8691,N_6159,N_6859);
or U8692 (N_8692,N_7485,N_7881);
or U8693 (N_8693,N_5467,N_5872);
or U8694 (N_8694,N_5590,N_7646);
xnor U8695 (N_8695,N_6265,N_6177);
and U8696 (N_8696,N_5436,N_4172);
or U8697 (N_8697,N_7595,N_6390);
or U8698 (N_8698,N_7975,N_4522);
and U8699 (N_8699,N_4857,N_4689);
or U8700 (N_8700,N_5301,N_6775);
nand U8701 (N_8701,N_4182,N_4770);
xor U8702 (N_8702,N_7027,N_7098);
and U8703 (N_8703,N_6264,N_6962);
or U8704 (N_8704,N_6143,N_7968);
or U8705 (N_8705,N_7572,N_6558);
nor U8706 (N_8706,N_6364,N_6807);
or U8707 (N_8707,N_7399,N_5591);
or U8708 (N_8708,N_7753,N_6510);
and U8709 (N_8709,N_4711,N_7310);
and U8710 (N_8710,N_5647,N_4230);
nor U8711 (N_8711,N_6688,N_5392);
or U8712 (N_8712,N_5331,N_5757);
or U8713 (N_8713,N_6701,N_5317);
nor U8714 (N_8714,N_7204,N_6053);
and U8715 (N_8715,N_6014,N_5032);
xor U8716 (N_8716,N_7489,N_4037);
and U8717 (N_8717,N_6507,N_6415);
xor U8718 (N_8718,N_5154,N_5005);
or U8719 (N_8719,N_6079,N_7007);
and U8720 (N_8720,N_6787,N_6076);
or U8721 (N_8721,N_4698,N_5158);
or U8722 (N_8722,N_4106,N_7357);
xnor U8723 (N_8723,N_6615,N_5788);
and U8724 (N_8724,N_5673,N_7122);
nor U8725 (N_8725,N_4887,N_4005);
or U8726 (N_8726,N_7323,N_6999);
or U8727 (N_8727,N_5994,N_6280);
and U8728 (N_8728,N_6684,N_7672);
nand U8729 (N_8729,N_6275,N_4835);
nand U8730 (N_8730,N_4380,N_6430);
nand U8731 (N_8731,N_5827,N_6105);
and U8732 (N_8732,N_4725,N_4569);
or U8733 (N_8733,N_6307,N_6131);
xor U8734 (N_8734,N_4620,N_4187);
nand U8735 (N_8735,N_5501,N_5618);
or U8736 (N_8736,N_4378,N_5427);
nor U8737 (N_8737,N_5087,N_4083);
or U8738 (N_8738,N_6051,N_7814);
and U8739 (N_8739,N_5122,N_6527);
or U8740 (N_8740,N_7673,N_6861);
nor U8741 (N_8741,N_5987,N_5617);
nor U8742 (N_8742,N_4229,N_5271);
nor U8743 (N_8743,N_7157,N_7525);
or U8744 (N_8744,N_6866,N_4697);
nor U8745 (N_8745,N_4548,N_5289);
and U8746 (N_8746,N_7728,N_7770);
nand U8747 (N_8747,N_7124,N_7092);
nor U8748 (N_8748,N_6917,N_6133);
nand U8749 (N_8749,N_7263,N_5531);
nor U8750 (N_8750,N_4914,N_4016);
or U8751 (N_8751,N_4912,N_5851);
nand U8752 (N_8752,N_5428,N_7386);
nand U8753 (N_8753,N_6136,N_5386);
and U8754 (N_8754,N_5008,N_5863);
and U8755 (N_8755,N_7930,N_5062);
nand U8756 (N_8756,N_6221,N_5067);
and U8757 (N_8757,N_6019,N_4688);
or U8758 (N_8758,N_4489,N_6130);
xnor U8759 (N_8759,N_4027,N_5864);
and U8760 (N_8760,N_4930,N_4746);
or U8761 (N_8761,N_4539,N_5056);
or U8762 (N_8762,N_4577,N_5972);
or U8763 (N_8763,N_7691,N_5424);
and U8764 (N_8764,N_7441,N_6270);
nand U8765 (N_8765,N_5897,N_5037);
nand U8766 (N_8766,N_7142,N_4070);
and U8767 (N_8767,N_7951,N_5441);
nand U8768 (N_8768,N_7089,N_4762);
nor U8769 (N_8769,N_6282,N_5908);
xnor U8770 (N_8770,N_4040,N_4558);
or U8771 (N_8771,N_6874,N_7118);
nand U8772 (N_8772,N_7491,N_6946);
nand U8773 (N_8773,N_4940,N_6326);
nor U8774 (N_8774,N_5073,N_7132);
nand U8775 (N_8775,N_5257,N_5389);
or U8776 (N_8776,N_7777,N_6827);
nand U8777 (N_8777,N_4023,N_4928);
or U8778 (N_8778,N_5368,N_7475);
nor U8779 (N_8779,N_5566,N_4972);
xor U8780 (N_8780,N_6022,N_7945);
and U8781 (N_8781,N_5779,N_6162);
or U8782 (N_8782,N_4743,N_4469);
and U8783 (N_8783,N_4058,N_7785);
or U8784 (N_8784,N_5559,N_7061);
nor U8785 (N_8785,N_7731,N_5310);
and U8786 (N_8786,N_7404,N_5861);
or U8787 (N_8787,N_7217,N_4906);
and U8788 (N_8788,N_7419,N_6400);
nand U8789 (N_8789,N_5358,N_5155);
and U8790 (N_8790,N_4350,N_7035);
nand U8791 (N_8791,N_4911,N_6573);
nor U8792 (N_8792,N_7904,N_4091);
nand U8793 (N_8793,N_4624,N_4880);
or U8794 (N_8794,N_7303,N_6038);
nand U8795 (N_8795,N_6698,N_6186);
nor U8796 (N_8796,N_5093,N_7898);
and U8797 (N_8797,N_4864,N_5762);
nand U8798 (N_8798,N_6749,N_7739);
or U8799 (N_8799,N_6391,N_7848);
nand U8800 (N_8800,N_7632,N_4096);
nand U8801 (N_8801,N_7147,N_5815);
nand U8802 (N_8802,N_5051,N_4551);
xor U8803 (N_8803,N_5592,N_6865);
nand U8804 (N_8804,N_6880,N_7751);
and U8805 (N_8805,N_4804,N_6841);
nand U8806 (N_8806,N_5172,N_5644);
or U8807 (N_8807,N_7470,N_4976);
and U8808 (N_8808,N_7827,N_5535);
nor U8809 (N_8809,N_7634,N_4206);
nand U8810 (N_8810,N_7763,N_7571);
and U8811 (N_8811,N_4510,N_4954);
and U8812 (N_8812,N_6598,N_7352);
and U8813 (N_8813,N_7176,N_5678);
and U8814 (N_8814,N_7702,N_4626);
nand U8815 (N_8815,N_4810,N_6365);
and U8816 (N_8816,N_6530,N_7180);
or U8817 (N_8817,N_6783,N_5128);
and U8818 (N_8818,N_4361,N_7003);
nand U8819 (N_8819,N_6170,N_6309);
xnor U8820 (N_8820,N_7214,N_4416);
nor U8821 (N_8821,N_6928,N_5195);
nor U8822 (N_8822,N_4756,N_7746);
nand U8823 (N_8823,N_5243,N_6786);
and U8824 (N_8824,N_4281,N_7875);
and U8825 (N_8825,N_7982,N_6867);
nand U8826 (N_8826,N_7480,N_7369);
nand U8827 (N_8827,N_4298,N_5578);
nand U8828 (N_8828,N_7021,N_6174);
or U8829 (N_8829,N_5835,N_4553);
and U8830 (N_8830,N_6726,N_4903);
or U8831 (N_8831,N_7426,N_5866);
and U8832 (N_8832,N_6199,N_6872);
or U8833 (N_8833,N_4331,N_6405);
nand U8834 (N_8834,N_4607,N_5845);
or U8835 (N_8835,N_7131,N_7567);
nand U8836 (N_8836,N_5679,N_5011);
and U8837 (N_8837,N_4455,N_7481);
nor U8838 (N_8838,N_7042,N_5491);
and U8839 (N_8839,N_7817,N_4457);
or U8840 (N_8840,N_5248,N_6625);
or U8841 (N_8841,N_7741,N_7230);
and U8842 (N_8842,N_6151,N_7194);
nor U8843 (N_8843,N_5928,N_5556);
or U8844 (N_8844,N_7888,N_5806);
nand U8845 (N_8845,N_6501,N_4433);
xnor U8846 (N_8846,N_4135,N_4840);
and U8847 (N_8847,N_5982,N_6488);
xor U8848 (N_8848,N_5308,N_5898);
or U8849 (N_8849,N_7320,N_6839);
nand U8850 (N_8850,N_7620,N_5834);
or U8851 (N_8851,N_4452,N_4454);
or U8852 (N_8852,N_4354,N_4701);
nand U8853 (N_8853,N_5579,N_6588);
and U8854 (N_8854,N_4965,N_5635);
xnor U8855 (N_8855,N_7371,N_4039);
nor U8856 (N_8856,N_4809,N_5071);
xnor U8857 (N_8857,N_4155,N_4530);
xor U8858 (N_8858,N_7615,N_7005);
nor U8859 (N_8859,N_6748,N_5288);
or U8860 (N_8860,N_5228,N_5760);
or U8861 (N_8861,N_5933,N_5752);
or U8862 (N_8862,N_7100,N_4269);
nor U8863 (N_8863,N_7037,N_5838);
xnor U8864 (N_8864,N_4936,N_5405);
or U8865 (N_8865,N_7134,N_6466);
or U8866 (N_8866,N_5973,N_6862);
nor U8867 (N_8867,N_4910,N_4334);
nand U8868 (N_8868,N_6298,N_7469);
nor U8869 (N_8869,N_5502,N_4797);
nor U8870 (N_8870,N_5181,N_4739);
nor U8871 (N_8871,N_5509,N_4164);
or U8872 (N_8872,N_6605,N_7034);
and U8873 (N_8873,N_4524,N_6563);
nand U8874 (N_8874,N_6146,N_5716);
and U8875 (N_8875,N_5216,N_4944);
nand U8876 (N_8876,N_4150,N_4851);
nor U8877 (N_8877,N_4395,N_7740);
nand U8878 (N_8878,N_4597,N_6208);
and U8879 (N_8879,N_5100,N_6313);
or U8880 (N_8880,N_4744,N_4432);
and U8881 (N_8881,N_4926,N_5180);
nand U8882 (N_8882,N_6227,N_7897);
and U8883 (N_8883,N_6303,N_4863);
xnor U8884 (N_8884,N_6941,N_4491);
nor U8885 (N_8885,N_7908,N_5924);
nand U8886 (N_8886,N_5024,N_5324);
or U8887 (N_8887,N_5239,N_7971);
or U8888 (N_8888,N_7237,N_5483);
nor U8889 (N_8889,N_6761,N_7148);
or U8890 (N_8890,N_7414,N_6472);
or U8891 (N_8891,N_6178,N_6623);
nor U8892 (N_8892,N_4596,N_5995);
xnor U8893 (N_8893,N_4501,N_6284);
or U8894 (N_8894,N_5980,N_4916);
nand U8895 (N_8895,N_4328,N_6992);
nor U8896 (N_8896,N_5223,N_7804);
nor U8897 (N_8897,N_4190,N_6073);
xor U8898 (N_8898,N_4422,N_5481);
nand U8899 (N_8899,N_6526,N_7415);
xor U8900 (N_8900,N_7797,N_4534);
or U8901 (N_8901,N_5425,N_7410);
nor U8902 (N_8902,N_5894,N_5300);
or U8903 (N_8903,N_7253,N_4450);
and U8904 (N_8904,N_4504,N_7060);
or U8905 (N_8905,N_7873,N_5156);
or U8906 (N_8906,N_7948,N_5484);
and U8907 (N_8907,N_5130,N_5858);
nand U8908 (N_8908,N_4989,N_6559);
nand U8909 (N_8909,N_5889,N_7758);
and U8910 (N_8910,N_7528,N_4383);
or U8911 (N_8911,N_4717,N_7190);
or U8912 (N_8912,N_7054,N_5802);
or U8913 (N_8913,N_4486,N_5512);
and U8914 (N_8914,N_7649,N_4813);
and U8915 (N_8915,N_6125,N_7720);
or U8916 (N_8916,N_4297,N_6655);
or U8917 (N_8917,N_4282,N_5391);
nor U8918 (N_8918,N_4853,N_6896);
nor U8919 (N_8919,N_6729,N_5311);
or U8920 (N_8920,N_7078,N_5319);
or U8921 (N_8921,N_6620,N_6565);
xor U8922 (N_8922,N_5586,N_7033);
or U8923 (N_8923,N_5036,N_5839);
or U8924 (N_8924,N_7925,N_6042);
or U8925 (N_8925,N_5084,N_5471);
xor U8926 (N_8926,N_4532,N_7436);
or U8927 (N_8927,N_5486,N_5595);
nor U8928 (N_8928,N_4990,N_6176);
xnor U8929 (N_8929,N_5508,N_4973);
nand U8930 (N_8930,N_4650,N_6736);
nor U8931 (N_8931,N_6524,N_7226);
or U8932 (N_8932,N_4310,N_7601);
nor U8933 (N_8933,N_7583,N_5229);
nand U8934 (N_8934,N_7425,N_7111);
or U8935 (N_8935,N_7213,N_5580);
nor U8936 (N_8936,N_7657,N_6086);
and U8937 (N_8937,N_6712,N_6912);
nand U8938 (N_8938,N_4886,N_5161);
xnor U8939 (N_8939,N_6320,N_4962);
nand U8940 (N_8940,N_5558,N_5103);
or U8941 (N_8941,N_4042,N_6440);
nand U8942 (N_8942,N_7612,N_4119);
nor U8943 (N_8943,N_4161,N_4829);
and U8944 (N_8944,N_6124,N_4901);
xor U8945 (N_8945,N_4578,N_4718);
nand U8946 (N_8946,N_4740,N_5101);
nor U8947 (N_8947,N_7405,N_7471);
or U8948 (N_8948,N_5664,N_7227);
nand U8949 (N_8949,N_7354,N_4488);
nor U8950 (N_8950,N_4211,N_6341);
nand U8951 (N_8951,N_7208,N_7468);
nand U8952 (N_8952,N_6249,N_4868);
or U8953 (N_8953,N_5120,N_5457);
or U8954 (N_8954,N_4516,N_4557);
nor U8955 (N_8955,N_4080,N_5879);
or U8956 (N_8956,N_7138,N_6092);
and U8957 (N_8957,N_7391,N_7302);
or U8958 (N_8958,N_7839,N_4821);
and U8959 (N_8959,N_5712,N_6109);
nor U8960 (N_8960,N_5539,N_6246);
or U8961 (N_8961,N_6347,N_7272);
xor U8962 (N_8962,N_4507,N_6401);
nor U8963 (N_8963,N_5680,N_4776);
or U8964 (N_8964,N_5906,N_6980);
nand U8965 (N_8965,N_4598,N_7101);
nand U8966 (N_8966,N_4052,N_4366);
nand U8967 (N_8967,N_4661,N_7311);
nand U8968 (N_8968,N_7822,N_7149);
nor U8969 (N_8969,N_6310,N_6194);
nand U8970 (N_8970,N_6953,N_5140);
nand U8971 (N_8971,N_7943,N_6889);
or U8972 (N_8972,N_4355,N_6368);
and U8973 (N_8973,N_4993,N_7860);
nand U8974 (N_8974,N_6788,N_5076);
nand U8975 (N_8975,N_7497,N_7141);
nor U8976 (N_8976,N_6743,N_4602);
xnor U8977 (N_8977,N_6490,N_5468);
or U8978 (N_8978,N_6431,N_4841);
nor U8979 (N_8979,N_6528,N_6976);
nor U8980 (N_8980,N_4121,N_4896);
and U8981 (N_8981,N_4389,N_4778);
nand U8982 (N_8982,N_4513,N_5728);
nor U8983 (N_8983,N_6594,N_4406);
and U8984 (N_8984,N_7862,N_5215);
nand U8985 (N_8985,N_7215,N_6838);
and U8986 (N_8986,N_6998,N_5044);
or U8987 (N_8987,N_5422,N_5725);
xor U8988 (N_8988,N_4605,N_5408);
nand U8989 (N_8989,N_6848,N_6561);
and U8990 (N_8990,N_4425,N_7799);
nor U8991 (N_8991,N_7106,N_6818);
or U8992 (N_8992,N_7108,N_5652);
or U8993 (N_8993,N_5853,N_5940);
or U8994 (N_8994,N_6108,N_6290);
nor U8995 (N_8995,N_4283,N_4858);
or U8996 (N_8996,N_6222,N_4339);
nor U8997 (N_8997,N_4838,N_4875);
nor U8998 (N_8998,N_6835,N_6044);
or U8999 (N_8999,N_5596,N_5165);
or U9000 (N_9000,N_7380,N_7637);
xnor U9001 (N_9001,N_6758,N_4343);
xnor U9002 (N_9002,N_7325,N_6741);
or U9003 (N_9003,N_6427,N_6189);
or U9004 (N_9004,N_4537,N_4924);
nand U9005 (N_9005,N_4665,N_5211);
and U9006 (N_9006,N_7501,N_6933);
nor U9007 (N_9007,N_6252,N_4736);
xor U9008 (N_9008,N_4141,N_7986);
nand U9009 (N_9009,N_7917,N_5709);
and U9010 (N_9010,N_4301,N_5476);
nand U9011 (N_9011,N_7642,N_6986);
nor U9012 (N_9012,N_6716,N_6450);
xor U9013 (N_9013,N_4373,N_7674);
and U9014 (N_9014,N_5628,N_6171);
nor U9015 (N_9015,N_5151,N_6013);
and U9016 (N_9016,N_4047,N_5742);
nand U9017 (N_9017,N_7838,N_5667);
xor U9018 (N_9018,N_4986,N_5798);
nor U9019 (N_9019,N_6074,N_4526);
nor U9020 (N_9020,N_5303,N_6045);
and U9021 (N_9021,N_6161,N_5472);
or U9022 (N_9022,N_4467,N_7744);
and U9023 (N_9023,N_6067,N_6491);
or U9024 (N_9024,N_4788,N_7461);
nand U9025 (N_9025,N_4782,N_7530);
or U9026 (N_9026,N_5903,N_7234);
nand U9027 (N_9027,N_4240,N_5072);
nor U9028 (N_9028,N_7343,N_5298);
nor U9029 (N_9029,N_5768,N_4726);
or U9030 (N_9030,N_5192,N_7990);
and U9031 (N_9031,N_5109,N_7179);
or U9032 (N_9032,N_5614,N_6529);
nor U9033 (N_9033,N_7667,N_6922);
or U9034 (N_9034,N_7887,N_6119);
nor U9035 (N_9035,N_6152,N_7462);
nand U9036 (N_9036,N_7393,N_4280);
and U9037 (N_9037,N_4825,N_6069);
or U9038 (N_9038,N_7663,N_4068);
or U9039 (N_9039,N_4806,N_7896);
xnor U9040 (N_9040,N_6345,N_4984);
nor U9041 (N_9041,N_6693,N_6808);
and U9042 (N_9042,N_6738,N_5105);
nand U9043 (N_9043,N_4695,N_7279);
xnor U9044 (N_9044,N_6328,N_5045);
or U9045 (N_9045,N_5816,N_5437);
and U9046 (N_9046,N_7949,N_5159);
or U9047 (N_9047,N_7289,N_5380);
or U9048 (N_9048,N_6654,N_6005);
or U9049 (N_9049,N_6540,N_7241);
nand U9050 (N_9050,N_5778,N_6627);
or U9051 (N_9051,N_6372,N_6757);
nor U9052 (N_9052,N_6640,N_4663);
or U9053 (N_9053,N_7322,N_7375);
and U9054 (N_9054,N_4682,N_7866);
nor U9055 (N_9055,N_7677,N_6774);
xnor U9056 (N_9056,N_5495,N_4509);
and U9057 (N_9057,N_5242,N_6158);
and U9058 (N_9058,N_6517,N_5541);
nand U9059 (N_9059,N_7125,N_7238);
nand U9060 (N_9060,N_5025,N_7959);
and U9061 (N_9061,N_5136,N_6935);
nand U9062 (N_9062,N_6667,N_6974);
and U9063 (N_9063,N_5143,N_6981);
or U9064 (N_9064,N_5251,N_4220);
or U9065 (N_9065,N_7466,N_5344);
and U9066 (N_9066,N_6048,N_6426);
nor U9067 (N_9067,N_6950,N_5584);
and U9068 (N_9068,N_5210,N_7365);
and U9069 (N_9069,N_5246,N_6637);
xnor U9070 (N_9070,N_7189,N_7490);
nand U9071 (N_9071,N_5698,N_4917);
nor U9072 (N_9072,N_5805,N_6777);
nor U9073 (N_9073,N_4377,N_6636);
xor U9074 (N_9074,N_5330,N_4120);
nand U9075 (N_9075,N_6344,N_4390);
and U9076 (N_9076,N_7257,N_7183);
nor U9077 (N_9077,N_5400,N_5115);
nor U9078 (N_9078,N_6870,N_5290);
or U9079 (N_9079,N_6997,N_5038);
nor U9080 (N_9080,N_4288,N_5797);
or U9081 (N_9081,N_4807,N_4036);
and U9082 (N_9082,N_7921,N_4760);
nand U9083 (N_9083,N_7809,N_7565);
nor U9084 (N_9084,N_4177,N_5458);
nand U9085 (N_9085,N_6120,N_7547);
or U9086 (N_9086,N_6148,N_6875);
or U9087 (N_9087,N_7174,N_7313);
or U9088 (N_9088,N_7987,N_4842);
xnor U9089 (N_9089,N_4724,N_6692);
or U9090 (N_9090,N_4204,N_6097);
xnor U9091 (N_9091,N_7353,N_6493);
nand U9092 (N_9092,N_6411,N_6459);
nand U9093 (N_9093,N_4974,N_6780);
or U9094 (N_9094,N_6498,N_5343);
and U9095 (N_9095,N_4978,N_5567);
xor U9096 (N_9096,N_4854,N_4019);
nor U9097 (N_9097,N_7254,N_7080);
nor U9098 (N_9098,N_7690,N_5607);
or U9099 (N_9099,N_6608,N_4642);
nor U9100 (N_9100,N_5771,N_5456);
and U9101 (N_9101,N_5121,N_6496);
nand U9102 (N_9102,N_5826,N_7594);
nand U9103 (N_9103,N_5399,N_4720);
and U9104 (N_9104,N_7538,N_6660);
and U9105 (N_9105,N_6675,N_4792);
nand U9106 (N_9106,N_6356,N_5279);
nand U9107 (N_9107,N_4787,N_6389);
nor U9108 (N_9108,N_5010,N_6497);
or U9109 (N_9109,N_4114,N_7645);
and U9110 (N_9110,N_5843,N_7370);
nand U9111 (N_9111,N_7072,N_6854);
xnor U9112 (N_9112,N_7438,N_6539);
nor U9113 (N_9113,N_4571,N_5594);
xnor U9114 (N_9114,N_7730,N_6759);
nor U9115 (N_9115,N_4819,N_6337);
nand U9116 (N_9116,N_4922,N_5329);
and U9117 (N_9117,N_6868,N_4587);
and U9118 (N_9118,N_5717,N_6024);
or U9119 (N_9119,N_7520,N_5751);
nand U9120 (N_9120,N_4981,N_5917);
nand U9121 (N_9121,N_7093,N_5547);
or U9122 (N_9122,N_6638,N_4441);
and U9123 (N_9123,N_6904,N_5876);
nor U9124 (N_9124,N_6532,N_7886);
and U9125 (N_9125,N_6134,N_5807);
nor U9126 (N_9126,N_5730,N_5703);
and U9127 (N_9127,N_7609,N_7197);
nand U9128 (N_9128,N_4592,N_6669);
nand U9129 (N_9129,N_7196,N_7790);
and U9130 (N_9130,N_6737,N_4137);
and U9131 (N_9131,N_7340,N_6191);
nor U9132 (N_9132,N_4649,N_5977);
or U9133 (N_9133,N_7505,N_4999);
or U9134 (N_9134,N_6085,N_7114);
and U9135 (N_9135,N_4167,N_7017);
nor U9136 (N_9136,N_5983,N_6274);
nor U9137 (N_9137,N_5267,N_7559);
or U9138 (N_9138,N_7264,N_5553);
nand U9139 (N_9139,N_7997,N_4194);
nand U9140 (N_9140,N_5953,N_6113);
and U9141 (N_9141,N_7246,N_6613);
and U9142 (N_9142,N_6647,N_6066);
nand U9143 (N_9143,N_7452,N_4555);
and U9144 (N_9144,N_7478,N_4348);
nor U9145 (N_9145,N_7899,N_5012);
and U9146 (N_9146,N_5477,N_7097);
xnor U9147 (N_9147,N_4239,N_7158);
nand U9148 (N_9148,N_7465,N_5862);
and U9149 (N_9149,N_7575,N_6665);
xor U9150 (N_9150,N_5993,N_5114);
nand U9151 (N_9151,N_7056,N_5654);
and U9152 (N_9152,N_5016,N_5421);
or U9153 (N_9153,N_7874,N_7852);
nor U9154 (N_9154,N_7117,N_4329);
and U9155 (N_9155,N_5684,N_5532);
or U9156 (N_9156,N_7300,N_4252);
nand U9157 (N_9157,N_4188,N_6312);
nor U9158 (N_9158,N_7504,N_7079);
nor U9159 (N_9159,N_6283,N_7619);
and U9160 (N_9160,N_4245,N_4250);
nand U9161 (N_9161,N_4275,N_5960);
nor U9162 (N_9162,N_7828,N_4259);
nor U9163 (N_9163,N_4565,N_4579);
nand U9164 (N_9164,N_5658,N_6257);
or U9165 (N_9165,N_7428,N_5642);
nor U9166 (N_9166,N_6267,N_4087);
or U9167 (N_9167,N_7362,N_4846);
xor U9168 (N_9168,N_4907,N_6080);
nand U9169 (N_9169,N_5413,N_7332);
nand U9170 (N_9170,N_5448,N_5686);
nor U9171 (N_9171,N_7249,N_5773);
and U9172 (N_9172,N_6055,N_7198);
nor U9173 (N_9173,N_6543,N_5849);
nand U9174 (N_9174,N_7981,N_4576);
or U9175 (N_9175,N_6574,N_4370);
nand U9176 (N_9176,N_6089,N_5273);
or U9177 (N_9177,N_5713,N_5327);
nand U9178 (N_9178,N_6409,N_7910);
nand U9179 (N_9179,N_5634,N_5446);
nand U9180 (N_9180,N_5627,N_5922);
nor U9181 (N_9181,N_5055,N_6699);
and U9182 (N_9182,N_6460,N_7939);
and U9183 (N_9183,N_7864,N_7389);
nor U9184 (N_9184,N_7892,N_7964);
or U9185 (N_9185,N_4883,N_7000);
xor U9186 (N_9186,N_7055,N_6182);
or U9187 (N_9187,N_5514,N_5538);
nand U9188 (N_9188,N_6920,N_4400);
and U9189 (N_9189,N_4061,N_7175);
and U9190 (N_9190,N_4011,N_6012);
or U9191 (N_9191,N_5204,N_5326);
nand U9192 (N_9192,N_7810,N_6732);
nor U9193 (N_9193,N_5689,N_7600);
nor U9194 (N_9194,N_6895,N_7019);
nand U9195 (N_9195,N_4267,N_6584);
or U9196 (N_9196,N_6725,N_7611);
nand U9197 (N_9197,N_5314,N_4908);
nor U9198 (N_9198,N_7726,N_7434);
nor U9199 (N_9199,N_6416,N_4111);
and U9200 (N_9200,N_5410,N_5046);
nor U9201 (N_9201,N_6659,N_6731);
or U9202 (N_9202,N_7578,N_6095);
or U9203 (N_9203,N_5402,N_4581);
nor U9204 (N_9204,N_6201,N_4585);
and U9205 (N_9205,N_6278,N_7689);
nand U9206 (N_9206,N_5198,N_5619);
and U9207 (N_9207,N_4967,N_7710);
nand U9208 (N_9208,N_6930,N_5199);
or U9209 (N_9209,N_4369,N_7579);
and U9210 (N_9210,N_6023,N_5283);
xor U9211 (N_9211,N_6373,N_7509);
nand U9212 (N_9212,N_6449,N_5206);
nand U9213 (N_9213,N_7644,N_5754);
nor U9214 (N_9214,N_5157,N_7902);
nand U9215 (N_9215,N_5035,N_5292);
or U9216 (N_9216,N_5857,N_6118);
nor U9217 (N_9217,N_6511,N_4209);
nor U9218 (N_9218,N_5470,N_6020);
xor U9219 (N_9219,N_5765,N_7482);
and U9220 (N_9220,N_7057,N_5030);
xnor U9221 (N_9221,N_6492,N_4656);
nor U9222 (N_9222,N_6599,N_6369);
nand U9223 (N_9223,N_6885,N_5341);
or U9224 (N_9224,N_6135,N_6340);
or U9225 (N_9225,N_4730,N_4951);
or U9226 (N_9226,N_6816,N_5790);
xnor U9227 (N_9227,N_4200,N_4015);
nor U9228 (N_9228,N_4174,N_5066);
nor U9229 (N_9229,N_6291,N_4678);
or U9230 (N_9230,N_4900,N_6708);
and U9231 (N_9231,N_6849,N_6768);
or U9232 (N_9232,N_4349,N_6718);
nand U9233 (N_9233,N_7235,N_4719);
and U9234 (N_9234,N_4487,N_7507);
and U9235 (N_9235,N_7590,N_4589);
nand U9236 (N_9236,N_7526,N_5697);
xnor U9237 (N_9237,N_7533,N_5743);
or U9238 (N_9238,N_7573,N_4438);
and U9239 (N_9239,N_4394,N_5490);
nand U9240 (N_9240,N_7477,N_5874);
nand U9241 (N_9241,N_4860,N_4327);
nand U9242 (N_9242,N_5576,N_7297);
and U9243 (N_9243,N_4518,N_7719);
and U9244 (N_9244,N_6016,N_4599);
and U9245 (N_9245,N_7411,N_4292);
nor U9246 (N_9246,N_5792,N_7894);
xor U9247 (N_9247,N_7582,N_6586);
nand U9248 (N_9248,N_6882,N_6437);
xor U9249 (N_9249,N_6403,N_7211);
or U9250 (N_9250,N_5054,N_5942);
or U9251 (N_9251,N_7792,N_6607);
or U9252 (N_9252,N_7734,N_7459);
and U9253 (N_9253,N_5497,N_5118);
nand U9254 (N_9254,N_6892,N_5609);
nand U9255 (N_9255,N_4671,N_7049);
xnor U9256 (N_9256,N_7499,N_4503);
or U9257 (N_9257,N_6566,N_6756);
or U9258 (N_9258,N_4198,N_7417);
nor U9259 (N_9259,N_5075,N_5240);
nand U9260 (N_9260,N_4226,N_4081);
nand U9261 (N_9261,N_4436,N_5320);
nor U9262 (N_9262,N_5787,N_4747);
or U9263 (N_9263,N_7178,N_7070);
nor U9264 (N_9264,N_5264,N_6181);
nand U9265 (N_9265,N_5034,N_6036);
or U9266 (N_9266,N_6297,N_4112);
and U9267 (N_9267,N_5297,N_4251);
nor U9268 (N_9268,N_5174,N_6486);
nand U9269 (N_9269,N_4078,N_7163);
xnor U9270 (N_9270,N_4302,N_7983);
nand U9271 (N_9271,N_4681,N_4434);
or U9272 (N_9272,N_7514,N_4470);
nand U9273 (N_9273,N_5226,N_7808);
nand U9274 (N_9274,N_7110,N_4633);
xnor U9275 (N_9275,N_5409,N_5557);
or U9276 (N_9276,N_4977,N_7395);
or U9277 (N_9277,N_6329,N_5739);
nor U9278 (N_9278,N_4938,N_6122);
or U9279 (N_9279,N_6513,N_4228);
nand U9280 (N_9280,N_7675,N_4471);
and U9281 (N_9281,N_7544,N_4248);
or U9282 (N_9282,N_5085,N_4303);
xor U9283 (N_9283,N_7316,N_7589);
nand U9284 (N_9284,N_6682,N_7068);
or U9285 (N_9285,N_6592,N_7455);
or U9286 (N_9286,N_4353,N_7063);
or U9287 (N_9287,N_4270,N_4499);
and U9288 (N_9288,N_5169,N_6845);
nor U9289 (N_9289,N_6811,N_7756);
nor U9290 (N_9290,N_4946,N_6940);
or U9291 (N_9291,N_7610,N_4996);
nand U9292 (N_9292,N_7094,N_5356);
xor U9293 (N_9293,N_4115,N_6139);
or U9294 (N_9294,N_7802,N_6407);
nand U9295 (N_9295,N_5969,N_6739);
and U9296 (N_9296,N_4193,N_6233);
xor U9297 (N_9297,N_7355,N_6436);
nand U9298 (N_9298,N_4876,N_6308);
and U9299 (N_9299,N_5944,N_6656);
nand U9300 (N_9300,N_5124,N_6434);
nor U9301 (N_9301,N_6195,N_4800);
nor U9302 (N_9302,N_7806,N_7448);
nor U9303 (N_9303,N_5474,N_7143);
nor U9304 (N_9304,N_6062,N_5304);
and U9305 (N_9305,N_7220,N_7351);
nand U9306 (N_9306,N_6661,N_4142);
and U9307 (N_9307,N_7605,N_4419);
nand U9308 (N_9308,N_6626,N_6634);
nor U9309 (N_9309,N_5939,N_7119);
nand U9310 (N_9310,N_6643,N_6294);
or U9311 (N_9311,N_4497,N_6523);
xnor U9312 (N_9312,N_5134,N_7317);
xor U9313 (N_9313,N_4265,N_5465);
or U9314 (N_9314,N_7772,N_4065);
nand U9315 (N_9315,N_4092,N_7191);
nand U9316 (N_9316,N_5104,N_7841);
and U9317 (N_9317,N_7926,N_7924);
xor U9318 (N_9318,N_7961,N_4478);
and U9319 (N_9319,N_6421,N_4738);
xnor U9320 (N_9320,N_6377,N_7240);
or U9321 (N_9321,N_5459,N_4563);
xor U9322 (N_9322,N_7081,N_5089);
xor U9323 (N_9323,N_5800,N_5254);
and U9324 (N_9324,N_5981,N_6676);
or U9325 (N_9325,N_4995,N_6043);
xnor U9326 (N_9326,N_5932,N_5018);
and U9327 (N_9327,N_5651,N_6944);
nand U9328 (N_9328,N_5573,N_5092);
or U9329 (N_9329,N_7783,N_6414);
or U9330 (N_9330,N_7281,N_7244);
nor U9331 (N_9331,N_6355,N_4375);
and U9332 (N_9332,N_5312,N_4030);
or U9333 (N_9333,N_5342,N_7512);
nor U9334 (N_9334,N_7685,N_4637);
and U9335 (N_9335,N_5622,N_6621);
and U9336 (N_9336,N_6234,N_5683);
xor U9337 (N_9337,N_5930,N_6703);
or U9338 (N_9338,N_4128,N_7536);
nand U9339 (N_9339,N_4741,N_7383);
and U9340 (N_9340,N_7126,N_5882);
and U9341 (N_9341,N_5549,N_5565);
or U9342 (N_9342,N_4843,N_4672);
and U9343 (N_9343,N_7635,N_4498);
or U9344 (N_9344,N_5886,N_6473);
nand U9345 (N_9345,N_4902,N_7735);
xnor U9346 (N_9346,N_4342,N_6007);
nor U9347 (N_9347,N_5636,N_5282);
nand U9348 (N_9348,N_7116,N_5498);
nand U9349 (N_9349,N_6099,N_6474);
and U9350 (N_9350,N_6366,N_6533);
xor U9351 (N_9351,N_6673,N_4437);
and U9352 (N_9352,N_5293,N_7655);
nor U9353 (N_9353,N_7915,N_7255);
nand U9354 (N_9354,N_7121,N_4664);
nand U9355 (N_9355,N_6315,N_4781);
and U9356 (N_9356,N_7156,N_5962);
nor U9357 (N_9357,N_6589,N_6696);
and U9358 (N_9358,N_5885,N_4003);
and U9359 (N_9359,N_5233,N_7969);
or U9360 (N_9360,N_5785,N_6037);
nor U9361 (N_9361,N_6374,N_6713);
or U9362 (N_9362,N_6856,N_7379);
nand U9363 (N_9363,N_6681,N_6078);
or U9364 (N_9364,N_7243,N_4009);
or U9365 (N_9365,N_7593,N_5931);
nor U9366 (N_9366,N_4430,N_7521);
or U9367 (N_9367,N_4795,N_6205);
or U9368 (N_9368,N_6481,N_4882);
nand U9369 (N_9369,N_5325,N_5004);
nand U9370 (N_9370,N_6668,N_5139);
nand U9371 (N_9371,N_6164,N_6833);
or U9372 (N_9372,N_5840,N_6030);
nand U9373 (N_9373,N_6226,N_4138);
nor U9374 (N_9374,N_6571,N_7793);
nand U9375 (N_9375,N_5729,N_4865);
and U9376 (N_9376,N_5443,N_4830);
and U9377 (N_9377,N_4116,N_6348);
xnor U9378 (N_9378,N_4026,N_4705);
nor U9379 (N_9379,N_4931,N_7789);
nor U9380 (N_9380,N_7938,N_4291);
nand U9381 (N_9381,N_6223,N_6973);
nor U9382 (N_9382,N_6689,N_5057);
and U9383 (N_9383,N_5079,N_5260);
and U9384 (N_9384,N_6596,N_7484);
xor U9385 (N_9385,N_5345,N_5372);
nand U9386 (N_9386,N_7400,N_6601);
or U9387 (N_9387,N_4170,N_5952);
nor U9388 (N_9388,N_4063,N_7145);
nand U9389 (N_9389,N_7105,N_7529);
or U9390 (N_9390,N_6296,N_5378);
and U9391 (N_9391,N_4893,N_6804);
nor U9392 (N_9392,N_7631,N_6417);
xnor U9393 (N_9393,N_6975,N_7233);
xor U9394 (N_9394,N_4412,N_5870);
or U9395 (N_9395,N_7210,N_6147);
and U9396 (N_9396,N_4987,N_5255);
and U9397 (N_9397,N_5753,N_4894);
nand U9398 (N_9398,N_4685,N_6907);
and U9399 (N_9399,N_6853,N_6671);
nand U9400 (N_9400,N_7151,N_5770);
and U9401 (N_9401,N_7965,N_4132);
and U9402 (N_9402,N_7972,N_7916);
and U9403 (N_9403,N_5061,N_7869);
nand U9404 (N_9404,N_5194,N_7222);
nor U9405 (N_9405,N_4261,N_4545);
nand U9406 (N_9406,N_7443,N_7773);
and U9407 (N_9407,N_4105,N_6192);
nor U9408 (N_9408,N_4628,N_5263);
nor U9409 (N_9409,N_4379,N_7818);
nor U9410 (N_9410,N_5274,N_6483);
or U9411 (N_9411,N_4643,N_6006);
nand U9412 (N_9412,N_4368,N_7967);
and U9413 (N_9413,N_7223,N_4224);
or U9414 (N_9414,N_4567,N_7704);
or U9415 (N_9415,N_4403,N_7767);
nand U9416 (N_9416,N_5097,N_4852);
or U9417 (N_9417,N_6611,N_5108);
xor U9418 (N_9418,N_6057,N_4253);
nand U9419 (N_9419,N_6101,N_4496);
or U9420 (N_9420,N_6244,N_6096);
nand U9421 (N_9421,N_6216,N_5844);
and U9422 (N_9422,N_5184,N_6467);
xnor U9423 (N_9423,N_5021,N_5489);
or U9424 (N_9424,N_7666,N_7984);
nand U9425 (N_9425,N_4502,N_6968);
nand U9426 (N_9426,N_6518,N_4621);
nand U9427 (N_9427,N_7779,N_4817);
and U9428 (N_9428,N_5937,N_5921);
and U9429 (N_9429,N_4258,N_5200);
nor U9430 (N_9430,N_6798,N_4731);
xor U9431 (N_9431,N_5203,N_6260);
nand U9432 (N_9432,N_7566,N_5452);
nand U9433 (N_9433,N_4523,N_6392);
nor U9434 (N_9434,N_7653,N_7433);
nand U9435 (N_9435,N_6059,N_6955);
and U9436 (N_9436,N_7778,N_4975);
or U9437 (N_9437,N_6990,N_5064);
nand U9438 (N_9438,N_6942,N_5918);
or U9439 (N_9439,N_6258,N_5735);
and U9440 (N_9440,N_4274,N_5706);
nor U9441 (N_9441,N_6302,N_5820);
and U9442 (N_9442,N_5976,N_6489);
xor U9443 (N_9443,N_7825,N_7980);
nor U9444 (N_9444,N_5395,N_4506);
or U9445 (N_9445,N_5720,N_7592);
and U9446 (N_9446,N_6384,N_6587);
nand U9447 (N_9447,N_6763,N_4971);
nor U9448 (N_9448,N_7680,N_5382);
nor U9449 (N_9449,N_4580,N_6908);
or U9450 (N_9450,N_6909,N_5852);
or U9451 (N_9451,N_7551,N_5266);
or U9452 (N_9452,N_5339,N_7184);
nor U9453 (N_9453,N_7555,N_4048);
nand U9454 (N_9454,N_5836,N_4699);
xor U9455 (N_9455,N_7811,N_6649);
xnor U9456 (N_9456,N_6228,N_7268);
nand U9457 (N_9457,N_4950,N_6994);
and U9458 (N_9458,N_4921,N_6033);
nor U9459 (N_9459,N_7011,N_6065);
nor U9460 (N_9460,N_7628,N_6657);
or U9461 (N_9461,N_6883,N_6800);
or U9462 (N_9462,N_4877,N_5904);
nor U9463 (N_9463,N_7298,N_4287);
or U9464 (N_9464,N_7807,N_5623);
nor U9465 (N_9465,N_6018,N_5193);
xor U9466 (N_9466,N_7483,N_4604);
and U9467 (N_9467,N_4299,N_7518);
nand U9468 (N_9468,N_4201,N_4793);
xor U9469 (N_9469,N_5123,N_6597);
and U9470 (N_9470,N_4546,N_5227);
nand U9471 (N_9471,N_6893,N_6242);
nor U9472 (N_9472,N_6531,N_5052);
or U9473 (N_9473,N_4286,N_6408);
and U9474 (N_9474,N_4356,N_6850);
nor U9475 (N_9475,N_7574,N_5653);
nand U9476 (N_9476,N_6009,N_5833);
nor U9477 (N_9477,N_5094,N_5214);
nand U9478 (N_9478,N_4004,N_7885);
nor U9479 (N_9479,N_4312,N_4632);
nor U9480 (N_9480,N_4722,N_4700);
or U9481 (N_9481,N_5328,N_4855);
and U9482 (N_9482,N_6577,N_6075);
nand U9483 (N_9483,N_7392,N_5896);
nand U9484 (N_9484,N_6484,N_6672);
and U9485 (N_9485,N_5970,N_6551);
nor U9486 (N_9486,N_6251,N_6516);
nand U9487 (N_9487,N_7966,N_7016);
and U9488 (N_9488,N_5023,N_6339);
and U9489 (N_9489,N_4603,N_4100);
or U9490 (N_9490,N_7878,N_4359);
xor U9491 (N_9491,N_5749,N_6305);
or U9492 (N_9492,N_4750,N_5645);
xor U9493 (N_9493,N_5220,N_4515);
nor U9494 (N_9494,N_6145,N_4764);
nor U9495 (N_9495,N_4391,N_5444);
nor U9496 (N_9496,N_4223,N_5313);
or U9497 (N_9497,N_5731,N_6241);
xor U9498 (N_9498,N_4710,N_5695);
and U9499 (N_9499,N_7510,N_4474);
and U9500 (N_9500,N_6468,N_4754);
nor U9501 (N_9501,N_4453,N_6966);
xor U9502 (N_9502,N_6985,N_5526);
or U9503 (N_9503,N_5926,N_4051);
nor U9504 (N_9504,N_6428,N_4326);
nand U9505 (N_9505,N_5711,N_5371);
nand U9506 (N_9506,N_5955,N_6160);
nor U9507 (N_9507,N_6936,N_5794);
xor U9508 (N_9508,N_5058,N_4595);
or U9509 (N_9509,N_6318,N_5984);
xnor U9510 (N_9510,N_5394,N_4242);
and U9511 (N_9511,N_7445,N_5630);
nor U9512 (N_9512,N_4423,N_6658);
xnor U9513 (N_9513,N_7976,N_7937);
nor U9514 (N_9514,N_5612,N_7193);
xor U9515 (N_9515,N_7695,N_5719);
nand U9516 (N_9516,N_4221,N_4963);
nor U9517 (N_9517,N_6375,N_4124);
nor U9518 (N_9518,N_5958,N_6879);
and U9519 (N_9519,N_4616,N_5429);
xnor U9520 (N_9520,N_6259,N_6901);
nand U9521 (N_9521,N_6554,N_6052);
nand U9522 (N_9522,N_4409,N_5127);
nor U9523 (N_9523,N_6977,N_5179);
or U9524 (N_9524,N_7164,N_7014);
and U9525 (N_9525,N_7761,N_7515);
or U9526 (N_9526,N_6911,N_7307);
and U9527 (N_9527,N_7069,N_5887);
xnor U9528 (N_9528,N_5029,N_6083);
nand U9529 (N_9529,N_7091,N_7700);
nor U9530 (N_9530,N_6697,N_6455);
or U9531 (N_9531,N_5360,N_4889);
and U9532 (N_9532,N_4278,N_4413);
and U9533 (N_9533,N_6361,N_5822);
or U9534 (N_9534,N_5801,N_6224);
or U9535 (N_9535,N_5966,N_4666);
nor U9536 (N_9536,N_7602,N_5551);
xor U9537 (N_9537,N_6685,N_6735);
and U9538 (N_9538,N_7186,N_5710);
nand U9539 (N_9539,N_6578,N_5336);
xnor U9540 (N_9540,N_7545,N_5620);
nor U9541 (N_9541,N_6958,N_7232);
nor U9542 (N_9542,N_5153,N_6142);
or U9543 (N_9543,N_4862,N_5523);
nor U9544 (N_9544,N_5648,N_5086);
xor U9545 (N_9545,N_6740,N_5253);
nor U9546 (N_9546,N_7519,N_5795);
or U9547 (N_9547,N_6070,N_5825);
nor U9548 (N_9548,N_6132,N_4007);
and U9549 (N_9549,N_4755,N_5417);
nand U9550 (N_9550,N_6680,N_5299);
and U9551 (N_9551,N_6487,N_5527);
or U9552 (N_9552,N_5971,N_4381);
or U9553 (N_9553,N_5610,N_4675);
and U9554 (N_9554,N_6711,N_6454);
nor U9555 (N_9555,N_7274,N_4404);
nand U9556 (N_9556,N_5133,N_4336);
and U9557 (N_9557,N_5261,N_7749);
nand U9558 (N_9558,N_4848,N_5828);
and U9559 (N_9559,N_7418,N_6444);
nand U9560 (N_9560,N_4694,N_4879);
nor U9561 (N_9561,N_4049,N_6581);
and U9562 (N_9562,N_7048,N_4561);
xor U9563 (N_9563,N_4968,N_4266);
or U9564 (N_9564,N_7457,N_5001);
nor U9565 (N_9565,N_7745,N_5946);
nor U9566 (N_9566,N_5218,N_5671);
or U9567 (N_9567,N_6169,N_4884);
or U9568 (N_9568,N_5106,N_4257);
xor U9569 (N_9569,N_4072,N_7136);
nand U9570 (N_9570,N_4617,N_7073);
or U9571 (N_9571,N_5761,N_4402);
nand U9572 (N_9572,N_4952,N_5447);
nand U9573 (N_9573,N_6961,N_4625);
nand U9574 (N_9574,N_5905,N_5823);
or U9575 (N_9575,N_4634,N_6795);
and U9576 (N_9576,N_7863,N_4317);
and U9577 (N_9577,N_7553,N_4505);
xor U9578 (N_9578,N_4885,N_5207);
or U9579 (N_9579,N_7075,N_5287);
nor U9580 (N_9580,N_4639,N_6629);
nand U9581 (N_9581,N_6399,N_6335);
nor U9582 (N_9582,N_7046,N_7816);
nand U9583 (N_9583,N_7344,N_5542);
nand U9584 (N_9584,N_6652,N_4559);
nor U9585 (N_9585,N_5377,N_4025);
nand U9586 (N_9586,N_5682,N_7914);
or U9587 (N_9587,N_6555,N_7301);
nor U9588 (N_9588,N_7597,N_4517);
nand U9589 (N_9589,N_4638,N_7913);
nand U9590 (N_9590,N_7876,N_4535);
and U9591 (N_9591,N_7558,N_7458);
nor U9592 (N_9592,N_4541,N_5676);
or U9593 (N_9593,N_4296,N_4780);
nor U9594 (N_9594,N_7795,N_7846);
nor U9595 (N_9595,N_7129,N_4046);
nor U9596 (N_9596,N_7423,N_5348);
xnor U9597 (N_9597,N_6207,N_6179);
nor U9598 (N_9598,N_6213,N_5059);
or U9599 (N_9599,N_4234,N_4646);
or U9600 (N_9600,N_4918,N_5646);
nor U9601 (N_9601,N_4758,N_7432);
nand U9602 (N_9602,N_5164,N_7868);
and U9603 (N_9603,N_4714,N_4676);
and U9604 (N_9604,N_7850,N_4086);
or U9605 (N_9605,N_4294,N_7670);
or U9606 (N_9606,N_7464,N_7598);
or U9607 (N_9607,N_4014,N_6137);
xor U9608 (N_9608,N_6918,N_7705);
xnor U9609 (N_9609,N_5758,N_7275);
nor U9610 (N_9610,N_7933,N_4673);
nor U9611 (N_9611,N_4751,N_7329);
nand U9612 (N_9612,N_6650,N_5026);
nor U9613 (N_9613,N_5615,N_5388);
nand U9614 (N_9614,N_6843,N_5451);
nor U9615 (N_9615,N_5575,N_4476);
nand U9616 (N_9616,N_4401,N_5406);
or U9617 (N_9617,N_5533,N_4927);
nor U9618 (N_9618,N_6949,N_7570);
nor U9619 (N_9619,N_4943,N_7338);
or U9620 (N_9620,N_7999,N_7376);
nor U9621 (N_9621,N_4318,N_4374);
nor U9622 (N_9622,N_7154,N_4823);
nor U9623 (N_9623,N_4983,N_7133);
and U9624 (N_9624,N_5354,N_5781);
nor U9625 (N_9625,N_4601,N_5323);
or U9626 (N_9626,N_6767,N_5252);
nand U9627 (N_9627,N_4363,N_6683);
or U9628 (N_9628,N_5587,N_5881);
nor U9629 (N_9629,N_5196,N_6412);
or U9630 (N_9630,N_4254,N_5347);
xor U9631 (N_9631,N_5691,N_7780);
nor U9632 (N_9632,N_6664,N_5764);
nor U9633 (N_9633,N_7723,N_7312);
nor U9634 (N_9634,N_6394,N_4166);
nor U9635 (N_9635,N_5393,N_4992);
nor U9636 (N_9636,N_6077,N_7309);
or U9637 (N_9637,N_6352,N_7523);
nand U9638 (N_9638,N_5902,N_7476);
nor U9639 (N_9639,N_7535,N_6386);
nor U9640 (N_9640,N_5418,N_4118);
or U9641 (N_9641,N_5146,N_5964);
xor U9642 (N_9642,N_5189,N_7447);
nor U9643 (N_9643,N_6453,N_7845);
or U9644 (N_9644,N_6766,N_4850);
and U9645 (N_9645,N_6190,N_5513);
or U9646 (N_9646,N_7762,N_7006);
xnor U9647 (N_9647,N_7348,N_7622);
or U9648 (N_9648,N_7979,N_6289);
xor U9649 (N_9649,N_5967,N_6722);
nand U9650 (N_9650,N_7295,N_6376);
nor U9651 (N_9651,N_5091,N_6461);
or U9652 (N_9652,N_6993,N_6536);
nand U9653 (N_9653,N_5564,N_7861);
and U9654 (N_9654,N_4098,N_5621);
nor U9655 (N_9655,N_6279,N_7010);
or U9656 (N_9656,N_4820,N_7071);
nor U9657 (N_9657,N_7947,N_4382);
xor U9658 (N_9658,N_5315,N_5968);
and U9659 (N_9659,N_6972,N_6003);
xor U9660 (N_9660,N_4873,N_5440);
and U9661 (N_9661,N_7508,N_5069);
nand U9662 (N_9662,N_5384,N_6572);
and U9663 (N_9663,N_7936,N_5296);
nor U9664 (N_9664,N_6570,N_4407);
nand U9665 (N_9665,N_4323,N_6269);
nor U9666 (N_9666,N_4512,N_7450);
xor U9667 (N_9667,N_7026,N_5453);
and U9668 (N_9668,N_6760,N_6742);
nor U9669 (N_9669,N_4871,N_7935);
or U9670 (N_9670,N_4941,N_7342);
or U9671 (N_9671,N_5374,N_6776);
or U9672 (N_9672,N_4411,N_6442);
nor U9673 (N_9673,N_4315,N_5346);
nand U9674 (N_9674,N_7333,N_7278);
nand U9675 (N_9675,N_7022,N_4344);
nand U9676 (N_9676,N_5589,N_6751);
nand U9677 (N_9677,N_5144,N_5920);
xor U9678 (N_9678,N_4816,N_6219);
and U9679 (N_9679,N_7713,N_4878);
xor U9680 (N_9680,N_5142,N_6971);
or U9681 (N_9681,N_5665,N_7336);
nor U9682 (N_9682,N_6959,N_7586);
and U9683 (N_9683,N_4108,N_6773);
and U9684 (N_9684,N_5167,N_6087);
xnor U9685 (N_9685,N_5493,N_5997);
and U9686 (N_9686,N_6188,N_5569);
or U9687 (N_9687,N_4157,N_6140);
or U9688 (N_9688,N_6886,N_4352);
xor U9689 (N_9689,N_4824,N_4466);
and U9690 (N_9690,N_7697,N_6061);
or U9691 (N_9691,N_5168,N_7684);
nand U9692 (N_9692,N_4001,N_7651);
xor U9693 (N_9693,N_6321,N_7560);
nor U9694 (N_9694,N_7577,N_5047);
or U9695 (N_9695,N_5492,N_7872);
or U9696 (N_9696,N_4439,N_6745);
nand U9697 (N_9697,N_5693,N_4093);
and U9698 (N_9698,N_7998,N_7492);
nor U9699 (N_9699,N_5796,N_4704);
nand U9700 (N_9700,N_5951,N_4145);
and U9701 (N_9701,N_6727,N_6035);
or U9702 (N_9702,N_4612,N_5522);
or U9703 (N_9703,N_7315,N_5681);
nand U9704 (N_9704,N_7038,N_4687);
or U9705 (N_9705,N_6630,N_4231);
xnor U9706 (N_9706,N_4056,N_6104);
or U9707 (N_9707,N_6720,N_6956);
nor U9708 (N_9708,N_4684,N_4622);
and U9709 (N_9709,N_4898,N_7162);
xor U9710 (N_9710,N_6770,N_7724);
or U9711 (N_9711,N_6989,N_6877);
and U9712 (N_9712,N_4464,N_4075);
xor U9713 (N_9713,N_4475,N_4008);
or U9714 (N_9714,N_7102,N_4260);
and U9715 (N_9715,N_6154,N_4834);
or U9716 (N_9716,N_5359,N_5775);
and U9717 (N_9717,N_4554,N_4777);
or U9718 (N_9718,N_6706,N_6622);
and U9719 (N_9719,N_6603,N_5450);
nand U9720 (N_9720,N_4891,N_5957);
nand U9721 (N_9721,N_5748,N_6855);
or U9722 (N_9722,N_7946,N_7929);
xor U9723 (N_9723,N_5217,N_5175);
nor U9724 (N_9724,N_4018,N_5631);
or U9725 (N_9725,N_4255,N_7473);
nor U9726 (N_9726,N_4881,N_4029);
nand U9727 (N_9727,N_6750,N_6830);
and U9728 (N_9728,N_5041,N_4959);
nand U9729 (N_9729,N_5333,N_4614);
nor U9730 (N_9730,N_7557,N_6225);
nor U9731 (N_9731,N_4171,N_7087);
nand U9732 (N_9732,N_7851,N_6651);
nor U9733 (N_9733,N_7717,N_5166);
and U9734 (N_9734,N_4465,N_4156);
and U9735 (N_9735,N_5837,N_6707);
and U9736 (N_9736,N_4189,N_4573);
nor U9737 (N_9737,N_5364,N_5480);
xor U9738 (N_9738,N_7659,N_7324);
nand U9739 (N_9739,N_7130,N_4000);
or U9740 (N_9740,N_6114,N_4997);
and U9741 (N_9741,N_7781,N_4424);
xor U9742 (N_9742,N_6733,N_6319);
or U9743 (N_9743,N_7503,N_6644);
and U9744 (N_9744,N_7879,N_7328);
and U9745 (N_9745,N_4293,N_6960);
nand U9746 (N_9746,N_4191,N_5943);
xnor U9747 (N_9747,N_5979,N_7290);
nand U9748 (N_9748,N_5112,N_5707);
nand U9749 (N_9749,N_4905,N_5511);
or U9750 (N_9750,N_4785,N_4966);
and U9751 (N_9751,N_4325,N_5603);
or U9752 (N_9752,N_7350,N_5911);
nand U9753 (N_9753,N_4479,N_7127);
xor U9754 (N_9754,N_5722,N_4970);
xor U9755 (N_9755,N_4044,N_4337);
nor U9756 (N_9756,N_4679,N_7952);
xor U9757 (N_9757,N_4360,N_7647);
nor U9758 (N_9758,N_6395,N_4948);
and U9759 (N_9759,N_5213,N_5415);
nor U9760 (N_9760,N_5875,N_7059);
xnor U9761 (N_9761,N_4583,N_7742);
xnor U9762 (N_9762,N_6560,N_4152);
nor U9763 (N_9763,N_6826,N_4847);
or U9764 (N_9764,N_4271,N_5352);
and U9765 (N_9765,N_7692,N_6888);
nand U9766 (N_9766,N_5461,N_5956);
or U9767 (N_9767,N_4659,N_5860);
xnor U9768 (N_9768,N_6247,N_5505);
or U9769 (N_9769,N_5608,N_7439);
and U9770 (N_9770,N_5947,N_4345);
xor U9771 (N_9771,N_7368,N_5640);
or U9772 (N_9772,N_7956,N_6556);
nand U9773 (N_9773,N_4549,N_5335);
xor U9774 (N_9774,N_5708,N_4615);
nor U9775 (N_9775,N_5517,N_5662);
nand U9776 (N_9776,N_6168,N_4610);
and U9777 (N_9777,N_6817,N_7599);
nor U9778 (N_9778,N_4033,N_4461);
and U9779 (N_9779,N_6235,N_6964);
and U9780 (N_9780,N_6771,N_6480);
nor U9781 (N_9781,N_5907,N_4256);
nand U9782 (N_9782,N_6211,N_5574);
nand U9783 (N_9783,N_6149,N_7532);
or U9784 (N_9784,N_7112,N_4192);
and U9785 (N_9785,N_7109,N_7912);
nor U9786 (N_9786,N_7681,N_6458);
nor U9787 (N_9787,N_7115,N_6579);
or U9788 (N_9788,N_7771,N_6752);
nor U9789 (N_9789,N_7722,N_4273);
nor U9790 (N_9790,N_5883,N_5783);
nor U9791 (N_9791,N_7748,N_5793);
or U9792 (N_9792,N_5185,N_4013);
and U9793 (N_9793,N_4032,N_5747);
nor U9794 (N_9794,N_6285,N_5307);
nand U9795 (N_9795,N_7580,N_4540);
nand U9796 (N_9796,N_5225,N_6056);
nor U9797 (N_9797,N_5734,N_4562);
or U9798 (N_9798,N_5633,N_7922);
or U9799 (N_9799,N_5482,N_6180);
nor U9800 (N_9800,N_4062,N_7319);
and U9801 (N_9801,N_7880,N_7025);
xor U9802 (N_9802,N_7002,N_7067);
or U9803 (N_9803,N_7766,N_7294);
or U9804 (N_9804,N_7472,N_7534);
nor U9805 (N_9805,N_5423,N_7384);
nand U9806 (N_9806,N_5455,N_4217);
nor U9807 (N_9807,N_6017,N_6477);
nand U9808 (N_9808,N_6631,N_6802);
nor U9809 (N_9809,N_4420,N_6582);
or U9810 (N_9810,N_6648,N_5494);
nor U9811 (N_9811,N_5401,N_7394);
xnor U9812 (N_9812,N_6690,N_4729);
or U9813 (N_9813,N_5639,N_5733);
nor U9814 (N_9814,N_6478,N_5923);
or U9815 (N_9815,N_6439,N_4045);
and U9816 (N_9816,N_6058,N_4692);
and U9817 (N_9817,N_5050,N_4305);
nand U9818 (N_9818,N_7012,N_6465);
or U9819 (N_9819,N_4693,N_6796);
nor U9820 (N_9820,N_4799,N_5420);
xnor U9821 (N_9821,N_4238,N_7668);
nand U9822 (N_9822,N_7095,N_6937);
nand U9823 (N_9823,N_4767,N_4384);
nand U9824 (N_9824,N_4608,N_6590);
nand U9825 (N_9825,N_5190,N_7625);
or U9826 (N_9826,N_7276,N_7385);
or U9827 (N_9827,N_5963,N_7030);
or U9828 (N_9828,N_6040,N_5366);
nand U9829 (N_9829,N_4828,N_4645);
nor U9830 (N_9830,N_5244,N_5985);
nand U9831 (N_9831,N_4774,N_5234);
or U9832 (N_9832,N_5624,N_5191);
nand U9833 (N_9833,N_6128,N_4791);
nor U9834 (N_9834,N_4570,N_4939);
nand U9835 (N_9835,N_5262,N_4801);
nor U9836 (N_9836,N_7305,N_5187);
nor U9837 (N_9837,N_5830,N_7940);
or U9838 (N_9838,N_5991,N_4151);
nand U9839 (N_9839,N_5013,N_6822);
nor U9840 (N_9840,N_5463,N_4715);
or U9841 (N_9841,N_7903,N_7160);
and U9842 (N_9842,N_7752,N_4263);
and U9843 (N_9843,N_7252,N_4732);
nor U9844 (N_9844,N_5039,N_6791);
nand U9845 (N_9845,N_7099,N_5824);
nor U9846 (N_9846,N_5040,N_6670);
nand U9847 (N_9847,N_6144,N_7171);
nor U9848 (N_9848,N_4123,N_5572);
or U9849 (N_9849,N_7330,N_6304);
nor U9850 (N_9850,N_5208,N_7865);
nor U9851 (N_9851,N_7604,N_4459);
nand U9852 (N_9852,N_7669,N_4125);
nand U9853 (N_9853,N_6210,N_5571);
nand U9854 (N_9854,N_7216,N_4988);
nand U9855 (N_9855,N_4289,N_6115);
nand U9856 (N_9856,N_6512,N_4867);
nor U9857 (N_9857,N_7540,N_4837);
xnor U9858 (N_9858,N_7754,N_6728);
or U9859 (N_9859,N_6508,N_6782);
xor U9860 (N_9860,N_6443,N_7527);
and U9861 (N_9861,N_7083,N_4845);
and U9862 (N_9862,N_4022,N_5774);
and U9863 (N_9863,N_6797,N_7835);
and U9864 (N_9864,N_5536,N_5690);
and U9865 (N_9865,N_4102,N_4606);
and U9866 (N_9866,N_7396,N_5277);
and U9867 (N_9867,N_4057,N_5014);
and U9868 (N_9868,N_4980,N_6910);
and U9869 (N_9869,N_4099,N_6957);
nor U9870 (N_9870,N_5247,N_5701);
or U9871 (N_9871,N_5949,N_5132);
nand U9872 (N_9872,N_4129,N_4276);
nor U9873 (N_9873,N_6825,N_5435);
or U9874 (N_9874,N_5473,N_7488);
and U9875 (N_9875,N_6525,N_5022);
or U9876 (N_9876,N_5107,N_7627);
nand U9877 (N_9877,N_5950,N_6004);
nor U9878 (N_9878,N_6793,N_4168);
nor U9879 (N_9879,N_5090,N_4097);
or U9880 (N_9880,N_7219,N_4386);
or U9881 (N_9881,N_4122,N_7139);
nand U9882 (N_9882,N_7890,N_4525);
xor U9883 (N_9883,N_4798,N_5383);
nor U9884 (N_9884,N_6002,N_5892);
or U9885 (N_9885,N_7977,N_6060);
xor U9886 (N_9886,N_6547,N_6857);
or U9887 (N_9887,N_7725,N_4444);
nand U9888 (N_9888,N_7495,N_6306);
and U9889 (N_9889,N_7463,N_4071);
nand U9890 (N_9890,N_6071,N_5349);
nand U9891 (N_9891,N_7339,N_5129);
or U9892 (N_9892,N_5276,N_7185);
and U9893 (N_9893,N_5561,N_7271);
nor U9894 (N_9894,N_4566,N_7537);
and U9895 (N_9895,N_6686,N_5927);
xnor U9896 (N_9896,N_7871,N_7456);
nor U9897 (N_9897,N_6255,N_7701);
or U9898 (N_9898,N_5919,N_6317);
or U9899 (N_9899,N_6616,N_7437);
nand U9900 (N_9900,N_6243,N_7549);
and U9901 (N_9901,N_6435,N_6418);
and U9902 (N_9902,N_6932,N_4655);
and U9903 (N_9903,N_6299,N_7044);
and U9904 (N_9904,N_7064,N_4575);
nand U9905 (N_9905,N_7413,N_7066);
or U9906 (N_9906,N_6214,N_5675);
nor U9907 (N_9907,N_7905,N_7787);
nor U9908 (N_9908,N_7776,N_6419);
nand U9909 (N_9909,N_6425,N_7403);
nor U9910 (N_9910,N_4448,N_5176);
or U9911 (N_9911,N_7041,N_5784);
or U9912 (N_9912,N_6379,N_7955);
nor U9913 (N_9913,N_7800,N_5570);
or U9914 (N_9914,N_7051,N_7550);
or U9915 (N_9915,N_6237,N_4761);
nand U9916 (N_9916,N_6383,N_6438);
or U9917 (N_9917,N_4786,N_7416);
or U9918 (N_9918,N_5702,N_4933);
nand U9919 (N_9919,N_5369,N_4594);
nor U9920 (N_9920,N_4985,N_6674);
nand U9921 (N_9921,N_6495,N_4073);
or U9922 (N_9922,N_4519,N_4920);
nand U9923 (N_9923,N_7008,N_4511);
nor U9924 (N_9924,N_6963,N_4619);
or U9925 (N_9925,N_7187,N_6050);
and U9926 (N_9926,N_5715,N_5149);
or U9927 (N_9927,N_7820,N_6639);
nand U9928 (N_9928,N_5499,N_4677);
or U9929 (N_9929,N_6858,N_5890);
nor U9930 (N_9930,N_6677,N_5744);
nand U9931 (N_9931,N_5375,N_7591);
xnor U9932 (N_9932,N_7269,N_5560);
xor U9933 (N_9933,N_4199,N_6281);
nand U9934 (N_9934,N_7076,N_7453);
or U9935 (N_9935,N_7883,N_4861);
nor U9936 (N_9936,N_5978,N_5756);
nor U9937 (N_9937,N_7633,N_7774);
xor U9938 (N_9938,N_6744,N_5426);
or U9939 (N_9939,N_6276,N_6353);
nor U9940 (N_9940,N_5241,N_4012);
nor U9941 (N_9941,N_4472,N_4272);
nor U9942 (N_9942,N_7652,N_5268);
and U9943 (N_9943,N_6747,N_4890);
or U9944 (N_9944,N_7165,N_5338);
nor U9945 (N_9945,N_4183,N_6354);
or U9946 (N_9946,N_5877,N_5235);
and U9947 (N_9947,N_5914,N_4733);
xnor U9948 (N_9948,N_6047,N_6847);
and U9949 (N_9949,N_7703,N_7236);
or U9950 (N_9950,N_4789,N_7248);
nand U9951 (N_9951,N_7388,N_4783);
or U9952 (N_9952,N_7364,N_4651);
nor U9953 (N_9953,N_6476,N_7496);
nand U9954 (N_9954,N_5746,N_4207);
nand U9955 (N_9955,N_7150,N_6635);
nor U9956 (N_9956,N_4002,N_4076);
xor U9957 (N_9957,N_4175,N_6801);
and U9958 (N_9958,N_4790,N_6273);
nor U9959 (N_9959,N_4335,N_5666);
or U9960 (N_9960,N_5600,N_7944);
and U9961 (N_9961,N_7335,N_5721);
nand U9962 (N_9962,N_7618,N_6166);
and U9963 (N_9963,N_5449,N_7522);
nor U9964 (N_9964,N_6126,N_7775);
or U9965 (N_9965,N_4542,N_6840);
xnor U9966 (N_9966,N_5884,N_7378);
or U9967 (N_9967,N_7397,N_5808);
nor U9968 (N_9968,N_7104,N_6268);
and U9969 (N_9969,N_7096,N_4771);
nor U9970 (N_9970,N_5789,N_7931);
nand U9971 (N_9971,N_4727,N_7251);
nor U9972 (N_9972,N_7660,N_5868);
nor U9973 (N_9973,N_5291,N_5006);
nor U9974 (N_9974,N_5411,N_5859);
and U9975 (N_9975,N_7363,N_6100);
nand U9976 (N_9976,N_4043,N_7716);
or U9977 (N_9977,N_5604,N_6218);
nand U9978 (N_9978,N_7506,N_7830);
nand U9979 (N_9979,N_4431,N_7334);
and U9980 (N_9980,N_6091,N_6286);
and U9981 (N_9981,N_6485,N_7747);
and U9982 (N_9982,N_7585,N_6923);
nand U9983 (N_9983,N_7387,N_7260);
and U9984 (N_9984,N_7358,N_4462);
nor U9985 (N_9985,N_4371,N_7177);
xnor U9986 (N_9986,N_5390,N_5941);
nand U9987 (N_9987,N_7554,N_7791);
and U9988 (N_9988,N_7024,N_7962);
and U9989 (N_9989,N_4713,N_4084);
and U9990 (N_9990,N_4415,N_7039);
xnor U9991 (N_9991,N_4184,N_4236);
nand U9992 (N_9992,N_4456,N_7228);
or U9993 (N_9993,N_7494,N_5286);
and U9994 (N_9994,N_5732,N_6864);
or U9995 (N_9995,N_4773,N_7085);
nor U9996 (N_9996,N_4176,N_7858);
or U9997 (N_9997,N_4919,N_7833);
nor U9998 (N_9998,N_6619,N_4769);
nand U9999 (N_9999,N_4017,N_5442);
and U10000 (N_10000,N_5113,N_7486);
or U10001 (N_10001,N_6691,N_4283);
or U10002 (N_10002,N_7112,N_5451);
and U10003 (N_10003,N_4256,N_4154);
or U10004 (N_10004,N_5598,N_5649);
nand U10005 (N_10005,N_6714,N_5637);
and U10006 (N_10006,N_7178,N_6379);
or U10007 (N_10007,N_4452,N_5794);
xor U10008 (N_10008,N_7599,N_5050);
or U10009 (N_10009,N_4334,N_5778);
or U10010 (N_10010,N_4531,N_6234);
or U10011 (N_10011,N_4937,N_7718);
xor U10012 (N_10012,N_4950,N_4758);
nand U10013 (N_10013,N_6398,N_6857);
and U10014 (N_10014,N_7924,N_4570);
nand U10015 (N_10015,N_4904,N_5313);
and U10016 (N_10016,N_5621,N_6370);
and U10017 (N_10017,N_5901,N_7410);
nand U10018 (N_10018,N_6859,N_4706);
or U10019 (N_10019,N_4979,N_5047);
nor U10020 (N_10020,N_4926,N_5419);
or U10021 (N_10021,N_6099,N_6787);
and U10022 (N_10022,N_5184,N_5121);
xnor U10023 (N_10023,N_6980,N_5568);
nand U10024 (N_10024,N_7458,N_6649);
or U10025 (N_10025,N_4528,N_7316);
nor U10026 (N_10026,N_5030,N_6539);
nand U10027 (N_10027,N_7314,N_4466);
nor U10028 (N_10028,N_4849,N_5617);
xor U10029 (N_10029,N_6546,N_6472);
or U10030 (N_10030,N_5759,N_5181);
and U10031 (N_10031,N_7666,N_7181);
xor U10032 (N_10032,N_7283,N_6423);
and U10033 (N_10033,N_6158,N_4264);
and U10034 (N_10034,N_7103,N_7713);
and U10035 (N_10035,N_4031,N_6499);
or U10036 (N_10036,N_7530,N_6035);
or U10037 (N_10037,N_4831,N_4272);
nor U10038 (N_10038,N_5672,N_7534);
nand U10039 (N_10039,N_5035,N_7694);
nor U10040 (N_10040,N_7641,N_6161);
nor U10041 (N_10041,N_5300,N_5243);
or U10042 (N_10042,N_7149,N_6787);
or U10043 (N_10043,N_7290,N_7345);
or U10044 (N_10044,N_7986,N_4679);
nor U10045 (N_10045,N_6454,N_6510);
nand U10046 (N_10046,N_6480,N_6531);
nor U10047 (N_10047,N_5058,N_4897);
or U10048 (N_10048,N_6163,N_6231);
nor U10049 (N_10049,N_4754,N_4688);
and U10050 (N_10050,N_7140,N_4699);
nor U10051 (N_10051,N_5225,N_6691);
nor U10052 (N_10052,N_7243,N_5761);
xor U10053 (N_10053,N_5311,N_7586);
and U10054 (N_10054,N_6099,N_5564);
or U10055 (N_10055,N_7176,N_7071);
or U10056 (N_10056,N_4915,N_5111);
and U10057 (N_10057,N_6610,N_6488);
nand U10058 (N_10058,N_5482,N_7333);
and U10059 (N_10059,N_4188,N_5302);
nand U10060 (N_10060,N_4954,N_5014);
and U10061 (N_10061,N_5411,N_5508);
and U10062 (N_10062,N_5231,N_4124);
or U10063 (N_10063,N_5147,N_7097);
and U10064 (N_10064,N_5634,N_4846);
or U10065 (N_10065,N_4032,N_6253);
or U10066 (N_10066,N_4715,N_4137);
xor U10067 (N_10067,N_5470,N_7937);
nor U10068 (N_10068,N_6684,N_6393);
or U10069 (N_10069,N_4903,N_4905);
and U10070 (N_10070,N_6825,N_6424);
and U10071 (N_10071,N_6344,N_5353);
nor U10072 (N_10072,N_7410,N_6180);
or U10073 (N_10073,N_4993,N_6959);
nand U10074 (N_10074,N_4272,N_6551);
or U10075 (N_10075,N_6846,N_6016);
nand U10076 (N_10076,N_6609,N_7080);
nand U10077 (N_10077,N_4793,N_5108);
nor U10078 (N_10078,N_7437,N_5665);
or U10079 (N_10079,N_4399,N_4790);
and U10080 (N_10080,N_5532,N_4919);
nand U10081 (N_10081,N_4304,N_4576);
and U10082 (N_10082,N_5717,N_7094);
or U10083 (N_10083,N_4872,N_6379);
nand U10084 (N_10084,N_5127,N_5250);
nor U10085 (N_10085,N_4225,N_4651);
and U10086 (N_10086,N_7391,N_4721);
xnor U10087 (N_10087,N_4311,N_5308);
or U10088 (N_10088,N_7415,N_7206);
nor U10089 (N_10089,N_6212,N_4521);
and U10090 (N_10090,N_4750,N_4414);
and U10091 (N_10091,N_7248,N_4578);
and U10092 (N_10092,N_4712,N_5909);
and U10093 (N_10093,N_7980,N_6147);
or U10094 (N_10094,N_7187,N_5643);
xor U10095 (N_10095,N_7168,N_5748);
nand U10096 (N_10096,N_4465,N_5537);
and U10097 (N_10097,N_4837,N_4663);
and U10098 (N_10098,N_7900,N_5170);
or U10099 (N_10099,N_5784,N_7692);
and U10100 (N_10100,N_5268,N_4959);
nand U10101 (N_10101,N_7058,N_5519);
nand U10102 (N_10102,N_5436,N_4939);
nand U10103 (N_10103,N_7451,N_4444);
or U10104 (N_10104,N_6150,N_4317);
and U10105 (N_10105,N_7826,N_6807);
nand U10106 (N_10106,N_6018,N_7092);
and U10107 (N_10107,N_4950,N_4148);
xnor U10108 (N_10108,N_5425,N_4121);
or U10109 (N_10109,N_4665,N_4547);
nor U10110 (N_10110,N_7138,N_4112);
or U10111 (N_10111,N_4015,N_5400);
or U10112 (N_10112,N_6035,N_4183);
or U10113 (N_10113,N_4084,N_6535);
xor U10114 (N_10114,N_4663,N_6943);
or U10115 (N_10115,N_6865,N_4233);
or U10116 (N_10116,N_7096,N_4168);
nor U10117 (N_10117,N_6896,N_7627);
nor U10118 (N_10118,N_5582,N_7465);
and U10119 (N_10119,N_5231,N_7386);
nor U10120 (N_10120,N_5915,N_4881);
nand U10121 (N_10121,N_4972,N_6062);
nor U10122 (N_10122,N_5890,N_6038);
and U10123 (N_10123,N_4491,N_6797);
and U10124 (N_10124,N_7159,N_7024);
or U10125 (N_10125,N_4815,N_4283);
or U10126 (N_10126,N_6573,N_6374);
xnor U10127 (N_10127,N_5717,N_6283);
nand U10128 (N_10128,N_5982,N_7318);
xor U10129 (N_10129,N_4225,N_4393);
nand U10130 (N_10130,N_4913,N_7379);
and U10131 (N_10131,N_4796,N_4252);
and U10132 (N_10132,N_4579,N_6609);
or U10133 (N_10133,N_7190,N_6208);
nand U10134 (N_10134,N_7380,N_5318);
nor U10135 (N_10135,N_5446,N_7729);
nor U10136 (N_10136,N_4081,N_7057);
nand U10137 (N_10137,N_6547,N_6824);
and U10138 (N_10138,N_6463,N_4907);
nand U10139 (N_10139,N_7485,N_7192);
nand U10140 (N_10140,N_7742,N_5171);
nand U10141 (N_10141,N_6823,N_5504);
nor U10142 (N_10142,N_4750,N_4130);
and U10143 (N_10143,N_6852,N_6550);
or U10144 (N_10144,N_6896,N_6747);
or U10145 (N_10145,N_7723,N_7167);
and U10146 (N_10146,N_4499,N_4644);
nand U10147 (N_10147,N_7395,N_7570);
nand U10148 (N_10148,N_7570,N_5940);
or U10149 (N_10149,N_7489,N_7055);
nand U10150 (N_10150,N_5190,N_7965);
and U10151 (N_10151,N_7520,N_5260);
nor U10152 (N_10152,N_5992,N_4094);
nand U10153 (N_10153,N_6788,N_4823);
nand U10154 (N_10154,N_7094,N_5262);
nor U10155 (N_10155,N_4753,N_5253);
nand U10156 (N_10156,N_6348,N_7605);
or U10157 (N_10157,N_4523,N_4656);
nor U10158 (N_10158,N_4023,N_6706);
or U10159 (N_10159,N_4519,N_6669);
nor U10160 (N_10160,N_7414,N_5664);
nand U10161 (N_10161,N_4854,N_7943);
nor U10162 (N_10162,N_7365,N_4522);
nand U10163 (N_10163,N_7864,N_5337);
nand U10164 (N_10164,N_6236,N_7890);
or U10165 (N_10165,N_7346,N_4555);
or U10166 (N_10166,N_7562,N_4768);
and U10167 (N_10167,N_6773,N_4095);
or U10168 (N_10168,N_4299,N_6975);
and U10169 (N_10169,N_5239,N_4346);
or U10170 (N_10170,N_7632,N_4361);
and U10171 (N_10171,N_6410,N_7293);
or U10172 (N_10172,N_4201,N_5410);
nor U10173 (N_10173,N_6513,N_7088);
nand U10174 (N_10174,N_4941,N_6398);
nor U10175 (N_10175,N_6031,N_6799);
nand U10176 (N_10176,N_5544,N_7667);
nor U10177 (N_10177,N_6099,N_5277);
nand U10178 (N_10178,N_4014,N_7442);
nor U10179 (N_10179,N_5354,N_4315);
and U10180 (N_10180,N_6381,N_4089);
or U10181 (N_10181,N_6184,N_5960);
and U10182 (N_10182,N_6993,N_4198);
nand U10183 (N_10183,N_6166,N_5656);
or U10184 (N_10184,N_5524,N_5218);
or U10185 (N_10185,N_4526,N_7300);
nor U10186 (N_10186,N_6260,N_4022);
nand U10187 (N_10187,N_5044,N_4066);
and U10188 (N_10188,N_4781,N_4600);
nand U10189 (N_10189,N_7024,N_7956);
and U10190 (N_10190,N_4372,N_5555);
nor U10191 (N_10191,N_5240,N_7701);
and U10192 (N_10192,N_4609,N_4554);
nor U10193 (N_10193,N_4469,N_6553);
nand U10194 (N_10194,N_7765,N_4414);
nand U10195 (N_10195,N_7636,N_5348);
and U10196 (N_10196,N_6200,N_7958);
or U10197 (N_10197,N_7565,N_5091);
xor U10198 (N_10198,N_4483,N_6380);
xor U10199 (N_10199,N_4781,N_6468);
or U10200 (N_10200,N_4939,N_6818);
nor U10201 (N_10201,N_4911,N_6557);
and U10202 (N_10202,N_6016,N_5722);
and U10203 (N_10203,N_4323,N_6652);
nor U10204 (N_10204,N_4322,N_5335);
xor U10205 (N_10205,N_5898,N_4714);
nor U10206 (N_10206,N_4630,N_4512);
xnor U10207 (N_10207,N_4501,N_4023);
or U10208 (N_10208,N_5491,N_5503);
or U10209 (N_10209,N_4534,N_6312);
xnor U10210 (N_10210,N_5234,N_6787);
or U10211 (N_10211,N_6544,N_7573);
or U10212 (N_10212,N_7420,N_6035);
or U10213 (N_10213,N_4723,N_5419);
nand U10214 (N_10214,N_7100,N_5553);
and U10215 (N_10215,N_5779,N_5217);
or U10216 (N_10216,N_6891,N_4289);
nor U10217 (N_10217,N_4574,N_4160);
nand U10218 (N_10218,N_7810,N_4525);
nand U10219 (N_10219,N_7540,N_6268);
nand U10220 (N_10220,N_7497,N_4349);
nor U10221 (N_10221,N_7218,N_6452);
or U10222 (N_10222,N_4538,N_7567);
nand U10223 (N_10223,N_4301,N_7252);
nor U10224 (N_10224,N_4534,N_6099);
or U10225 (N_10225,N_4682,N_4766);
nand U10226 (N_10226,N_6031,N_7785);
or U10227 (N_10227,N_6641,N_6483);
or U10228 (N_10228,N_7064,N_7124);
nor U10229 (N_10229,N_6464,N_4602);
nor U10230 (N_10230,N_6901,N_7642);
or U10231 (N_10231,N_5735,N_5489);
xnor U10232 (N_10232,N_4352,N_5415);
and U10233 (N_10233,N_4515,N_5898);
and U10234 (N_10234,N_5418,N_5762);
and U10235 (N_10235,N_6409,N_6973);
or U10236 (N_10236,N_5052,N_5663);
nor U10237 (N_10237,N_4836,N_6224);
and U10238 (N_10238,N_6306,N_5160);
nand U10239 (N_10239,N_6126,N_5864);
or U10240 (N_10240,N_6633,N_6814);
or U10241 (N_10241,N_4328,N_7811);
nor U10242 (N_10242,N_7335,N_5458);
nor U10243 (N_10243,N_7773,N_6822);
and U10244 (N_10244,N_5690,N_6221);
or U10245 (N_10245,N_4899,N_6911);
or U10246 (N_10246,N_7520,N_7046);
or U10247 (N_10247,N_4768,N_5579);
and U10248 (N_10248,N_5123,N_5784);
and U10249 (N_10249,N_4599,N_4698);
nand U10250 (N_10250,N_7910,N_5359);
nand U10251 (N_10251,N_5147,N_7209);
and U10252 (N_10252,N_5698,N_4120);
and U10253 (N_10253,N_7325,N_6489);
and U10254 (N_10254,N_6144,N_4426);
nand U10255 (N_10255,N_5783,N_7387);
or U10256 (N_10256,N_5233,N_4535);
nor U10257 (N_10257,N_6456,N_5466);
xor U10258 (N_10258,N_7719,N_7250);
nor U10259 (N_10259,N_5423,N_6284);
and U10260 (N_10260,N_6693,N_5210);
and U10261 (N_10261,N_7447,N_4767);
or U10262 (N_10262,N_7440,N_4570);
and U10263 (N_10263,N_6683,N_4859);
nand U10264 (N_10264,N_5623,N_6822);
nand U10265 (N_10265,N_4094,N_4305);
nor U10266 (N_10266,N_4505,N_4107);
nor U10267 (N_10267,N_6857,N_4399);
and U10268 (N_10268,N_5094,N_6407);
nand U10269 (N_10269,N_6445,N_6780);
and U10270 (N_10270,N_7096,N_7365);
and U10271 (N_10271,N_4375,N_4646);
and U10272 (N_10272,N_5938,N_7287);
nand U10273 (N_10273,N_4300,N_6509);
nand U10274 (N_10274,N_6748,N_7467);
or U10275 (N_10275,N_6479,N_7241);
and U10276 (N_10276,N_5076,N_7490);
or U10277 (N_10277,N_7291,N_7300);
xor U10278 (N_10278,N_6944,N_7539);
nor U10279 (N_10279,N_6651,N_4445);
xor U10280 (N_10280,N_4766,N_5205);
or U10281 (N_10281,N_4314,N_6513);
and U10282 (N_10282,N_4265,N_5174);
xnor U10283 (N_10283,N_6213,N_4473);
and U10284 (N_10284,N_7528,N_5094);
and U10285 (N_10285,N_6772,N_6383);
and U10286 (N_10286,N_4418,N_6231);
and U10287 (N_10287,N_6410,N_5420);
and U10288 (N_10288,N_4692,N_4936);
nand U10289 (N_10289,N_4672,N_4122);
nand U10290 (N_10290,N_7597,N_5344);
xor U10291 (N_10291,N_7123,N_7411);
nand U10292 (N_10292,N_5405,N_4986);
xnor U10293 (N_10293,N_5865,N_6651);
nand U10294 (N_10294,N_6984,N_5691);
or U10295 (N_10295,N_7483,N_5880);
nor U10296 (N_10296,N_4900,N_4794);
or U10297 (N_10297,N_6961,N_4496);
nor U10298 (N_10298,N_4615,N_5455);
nor U10299 (N_10299,N_6246,N_4973);
nand U10300 (N_10300,N_5328,N_6791);
or U10301 (N_10301,N_7883,N_7707);
xor U10302 (N_10302,N_6261,N_4626);
and U10303 (N_10303,N_4620,N_7377);
and U10304 (N_10304,N_5327,N_4871);
nand U10305 (N_10305,N_4366,N_5320);
nand U10306 (N_10306,N_6584,N_6769);
nand U10307 (N_10307,N_6271,N_5742);
nand U10308 (N_10308,N_4314,N_6595);
nand U10309 (N_10309,N_4655,N_7945);
or U10310 (N_10310,N_6824,N_5894);
and U10311 (N_10311,N_5872,N_6263);
nor U10312 (N_10312,N_4173,N_4259);
nand U10313 (N_10313,N_5658,N_7903);
xnor U10314 (N_10314,N_7401,N_5192);
and U10315 (N_10315,N_6101,N_7971);
or U10316 (N_10316,N_5588,N_5538);
or U10317 (N_10317,N_7598,N_7619);
and U10318 (N_10318,N_6422,N_6010);
or U10319 (N_10319,N_5652,N_4815);
nand U10320 (N_10320,N_4518,N_6748);
or U10321 (N_10321,N_4549,N_4633);
xnor U10322 (N_10322,N_7752,N_6182);
nand U10323 (N_10323,N_4718,N_7715);
or U10324 (N_10324,N_7846,N_5482);
or U10325 (N_10325,N_7493,N_4529);
or U10326 (N_10326,N_6256,N_7182);
nor U10327 (N_10327,N_4067,N_5485);
xor U10328 (N_10328,N_6705,N_4243);
nor U10329 (N_10329,N_7644,N_5513);
xnor U10330 (N_10330,N_7414,N_5280);
nor U10331 (N_10331,N_5069,N_6631);
and U10332 (N_10332,N_6004,N_5841);
nor U10333 (N_10333,N_7337,N_4717);
nor U10334 (N_10334,N_4106,N_4858);
and U10335 (N_10335,N_5894,N_4532);
nand U10336 (N_10336,N_4521,N_6051);
nor U10337 (N_10337,N_5214,N_4010);
or U10338 (N_10338,N_7131,N_7053);
xor U10339 (N_10339,N_7987,N_7893);
nor U10340 (N_10340,N_6087,N_7233);
nor U10341 (N_10341,N_6966,N_5901);
nor U10342 (N_10342,N_5314,N_6910);
and U10343 (N_10343,N_5055,N_4766);
nor U10344 (N_10344,N_7904,N_7308);
and U10345 (N_10345,N_7785,N_6180);
nor U10346 (N_10346,N_4930,N_4605);
and U10347 (N_10347,N_4696,N_4744);
and U10348 (N_10348,N_5550,N_4276);
nor U10349 (N_10349,N_6078,N_6487);
nand U10350 (N_10350,N_6179,N_4033);
and U10351 (N_10351,N_7294,N_7061);
nand U10352 (N_10352,N_4955,N_6722);
and U10353 (N_10353,N_6954,N_4862);
nand U10354 (N_10354,N_4572,N_7451);
nand U10355 (N_10355,N_6714,N_4766);
nand U10356 (N_10356,N_5752,N_4385);
and U10357 (N_10357,N_5585,N_4609);
or U10358 (N_10358,N_5348,N_5854);
and U10359 (N_10359,N_6157,N_6847);
nor U10360 (N_10360,N_4428,N_4784);
and U10361 (N_10361,N_6731,N_5970);
and U10362 (N_10362,N_7415,N_5584);
nor U10363 (N_10363,N_4251,N_6016);
or U10364 (N_10364,N_4267,N_5670);
nand U10365 (N_10365,N_6975,N_7590);
or U10366 (N_10366,N_4936,N_4815);
or U10367 (N_10367,N_7708,N_7463);
or U10368 (N_10368,N_4710,N_5711);
and U10369 (N_10369,N_6477,N_4203);
xnor U10370 (N_10370,N_6576,N_4258);
nand U10371 (N_10371,N_7193,N_6587);
and U10372 (N_10372,N_7759,N_7614);
and U10373 (N_10373,N_7732,N_7283);
nor U10374 (N_10374,N_5933,N_6914);
nand U10375 (N_10375,N_4180,N_6349);
xnor U10376 (N_10376,N_7546,N_4260);
xor U10377 (N_10377,N_7155,N_6051);
nand U10378 (N_10378,N_7215,N_6586);
or U10379 (N_10379,N_7363,N_7083);
nand U10380 (N_10380,N_4037,N_7381);
nand U10381 (N_10381,N_5814,N_6415);
and U10382 (N_10382,N_5247,N_4395);
xnor U10383 (N_10383,N_7197,N_4338);
nand U10384 (N_10384,N_5995,N_4175);
xor U10385 (N_10385,N_6057,N_4680);
or U10386 (N_10386,N_5027,N_4033);
or U10387 (N_10387,N_5124,N_7481);
and U10388 (N_10388,N_4768,N_6110);
and U10389 (N_10389,N_4419,N_4774);
and U10390 (N_10390,N_7109,N_5250);
and U10391 (N_10391,N_4303,N_5363);
nor U10392 (N_10392,N_5071,N_5275);
nand U10393 (N_10393,N_6960,N_5849);
and U10394 (N_10394,N_7104,N_7270);
and U10395 (N_10395,N_4961,N_6921);
nand U10396 (N_10396,N_7353,N_5539);
nand U10397 (N_10397,N_6993,N_4782);
and U10398 (N_10398,N_7215,N_7545);
and U10399 (N_10399,N_7314,N_6541);
or U10400 (N_10400,N_4231,N_4874);
or U10401 (N_10401,N_6187,N_5829);
nor U10402 (N_10402,N_7981,N_4772);
nand U10403 (N_10403,N_4487,N_4270);
and U10404 (N_10404,N_4237,N_6290);
xor U10405 (N_10405,N_4220,N_6656);
nand U10406 (N_10406,N_6195,N_4622);
xnor U10407 (N_10407,N_6559,N_7755);
and U10408 (N_10408,N_6641,N_6987);
and U10409 (N_10409,N_7527,N_5383);
xor U10410 (N_10410,N_7790,N_4665);
nand U10411 (N_10411,N_4204,N_4252);
or U10412 (N_10412,N_6341,N_7608);
xor U10413 (N_10413,N_4705,N_7347);
and U10414 (N_10414,N_4131,N_5887);
or U10415 (N_10415,N_6426,N_6044);
nand U10416 (N_10416,N_7067,N_7327);
nand U10417 (N_10417,N_6326,N_4042);
nand U10418 (N_10418,N_4673,N_6793);
nand U10419 (N_10419,N_5006,N_6925);
nor U10420 (N_10420,N_7939,N_6643);
nand U10421 (N_10421,N_6305,N_6239);
and U10422 (N_10422,N_7397,N_4388);
xor U10423 (N_10423,N_7118,N_4413);
and U10424 (N_10424,N_5204,N_7442);
nor U10425 (N_10425,N_5670,N_5856);
and U10426 (N_10426,N_5240,N_7826);
nand U10427 (N_10427,N_4750,N_4214);
nand U10428 (N_10428,N_6899,N_5717);
and U10429 (N_10429,N_7627,N_7403);
nand U10430 (N_10430,N_5689,N_5730);
or U10431 (N_10431,N_6559,N_4936);
or U10432 (N_10432,N_7529,N_5332);
nor U10433 (N_10433,N_7114,N_7400);
or U10434 (N_10434,N_5428,N_7025);
nand U10435 (N_10435,N_6247,N_4537);
nand U10436 (N_10436,N_4026,N_6381);
and U10437 (N_10437,N_6273,N_5169);
nand U10438 (N_10438,N_4356,N_5703);
or U10439 (N_10439,N_5103,N_4466);
nor U10440 (N_10440,N_6170,N_7483);
nand U10441 (N_10441,N_6762,N_4931);
and U10442 (N_10442,N_7237,N_5565);
xnor U10443 (N_10443,N_4558,N_4154);
nand U10444 (N_10444,N_4356,N_7958);
and U10445 (N_10445,N_7807,N_7624);
nor U10446 (N_10446,N_6668,N_6608);
and U10447 (N_10447,N_7353,N_4475);
and U10448 (N_10448,N_7354,N_7234);
nor U10449 (N_10449,N_5951,N_7030);
and U10450 (N_10450,N_7786,N_5671);
nor U10451 (N_10451,N_6610,N_7685);
and U10452 (N_10452,N_5987,N_7121);
and U10453 (N_10453,N_6588,N_5699);
or U10454 (N_10454,N_5826,N_6561);
and U10455 (N_10455,N_4155,N_7338);
nand U10456 (N_10456,N_5277,N_5947);
nor U10457 (N_10457,N_4720,N_7710);
xnor U10458 (N_10458,N_4109,N_5929);
nand U10459 (N_10459,N_5287,N_5041);
nor U10460 (N_10460,N_7405,N_4160);
or U10461 (N_10461,N_6142,N_4409);
nand U10462 (N_10462,N_4123,N_4085);
and U10463 (N_10463,N_7084,N_5805);
and U10464 (N_10464,N_4830,N_4575);
nor U10465 (N_10465,N_6666,N_6474);
or U10466 (N_10466,N_4549,N_4335);
nor U10467 (N_10467,N_5146,N_7662);
and U10468 (N_10468,N_7518,N_5323);
nand U10469 (N_10469,N_5870,N_6356);
xor U10470 (N_10470,N_5586,N_6966);
nor U10471 (N_10471,N_4094,N_5421);
nand U10472 (N_10472,N_5236,N_4434);
nor U10473 (N_10473,N_7605,N_4901);
and U10474 (N_10474,N_4348,N_4546);
nor U10475 (N_10475,N_5163,N_7084);
nand U10476 (N_10476,N_5901,N_6302);
and U10477 (N_10477,N_4350,N_5504);
nand U10478 (N_10478,N_7194,N_6908);
and U10479 (N_10479,N_4535,N_7965);
nand U10480 (N_10480,N_6810,N_5401);
nor U10481 (N_10481,N_4534,N_5722);
xnor U10482 (N_10482,N_7524,N_4251);
nand U10483 (N_10483,N_6589,N_5685);
nor U10484 (N_10484,N_5115,N_7263);
xnor U10485 (N_10485,N_4468,N_6685);
and U10486 (N_10486,N_7571,N_4355);
nor U10487 (N_10487,N_4151,N_6317);
and U10488 (N_10488,N_6663,N_6730);
nor U10489 (N_10489,N_7528,N_7446);
nand U10490 (N_10490,N_4702,N_4513);
xor U10491 (N_10491,N_7765,N_6014);
nor U10492 (N_10492,N_5419,N_6196);
and U10493 (N_10493,N_7890,N_5451);
nor U10494 (N_10494,N_7780,N_7450);
and U10495 (N_10495,N_4965,N_5865);
or U10496 (N_10496,N_5764,N_7369);
and U10497 (N_10497,N_5829,N_4987);
xnor U10498 (N_10498,N_7971,N_7698);
xor U10499 (N_10499,N_4054,N_7018);
nand U10500 (N_10500,N_7701,N_6672);
nor U10501 (N_10501,N_7451,N_7650);
nor U10502 (N_10502,N_7053,N_4268);
nor U10503 (N_10503,N_4936,N_5366);
nor U10504 (N_10504,N_4594,N_6880);
nor U10505 (N_10505,N_4588,N_6452);
nor U10506 (N_10506,N_6658,N_4178);
nand U10507 (N_10507,N_6915,N_7046);
xor U10508 (N_10508,N_4240,N_5084);
nor U10509 (N_10509,N_4679,N_4350);
nand U10510 (N_10510,N_4058,N_6629);
nand U10511 (N_10511,N_7536,N_5643);
nand U10512 (N_10512,N_7724,N_6582);
nor U10513 (N_10513,N_4234,N_7474);
and U10514 (N_10514,N_5712,N_7413);
nand U10515 (N_10515,N_5784,N_6099);
and U10516 (N_10516,N_4422,N_7425);
and U10517 (N_10517,N_4461,N_4458);
nand U10518 (N_10518,N_6315,N_5950);
nand U10519 (N_10519,N_5749,N_7776);
or U10520 (N_10520,N_7072,N_4891);
nand U10521 (N_10521,N_4538,N_6759);
or U10522 (N_10522,N_6319,N_7876);
nor U10523 (N_10523,N_7970,N_7957);
nand U10524 (N_10524,N_6694,N_4066);
nand U10525 (N_10525,N_4576,N_5086);
nand U10526 (N_10526,N_4223,N_6852);
and U10527 (N_10527,N_5551,N_5104);
nand U10528 (N_10528,N_4007,N_6749);
nand U10529 (N_10529,N_5193,N_5267);
nand U10530 (N_10530,N_5696,N_6155);
nand U10531 (N_10531,N_7711,N_6724);
xnor U10532 (N_10532,N_5330,N_5704);
nor U10533 (N_10533,N_5747,N_5484);
nor U10534 (N_10534,N_7689,N_7374);
or U10535 (N_10535,N_4708,N_7801);
and U10536 (N_10536,N_4441,N_7766);
and U10537 (N_10537,N_4557,N_5535);
nand U10538 (N_10538,N_4694,N_7541);
nor U10539 (N_10539,N_5646,N_5506);
or U10540 (N_10540,N_7838,N_5657);
nor U10541 (N_10541,N_4358,N_7013);
and U10542 (N_10542,N_5725,N_7634);
and U10543 (N_10543,N_7572,N_5380);
and U10544 (N_10544,N_4031,N_7507);
and U10545 (N_10545,N_4879,N_6192);
and U10546 (N_10546,N_6874,N_6148);
xnor U10547 (N_10547,N_6289,N_7288);
xor U10548 (N_10548,N_6089,N_6346);
nor U10549 (N_10549,N_4528,N_7943);
or U10550 (N_10550,N_7418,N_7847);
or U10551 (N_10551,N_5108,N_4283);
and U10552 (N_10552,N_5210,N_4279);
nor U10553 (N_10553,N_4020,N_4072);
and U10554 (N_10554,N_5941,N_5056);
or U10555 (N_10555,N_7819,N_4111);
nand U10556 (N_10556,N_5520,N_7512);
or U10557 (N_10557,N_7162,N_5850);
and U10558 (N_10558,N_7046,N_4495);
nand U10559 (N_10559,N_4412,N_7349);
and U10560 (N_10560,N_5649,N_7480);
nor U10561 (N_10561,N_6143,N_5084);
nor U10562 (N_10562,N_6429,N_5033);
and U10563 (N_10563,N_4326,N_7141);
nor U10564 (N_10564,N_6562,N_4495);
nand U10565 (N_10565,N_7314,N_5301);
xor U10566 (N_10566,N_4184,N_5427);
nor U10567 (N_10567,N_5623,N_5762);
or U10568 (N_10568,N_6006,N_5111);
and U10569 (N_10569,N_6617,N_5556);
xor U10570 (N_10570,N_4759,N_4065);
xor U10571 (N_10571,N_7247,N_4983);
and U10572 (N_10572,N_7147,N_6504);
xor U10573 (N_10573,N_7857,N_5285);
nand U10574 (N_10574,N_7915,N_6711);
and U10575 (N_10575,N_5015,N_7386);
or U10576 (N_10576,N_7569,N_6945);
or U10577 (N_10577,N_6407,N_4455);
and U10578 (N_10578,N_7363,N_6181);
xor U10579 (N_10579,N_5959,N_5063);
or U10580 (N_10580,N_6525,N_4961);
nand U10581 (N_10581,N_4931,N_4922);
nand U10582 (N_10582,N_4689,N_4825);
nor U10583 (N_10583,N_5183,N_5573);
and U10584 (N_10584,N_7135,N_4239);
or U10585 (N_10585,N_5438,N_7883);
or U10586 (N_10586,N_4172,N_5277);
nor U10587 (N_10587,N_4188,N_6906);
nand U10588 (N_10588,N_6477,N_5814);
xor U10589 (N_10589,N_5596,N_4041);
nand U10590 (N_10590,N_5880,N_6816);
nand U10591 (N_10591,N_6442,N_5813);
and U10592 (N_10592,N_6540,N_4352);
nand U10593 (N_10593,N_4457,N_6915);
nand U10594 (N_10594,N_4749,N_5949);
or U10595 (N_10595,N_4093,N_7131);
or U10596 (N_10596,N_6761,N_6369);
nand U10597 (N_10597,N_4983,N_6247);
nor U10598 (N_10598,N_6796,N_5254);
nand U10599 (N_10599,N_6366,N_5443);
nor U10600 (N_10600,N_4680,N_7562);
nand U10601 (N_10601,N_6426,N_6027);
xor U10602 (N_10602,N_4052,N_7107);
nor U10603 (N_10603,N_7560,N_7247);
or U10604 (N_10604,N_7481,N_7840);
nand U10605 (N_10605,N_4261,N_5061);
nand U10606 (N_10606,N_5917,N_6369);
xnor U10607 (N_10607,N_5531,N_6353);
and U10608 (N_10608,N_5372,N_5677);
xor U10609 (N_10609,N_4366,N_4250);
nand U10610 (N_10610,N_5750,N_6113);
or U10611 (N_10611,N_6046,N_4031);
and U10612 (N_10612,N_6628,N_6784);
or U10613 (N_10613,N_6912,N_4416);
nor U10614 (N_10614,N_5227,N_7102);
and U10615 (N_10615,N_4676,N_4994);
nor U10616 (N_10616,N_5782,N_4428);
or U10617 (N_10617,N_7031,N_6756);
nand U10618 (N_10618,N_4238,N_4988);
nor U10619 (N_10619,N_4623,N_5915);
or U10620 (N_10620,N_7073,N_6591);
or U10621 (N_10621,N_7262,N_4184);
nand U10622 (N_10622,N_6597,N_6157);
and U10623 (N_10623,N_6959,N_5640);
xnor U10624 (N_10624,N_5926,N_5799);
nand U10625 (N_10625,N_4366,N_6149);
or U10626 (N_10626,N_5392,N_4230);
or U10627 (N_10627,N_7977,N_7855);
or U10628 (N_10628,N_5459,N_4883);
nor U10629 (N_10629,N_6768,N_4171);
xor U10630 (N_10630,N_7800,N_7734);
or U10631 (N_10631,N_7364,N_5895);
nand U10632 (N_10632,N_4092,N_6125);
and U10633 (N_10633,N_4337,N_4451);
nand U10634 (N_10634,N_7590,N_4241);
or U10635 (N_10635,N_6954,N_4710);
nand U10636 (N_10636,N_6760,N_6614);
nor U10637 (N_10637,N_5545,N_4228);
xnor U10638 (N_10638,N_7176,N_7163);
and U10639 (N_10639,N_4888,N_5258);
nor U10640 (N_10640,N_7623,N_7904);
nand U10641 (N_10641,N_4326,N_7424);
nor U10642 (N_10642,N_5086,N_5612);
or U10643 (N_10643,N_7415,N_4008);
and U10644 (N_10644,N_4195,N_7292);
or U10645 (N_10645,N_7339,N_6903);
or U10646 (N_10646,N_4593,N_7069);
and U10647 (N_10647,N_4809,N_6773);
nand U10648 (N_10648,N_7703,N_5415);
nand U10649 (N_10649,N_7686,N_6750);
or U10650 (N_10650,N_7163,N_5565);
and U10651 (N_10651,N_7477,N_4636);
or U10652 (N_10652,N_4995,N_6413);
nor U10653 (N_10653,N_6417,N_5580);
or U10654 (N_10654,N_6757,N_4211);
nand U10655 (N_10655,N_5738,N_6694);
or U10656 (N_10656,N_6359,N_7266);
nand U10657 (N_10657,N_4295,N_5258);
and U10658 (N_10658,N_5092,N_4966);
nand U10659 (N_10659,N_4647,N_7519);
nor U10660 (N_10660,N_5589,N_4181);
or U10661 (N_10661,N_7723,N_7147);
or U10662 (N_10662,N_4061,N_7185);
or U10663 (N_10663,N_6985,N_6523);
or U10664 (N_10664,N_4088,N_4119);
and U10665 (N_10665,N_7520,N_5406);
or U10666 (N_10666,N_5981,N_7623);
and U10667 (N_10667,N_5002,N_5492);
nor U10668 (N_10668,N_4508,N_5805);
and U10669 (N_10669,N_4928,N_4472);
xnor U10670 (N_10670,N_6325,N_7522);
and U10671 (N_10671,N_7223,N_4400);
nor U10672 (N_10672,N_5569,N_6025);
nand U10673 (N_10673,N_5721,N_4293);
nor U10674 (N_10674,N_6037,N_6631);
nand U10675 (N_10675,N_6535,N_7855);
nor U10676 (N_10676,N_6435,N_5111);
nand U10677 (N_10677,N_6895,N_4253);
xnor U10678 (N_10678,N_4372,N_7492);
xor U10679 (N_10679,N_7745,N_6320);
nand U10680 (N_10680,N_7069,N_6289);
or U10681 (N_10681,N_4411,N_7315);
and U10682 (N_10682,N_5458,N_7191);
or U10683 (N_10683,N_4846,N_5359);
nor U10684 (N_10684,N_6485,N_5703);
or U10685 (N_10685,N_7912,N_6949);
or U10686 (N_10686,N_5953,N_7220);
nor U10687 (N_10687,N_5712,N_4787);
and U10688 (N_10688,N_5968,N_5136);
nor U10689 (N_10689,N_7874,N_4816);
nand U10690 (N_10690,N_5972,N_5445);
or U10691 (N_10691,N_5053,N_6915);
or U10692 (N_10692,N_5685,N_7657);
nand U10693 (N_10693,N_6184,N_7629);
nand U10694 (N_10694,N_4512,N_7742);
nor U10695 (N_10695,N_7807,N_5720);
xnor U10696 (N_10696,N_6066,N_5283);
or U10697 (N_10697,N_4628,N_5260);
nor U10698 (N_10698,N_5165,N_5055);
and U10699 (N_10699,N_4882,N_6682);
nand U10700 (N_10700,N_6082,N_4978);
nand U10701 (N_10701,N_4160,N_4307);
or U10702 (N_10702,N_6111,N_5675);
xnor U10703 (N_10703,N_4389,N_5890);
xnor U10704 (N_10704,N_4030,N_5763);
nor U10705 (N_10705,N_4454,N_6591);
nor U10706 (N_10706,N_6100,N_7052);
nand U10707 (N_10707,N_6924,N_7880);
nor U10708 (N_10708,N_7159,N_6617);
or U10709 (N_10709,N_6574,N_6679);
and U10710 (N_10710,N_4463,N_7106);
or U10711 (N_10711,N_6837,N_5538);
nor U10712 (N_10712,N_6774,N_6827);
nor U10713 (N_10713,N_7163,N_6530);
or U10714 (N_10714,N_6698,N_4005);
or U10715 (N_10715,N_5242,N_6966);
and U10716 (N_10716,N_6381,N_7374);
nand U10717 (N_10717,N_4589,N_4320);
xor U10718 (N_10718,N_6520,N_6355);
nand U10719 (N_10719,N_7516,N_4658);
or U10720 (N_10720,N_4841,N_7455);
or U10721 (N_10721,N_6391,N_5320);
nor U10722 (N_10722,N_5337,N_4354);
nor U10723 (N_10723,N_7429,N_6071);
nor U10724 (N_10724,N_5877,N_6161);
and U10725 (N_10725,N_7259,N_4010);
or U10726 (N_10726,N_6592,N_6457);
nand U10727 (N_10727,N_5106,N_7095);
or U10728 (N_10728,N_5632,N_7023);
nor U10729 (N_10729,N_7939,N_7143);
nor U10730 (N_10730,N_4107,N_6183);
or U10731 (N_10731,N_7627,N_4061);
and U10732 (N_10732,N_5688,N_7108);
nand U10733 (N_10733,N_5548,N_4283);
xor U10734 (N_10734,N_5526,N_5784);
and U10735 (N_10735,N_7442,N_5186);
and U10736 (N_10736,N_6847,N_6134);
nor U10737 (N_10737,N_7227,N_6994);
or U10738 (N_10738,N_5420,N_6574);
xor U10739 (N_10739,N_6060,N_7472);
or U10740 (N_10740,N_5934,N_5990);
nor U10741 (N_10741,N_4605,N_6980);
xnor U10742 (N_10742,N_7089,N_4590);
or U10743 (N_10743,N_6431,N_4574);
or U10744 (N_10744,N_4617,N_4641);
or U10745 (N_10745,N_7986,N_6027);
nor U10746 (N_10746,N_6049,N_7792);
or U10747 (N_10747,N_6836,N_5523);
nand U10748 (N_10748,N_4354,N_7436);
nor U10749 (N_10749,N_6235,N_5586);
nor U10750 (N_10750,N_5348,N_4334);
or U10751 (N_10751,N_4098,N_4534);
xor U10752 (N_10752,N_7048,N_4490);
and U10753 (N_10753,N_5452,N_6404);
or U10754 (N_10754,N_6858,N_6777);
or U10755 (N_10755,N_6773,N_5369);
and U10756 (N_10756,N_5572,N_5564);
xor U10757 (N_10757,N_4073,N_5835);
and U10758 (N_10758,N_7218,N_4976);
xnor U10759 (N_10759,N_4468,N_4242);
and U10760 (N_10760,N_6916,N_4044);
or U10761 (N_10761,N_5505,N_4419);
or U10762 (N_10762,N_4218,N_5827);
nor U10763 (N_10763,N_7101,N_7046);
or U10764 (N_10764,N_4508,N_6588);
or U10765 (N_10765,N_6044,N_4736);
or U10766 (N_10766,N_5777,N_6546);
nor U10767 (N_10767,N_6750,N_7368);
nand U10768 (N_10768,N_7365,N_4102);
and U10769 (N_10769,N_6267,N_4241);
and U10770 (N_10770,N_4611,N_5194);
nand U10771 (N_10771,N_4215,N_5025);
nor U10772 (N_10772,N_5041,N_7042);
nor U10773 (N_10773,N_6640,N_5866);
and U10774 (N_10774,N_6217,N_4384);
and U10775 (N_10775,N_7402,N_5403);
nor U10776 (N_10776,N_7453,N_6638);
and U10777 (N_10777,N_7065,N_7490);
nor U10778 (N_10778,N_5510,N_4684);
nor U10779 (N_10779,N_4153,N_5351);
or U10780 (N_10780,N_4353,N_6728);
nor U10781 (N_10781,N_7988,N_6643);
nor U10782 (N_10782,N_7140,N_4943);
nand U10783 (N_10783,N_5046,N_4190);
nand U10784 (N_10784,N_6941,N_4538);
nor U10785 (N_10785,N_7486,N_6910);
and U10786 (N_10786,N_6578,N_5654);
and U10787 (N_10787,N_7929,N_6637);
or U10788 (N_10788,N_4881,N_5271);
and U10789 (N_10789,N_7639,N_4986);
xnor U10790 (N_10790,N_6726,N_5667);
or U10791 (N_10791,N_4919,N_5320);
nand U10792 (N_10792,N_7438,N_7498);
nand U10793 (N_10793,N_7952,N_5474);
nand U10794 (N_10794,N_5582,N_6903);
or U10795 (N_10795,N_5917,N_6954);
nand U10796 (N_10796,N_6341,N_6752);
xnor U10797 (N_10797,N_6572,N_6264);
nand U10798 (N_10798,N_6261,N_7184);
nor U10799 (N_10799,N_6372,N_7578);
xnor U10800 (N_10800,N_5795,N_5097);
nand U10801 (N_10801,N_4079,N_4977);
xor U10802 (N_10802,N_5224,N_5437);
nor U10803 (N_10803,N_6925,N_4009);
and U10804 (N_10804,N_7157,N_4623);
and U10805 (N_10805,N_7179,N_5550);
and U10806 (N_10806,N_7808,N_5512);
or U10807 (N_10807,N_5338,N_6252);
and U10808 (N_10808,N_6756,N_4315);
and U10809 (N_10809,N_4871,N_5537);
xor U10810 (N_10810,N_5888,N_7490);
nor U10811 (N_10811,N_5384,N_5640);
or U10812 (N_10812,N_5215,N_6785);
xor U10813 (N_10813,N_5424,N_7293);
nor U10814 (N_10814,N_4406,N_5500);
nand U10815 (N_10815,N_6067,N_5380);
nor U10816 (N_10816,N_6377,N_6370);
nand U10817 (N_10817,N_5035,N_7310);
and U10818 (N_10818,N_4695,N_7595);
and U10819 (N_10819,N_5312,N_4188);
nand U10820 (N_10820,N_4985,N_4648);
nor U10821 (N_10821,N_6769,N_4525);
xor U10822 (N_10822,N_6982,N_6572);
nor U10823 (N_10823,N_4471,N_4358);
or U10824 (N_10824,N_4698,N_5030);
and U10825 (N_10825,N_4209,N_5983);
nor U10826 (N_10826,N_5363,N_4404);
nand U10827 (N_10827,N_5396,N_4572);
nor U10828 (N_10828,N_6124,N_5383);
and U10829 (N_10829,N_4426,N_6265);
nor U10830 (N_10830,N_4636,N_6974);
nand U10831 (N_10831,N_4410,N_4479);
and U10832 (N_10832,N_6186,N_7649);
and U10833 (N_10833,N_5176,N_5174);
nor U10834 (N_10834,N_7249,N_4079);
or U10835 (N_10835,N_5122,N_6776);
nor U10836 (N_10836,N_4868,N_4980);
and U10837 (N_10837,N_4725,N_5870);
nor U10838 (N_10838,N_4203,N_5812);
nor U10839 (N_10839,N_7845,N_5132);
xor U10840 (N_10840,N_7694,N_7177);
and U10841 (N_10841,N_7731,N_6738);
or U10842 (N_10842,N_7715,N_5592);
or U10843 (N_10843,N_5050,N_7873);
and U10844 (N_10844,N_4880,N_6772);
and U10845 (N_10845,N_4887,N_4166);
or U10846 (N_10846,N_6306,N_5883);
nand U10847 (N_10847,N_7418,N_4116);
and U10848 (N_10848,N_5579,N_4647);
nor U10849 (N_10849,N_5089,N_4012);
and U10850 (N_10850,N_6469,N_4799);
nor U10851 (N_10851,N_7907,N_7847);
or U10852 (N_10852,N_6515,N_7582);
nand U10853 (N_10853,N_7410,N_6353);
nand U10854 (N_10854,N_5841,N_4764);
nor U10855 (N_10855,N_5495,N_6615);
nand U10856 (N_10856,N_6253,N_6073);
xor U10857 (N_10857,N_5976,N_6095);
nand U10858 (N_10858,N_4922,N_6542);
nor U10859 (N_10859,N_6739,N_4618);
or U10860 (N_10860,N_6795,N_4614);
nor U10861 (N_10861,N_5520,N_4056);
and U10862 (N_10862,N_7922,N_7888);
nor U10863 (N_10863,N_7925,N_6770);
and U10864 (N_10864,N_5105,N_7434);
or U10865 (N_10865,N_7495,N_6929);
and U10866 (N_10866,N_4945,N_5796);
or U10867 (N_10867,N_4594,N_4738);
nand U10868 (N_10868,N_5044,N_6355);
and U10869 (N_10869,N_5137,N_5208);
nor U10870 (N_10870,N_4356,N_7381);
nand U10871 (N_10871,N_6705,N_4246);
or U10872 (N_10872,N_5109,N_4271);
nand U10873 (N_10873,N_4893,N_4079);
or U10874 (N_10874,N_5536,N_7439);
nand U10875 (N_10875,N_5159,N_6944);
nor U10876 (N_10876,N_5653,N_6765);
nor U10877 (N_10877,N_5988,N_6452);
nand U10878 (N_10878,N_5293,N_5229);
nand U10879 (N_10879,N_4958,N_7246);
nand U10880 (N_10880,N_7804,N_5732);
nand U10881 (N_10881,N_5029,N_4827);
nand U10882 (N_10882,N_6048,N_6298);
and U10883 (N_10883,N_7253,N_5448);
nor U10884 (N_10884,N_6433,N_4179);
xnor U10885 (N_10885,N_7067,N_5396);
nor U10886 (N_10886,N_4298,N_5855);
or U10887 (N_10887,N_6800,N_5651);
or U10888 (N_10888,N_4271,N_6117);
nor U10889 (N_10889,N_6202,N_7449);
xor U10890 (N_10890,N_5193,N_7477);
nand U10891 (N_10891,N_6963,N_7955);
nor U10892 (N_10892,N_7398,N_4197);
nand U10893 (N_10893,N_6222,N_7856);
or U10894 (N_10894,N_5895,N_6607);
nor U10895 (N_10895,N_4737,N_7733);
nor U10896 (N_10896,N_6942,N_6299);
nand U10897 (N_10897,N_5828,N_5379);
nor U10898 (N_10898,N_4530,N_7260);
xor U10899 (N_10899,N_7392,N_6921);
nand U10900 (N_10900,N_4695,N_5308);
nor U10901 (N_10901,N_4625,N_5494);
nand U10902 (N_10902,N_7641,N_5212);
nand U10903 (N_10903,N_6615,N_4467);
and U10904 (N_10904,N_6149,N_4804);
nand U10905 (N_10905,N_5746,N_4739);
nand U10906 (N_10906,N_7342,N_5568);
and U10907 (N_10907,N_4957,N_4534);
nand U10908 (N_10908,N_4585,N_7947);
and U10909 (N_10909,N_6434,N_4489);
and U10910 (N_10910,N_7913,N_6212);
and U10911 (N_10911,N_4819,N_4856);
and U10912 (N_10912,N_6984,N_6986);
or U10913 (N_10913,N_6313,N_6572);
or U10914 (N_10914,N_5848,N_5037);
nor U10915 (N_10915,N_6539,N_4915);
or U10916 (N_10916,N_6569,N_5718);
or U10917 (N_10917,N_5465,N_6728);
nor U10918 (N_10918,N_6749,N_6400);
nand U10919 (N_10919,N_4294,N_4293);
and U10920 (N_10920,N_5092,N_4702);
xnor U10921 (N_10921,N_5342,N_4755);
xor U10922 (N_10922,N_6676,N_4348);
or U10923 (N_10923,N_4454,N_6249);
xor U10924 (N_10924,N_6744,N_4662);
or U10925 (N_10925,N_4457,N_7934);
xor U10926 (N_10926,N_5733,N_6861);
nand U10927 (N_10927,N_6036,N_7031);
xor U10928 (N_10928,N_4999,N_6725);
xnor U10929 (N_10929,N_4976,N_6102);
or U10930 (N_10930,N_6453,N_6065);
xor U10931 (N_10931,N_4172,N_4631);
or U10932 (N_10932,N_4840,N_6544);
nor U10933 (N_10933,N_7328,N_6137);
nor U10934 (N_10934,N_7867,N_6453);
and U10935 (N_10935,N_7707,N_4267);
or U10936 (N_10936,N_4211,N_6399);
or U10937 (N_10937,N_7915,N_5764);
or U10938 (N_10938,N_6520,N_6370);
nand U10939 (N_10939,N_7924,N_6959);
xor U10940 (N_10940,N_6078,N_6203);
nand U10941 (N_10941,N_7728,N_6508);
nor U10942 (N_10942,N_4580,N_4560);
nor U10943 (N_10943,N_6256,N_4895);
nand U10944 (N_10944,N_5628,N_4863);
or U10945 (N_10945,N_5066,N_6557);
or U10946 (N_10946,N_5436,N_4416);
nand U10947 (N_10947,N_6278,N_7352);
nand U10948 (N_10948,N_4464,N_7734);
or U10949 (N_10949,N_7968,N_4278);
and U10950 (N_10950,N_7192,N_5567);
or U10951 (N_10951,N_5864,N_6615);
nor U10952 (N_10952,N_7594,N_7451);
nor U10953 (N_10953,N_6115,N_5663);
nor U10954 (N_10954,N_6196,N_5644);
nor U10955 (N_10955,N_7869,N_5366);
nand U10956 (N_10956,N_7422,N_4505);
nand U10957 (N_10957,N_6817,N_7170);
nor U10958 (N_10958,N_4354,N_4103);
nor U10959 (N_10959,N_4206,N_5198);
nor U10960 (N_10960,N_5979,N_7904);
nand U10961 (N_10961,N_4452,N_4244);
or U10962 (N_10962,N_6232,N_6491);
nor U10963 (N_10963,N_4099,N_5764);
or U10964 (N_10964,N_7471,N_4037);
and U10965 (N_10965,N_5629,N_7762);
xnor U10966 (N_10966,N_5884,N_4087);
nand U10967 (N_10967,N_5185,N_7491);
xnor U10968 (N_10968,N_5665,N_4657);
and U10969 (N_10969,N_7722,N_5669);
or U10970 (N_10970,N_7196,N_4979);
and U10971 (N_10971,N_4984,N_5206);
and U10972 (N_10972,N_4534,N_7713);
nand U10973 (N_10973,N_4538,N_4236);
nand U10974 (N_10974,N_7565,N_7677);
and U10975 (N_10975,N_5975,N_7445);
and U10976 (N_10976,N_6631,N_4817);
and U10977 (N_10977,N_7146,N_6342);
nor U10978 (N_10978,N_6579,N_6513);
or U10979 (N_10979,N_7002,N_5575);
and U10980 (N_10980,N_6536,N_4695);
nand U10981 (N_10981,N_5445,N_7718);
or U10982 (N_10982,N_6551,N_6977);
nand U10983 (N_10983,N_6840,N_7619);
nand U10984 (N_10984,N_4267,N_5305);
and U10985 (N_10985,N_6732,N_7089);
and U10986 (N_10986,N_7970,N_7891);
or U10987 (N_10987,N_5893,N_7400);
and U10988 (N_10988,N_5215,N_4678);
xor U10989 (N_10989,N_4031,N_5431);
xor U10990 (N_10990,N_7784,N_7586);
or U10991 (N_10991,N_5732,N_7208);
and U10992 (N_10992,N_4951,N_7545);
xor U10993 (N_10993,N_7065,N_5068);
xnor U10994 (N_10994,N_5406,N_5263);
or U10995 (N_10995,N_4976,N_5219);
nor U10996 (N_10996,N_7529,N_6904);
or U10997 (N_10997,N_5358,N_4105);
and U10998 (N_10998,N_4712,N_5573);
nand U10999 (N_10999,N_6591,N_6786);
nor U11000 (N_11000,N_4619,N_7940);
and U11001 (N_11001,N_5881,N_5840);
xor U11002 (N_11002,N_4432,N_6632);
nand U11003 (N_11003,N_6610,N_6429);
and U11004 (N_11004,N_7062,N_4474);
and U11005 (N_11005,N_6913,N_6783);
and U11006 (N_11006,N_6550,N_6767);
and U11007 (N_11007,N_6045,N_5669);
and U11008 (N_11008,N_6961,N_4485);
nand U11009 (N_11009,N_5114,N_5649);
xnor U11010 (N_11010,N_6476,N_5030);
and U11011 (N_11011,N_5613,N_5565);
nor U11012 (N_11012,N_6257,N_7254);
nor U11013 (N_11013,N_7443,N_4660);
or U11014 (N_11014,N_5028,N_5723);
nand U11015 (N_11015,N_4893,N_4335);
or U11016 (N_11016,N_4475,N_4716);
nor U11017 (N_11017,N_6993,N_7958);
or U11018 (N_11018,N_7448,N_4362);
nor U11019 (N_11019,N_5408,N_5473);
nor U11020 (N_11020,N_7627,N_4847);
and U11021 (N_11021,N_6992,N_6412);
nor U11022 (N_11022,N_6402,N_5431);
nor U11023 (N_11023,N_7411,N_6135);
nor U11024 (N_11024,N_4954,N_4605);
nand U11025 (N_11025,N_4829,N_7166);
nand U11026 (N_11026,N_6068,N_5649);
and U11027 (N_11027,N_5827,N_6718);
and U11028 (N_11028,N_6197,N_4562);
xor U11029 (N_11029,N_5686,N_6783);
nor U11030 (N_11030,N_6200,N_7456);
nor U11031 (N_11031,N_5848,N_5846);
or U11032 (N_11032,N_4548,N_4891);
nand U11033 (N_11033,N_6332,N_4865);
and U11034 (N_11034,N_5452,N_7683);
nor U11035 (N_11035,N_7772,N_7918);
nand U11036 (N_11036,N_7604,N_5094);
nand U11037 (N_11037,N_7229,N_4981);
nor U11038 (N_11038,N_7770,N_4627);
and U11039 (N_11039,N_6117,N_6292);
nor U11040 (N_11040,N_7308,N_7417);
and U11041 (N_11041,N_7100,N_5037);
nand U11042 (N_11042,N_7800,N_5603);
nor U11043 (N_11043,N_5229,N_4077);
nand U11044 (N_11044,N_6058,N_5933);
nor U11045 (N_11045,N_4282,N_6042);
nor U11046 (N_11046,N_5256,N_7962);
and U11047 (N_11047,N_5742,N_6447);
nand U11048 (N_11048,N_4776,N_4147);
and U11049 (N_11049,N_7389,N_6054);
nor U11050 (N_11050,N_4061,N_6102);
nand U11051 (N_11051,N_4585,N_7467);
nor U11052 (N_11052,N_5853,N_4836);
and U11053 (N_11053,N_7913,N_6098);
nor U11054 (N_11054,N_7830,N_6820);
nor U11055 (N_11055,N_5364,N_7391);
and U11056 (N_11056,N_6844,N_5961);
and U11057 (N_11057,N_4745,N_7880);
and U11058 (N_11058,N_5766,N_4930);
xnor U11059 (N_11059,N_4654,N_4777);
or U11060 (N_11060,N_5916,N_7915);
xor U11061 (N_11061,N_6043,N_5644);
xnor U11062 (N_11062,N_4497,N_4123);
nand U11063 (N_11063,N_6783,N_5875);
nand U11064 (N_11064,N_4357,N_7734);
and U11065 (N_11065,N_5320,N_7443);
xor U11066 (N_11066,N_6088,N_6857);
and U11067 (N_11067,N_4797,N_4851);
xnor U11068 (N_11068,N_4612,N_7965);
and U11069 (N_11069,N_7657,N_6593);
nor U11070 (N_11070,N_5931,N_6316);
and U11071 (N_11071,N_6341,N_4350);
nand U11072 (N_11072,N_7760,N_4431);
nand U11073 (N_11073,N_5045,N_5197);
nor U11074 (N_11074,N_6927,N_5024);
or U11075 (N_11075,N_6129,N_4788);
nand U11076 (N_11076,N_5445,N_5826);
nand U11077 (N_11077,N_5482,N_5716);
xor U11078 (N_11078,N_6764,N_7678);
nor U11079 (N_11079,N_4428,N_5617);
xnor U11080 (N_11080,N_4559,N_6201);
or U11081 (N_11081,N_7202,N_4788);
nor U11082 (N_11082,N_5871,N_6667);
and U11083 (N_11083,N_6317,N_5455);
and U11084 (N_11084,N_4542,N_7544);
nand U11085 (N_11085,N_5269,N_5533);
nor U11086 (N_11086,N_7583,N_6644);
and U11087 (N_11087,N_6717,N_6759);
or U11088 (N_11088,N_5872,N_5788);
and U11089 (N_11089,N_7357,N_5833);
nor U11090 (N_11090,N_6123,N_7170);
nor U11091 (N_11091,N_7763,N_4942);
nand U11092 (N_11092,N_6972,N_7683);
or U11093 (N_11093,N_4081,N_7795);
and U11094 (N_11094,N_5896,N_7581);
xnor U11095 (N_11095,N_6174,N_5831);
and U11096 (N_11096,N_4488,N_7401);
and U11097 (N_11097,N_6528,N_4558);
or U11098 (N_11098,N_4129,N_7045);
or U11099 (N_11099,N_6807,N_7365);
or U11100 (N_11100,N_6589,N_5808);
xnor U11101 (N_11101,N_4070,N_5601);
and U11102 (N_11102,N_5560,N_6246);
nor U11103 (N_11103,N_5062,N_4479);
or U11104 (N_11104,N_7187,N_4091);
nor U11105 (N_11105,N_4561,N_6278);
nand U11106 (N_11106,N_4557,N_7224);
nor U11107 (N_11107,N_7104,N_7854);
nand U11108 (N_11108,N_5256,N_4448);
nand U11109 (N_11109,N_5188,N_5554);
nand U11110 (N_11110,N_7082,N_4140);
or U11111 (N_11111,N_5513,N_5592);
nand U11112 (N_11112,N_4286,N_5099);
or U11113 (N_11113,N_4747,N_6053);
nor U11114 (N_11114,N_4369,N_5461);
or U11115 (N_11115,N_4270,N_5963);
or U11116 (N_11116,N_5966,N_7565);
or U11117 (N_11117,N_5484,N_6328);
or U11118 (N_11118,N_5233,N_4813);
or U11119 (N_11119,N_6891,N_5168);
nor U11120 (N_11120,N_7799,N_4860);
nand U11121 (N_11121,N_5263,N_7145);
nor U11122 (N_11122,N_4277,N_4590);
or U11123 (N_11123,N_7871,N_4419);
nand U11124 (N_11124,N_7510,N_4557);
or U11125 (N_11125,N_5114,N_7932);
or U11126 (N_11126,N_5650,N_4871);
and U11127 (N_11127,N_4425,N_7212);
nand U11128 (N_11128,N_7565,N_7101);
xor U11129 (N_11129,N_7105,N_5290);
nor U11130 (N_11130,N_6660,N_5117);
and U11131 (N_11131,N_6880,N_6147);
or U11132 (N_11132,N_5986,N_7075);
and U11133 (N_11133,N_6351,N_4830);
or U11134 (N_11134,N_5400,N_5777);
nor U11135 (N_11135,N_7798,N_7859);
nor U11136 (N_11136,N_7197,N_6247);
nand U11137 (N_11137,N_5714,N_4092);
or U11138 (N_11138,N_4099,N_4383);
and U11139 (N_11139,N_6863,N_6920);
and U11140 (N_11140,N_5669,N_4919);
or U11141 (N_11141,N_4759,N_7203);
nand U11142 (N_11142,N_4419,N_6262);
or U11143 (N_11143,N_4117,N_5949);
xor U11144 (N_11144,N_6759,N_7508);
xor U11145 (N_11145,N_6312,N_6845);
xor U11146 (N_11146,N_6156,N_7143);
nor U11147 (N_11147,N_6085,N_5490);
nor U11148 (N_11148,N_5679,N_4215);
nand U11149 (N_11149,N_4563,N_6306);
xnor U11150 (N_11150,N_7341,N_7435);
or U11151 (N_11151,N_4721,N_4869);
nor U11152 (N_11152,N_5320,N_4537);
nand U11153 (N_11153,N_7879,N_6362);
and U11154 (N_11154,N_6389,N_7489);
and U11155 (N_11155,N_7146,N_4059);
and U11156 (N_11156,N_7336,N_4262);
nand U11157 (N_11157,N_5652,N_5075);
nand U11158 (N_11158,N_5112,N_4259);
or U11159 (N_11159,N_4046,N_4036);
or U11160 (N_11160,N_7110,N_5693);
or U11161 (N_11161,N_4759,N_6707);
nor U11162 (N_11162,N_5743,N_4033);
and U11163 (N_11163,N_5807,N_4401);
xor U11164 (N_11164,N_6292,N_7858);
xnor U11165 (N_11165,N_6303,N_5360);
and U11166 (N_11166,N_6162,N_6152);
xnor U11167 (N_11167,N_4575,N_5919);
and U11168 (N_11168,N_5697,N_4295);
xor U11169 (N_11169,N_6709,N_6061);
and U11170 (N_11170,N_7605,N_6769);
and U11171 (N_11171,N_6607,N_5255);
xor U11172 (N_11172,N_6798,N_6263);
nor U11173 (N_11173,N_5442,N_4869);
and U11174 (N_11174,N_4716,N_5068);
and U11175 (N_11175,N_4227,N_4838);
nor U11176 (N_11176,N_6584,N_6770);
or U11177 (N_11177,N_7701,N_7518);
nand U11178 (N_11178,N_7789,N_7906);
nor U11179 (N_11179,N_5650,N_4900);
and U11180 (N_11180,N_4887,N_4225);
and U11181 (N_11181,N_6853,N_4996);
and U11182 (N_11182,N_7620,N_6604);
and U11183 (N_11183,N_6183,N_7987);
and U11184 (N_11184,N_6443,N_5347);
nor U11185 (N_11185,N_7581,N_7210);
and U11186 (N_11186,N_4651,N_5541);
or U11187 (N_11187,N_7910,N_4068);
nand U11188 (N_11188,N_7486,N_4516);
and U11189 (N_11189,N_7410,N_6755);
or U11190 (N_11190,N_6686,N_7984);
or U11191 (N_11191,N_4482,N_6330);
and U11192 (N_11192,N_7870,N_7066);
nand U11193 (N_11193,N_4217,N_5163);
and U11194 (N_11194,N_5392,N_7828);
or U11195 (N_11195,N_6375,N_5611);
nor U11196 (N_11196,N_6367,N_5177);
or U11197 (N_11197,N_5812,N_5573);
and U11198 (N_11198,N_4135,N_5972);
and U11199 (N_11199,N_5144,N_6685);
nor U11200 (N_11200,N_6608,N_5290);
nor U11201 (N_11201,N_5122,N_5568);
nand U11202 (N_11202,N_6738,N_4117);
xnor U11203 (N_11203,N_4224,N_5198);
or U11204 (N_11204,N_7480,N_5981);
and U11205 (N_11205,N_6150,N_4804);
or U11206 (N_11206,N_4459,N_4223);
xnor U11207 (N_11207,N_4001,N_5339);
or U11208 (N_11208,N_7983,N_4884);
or U11209 (N_11209,N_5034,N_6414);
xor U11210 (N_11210,N_5219,N_4148);
and U11211 (N_11211,N_6001,N_7210);
and U11212 (N_11212,N_7865,N_4631);
and U11213 (N_11213,N_6301,N_4770);
nand U11214 (N_11214,N_7360,N_7436);
and U11215 (N_11215,N_4680,N_4080);
nand U11216 (N_11216,N_7617,N_5311);
or U11217 (N_11217,N_7528,N_6626);
and U11218 (N_11218,N_4502,N_4522);
or U11219 (N_11219,N_7553,N_6014);
nor U11220 (N_11220,N_7199,N_5076);
xor U11221 (N_11221,N_7928,N_7874);
and U11222 (N_11222,N_5161,N_7504);
nor U11223 (N_11223,N_6576,N_4978);
nand U11224 (N_11224,N_7997,N_4670);
xor U11225 (N_11225,N_5907,N_7646);
and U11226 (N_11226,N_6797,N_5428);
and U11227 (N_11227,N_7842,N_5091);
xnor U11228 (N_11228,N_7000,N_7315);
or U11229 (N_11229,N_4110,N_6552);
nor U11230 (N_11230,N_6727,N_5077);
nand U11231 (N_11231,N_6631,N_7834);
nor U11232 (N_11232,N_6526,N_5834);
or U11233 (N_11233,N_7783,N_5873);
and U11234 (N_11234,N_4602,N_5900);
and U11235 (N_11235,N_6762,N_7941);
nand U11236 (N_11236,N_4353,N_4120);
and U11237 (N_11237,N_7755,N_6879);
and U11238 (N_11238,N_6855,N_6153);
nor U11239 (N_11239,N_4107,N_5204);
nand U11240 (N_11240,N_7998,N_4650);
or U11241 (N_11241,N_4460,N_6268);
and U11242 (N_11242,N_5626,N_5480);
or U11243 (N_11243,N_4832,N_5354);
and U11244 (N_11244,N_4932,N_4041);
nor U11245 (N_11245,N_7199,N_6152);
nand U11246 (N_11246,N_7330,N_4006);
xnor U11247 (N_11247,N_5743,N_4319);
or U11248 (N_11248,N_7913,N_4218);
nand U11249 (N_11249,N_6190,N_7962);
nor U11250 (N_11250,N_5863,N_4178);
or U11251 (N_11251,N_6542,N_4405);
and U11252 (N_11252,N_6850,N_6940);
nor U11253 (N_11253,N_6894,N_6657);
xnor U11254 (N_11254,N_6355,N_4717);
or U11255 (N_11255,N_5702,N_4709);
xor U11256 (N_11256,N_6654,N_6565);
nand U11257 (N_11257,N_7761,N_5179);
nor U11258 (N_11258,N_4710,N_4800);
nor U11259 (N_11259,N_4990,N_7808);
nand U11260 (N_11260,N_5357,N_5190);
or U11261 (N_11261,N_7085,N_7487);
xor U11262 (N_11262,N_7661,N_7624);
nand U11263 (N_11263,N_7309,N_5851);
and U11264 (N_11264,N_5145,N_6564);
or U11265 (N_11265,N_7560,N_7786);
nand U11266 (N_11266,N_7418,N_5455);
nand U11267 (N_11267,N_5996,N_7616);
nand U11268 (N_11268,N_6608,N_6995);
nand U11269 (N_11269,N_6435,N_6183);
nor U11270 (N_11270,N_5824,N_6051);
nor U11271 (N_11271,N_5909,N_6931);
and U11272 (N_11272,N_7301,N_7887);
or U11273 (N_11273,N_6677,N_6717);
and U11274 (N_11274,N_5461,N_7893);
nor U11275 (N_11275,N_4023,N_4245);
nor U11276 (N_11276,N_6346,N_7018);
nor U11277 (N_11277,N_6629,N_5805);
or U11278 (N_11278,N_7777,N_4281);
nand U11279 (N_11279,N_5648,N_7702);
xor U11280 (N_11280,N_7279,N_5068);
or U11281 (N_11281,N_4197,N_7189);
xnor U11282 (N_11282,N_4366,N_6710);
or U11283 (N_11283,N_5932,N_6278);
or U11284 (N_11284,N_7016,N_4919);
or U11285 (N_11285,N_7784,N_7562);
and U11286 (N_11286,N_7238,N_5159);
or U11287 (N_11287,N_4026,N_4014);
nand U11288 (N_11288,N_6568,N_7986);
and U11289 (N_11289,N_7915,N_4467);
xor U11290 (N_11290,N_7908,N_6016);
nand U11291 (N_11291,N_5394,N_4597);
or U11292 (N_11292,N_4640,N_4688);
or U11293 (N_11293,N_4694,N_7298);
nand U11294 (N_11294,N_7645,N_4818);
and U11295 (N_11295,N_5264,N_6676);
nand U11296 (N_11296,N_5814,N_5090);
and U11297 (N_11297,N_6722,N_6182);
or U11298 (N_11298,N_4821,N_7279);
and U11299 (N_11299,N_5249,N_4451);
xnor U11300 (N_11300,N_5625,N_5578);
nand U11301 (N_11301,N_6378,N_4373);
nand U11302 (N_11302,N_4766,N_5247);
nor U11303 (N_11303,N_6283,N_5011);
or U11304 (N_11304,N_5705,N_6548);
or U11305 (N_11305,N_4869,N_4205);
nor U11306 (N_11306,N_4747,N_5074);
xnor U11307 (N_11307,N_7479,N_4444);
and U11308 (N_11308,N_5329,N_6889);
and U11309 (N_11309,N_7606,N_7162);
and U11310 (N_11310,N_7438,N_5990);
nand U11311 (N_11311,N_6435,N_4689);
or U11312 (N_11312,N_5116,N_6066);
and U11313 (N_11313,N_6070,N_6577);
or U11314 (N_11314,N_7301,N_7334);
xor U11315 (N_11315,N_4983,N_5699);
nand U11316 (N_11316,N_6405,N_6152);
nand U11317 (N_11317,N_6272,N_5916);
and U11318 (N_11318,N_5524,N_7995);
and U11319 (N_11319,N_5452,N_7603);
or U11320 (N_11320,N_6055,N_7122);
and U11321 (N_11321,N_7053,N_6555);
and U11322 (N_11322,N_5869,N_6974);
nor U11323 (N_11323,N_5588,N_6948);
nand U11324 (N_11324,N_4337,N_4459);
xor U11325 (N_11325,N_7924,N_4204);
nor U11326 (N_11326,N_5578,N_6011);
or U11327 (N_11327,N_5203,N_6106);
xnor U11328 (N_11328,N_4065,N_6496);
or U11329 (N_11329,N_5788,N_6595);
and U11330 (N_11330,N_6047,N_7078);
and U11331 (N_11331,N_7421,N_5973);
nand U11332 (N_11332,N_7515,N_6812);
and U11333 (N_11333,N_6966,N_6375);
nand U11334 (N_11334,N_5369,N_4781);
nand U11335 (N_11335,N_6144,N_4032);
nor U11336 (N_11336,N_4480,N_6846);
nand U11337 (N_11337,N_5987,N_7985);
xor U11338 (N_11338,N_7151,N_5321);
nand U11339 (N_11339,N_6021,N_6723);
nand U11340 (N_11340,N_4366,N_6289);
xnor U11341 (N_11341,N_7818,N_6646);
and U11342 (N_11342,N_5343,N_7852);
nor U11343 (N_11343,N_4083,N_7533);
and U11344 (N_11344,N_5167,N_7469);
nand U11345 (N_11345,N_7170,N_6887);
and U11346 (N_11346,N_7414,N_5544);
and U11347 (N_11347,N_7542,N_4351);
and U11348 (N_11348,N_6134,N_4378);
and U11349 (N_11349,N_4437,N_5654);
or U11350 (N_11350,N_6732,N_6794);
and U11351 (N_11351,N_4878,N_6539);
nand U11352 (N_11352,N_4027,N_7385);
nor U11353 (N_11353,N_4070,N_4795);
nand U11354 (N_11354,N_5792,N_6222);
or U11355 (N_11355,N_7374,N_5072);
or U11356 (N_11356,N_4010,N_5029);
and U11357 (N_11357,N_4840,N_6819);
nand U11358 (N_11358,N_5606,N_5425);
and U11359 (N_11359,N_4387,N_4482);
nor U11360 (N_11360,N_7235,N_7770);
nand U11361 (N_11361,N_7827,N_7950);
nor U11362 (N_11362,N_7261,N_7609);
xor U11363 (N_11363,N_4049,N_6787);
nor U11364 (N_11364,N_7350,N_7793);
nand U11365 (N_11365,N_4197,N_6836);
and U11366 (N_11366,N_7764,N_5943);
nor U11367 (N_11367,N_7272,N_4821);
nor U11368 (N_11368,N_4297,N_7950);
and U11369 (N_11369,N_7063,N_7090);
and U11370 (N_11370,N_4451,N_7541);
or U11371 (N_11371,N_6450,N_5920);
and U11372 (N_11372,N_5606,N_7507);
xnor U11373 (N_11373,N_4119,N_4691);
and U11374 (N_11374,N_5807,N_6933);
or U11375 (N_11375,N_6898,N_5408);
xnor U11376 (N_11376,N_5681,N_4927);
nor U11377 (N_11377,N_4737,N_5046);
or U11378 (N_11378,N_4498,N_6991);
and U11379 (N_11379,N_4776,N_5010);
and U11380 (N_11380,N_6572,N_7843);
xnor U11381 (N_11381,N_6291,N_7688);
nand U11382 (N_11382,N_7613,N_4911);
or U11383 (N_11383,N_7915,N_4364);
nor U11384 (N_11384,N_5603,N_4089);
nand U11385 (N_11385,N_5229,N_5457);
or U11386 (N_11386,N_4408,N_7935);
xor U11387 (N_11387,N_7652,N_5746);
nor U11388 (N_11388,N_7532,N_5220);
or U11389 (N_11389,N_6870,N_5920);
nor U11390 (N_11390,N_7921,N_4711);
nor U11391 (N_11391,N_6065,N_6851);
nand U11392 (N_11392,N_6545,N_4997);
or U11393 (N_11393,N_4823,N_6822);
nor U11394 (N_11394,N_6197,N_5649);
nor U11395 (N_11395,N_7535,N_7382);
and U11396 (N_11396,N_4036,N_7445);
nand U11397 (N_11397,N_6915,N_4839);
or U11398 (N_11398,N_4387,N_4332);
nor U11399 (N_11399,N_7986,N_6572);
or U11400 (N_11400,N_4544,N_4342);
and U11401 (N_11401,N_6585,N_5763);
or U11402 (N_11402,N_7164,N_6796);
nand U11403 (N_11403,N_7342,N_7691);
nor U11404 (N_11404,N_7627,N_7197);
nand U11405 (N_11405,N_6283,N_5400);
and U11406 (N_11406,N_6389,N_4561);
or U11407 (N_11407,N_4946,N_5286);
nand U11408 (N_11408,N_4313,N_5604);
nand U11409 (N_11409,N_7018,N_4296);
or U11410 (N_11410,N_5094,N_4211);
and U11411 (N_11411,N_5659,N_5078);
xnor U11412 (N_11412,N_7469,N_6334);
and U11413 (N_11413,N_5635,N_4720);
nand U11414 (N_11414,N_7030,N_4743);
nand U11415 (N_11415,N_4222,N_5596);
and U11416 (N_11416,N_7318,N_5895);
nor U11417 (N_11417,N_7938,N_7580);
xnor U11418 (N_11418,N_4291,N_7068);
xnor U11419 (N_11419,N_4832,N_5690);
or U11420 (N_11420,N_6931,N_6299);
nand U11421 (N_11421,N_6082,N_6975);
and U11422 (N_11422,N_4906,N_7410);
and U11423 (N_11423,N_4138,N_6363);
or U11424 (N_11424,N_7814,N_4010);
and U11425 (N_11425,N_7641,N_7674);
nor U11426 (N_11426,N_7079,N_5708);
nor U11427 (N_11427,N_6867,N_4928);
or U11428 (N_11428,N_7366,N_6494);
or U11429 (N_11429,N_7954,N_5919);
nor U11430 (N_11430,N_4340,N_6780);
or U11431 (N_11431,N_7262,N_4109);
nand U11432 (N_11432,N_7379,N_4958);
nor U11433 (N_11433,N_7082,N_6454);
and U11434 (N_11434,N_4080,N_4302);
nor U11435 (N_11435,N_4914,N_4253);
nand U11436 (N_11436,N_7767,N_7319);
nor U11437 (N_11437,N_6827,N_5347);
or U11438 (N_11438,N_7380,N_6550);
or U11439 (N_11439,N_6384,N_7027);
xnor U11440 (N_11440,N_6811,N_4147);
nor U11441 (N_11441,N_4598,N_7652);
and U11442 (N_11442,N_7988,N_4705);
nand U11443 (N_11443,N_6224,N_4120);
nor U11444 (N_11444,N_5466,N_4873);
nor U11445 (N_11445,N_4671,N_6326);
nor U11446 (N_11446,N_5974,N_5036);
or U11447 (N_11447,N_4049,N_5351);
and U11448 (N_11448,N_4633,N_5135);
or U11449 (N_11449,N_7664,N_5912);
nor U11450 (N_11450,N_7819,N_5783);
or U11451 (N_11451,N_4581,N_4593);
xnor U11452 (N_11452,N_5299,N_4484);
and U11453 (N_11453,N_4762,N_4826);
nor U11454 (N_11454,N_4338,N_7712);
xnor U11455 (N_11455,N_4402,N_6752);
nand U11456 (N_11456,N_6910,N_4914);
nand U11457 (N_11457,N_5999,N_4220);
nor U11458 (N_11458,N_4512,N_7236);
nor U11459 (N_11459,N_6379,N_6610);
xor U11460 (N_11460,N_4100,N_5407);
and U11461 (N_11461,N_4850,N_5610);
or U11462 (N_11462,N_5423,N_6440);
nor U11463 (N_11463,N_4425,N_7302);
nand U11464 (N_11464,N_5871,N_7458);
and U11465 (N_11465,N_5360,N_5953);
or U11466 (N_11466,N_6802,N_6128);
nand U11467 (N_11467,N_5266,N_7422);
nand U11468 (N_11468,N_6161,N_6475);
nand U11469 (N_11469,N_7529,N_7502);
and U11470 (N_11470,N_6977,N_4663);
or U11471 (N_11471,N_7312,N_4684);
nor U11472 (N_11472,N_5719,N_5399);
nand U11473 (N_11473,N_6578,N_4639);
and U11474 (N_11474,N_6890,N_5064);
or U11475 (N_11475,N_7659,N_4169);
xnor U11476 (N_11476,N_4300,N_5800);
and U11477 (N_11477,N_4655,N_4716);
and U11478 (N_11478,N_5157,N_7204);
or U11479 (N_11479,N_4565,N_6186);
nand U11480 (N_11480,N_6384,N_6984);
nor U11481 (N_11481,N_5318,N_5019);
or U11482 (N_11482,N_6958,N_5833);
or U11483 (N_11483,N_4334,N_4728);
nor U11484 (N_11484,N_5306,N_5047);
and U11485 (N_11485,N_7164,N_5618);
or U11486 (N_11486,N_6393,N_4797);
nor U11487 (N_11487,N_5722,N_7315);
nor U11488 (N_11488,N_6007,N_5587);
xnor U11489 (N_11489,N_6078,N_4534);
nor U11490 (N_11490,N_6806,N_6650);
nand U11491 (N_11491,N_5830,N_6727);
nand U11492 (N_11492,N_5271,N_5046);
and U11493 (N_11493,N_6965,N_5550);
nand U11494 (N_11494,N_6633,N_4462);
or U11495 (N_11495,N_6536,N_6964);
or U11496 (N_11496,N_5988,N_4304);
or U11497 (N_11497,N_6918,N_6481);
or U11498 (N_11498,N_5832,N_6982);
and U11499 (N_11499,N_4432,N_7627);
or U11500 (N_11500,N_7568,N_6082);
or U11501 (N_11501,N_5649,N_6104);
and U11502 (N_11502,N_6748,N_6501);
nor U11503 (N_11503,N_6944,N_7967);
xor U11504 (N_11504,N_5957,N_6557);
nand U11505 (N_11505,N_7452,N_5193);
nor U11506 (N_11506,N_4095,N_5662);
nand U11507 (N_11507,N_6565,N_6877);
nor U11508 (N_11508,N_7620,N_7142);
nand U11509 (N_11509,N_5734,N_6422);
or U11510 (N_11510,N_7838,N_6284);
nand U11511 (N_11511,N_6828,N_6111);
or U11512 (N_11512,N_4446,N_5782);
nand U11513 (N_11513,N_7874,N_5419);
and U11514 (N_11514,N_5326,N_7666);
nand U11515 (N_11515,N_4041,N_5044);
nand U11516 (N_11516,N_5181,N_5108);
nor U11517 (N_11517,N_4404,N_5782);
and U11518 (N_11518,N_5973,N_4386);
or U11519 (N_11519,N_6284,N_7289);
nand U11520 (N_11520,N_6282,N_6150);
or U11521 (N_11521,N_5412,N_6760);
and U11522 (N_11522,N_4660,N_7532);
and U11523 (N_11523,N_4798,N_4022);
nand U11524 (N_11524,N_5405,N_5145);
nor U11525 (N_11525,N_6593,N_6552);
nor U11526 (N_11526,N_7704,N_6963);
and U11527 (N_11527,N_5413,N_4881);
and U11528 (N_11528,N_5925,N_4967);
nor U11529 (N_11529,N_4188,N_5579);
or U11530 (N_11530,N_5727,N_5386);
nor U11531 (N_11531,N_6989,N_5318);
or U11532 (N_11532,N_5882,N_6967);
nand U11533 (N_11533,N_4276,N_4299);
and U11534 (N_11534,N_7482,N_5734);
or U11535 (N_11535,N_4698,N_5693);
xnor U11536 (N_11536,N_6479,N_5137);
or U11537 (N_11537,N_4744,N_6283);
nand U11538 (N_11538,N_5224,N_7919);
and U11539 (N_11539,N_6826,N_4651);
and U11540 (N_11540,N_5832,N_7593);
or U11541 (N_11541,N_5528,N_6767);
and U11542 (N_11542,N_5957,N_6088);
or U11543 (N_11543,N_6106,N_4083);
nand U11544 (N_11544,N_4982,N_5544);
nand U11545 (N_11545,N_6617,N_4600);
nand U11546 (N_11546,N_7311,N_4186);
nor U11547 (N_11547,N_6990,N_5665);
nor U11548 (N_11548,N_7932,N_7538);
or U11549 (N_11549,N_5665,N_4433);
and U11550 (N_11550,N_6347,N_5087);
nand U11551 (N_11551,N_7962,N_7102);
or U11552 (N_11552,N_6873,N_6373);
and U11553 (N_11553,N_4025,N_6589);
or U11554 (N_11554,N_4170,N_5747);
or U11555 (N_11555,N_6677,N_7113);
or U11556 (N_11556,N_5601,N_5252);
nand U11557 (N_11557,N_6592,N_4770);
nor U11558 (N_11558,N_6146,N_5007);
xnor U11559 (N_11559,N_6353,N_4382);
nor U11560 (N_11560,N_7985,N_5323);
nor U11561 (N_11561,N_6547,N_5018);
xor U11562 (N_11562,N_7920,N_7021);
nor U11563 (N_11563,N_6201,N_5245);
nand U11564 (N_11564,N_6897,N_5756);
or U11565 (N_11565,N_4518,N_7201);
or U11566 (N_11566,N_5069,N_7627);
or U11567 (N_11567,N_7432,N_6425);
and U11568 (N_11568,N_7249,N_5370);
nor U11569 (N_11569,N_4862,N_4420);
nor U11570 (N_11570,N_4335,N_5761);
nand U11571 (N_11571,N_7111,N_4874);
or U11572 (N_11572,N_6735,N_7480);
xor U11573 (N_11573,N_6144,N_5621);
and U11574 (N_11574,N_6808,N_4443);
and U11575 (N_11575,N_5379,N_5137);
nand U11576 (N_11576,N_5256,N_5653);
and U11577 (N_11577,N_5818,N_6578);
nor U11578 (N_11578,N_5153,N_6407);
or U11579 (N_11579,N_4596,N_6608);
nor U11580 (N_11580,N_6364,N_5670);
nand U11581 (N_11581,N_7024,N_5096);
nor U11582 (N_11582,N_6744,N_6278);
and U11583 (N_11583,N_4147,N_6645);
xor U11584 (N_11584,N_5586,N_7510);
nand U11585 (N_11585,N_7654,N_5675);
and U11586 (N_11586,N_7236,N_7241);
or U11587 (N_11587,N_7318,N_5579);
nor U11588 (N_11588,N_6207,N_7123);
and U11589 (N_11589,N_6836,N_4602);
and U11590 (N_11590,N_5265,N_4878);
nor U11591 (N_11591,N_7536,N_4523);
nor U11592 (N_11592,N_4672,N_6526);
nand U11593 (N_11593,N_6994,N_5179);
nand U11594 (N_11594,N_6858,N_6004);
nor U11595 (N_11595,N_4768,N_4034);
nor U11596 (N_11596,N_4005,N_7747);
and U11597 (N_11597,N_5448,N_4224);
and U11598 (N_11598,N_6563,N_4140);
nor U11599 (N_11599,N_5347,N_6812);
xnor U11600 (N_11600,N_5017,N_7793);
nor U11601 (N_11601,N_7703,N_4873);
nand U11602 (N_11602,N_6865,N_5268);
nor U11603 (N_11603,N_5632,N_6561);
or U11604 (N_11604,N_5578,N_7057);
nand U11605 (N_11605,N_6716,N_4471);
and U11606 (N_11606,N_7043,N_7105);
nand U11607 (N_11607,N_4334,N_6213);
and U11608 (N_11608,N_6072,N_7349);
nand U11609 (N_11609,N_6344,N_4875);
nand U11610 (N_11610,N_5976,N_5772);
nor U11611 (N_11611,N_7078,N_6475);
nand U11612 (N_11612,N_6614,N_6309);
nand U11613 (N_11613,N_6946,N_6504);
and U11614 (N_11614,N_7979,N_6117);
or U11615 (N_11615,N_6190,N_6489);
nand U11616 (N_11616,N_7767,N_5204);
xor U11617 (N_11617,N_4591,N_7822);
nor U11618 (N_11618,N_5257,N_4630);
xnor U11619 (N_11619,N_6593,N_5869);
nand U11620 (N_11620,N_5799,N_4414);
nor U11621 (N_11621,N_5571,N_7645);
nand U11622 (N_11622,N_4897,N_6171);
nand U11623 (N_11623,N_7311,N_4559);
or U11624 (N_11624,N_7925,N_5548);
or U11625 (N_11625,N_4422,N_7934);
and U11626 (N_11626,N_6996,N_6222);
nor U11627 (N_11627,N_7054,N_7002);
and U11628 (N_11628,N_7731,N_5778);
xor U11629 (N_11629,N_6309,N_4608);
and U11630 (N_11630,N_5557,N_5941);
xnor U11631 (N_11631,N_6560,N_4457);
and U11632 (N_11632,N_5091,N_6521);
nor U11633 (N_11633,N_6437,N_5680);
nor U11634 (N_11634,N_4715,N_6135);
nor U11635 (N_11635,N_5526,N_6136);
and U11636 (N_11636,N_6125,N_5406);
nor U11637 (N_11637,N_6249,N_4693);
nor U11638 (N_11638,N_5131,N_5210);
nor U11639 (N_11639,N_4248,N_5171);
nand U11640 (N_11640,N_4747,N_6291);
or U11641 (N_11641,N_6248,N_7560);
nand U11642 (N_11642,N_6332,N_4055);
and U11643 (N_11643,N_7534,N_6320);
and U11644 (N_11644,N_4946,N_6117);
nor U11645 (N_11645,N_6169,N_6569);
or U11646 (N_11646,N_5136,N_6424);
nor U11647 (N_11647,N_5576,N_4945);
nor U11648 (N_11648,N_4723,N_5068);
nand U11649 (N_11649,N_6906,N_7069);
and U11650 (N_11650,N_6438,N_5860);
nand U11651 (N_11651,N_6245,N_7863);
nor U11652 (N_11652,N_6857,N_6027);
and U11653 (N_11653,N_4182,N_6212);
or U11654 (N_11654,N_5283,N_7465);
nand U11655 (N_11655,N_7239,N_5203);
nand U11656 (N_11656,N_6239,N_4916);
or U11657 (N_11657,N_7357,N_5011);
nand U11658 (N_11658,N_7830,N_5377);
nor U11659 (N_11659,N_6629,N_5387);
and U11660 (N_11660,N_7676,N_6614);
and U11661 (N_11661,N_5487,N_6261);
xor U11662 (N_11662,N_5874,N_4088);
or U11663 (N_11663,N_7759,N_6179);
nand U11664 (N_11664,N_6281,N_4092);
and U11665 (N_11665,N_7708,N_7799);
nand U11666 (N_11666,N_7983,N_6692);
xor U11667 (N_11667,N_6091,N_4767);
nor U11668 (N_11668,N_5027,N_5449);
and U11669 (N_11669,N_5210,N_6088);
and U11670 (N_11670,N_7747,N_5535);
nand U11671 (N_11671,N_7080,N_4825);
nor U11672 (N_11672,N_7893,N_6581);
nor U11673 (N_11673,N_6255,N_6534);
nor U11674 (N_11674,N_4961,N_6976);
or U11675 (N_11675,N_4530,N_4494);
xnor U11676 (N_11676,N_5887,N_5640);
nand U11677 (N_11677,N_4005,N_4426);
xor U11678 (N_11678,N_5060,N_4161);
xor U11679 (N_11679,N_5758,N_4918);
and U11680 (N_11680,N_7786,N_6010);
nand U11681 (N_11681,N_5831,N_5513);
nor U11682 (N_11682,N_4170,N_4132);
nor U11683 (N_11683,N_4010,N_7639);
nand U11684 (N_11684,N_4260,N_7793);
and U11685 (N_11685,N_5423,N_4374);
nor U11686 (N_11686,N_6027,N_5876);
nand U11687 (N_11687,N_6554,N_5963);
xnor U11688 (N_11688,N_5142,N_4209);
nand U11689 (N_11689,N_5051,N_7078);
nor U11690 (N_11690,N_5012,N_7356);
or U11691 (N_11691,N_6116,N_7194);
nor U11692 (N_11692,N_4312,N_4067);
nand U11693 (N_11693,N_6228,N_4645);
xor U11694 (N_11694,N_6971,N_5709);
xnor U11695 (N_11695,N_6652,N_7050);
nand U11696 (N_11696,N_6281,N_7151);
and U11697 (N_11697,N_4864,N_5589);
or U11698 (N_11698,N_4848,N_5518);
nor U11699 (N_11699,N_4041,N_4326);
xnor U11700 (N_11700,N_6438,N_7668);
nand U11701 (N_11701,N_5722,N_5397);
nor U11702 (N_11702,N_7021,N_4227);
or U11703 (N_11703,N_4312,N_5228);
or U11704 (N_11704,N_7589,N_6911);
nor U11705 (N_11705,N_5306,N_4435);
nand U11706 (N_11706,N_4703,N_6732);
and U11707 (N_11707,N_6402,N_7458);
nor U11708 (N_11708,N_5644,N_7838);
and U11709 (N_11709,N_4605,N_6392);
nor U11710 (N_11710,N_5341,N_7505);
nand U11711 (N_11711,N_4393,N_4165);
xnor U11712 (N_11712,N_4679,N_4170);
or U11713 (N_11713,N_7695,N_5904);
nand U11714 (N_11714,N_5986,N_6650);
or U11715 (N_11715,N_4306,N_6171);
nand U11716 (N_11716,N_4609,N_7690);
nand U11717 (N_11717,N_4388,N_7736);
xor U11718 (N_11718,N_6994,N_6628);
nand U11719 (N_11719,N_7099,N_7415);
nor U11720 (N_11720,N_7502,N_4029);
xor U11721 (N_11721,N_6155,N_4925);
or U11722 (N_11722,N_4555,N_5019);
or U11723 (N_11723,N_7581,N_5345);
and U11724 (N_11724,N_6825,N_7675);
nand U11725 (N_11725,N_7165,N_7229);
or U11726 (N_11726,N_7407,N_4735);
nor U11727 (N_11727,N_4751,N_6836);
nor U11728 (N_11728,N_6957,N_7586);
nor U11729 (N_11729,N_6006,N_7157);
nand U11730 (N_11730,N_5428,N_6483);
and U11731 (N_11731,N_4942,N_4099);
or U11732 (N_11732,N_7481,N_4408);
xor U11733 (N_11733,N_6967,N_7739);
xor U11734 (N_11734,N_7464,N_5543);
nand U11735 (N_11735,N_5597,N_7073);
or U11736 (N_11736,N_5983,N_7619);
nand U11737 (N_11737,N_4343,N_6119);
xnor U11738 (N_11738,N_7183,N_6615);
nand U11739 (N_11739,N_4461,N_7729);
or U11740 (N_11740,N_4360,N_6625);
and U11741 (N_11741,N_7394,N_4226);
nand U11742 (N_11742,N_7604,N_7219);
nand U11743 (N_11743,N_5980,N_5137);
or U11744 (N_11744,N_6875,N_7766);
and U11745 (N_11745,N_6668,N_6527);
xor U11746 (N_11746,N_6395,N_6288);
nor U11747 (N_11747,N_5193,N_4754);
xnor U11748 (N_11748,N_7434,N_5185);
nor U11749 (N_11749,N_6866,N_6980);
and U11750 (N_11750,N_6918,N_7910);
or U11751 (N_11751,N_4164,N_6427);
and U11752 (N_11752,N_5935,N_6529);
nor U11753 (N_11753,N_7770,N_6002);
and U11754 (N_11754,N_7948,N_7133);
nor U11755 (N_11755,N_5301,N_4416);
nand U11756 (N_11756,N_7586,N_6264);
nand U11757 (N_11757,N_7542,N_6476);
or U11758 (N_11758,N_7646,N_6129);
nor U11759 (N_11759,N_7478,N_4916);
or U11760 (N_11760,N_5841,N_5585);
and U11761 (N_11761,N_4309,N_5450);
nor U11762 (N_11762,N_4682,N_4979);
nor U11763 (N_11763,N_6040,N_7656);
nor U11764 (N_11764,N_4983,N_5927);
or U11765 (N_11765,N_6811,N_5281);
nor U11766 (N_11766,N_4345,N_4499);
or U11767 (N_11767,N_7761,N_4956);
and U11768 (N_11768,N_4892,N_7181);
and U11769 (N_11769,N_5717,N_7383);
and U11770 (N_11770,N_7082,N_4608);
or U11771 (N_11771,N_4096,N_5643);
or U11772 (N_11772,N_5088,N_7017);
and U11773 (N_11773,N_4091,N_7576);
nor U11774 (N_11774,N_5140,N_7200);
nor U11775 (N_11775,N_4729,N_4348);
and U11776 (N_11776,N_7506,N_5553);
nor U11777 (N_11777,N_7975,N_4859);
nor U11778 (N_11778,N_5011,N_4088);
and U11779 (N_11779,N_7245,N_6698);
nand U11780 (N_11780,N_5758,N_4778);
nand U11781 (N_11781,N_6686,N_4269);
and U11782 (N_11782,N_4677,N_4963);
nor U11783 (N_11783,N_6247,N_5095);
xor U11784 (N_11784,N_6223,N_7189);
nand U11785 (N_11785,N_7253,N_4509);
nand U11786 (N_11786,N_5280,N_7477);
and U11787 (N_11787,N_4165,N_7200);
and U11788 (N_11788,N_6221,N_5339);
nand U11789 (N_11789,N_4575,N_7466);
and U11790 (N_11790,N_6567,N_6120);
or U11791 (N_11791,N_6788,N_5023);
nor U11792 (N_11792,N_6488,N_4560);
nand U11793 (N_11793,N_6008,N_5664);
nand U11794 (N_11794,N_5484,N_7152);
nand U11795 (N_11795,N_6462,N_6597);
or U11796 (N_11796,N_6991,N_7761);
nor U11797 (N_11797,N_4317,N_5547);
xnor U11798 (N_11798,N_4993,N_7183);
nor U11799 (N_11799,N_7495,N_7378);
or U11800 (N_11800,N_7001,N_7195);
and U11801 (N_11801,N_4991,N_4511);
or U11802 (N_11802,N_6948,N_4956);
or U11803 (N_11803,N_7462,N_7836);
nor U11804 (N_11804,N_5249,N_7401);
xnor U11805 (N_11805,N_4844,N_6728);
nor U11806 (N_11806,N_5951,N_7134);
nor U11807 (N_11807,N_7659,N_7028);
nand U11808 (N_11808,N_4723,N_7607);
nand U11809 (N_11809,N_4262,N_4525);
nand U11810 (N_11810,N_6999,N_4586);
nand U11811 (N_11811,N_4188,N_4494);
nor U11812 (N_11812,N_7827,N_5215);
nor U11813 (N_11813,N_7699,N_6915);
and U11814 (N_11814,N_4524,N_6589);
nand U11815 (N_11815,N_6178,N_7853);
and U11816 (N_11816,N_4529,N_7344);
and U11817 (N_11817,N_4034,N_6817);
or U11818 (N_11818,N_7540,N_4073);
nor U11819 (N_11819,N_5673,N_5569);
nor U11820 (N_11820,N_6944,N_6108);
and U11821 (N_11821,N_5738,N_5287);
nor U11822 (N_11822,N_5510,N_7517);
nand U11823 (N_11823,N_6106,N_7269);
and U11824 (N_11824,N_5680,N_7126);
nand U11825 (N_11825,N_5052,N_7441);
and U11826 (N_11826,N_5420,N_5424);
nor U11827 (N_11827,N_6411,N_4282);
and U11828 (N_11828,N_7223,N_7408);
nand U11829 (N_11829,N_4836,N_4421);
nand U11830 (N_11830,N_6556,N_6815);
nor U11831 (N_11831,N_7361,N_4575);
nor U11832 (N_11832,N_7441,N_6061);
xnor U11833 (N_11833,N_4678,N_4656);
or U11834 (N_11834,N_4218,N_4128);
or U11835 (N_11835,N_4461,N_7024);
nand U11836 (N_11836,N_4848,N_7043);
nand U11837 (N_11837,N_5521,N_4235);
nor U11838 (N_11838,N_5067,N_5705);
nor U11839 (N_11839,N_7061,N_6159);
nand U11840 (N_11840,N_7108,N_5147);
xnor U11841 (N_11841,N_5425,N_4592);
or U11842 (N_11842,N_5415,N_5351);
nor U11843 (N_11843,N_7748,N_6380);
nand U11844 (N_11844,N_6975,N_6815);
nand U11845 (N_11845,N_5497,N_5891);
and U11846 (N_11846,N_6510,N_6919);
and U11847 (N_11847,N_4240,N_7725);
nand U11848 (N_11848,N_5199,N_6127);
nand U11849 (N_11849,N_4406,N_5149);
or U11850 (N_11850,N_7587,N_7250);
and U11851 (N_11851,N_4930,N_5492);
nand U11852 (N_11852,N_5764,N_4375);
nand U11853 (N_11853,N_7752,N_6925);
nand U11854 (N_11854,N_5172,N_4576);
nand U11855 (N_11855,N_6730,N_4538);
nand U11856 (N_11856,N_6535,N_4151);
and U11857 (N_11857,N_5671,N_6104);
or U11858 (N_11858,N_4877,N_6079);
and U11859 (N_11859,N_5725,N_6016);
nor U11860 (N_11860,N_4831,N_5140);
or U11861 (N_11861,N_5826,N_6781);
or U11862 (N_11862,N_6105,N_6539);
nor U11863 (N_11863,N_6965,N_5460);
and U11864 (N_11864,N_5796,N_5501);
nor U11865 (N_11865,N_7079,N_7217);
and U11866 (N_11866,N_5668,N_4740);
and U11867 (N_11867,N_6035,N_4290);
and U11868 (N_11868,N_4325,N_4732);
or U11869 (N_11869,N_6935,N_5724);
nor U11870 (N_11870,N_5307,N_7936);
nand U11871 (N_11871,N_4960,N_4854);
and U11872 (N_11872,N_7539,N_4098);
nand U11873 (N_11873,N_7963,N_4070);
and U11874 (N_11874,N_4122,N_7863);
and U11875 (N_11875,N_5409,N_5865);
and U11876 (N_11876,N_4414,N_7326);
nand U11877 (N_11877,N_5659,N_4399);
nor U11878 (N_11878,N_6681,N_6934);
xnor U11879 (N_11879,N_6198,N_7908);
nor U11880 (N_11880,N_5607,N_6104);
nor U11881 (N_11881,N_5425,N_6711);
or U11882 (N_11882,N_5863,N_5120);
or U11883 (N_11883,N_6229,N_5263);
or U11884 (N_11884,N_4731,N_6003);
nor U11885 (N_11885,N_4821,N_6046);
and U11886 (N_11886,N_6401,N_4377);
or U11887 (N_11887,N_7564,N_7499);
nor U11888 (N_11888,N_5363,N_5543);
or U11889 (N_11889,N_6351,N_4720);
nand U11890 (N_11890,N_5692,N_4337);
or U11891 (N_11891,N_7057,N_5194);
nand U11892 (N_11892,N_7317,N_4624);
nor U11893 (N_11893,N_6746,N_4203);
nor U11894 (N_11894,N_4755,N_6192);
or U11895 (N_11895,N_5771,N_4182);
nand U11896 (N_11896,N_5886,N_6604);
and U11897 (N_11897,N_6287,N_6020);
or U11898 (N_11898,N_6457,N_6982);
nand U11899 (N_11899,N_4297,N_5719);
nor U11900 (N_11900,N_4786,N_6438);
nand U11901 (N_11901,N_7280,N_4751);
xor U11902 (N_11902,N_6529,N_4086);
or U11903 (N_11903,N_4479,N_6091);
nand U11904 (N_11904,N_7010,N_5871);
and U11905 (N_11905,N_6741,N_5993);
and U11906 (N_11906,N_6808,N_4038);
nand U11907 (N_11907,N_5577,N_6691);
xnor U11908 (N_11908,N_5710,N_6109);
xnor U11909 (N_11909,N_5699,N_6881);
or U11910 (N_11910,N_6049,N_6084);
or U11911 (N_11911,N_5257,N_4749);
xnor U11912 (N_11912,N_5605,N_4009);
xnor U11913 (N_11913,N_7226,N_5245);
nor U11914 (N_11914,N_4068,N_4870);
or U11915 (N_11915,N_5921,N_6559);
or U11916 (N_11916,N_4749,N_6793);
nand U11917 (N_11917,N_6896,N_7573);
or U11918 (N_11918,N_5099,N_6012);
and U11919 (N_11919,N_4367,N_5829);
nor U11920 (N_11920,N_4367,N_4252);
and U11921 (N_11921,N_4703,N_6667);
and U11922 (N_11922,N_6135,N_6638);
nand U11923 (N_11923,N_7808,N_7331);
and U11924 (N_11924,N_6245,N_7200);
or U11925 (N_11925,N_7389,N_5210);
nand U11926 (N_11926,N_6879,N_7899);
and U11927 (N_11927,N_5364,N_4143);
nor U11928 (N_11928,N_6855,N_5429);
xor U11929 (N_11929,N_6179,N_5834);
nand U11930 (N_11930,N_5976,N_4661);
or U11931 (N_11931,N_5302,N_6424);
or U11932 (N_11932,N_7763,N_5981);
nand U11933 (N_11933,N_6015,N_4460);
nor U11934 (N_11934,N_4835,N_7064);
or U11935 (N_11935,N_7934,N_7476);
nand U11936 (N_11936,N_7205,N_5027);
or U11937 (N_11937,N_5368,N_7721);
nand U11938 (N_11938,N_7769,N_4982);
xor U11939 (N_11939,N_5281,N_7334);
or U11940 (N_11940,N_5778,N_6494);
nor U11941 (N_11941,N_4219,N_4415);
nand U11942 (N_11942,N_6171,N_5044);
xnor U11943 (N_11943,N_6330,N_7531);
and U11944 (N_11944,N_5744,N_4552);
nand U11945 (N_11945,N_5104,N_6434);
nor U11946 (N_11946,N_6110,N_4397);
xnor U11947 (N_11947,N_4700,N_7117);
nand U11948 (N_11948,N_4407,N_5761);
nor U11949 (N_11949,N_7064,N_6700);
nor U11950 (N_11950,N_6568,N_7638);
nor U11951 (N_11951,N_7357,N_6492);
and U11952 (N_11952,N_5526,N_6601);
nor U11953 (N_11953,N_7943,N_5957);
or U11954 (N_11954,N_4663,N_5979);
or U11955 (N_11955,N_4856,N_6538);
nor U11956 (N_11956,N_5142,N_5397);
or U11957 (N_11957,N_7876,N_6628);
nand U11958 (N_11958,N_5574,N_7210);
and U11959 (N_11959,N_4378,N_6532);
nand U11960 (N_11960,N_7991,N_7039);
or U11961 (N_11961,N_6913,N_4366);
nand U11962 (N_11962,N_7838,N_6396);
nand U11963 (N_11963,N_5886,N_5692);
nand U11964 (N_11964,N_6584,N_6083);
xor U11965 (N_11965,N_7592,N_6995);
nand U11966 (N_11966,N_4719,N_6851);
or U11967 (N_11967,N_4538,N_5751);
nor U11968 (N_11968,N_5733,N_6025);
nor U11969 (N_11969,N_4019,N_4526);
nor U11970 (N_11970,N_5681,N_5893);
and U11971 (N_11971,N_5693,N_4218);
nor U11972 (N_11972,N_5341,N_6476);
or U11973 (N_11973,N_4078,N_5724);
and U11974 (N_11974,N_5637,N_4122);
nand U11975 (N_11975,N_4205,N_6146);
or U11976 (N_11976,N_5562,N_5399);
nor U11977 (N_11977,N_5300,N_4043);
and U11978 (N_11978,N_6919,N_5875);
nor U11979 (N_11979,N_4644,N_4284);
or U11980 (N_11980,N_7207,N_4113);
xnor U11981 (N_11981,N_4375,N_7854);
nor U11982 (N_11982,N_4761,N_4027);
or U11983 (N_11983,N_7665,N_6322);
xnor U11984 (N_11984,N_4990,N_4460);
nand U11985 (N_11985,N_5657,N_4488);
nand U11986 (N_11986,N_5394,N_5641);
and U11987 (N_11987,N_6589,N_4427);
xnor U11988 (N_11988,N_6536,N_4431);
nand U11989 (N_11989,N_7319,N_7408);
nand U11990 (N_11990,N_5750,N_5372);
or U11991 (N_11991,N_6963,N_4237);
or U11992 (N_11992,N_7263,N_5709);
and U11993 (N_11993,N_6894,N_4834);
nor U11994 (N_11994,N_5273,N_5313);
nor U11995 (N_11995,N_6344,N_4152);
nor U11996 (N_11996,N_7317,N_4505);
nor U11997 (N_11997,N_4879,N_5837);
or U11998 (N_11998,N_4786,N_5387);
nand U11999 (N_11999,N_5911,N_4091);
nor U12000 (N_12000,N_8562,N_10428);
nand U12001 (N_12001,N_10839,N_11307);
and U12002 (N_12002,N_11302,N_11898);
nand U12003 (N_12003,N_8383,N_11842);
nor U12004 (N_12004,N_9547,N_8175);
and U12005 (N_12005,N_11888,N_11615);
nor U12006 (N_12006,N_8049,N_8745);
nand U12007 (N_12007,N_8209,N_11289);
nor U12008 (N_12008,N_10323,N_11740);
and U12009 (N_12009,N_8493,N_8803);
and U12010 (N_12010,N_8067,N_10707);
or U12011 (N_12011,N_8083,N_9945);
or U12012 (N_12012,N_10715,N_9364);
nor U12013 (N_12013,N_8201,N_8916);
and U12014 (N_12014,N_9005,N_9567);
and U12015 (N_12015,N_8579,N_9085);
xor U12016 (N_12016,N_11745,N_8038);
nor U12017 (N_12017,N_8110,N_10612);
or U12018 (N_12018,N_11677,N_8690);
nor U12019 (N_12019,N_11896,N_8819);
and U12020 (N_12020,N_8400,N_11381);
or U12021 (N_12021,N_8364,N_9862);
and U12022 (N_12022,N_8739,N_9358);
or U12023 (N_12023,N_11702,N_11216);
nor U12024 (N_12024,N_11061,N_11553);
or U12025 (N_12025,N_9150,N_8806);
nor U12026 (N_12026,N_8511,N_11574);
and U12027 (N_12027,N_11732,N_9522);
nor U12028 (N_12028,N_9981,N_8069);
and U12029 (N_12029,N_9561,N_11090);
or U12030 (N_12030,N_10792,N_11194);
nand U12031 (N_12031,N_10892,N_11271);
nand U12032 (N_12032,N_10972,N_10821);
nor U12033 (N_12033,N_10631,N_9394);
and U12034 (N_12034,N_8299,N_8642);
or U12035 (N_12035,N_9184,N_11037);
and U12036 (N_12036,N_9823,N_10077);
nand U12037 (N_12037,N_8312,N_8677);
nand U12038 (N_12038,N_8661,N_11407);
and U12039 (N_12039,N_9069,N_8646);
xnor U12040 (N_12040,N_10220,N_8024);
nor U12041 (N_12041,N_10257,N_9391);
nor U12042 (N_12042,N_10653,N_10749);
nand U12043 (N_12043,N_10879,N_10360);
or U12044 (N_12044,N_8010,N_10615);
and U12045 (N_12045,N_11914,N_8102);
or U12046 (N_12046,N_8007,N_11817);
or U12047 (N_12047,N_10090,N_10194);
nor U12048 (N_12048,N_10663,N_11211);
and U12049 (N_12049,N_9172,N_9185);
nand U12050 (N_12050,N_9271,N_10589);
or U12051 (N_12051,N_8023,N_11601);
or U12052 (N_12052,N_11573,N_11365);
or U12053 (N_12053,N_10001,N_10730);
nand U12054 (N_12054,N_8870,N_9385);
or U12055 (N_12055,N_10989,N_11959);
nor U12056 (N_12056,N_10401,N_9625);
nand U12057 (N_12057,N_10162,N_10561);
and U12058 (N_12058,N_10945,N_11242);
and U12059 (N_12059,N_9837,N_9633);
nand U12060 (N_12060,N_11921,N_9768);
or U12061 (N_12061,N_11186,N_9867);
or U12062 (N_12062,N_10777,N_11619);
or U12063 (N_12063,N_10270,N_10207);
nor U12064 (N_12064,N_10051,N_9194);
nand U12065 (N_12065,N_8073,N_8292);
and U12066 (N_12066,N_8471,N_9556);
or U12067 (N_12067,N_10539,N_8785);
nand U12068 (N_12068,N_11255,N_11383);
and U12069 (N_12069,N_9995,N_11296);
nor U12070 (N_12070,N_10126,N_9550);
and U12071 (N_12071,N_9415,N_10294);
and U12072 (N_12072,N_9666,N_10487);
xnor U12073 (N_12073,N_11934,N_9896);
nand U12074 (N_12074,N_9767,N_10180);
nor U12075 (N_12075,N_8713,N_10837);
and U12076 (N_12076,N_10074,N_8191);
xnor U12077 (N_12077,N_10130,N_8875);
or U12078 (N_12078,N_8027,N_9379);
xnor U12079 (N_12079,N_9505,N_8627);
or U12080 (N_12080,N_10228,N_11026);
xnor U12081 (N_12081,N_9730,N_11418);
and U12082 (N_12082,N_11179,N_9694);
xor U12083 (N_12083,N_9738,N_10702);
nor U12084 (N_12084,N_9611,N_9652);
xnor U12085 (N_12085,N_10720,N_10629);
xor U12086 (N_12086,N_8135,N_9779);
nand U12087 (N_12087,N_9451,N_10622);
xnor U12088 (N_12088,N_11110,N_8938);
nor U12089 (N_12089,N_9475,N_10408);
or U12090 (N_12090,N_8177,N_11968);
nor U12091 (N_12091,N_10606,N_8587);
nand U12092 (N_12092,N_10928,N_10475);
nand U12093 (N_12093,N_10915,N_8626);
and U12094 (N_12094,N_10661,N_9487);
and U12095 (N_12095,N_9039,N_10826);
or U12096 (N_12096,N_8431,N_11457);
or U12097 (N_12097,N_11355,N_10829);
nor U12098 (N_12098,N_11164,N_11741);
and U12099 (N_12099,N_8176,N_10277);
and U12100 (N_12100,N_9283,N_9885);
nor U12101 (N_12101,N_9196,N_8322);
nor U12102 (N_12102,N_10003,N_11710);
nand U12103 (N_12103,N_9711,N_10882);
and U12104 (N_12104,N_11685,N_10050);
or U12105 (N_12105,N_9168,N_10183);
nand U12106 (N_12106,N_8995,N_8205);
nor U12107 (N_12107,N_8347,N_8898);
or U12108 (N_12108,N_11718,N_11534);
nor U12109 (N_12109,N_10350,N_10549);
nand U12110 (N_12110,N_8470,N_8267);
and U12111 (N_12111,N_8143,N_10040);
nand U12112 (N_12112,N_11071,N_11017);
or U12113 (N_12113,N_8638,N_9020);
nand U12114 (N_12114,N_11929,N_10271);
nand U12115 (N_12115,N_10044,N_10933);
nor U12116 (N_12116,N_9850,N_11637);
or U12117 (N_12117,N_8540,N_11562);
nor U12118 (N_12118,N_9372,N_9340);
nand U12119 (N_12119,N_11111,N_9077);
nor U12120 (N_12120,N_10054,N_8340);
nor U12121 (N_12121,N_8577,N_11473);
nand U12122 (N_12122,N_11297,N_10112);
nor U12123 (N_12123,N_9059,N_8265);
or U12124 (N_12124,N_9788,N_9965);
or U12125 (N_12125,N_11020,N_11221);
nor U12126 (N_12126,N_10801,N_10555);
and U12127 (N_12127,N_8260,N_9435);
and U12128 (N_12128,N_8419,N_10354);
nand U12129 (N_12129,N_10480,N_8127);
and U12130 (N_12130,N_8824,N_11235);
or U12131 (N_12131,N_8883,N_8769);
and U12132 (N_12132,N_8757,N_10802);
and U12133 (N_12133,N_10202,N_9319);
xor U12134 (N_12134,N_9784,N_9247);
and U12135 (N_12135,N_11832,N_9672);
nand U12136 (N_12136,N_10156,N_8122);
nand U12137 (N_12137,N_11756,N_9496);
or U12138 (N_12138,N_11963,N_10708);
or U12139 (N_12139,N_8932,N_10380);
nor U12140 (N_12140,N_10466,N_10049);
and U12141 (N_12141,N_11816,N_10227);
nor U12142 (N_12142,N_9881,N_9317);
nor U12143 (N_12143,N_10426,N_11635);
and U12144 (N_12144,N_10514,N_8277);
and U12145 (N_12145,N_11632,N_8963);
nand U12146 (N_12146,N_10157,N_9038);
nor U12147 (N_12147,N_9064,N_8245);
and U12148 (N_12148,N_9783,N_11316);
nand U12149 (N_12149,N_9448,N_11197);
or U12150 (N_12150,N_10823,N_8615);
or U12151 (N_12151,N_9124,N_10610);
nor U12152 (N_12152,N_8231,N_11147);
nor U12153 (N_12153,N_10682,N_11156);
or U12154 (N_12154,N_10951,N_11638);
or U12155 (N_12155,N_10969,N_9143);
xnor U12156 (N_12156,N_8278,N_11446);
xnor U12157 (N_12157,N_11341,N_10973);
and U12158 (N_12158,N_9275,N_10290);
and U12159 (N_12159,N_8141,N_10109);
and U12160 (N_12160,N_8228,N_9929);
nand U12161 (N_12161,N_9032,N_10313);
nor U12162 (N_12162,N_9417,N_11466);
nor U12163 (N_12163,N_9467,N_9597);
and U12164 (N_12164,N_8940,N_9442);
and U12165 (N_12165,N_11137,N_8915);
or U12166 (N_12166,N_10656,N_10816);
nand U12167 (N_12167,N_9203,N_8199);
and U12168 (N_12168,N_9015,N_10326);
or U12169 (N_12169,N_11516,N_11919);
and U12170 (N_12170,N_8149,N_8697);
nor U12171 (N_12171,N_8094,N_9100);
nor U12172 (N_12172,N_9764,N_10926);
nor U12173 (N_12173,N_8728,N_9957);
nand U12174 (N_12174,N_9277,N_9373);
nor U12175 (N_12175,N_10287,N_8391);
or U12176 (N_12176,N_11041,N_9637);
or U12177 (N_12177,N_8331,N_10192);
nand U12178 (N_12178,N_10073,N_10925);
nor U12179 (N_12179,N_10693,N_9424);
and U12180 (N_12180,N_9987,N_10120);
xor U12181 (N_12181,N_9648,N_9916);
xor U12182 (N_12182,N_11973,N_10931);
nand U12183 (N_12183,N_8050,N_11541);
and U12184 (N_12184,N_10255,N_8575);
nand U12185 (N_12185,N_11441,N_10734);
nand U12186 (N_12186,N_11392,N_9169);
nor U12187 (N_12187,N_9350,N_8976);
nand U12188 (N_12188,N_11445,N_11547);
or U12189 (N_12189,N_11577,N_11944);
or U12190 (N_12190,N_9618,N_8537);
nor U12191 (N_12191,N_11421,N_8968);
nor U12192 (N_12192,N_10543,N_10453);
and U12193 (N_12193,N_10784,N_8681);
or U12194 (N_12194,N_11317,N_9634);
nand U12195 (N_12195,N_9743,N_11356);
nor U12196 (N_12196,N_8287,N_11662);
nand U12197 (N_12197,N_10022,N_11904);
or U12198 (N_12198,N_9873,N_8145);
nor U12199 (N_12199,N_9289,N_8255);
and U12200 (N_12200,N_9800,N_9164);
nand U12201 (N_12201,N_8480,N_11335);
nand U12202 (N_12202,N_8783,N_11893);
or U12203 (N_12203,N_11546,N_9432);
nand U12204 (N_12204,N_8807,N_11395);
and U12205 (N_12205,N_8885,N_10031);
nand U12206 (N_12206,N_8780,N_10011);
or U12207 (N_12207,N_10813,N_8495);
and U12208 (N_12208,N_11862,N_9534);
or U12209 (N_12209,N_9182,N_8812);
nand U12210 (N_12210,N_10534,N_8192);
and U12211 (N_12211,N_10705,N_9986);
or U12212 (N_12212,N_9586,N_8773);
nand U12213 (N_12213,N_10714,N_9845);
and U12214 (N_12214,N_10504,N_8653);
nand U12215 (N_12215,N_11788,N_10143);
or U12216 (N_12216,N_8309,N_10358);
nand U12217 (N_12217,N_8483,N_8256);
nand U12218 (N_12218,N_8695,N_8658);
xor U12219 (N_12219,N_9132,N_10528);
nand U12220 (N_12220,N_8893,N_11412);
nand U12221 (N_12221,N_9230,N_11048);
nor U12222 (N_12222,N_9361,N_8125);
nand U12223 (N_12223,N_11823,N_10413);
and U12224 (N_12224,N_8925,N_8830);
xor U12225 (N_12225,N_9501,N_10761);
and U12226 (N_12226,N_10893,N_10794);
or U12227 (N_12227,N_11848,N_11592);
xor U12228 (N_12228,N_8270,N_11042);
and U12229 (N_12229,N_8148,N_11604);
and U12230 (N_12230,N_11537,N_8787);
and U12231 (N_12231,N_11782,N_8999);
nand U12232 (N_12232,N_8468,N_11985);
xnor U12233 (N_12233,N_11419,N_8107);
xor U12234 (N_12234,N_10121,N_10754);
or U12235 (N_12235,N_8252,N_11626);
nand U12236 (N_12236,N_11520,N_10852);
nor U12237 (N_12237,N_9994,N_10786);
or U12238 (N_12238,N_11792,N_8283);
nor U12239 (N_12239,N_11172,N_9426);
nand U12240 (N_12240,N_8703,N_8451);
nand U12241 (N_12241,N_8836,N_11285);
xor U12242 (N_12242,N_9693,N_11451);
or U12243 (N_12243,N_10075,N_11845);
nor U12244 (N_12244,N_10778,N_8159);
or U12245 (N_12245,N_10377,N_11915);
xnor U12246 (N_12246,N_9046,N_9927);
nor U12247 (N_12247,N_9389,N_9831);
nor U12248 (N_12248,N_11762,N_11748);
and U12249 (N_12249,N_9892,N_9944);
and U12250 (N_12250,N_8801,N_10519);
nand U12251 (N_12251,N_10958,N_11545);
xnor U12252 (N_12252,N_10787,N_11493);
nor U12253 (N_12253,N_10348,N_8696);
xnor U12254 (N_12254,N_11183,N_10678);
nand U12255 (N_12255,N_8254,N_11855);
or U12256 (N_12256,N_11807,N_11349);
nand U12257 (N_12257,N_9369,N_9211);
nand U12258 (N_12258,N_11487,N_11723);
or U12259 (N_12259,N_10566,N_11393);
and U12260 (N_12260,N_9325,N_9096);
or U12261 (N_12261,N_9812,N_10435);
nand U12262 (N_12262,N_10764,N_9639);
xnor U12263 (N_12263,N_11170,N_10814);
nand U12264 (N_12264,N_10694,N_10752);
or U12265 (N_12265,N_11686,N_11288);
nand U12266 (N_12266,N_8363,N_8965);
nor U12267 (N_12267,N_9977,N_8742);
nand U12268 (N_12268,N_9197,N_10799);
nand U12269 (N_12269,N_9004,N_8591);
xor U12270 (N_12270,N_9623,N_8913);
and U12271 (N_12271,N_10230,N_9327);
nor U12272 (N_12272,N_11687,N_8202);
xnor U12273 (N_12273,N_10310,N_9596);
nor U12274 (N_12274,N_8058,N_8947);
nor U12275 (N_12275,N_9701,N_10060);
nand U12276 (N_12276,N_10991,N_11818);
nand U12277 (N_12277,N_11498,N_9330);
or U12278 (N_12278,N_9744,N_8794);
nand U12279 (N_12279,N_9688,N_9753);
nor U12280 (N_12280,N_11759,N_8154);
nor U12281 (N_12281,N_8565,N_9569);
nor U12282 (N_12282,N_11222,N_10770);
nor U12283 (N_12283,N_10918,N_10043);
xnor U12284 (N_12284,N_11861,N_11863);
and U12285 (N_12285,N_8590,N_11225);
and U12286 (N_12286,N_11808,N_8517);
xnor U12287 (N_12287,N_8381,N_11865);
nor U12288 (N_12288,N_9459,N_8662);
nor U12289 (N_12289,N_10195,N_11245);
nor U12290 (N_12290,N_8505,N_11113);
or U12291 (N_12291,N_8776,N_11034);
and U12292 (N_12292,N_11377,N_8799);
nand U12293 (N_12293,N_8025,N_9161);
and U12294 (N_12294,N_10009,N_8546);
and U12295 (N_12295,N_8499,N_8693);
nand U12296 (N_12296,N_11167,N_10221);
or U12297 (N_12297,N_9708,N_8421);
or U12298 (N_12298,N_11151,N_10501);
xor U12299 (N_12299,N_11091,N_11841);
or U12300 (N_12300,N_10138,N_11883);
nor U12301 (N_12301,N_9401,N_9139);
nor U12302 (N_12302,N_11187,N_10941);
xnor U12303 (N_12303,N_10979,N_11521);
xor U12304 (N_12304,N_8042,N_10654);
nand U12305 (N_12305,N_11836,N_11324);
nand U12306 (N_12306,N_9563,N_10330);
nor U12307 (N_12307,N_8525,N_8153);
and U12308 (N_12308,N_10507,N_9771);
nand U12309 (N_12309,N_10647,N_8046);
and U12310 (N_12310,N_8712,N_11301);
or U12311 (N_12311,N_11483,N_9117);
or U12312 (N_12312,N_10311,N_9638);
nand U12313 (N_12313,N_10096,N_9212);
nand U12314 (N_12314,N_9375,N_9436);
nor U12315 (N_12315,N_11918,N_10888);
and U12316 (N_12316,N_8303,N_10545);
nand U12317 (N_12317,N_9932,N_10669);
nor U12318 (N_12318,N_8726,N_10745);
and U12319 (N_12319,N_11875,N_11882);
or U12320 (N_12320,N_11767,N_9853);
nor U12321 (N_12321,N_9109,N_10586);
nor U12322 (N_12322,N_9199,N_11007);
and U12323 (N_12323,N_10057,N_11797);
nand U12324 (N_12324,N_10524,N_9393);
or U12325 (N_12325,N_8365,N_10414);
nor U12326 (N_12326,N_9642,N_9519);
or U12327 (N_12327,N_8438,N_10847);
or U12328 (N_12328,N_10964,N_8752);
nand U12329 (N_12329,N_10437,N_11103);
nand U12330 (N_12330,N_10151,N_10097);
nor U12331 (N_12331,N_9195,N_10342);
and U12332 (N_12332,N_9912,N_10505);
xnor U12333 (N_12333,N_10424,N_9173);
and U12334 (N_12334,N_9984,N_11424);
and U12335 (N_12335,N_10278,N_9595);
nand U12336 (N_12336,N_10399,N_8133);
nor U12337 (N_12337,N_9572,N_8571);
nand U12338 (N_12338,N_8911,N_9683);
or U12339 (N_12339,N_10667,N_8092);
or U12340 (N_12340,N_11540,N_8761);
and U12341 (N_12341,N_9508,N_10223);
nor U12342 (N_12342,N_11663,N_10869);
or U12343 (N_12343,N_9515,N_8137);
and U12344 (N_12344,N_9802,N_8814);
or U12345 (N_12345,N_11485,N_10738);
or U12346 (N_12346,N_10851,N_10478);
nor U12347 (N_12347,N_9750,N_9910);
nor U12348 (N_12348,N_8409,N_8311);
nor U12349 (N_12349,N_10594,N_10580);
and U12350 (N_12350,N_9209,N_10037);
nor U12351 (N_12351,N_8991,N_8142);
nor U12352 (N_12352,N_11484,N_10027);
nand U12353 (N_12353,N_11423,N_9162);
nand U12354 (N_12354,N_9244,N_11065);
and U12355 (N_12355,N_9461,N_10412);
nand U12356 (N_12356,N_8881,N_10637);
nand U12357 (N_12357,N_11295,N_10264);
nand U12358 (N_12358,N_10425,N_10870);
xor U12359 (N_12359,N_9838,N_9962);
nor U12360 (N_12360,N_10966,N_9263);
or U12361 (N_12361,N_9815,N_11202);
nand U12362 (N_12362,N_10857,N_11195);
or U12363 (N_12363,N_11112,N_10476);
and U12364 (N_12364,N_10692,N_11608);
nand U12365 (N_12365,N_8820,N_8194);
and U12366 (N_12366,N_10321,N_11426);
nand U12367 (N_12367,N_11001,N_8657);
xor U12368 (N_12368,N_8632,N_8542);
and U12369 (N_12369,N_11874,N_10703);
and U12370 (N_12370,N_10258,N_11913);
and U12371 (N_12371,N_8279,N_8047);
or U12372 (N_12372,N_10760,N_11389);
nor U12373 (N_12373,N_9051,N_11347);
nor U12374 (N_12374,N_11277,N_8111);
and U12375 (N_12375,N_11051,N_11434);
nand U12376 (N_12376,N_10249,N_8620);
and U12377 (N_12377,N_11531,N_11881);
xnor U12378 (N_12378,N_9599,N_9616);
or U12379 (N_12379,N_9719,N_8119);
nand U12380 (N_12380,N_10559,N_10884);
and U12381 (N_12381,N_9759,N_11858);
and U12382 (N_12382,N_11612,N_8321);
and U12383 (N_12383,N_10325,N_9359);
and U12384 (N_12384,N_10970,N_11384);
and U12385 (N_12385,N_9449,N_8942);
xnor U12386 (N_12386,N_11085,N_8478);
or U12387 (N_12387,N_9687,N_9801);
and U12388 (N_12388,N_11074,N_11139);
and U12389 (N_12389,N_9233,N_8760);
xor U12390 (N_12390,N_9741,N_8041);
or U12391 (N_12391,N_8541,N_11060);
or U12392 (N_12392,N_9159,N_9329);
and U12393 (N_12393,N_8235,N_11639);
nand U12394 (N_12394,N_8977,N_8293);
xnor U12395 (N_12395,N_8090,N_10046);
nor U12396 (N_12396,N_11370,N_10184);
or U12397 (N_12397,N_9691,N_11857);
nand U12398 (N_12398,N_11359,N_8264);
or U12399 (N_12399,N_9446,N_8339);
or U12400 (N_12400,N_9260,N_11430);
nand U12401 (N_12401,N_10309,N_10853);
nand U12402 (N_12402,N_11161,N_10990);
or U12403 (N_12403,N_8707,N_8956);
nor U12404 (N_12404,N_10621,N_10393);
nand U12405 (N_12405,N_8692,N_11429);
nand U12406 (N_12406,N_9560,N_9057);
and U12407 (N_12407,N_8220,N_11990);
nand U12408 (N_12408,N_11180,N_10176);
and U12409 (N_12409,N_9494,N_11337);
nor U12410 (N_12410,N_10938,N_10080);
nor U12411 (N_12411,N_9308,N_10082);
and U12412 (N_12412,N_9681,N_9499);
or U12413 (N_12413,N_10601,N_10616);
nor U12414 (N_12414,N_10627,N_11021);
nand U12415 (N_12415,N_10021,N_9651);
and U12416 (N_12416,N_11331,N_11709);
nand U12417 (N_12417,N_10626,N_11099);
and U12418 (N_12418,N_9092,N_10307);
nor U12419 (N_12419,N_10704,N_11079);
nand U12420 (N_12420,N_10141,N_10334);
or U12421 (N_12421,N_8221,N_11596);
xor U12422 (N_12422,N_9980,N_9528);
nor U12423 (N_12423,N_10876,N_9861);
or U12424 (N_12424,N_10535,N_9624);
nand U12425 (N_12425,N_11239,N_10827);
or U12426 (N_12426,N_10836,N_9114);
and U12427 (N_12427,N_9982,N_8621);
xnor U12428 (N_12428,N_11224,N_11645);
xor U12429 (N_12429,N_10206,N_8986);
nor U12430 (N_12430,N_10091,N_8497);
or U12431 (N_12431,N_10458,N_11565);
or U12432 (N_12432,N_9183,N_9050);
nor U12433 (N_12433,N_10685,N_9431);
nor U12434 (N_12434,N_9754,N_8866);
xor U12435 (N_12435,N_8847,N_9405);
and U12436 (N_12436,N_11654,N_11728);
and U12437 (N_12437,N_11515,N_9570);
nor U12438 (N_12438,N_10541,N_11804);
nand U12439 (N_12439,N_11542,N_11977);
xnor U12440 (N_12440,N_11958,N_8320);
and U12441 (N_12441,N_9761,N_11503);
nand U12442 (N_12442,N_9419,N_11850);
nand U12443 (N_12443,N_11045,N_11506);
nand U12444 (N_12444,N_11631,N_9574);
or U12445 (N_12445,N_10806,N_10758);
nor U12446 (N_12446,N_9964,N_11734);
nand U12447 (N_12447,N_11621,N_9052);
nor U12448 (N_12448,N_8648,N_9452);
nor U12449 (N_12449,N_9579,N_8759);
or U12450 (N_12450,N_9834,N_8490);
nor U12451 (N_12451,N_8345,N_9664);
and U12452 (N_12452,N_9993,N_9493);
or U12453 (N_12453,N_10256,N_11189);
nor U12454 (N_12454,N_10133,N_10473);
and U12455 (N_12455,N_11587,N_11784);
nor U12456 (N_12456,N_9931,N_8068);
nand U12457 (N_12457,N_9841,N_10547);
nor U12458 (N_12458,N_11084,N_10674);
nor U12459 (N_12459,N_9707,N_9121);
or U12460 (N_12460,N_9696,N_9306);
and U12461 (N_12461,N_11838,N_11396);
nand U12462 (N_12462,N_10628,N_11076);
and U12463 (N_12463,N_8064,N_8348);
and U12464 (N_12464,N_9757,N_9108);
and U12465 (N_12465,N_9001,N_8226);
xnor U12466 (N_12466,N_9923,N_8334);
or U12467 (N_12467,N_11291,N_9816);
nand U12468 (N_12468,N_10581,N_11941);
nor U12469 (N_12469,N_8933,N_10546);
and U12470 (N_12470,N_8433,N_8640);
or U12471 (N_12471,N_9665,N_11764);
nor U12472 (N_12472,N_8130,N_11124);
nor U12473 (N_12473,N_10525,N_10762);
nand U12474 (N_12474,N_10482,N_9526);
or U12475 (N_12475,N_8573,N_11131);
xor U12476 (N_12476,N_10772,N_8605);
nand U12477 (N_12477,N_9354,N_10000);
and U12478 (N_12478,N_8132,N_8411);
nor U12479 (N_12479,N_11984,N_11476);
nand U12480 (N_12480,N_11906,N_11098);
and U12481 (N_12481,N_9805,N_8997);
nor U12482 (N_12482,N_11877,N_9054);
nand U12483 (N_12483,N_8060,N_9456);
nor U12484 (N_12484,N_9933,N_10676);
nand U12485 (N_12485,N_10187,N_10910);
nor U12486 (N_12486,N_8269,N_11438);
or U12487 (N_12487,N_11829,N_8634);
nor U12488 (N_12488,N_11125,N_8652);
nand U12489 (N_12489,N_9631,N_9992);
or U12490 (N_12490,N_10681,N_8556);
nor U12491 (N_12491,N_11583,N_9430);
or U12492 (N_12492,N_10898,N_10630);
nand U12493 (N_12493,N_9453,N_10998);
and U12494 (N_12494,N_11217,N_9617);
and U12495 (N_12495,N_11625,N_11092);
or U12496 (N_12496,N_11554,N_9825);
nor U12497 (N_12497,N_9903,N_9378);
and U12498 (N_12498,N_10824,N_8899);
and U12499 (N_12499,N_11063,N_9236);
and U12500 (N_12500,N_9068,N_8670);
nor U12501 (N_12501,N_10240,N_9103);
and U12502 (N_12502,N_10613,N_9882);
or U12503 (N_12503,N_9905,N_10332);
or U12504 (N_12504,N_11514,N_11971);
xor U12505 (N_12505,N_8357,N_11907);
and U12506 (N_12506,N_10241,N_11097);
or U12507 (N_12507,N_9101,N_11561);
nor U12508 (N_12508,N_9857,N_8817);
nor U12509 (N_12509,N_11265,N_8518);
or U12510 (N_12510,N_11168,N_11489);
or U12511 (N_12511,N_8210,N_8301);
nand U12512 (N_12512,N_11589,N_11966);
xor U12513 (N_12513,N_8998,N_9581);
nand U12514 (N_12514,N_10265,N_8237);
nor U12515 (N_12515,N_11724,N_9975);
or U12516 (N_12516,N_9074,N_11385);
nand U12517 (N_12517,N_11130,N_8376);
or U12518 (N_12518,N_10523,N_9355);
xor U12519 (N_12519,N_11974,N_10607);
and U12520 (N_12520,N_9060,N_8981);
nand U12521 (N_12521,N_8660,N_8437);
nor U12522 (N_12522,N_11775,N_9474);
nand U12523 (N_12523,N_8765,N_10842);
nand U12524 (N_12524,N_11155,N_9615);
xor U12525 (N_12525,N_9868,N_11880);
nand U12526 (N_12526,N_10804,N_9469);
nor U12527 (N_12527,N_11144,N_9368);
nand U12528 (N_12528,N_11570,N_8002);
nand U12529 (N_12529,N_9402,N_9486);
and U12530 (N_12530,N_9017,N_11134);
xnor U12531 (N_12531,N_11715,N_10118);
or U12532 (N_12532,N_8197,N_9371);
and U12533 (N_12533,N_11119,N_8514);
or U12534 (N_12534,N_9049,N_9504);
nor U12535 (N_12535,N_10268,N_10585);
xor U12536 (N_12536,N_9062,N_10160);
or U12537 (N_12537,N_11834,N_11176);
nand U12538 (N_12538,N_10530,N_10282);
nor U12539 (N_12539,N_11117,N_10527);
xor U12540 (N_12540,N_11142,N_9590);
nand U12541 (N_12541,N_11089,N_11082);
nor U12542 (N_12542,N_9175,N_8912);
or U12543 (N_12543,N_10374,N_11800);
or U12544 (N_12544,N_8843,N_9473);
nor U12545 (N_12545,N_8949,N_11388);
nand U12546 (N_12546,N_10409,N_9082);
nor U12547 (N_12547,N_9351,N_8921);
nand U12548 (N_12548,N_8351,N_10395);
nor U12549 (N_12549,N_11864,N_8212);
nand U12550 (N_12550,N_11970,N_9208);
nor U12551 (N_12551,N_10197,N_8498);
or U12552 (N_12552,N_10666,N_10315);
and U12553 (N_12553,N_8926,N_8834);
and U12554 (N_12554,N_10253,N_10340);
xor U12555 (N_12555,N_10683,N_10689);
or U12556 (N_12556,N_8896,N_9799);
or U12557 (N_12557,N_8521,N_8844);
nor U12558 (N_12558,N_8667,N_10235);
and U12559 (N_12559,N_11744,N_9307);
and U12560 (N_12560,N_10569,N_10822);
nand U12561 (N_12561,N_8275,N_11086);
and U12562 (N_12562,N_9773,N_9978);
or U12563 (N_12563,N_8342,N_9188);
nand U12564 (N_12564,N_11622,N_11681);
or U12565 (N_12565,N_11640,N_11999);
or U12566 (N_12566,N_9097,N_11928);
nand U12567 (N_12567,N_8530,N_9548);
nor U12568 (N_12568,N_8624,N_11093);
and U12569 (N_12569,N_10140,N_8552);
and U12570 (N_12570,N_10696,N_9938);
nor U12571 (N_12571,N_9774,N_9552);
nand U12572 (N_12572,N_8716,N_11922);
nor U12573 (N_12573,N_11617,N_8371);
xor U12574 (N_12574,N_11598,N_11252);
xnor U12575 (N_12575,N_10573,N_11591);
nand U12576 (N_12576,N_9635,N_8871);
or U12577 (N_12577,N_8032,N_10443);
nand U12578 (N_12578,N_9710,N_9089);
nand U12579 (N_12579,N_9673,N_10485);
or U12580 (N_12580,N_8464,N_9663);
nor U12581 (N_12581,N_8475,N_8503);
and U12582 (N_12582,N_8884,N_8496);
or U12583 (N_12583,N_11468,N_9290);
and U12584 (N_12584,N_11866,N_11752);
nand U12585 (N_12585,N_10550,N_11499);
and U12586 (N_12586,N_10089,N_11286);
xnor U12587 (N_12587,N_8816,N_11126);
nand U12588 (N_12588,N_9029,N_9243);
and U12589 (N_12589,N_10298,N_8258);
and U12590 (N_12590,N_9295,N_9016);
nor U12591 (N_12591,N_9827,N_11054);
and U12592 (N_12592,N_10724,N_11140);
nor U12593 (N_12593,N_9261,N_8399);
nand U12594 (N_12594,N_8833,N_10913);
nand U12595 (N_12595,N_10564,N_10439);
nand U12596 (N_12596,N_8098,N_10106);
nor U12597 (N_12597,N_8402,N_9626);
nor U12598 (N_12598,N_11357,N_10643);
or U12599 (N_12599,N_10078,N_8786);
or U12600 (N_12600,N_11967,N_10247);
nand U12601 (N_12601,N_10376,N_8248);
or U12602 (N_12602,N_9760,N_11939);
and U12603 (N_12603,N_10285,N_9488);
nor U12604 (N_12604,N_10150,N_9942);
nor U12605 (N_12605,N_10381,N_9809);
nor U12606 (N_12606,N_10333,N_10403);
or U12607 (N_12607,N_9509,N_8481);
and U12608 (N_12608,N_11641,N_8647);
nand U12609 (N_12609,N_11600,N_9549);
nand U12610 (N_12610,N_9785,N_10099);
and U12611 (N_12611,N_11293,N_8725);
xnor U12612 (N_12612,N_8453,N_9983);
or U12613 (N_12613,N_11132,N_9344);
nand U12614 (N_12614,N_9135,N_8121);
nand U12615 (N_12615,N_11696,N_11870);
and U12616 (N_12616,N_10385,N_9680);
nor U12617 (N_12617,N_9471,N_11673);
nor U12618 (N_12618,N_11031,N_9298);
nand U12619 (N_12619,N_10557,N_11214);
nor U12620 (N_12620,N_10145,N_8936);
and U12621 (N_12621,N_8604,N_8778);
nand U12622 (N_12622,N_10675,N_10551);
nor U12623 (N_12623,N_10243,N_11366);
nand U12624 (N_12624,N_11853,N_8388);
nor U12625 (N_12625,N_11610,N_10384);
or U12626 (N_12626,N_8508,N_9104);
nand U12627 (N_12627,N_9217,N_8581);
nand U12628 (N_12628,N_10166,N_10301);
nor U12629 (N_12629,N_9535,N_8813);
nor U12630 (N_12630,N_9272,N_9353);
or U12631 (N_12631,N_11432,N_8280);
or U12632 (N_12632,N_8970,N_10763);
or U12633 (N_12633,N_8014,N_9591);
nand U12634 (N_12634,N_9541,N_10274);
xor U12635 (N_12635,N_9894,N_10831);
nand U12636 (N_12636,N_9888,N_9630);
and U12637 (N_12637,N_9860,N_11785);
nand U12638 (N_12638,N_10963,N_10742);
and U12639 (N_12639,N_8733,N_10319);
or U12640 (N_12640,N_8003,N_9377);
or U12641 (N_12641,N_9575,N_10880);
nand U12642 (N_12642,N_10185,N_11015);
nand U12643 (N_12643,N_8996,N_10338);
and U12644 (N_12644,N_8117,N_10825);
nor U12645 (N_12645,N_9669,N_11078);
xor U12646 (N_12646,N_10502,N_9420);
nand U12647 (N_12647,N_9545,N_10756);
nand U12648 (N_12648,N_8584,N_9846);
xor U12649 (N_12649,N_9292,N_11680);
nor U12650 (N_12650,N_9397,N_10727);
or U12651 (N_12651,N_9973,N_9177);
nor U12652 (N_12652,N_8569,N_11330);
or U12653 (N_12653,N_9811,N_9676);
or U12654 (N_12654,N_8729,N_9346);
nand U12655 (N_12655,N_10172,N_10467);
nand U12656 (N_12656,N_11802,N_10496);
nand U12657 (N_12657,N_11232,N_8456);
xnor U12658 (N_12658,N_8694,N_9914);
or U12659 (N_12659,N_8375,N_8355);
and U12660 (N_12660,N_9830,N_10122);
and U12661 (N_12661,N_10903,N_10747);
nand U12662 (N_12662,N_8238,N_10262);
and U12663 (N_12663,N_11315,N_11399);
nand U12664 (N_12664,N_8862,N_11548);
or U12665 (N_12665,N_9679,N_10544);
and U12666 (N_12666,N_11878,N_11975);
or U12667 (N_12667,N_9536,N_9922);
nand U12668 (N_12668,N_9153,N_8186);
nand U12669 (N_12669,N_9692,N_9048);
nand U12670 (N_12670,N_8346,N_11024);
nor U12671 (N_12671,N_10583,N_10679);
xnor U12672 (N_12672,N_10224,N_8180);
or U12673 (N_12673,N_10098,N_11449);
nor U12674 (N_12674,N_9406,N_9943);
or U12675 (N_12675,N_11783,N_9134);
nand U12676 (N_12676,N_8934,N_10602);
nor U12677 (N_12677,N_9998,N_10019);
and U12678 (N_12678,N_8930,N_11924);
or U12679 (N_12679,N_11544,N_11753);
or U12680 (N_12680,N_10026,N_10901);
nor U12681 (N_12681,N_9592,N_10303);
and U12682 (N_12682,N_11254,N_8244);
nor U12683 (N_12683,N_8013,N_8606);
and U12684 (N_12684,N_9558,N_11191);
and U12685 (N_12685,N_8631,N_9160);
nor U12686 (N_12686,N_9427,N_9416);
or U12687 (N_12687,N_8394,N_10993);
and U12688 (N_12688,N_8294,N_10906);
nand U12689 (N_12689,N_9958,N_10053);
nand U12690 (N_12690,N_11805,N_10618);
or U12691 (N_12691,N_8878,N_10978);
nor U12692 (N_12692,N_11066,N_10238);
or U12693 (N_12693,N_9842,N_8868);
or U12694 (N_12694,N_8045,N_9969);
or U12695 (N_12695,N_8849,N_9775);
nand U12696 (N_12696,N_9913,N_9546);
or U12697 (N_12697,N_11259,N_11372);
nand U12698 (N_12698,N_9758,N_11828);
nand U12699 (N_12699,N_9287,N_11083);
nor U12700 (N_12700,N_8608,N_8727);
or U12701 (N_12701,N_10104,N_8572);
nor U12702 (N_12702,N_10868,N_9086);
nor U12703 (N_12703,N_10862,N_8048);
nand U12704 (N_12704,N_11411,N_8952);
and U12705 (N_12705,N_11397,N_8570);
nand U12706 (N_12706,N_11153,N_10582);
nor U12707 (N_12707,N_10186,N_9131);
nand U12708 (N_12708,N_11795,N_9970);
nand U12709 (N_12709,N_9803,N_10855);
nor U12710 (N_12710,N_9840,N_11229);
nor U12711 (N_12711,N_11781,N_10861);
or U12712 (N_12712,N_11181,N_9305);
and U12713 (N_12713,N_8535,N_11100);
and U12714 (N_12714,N_9876,N_9439);
or U12715 (N_12715,N_8583,N_9067);
nor U12716 (N_12716,N_10095,N_11022);
and U12717 (N_12717,N_11607,N_8352);
nand U12718 (N_12718,N_9266,N_10318);
and U12719 (N_12719,N_10005,N_8116);
and U12720 (N_12720,N_10367,N_8564);
nor U12721 (N_12721,N_10175,N_10463);
or U12722 (N_12722,N_9403,N_10733);
nand U12723 (N_12723,N_9529,N_11509);
or U12724 (N_12724,N_9990,N_11358);
or U12725 (N_12725,N_10038,N_9608);
or U12726 (N_12726,N_8129,N_11666);
nor U12727 (N_12727,N_11892,N_10518);
nor U12728 (N_12728,N_10201,N_10378);
or U12729 (N_12729,N_9926,N_9739);
or U12730 (N_12730,N_9513,N_9187);
xor U12731 (N_12731,N_8740,N_8085);
nand U12732 (N_12732,N_11488,N_9619);
xnor U12733 (N_12733,N_11025,N_11081);
or U12734 (N_12734,N_9510,N_11743);
nand U12735 (N_12735,N_9690,N_10687);
xor U12736 (N_12736,N_9098,N_10028);
nand U12737 (N_12737,N_8860,N_8971);
nor U12738 (N_12738,N_11993,N_11129);
and U12739 (N_12739,N_10620,N_9365);
nor U12740 (N_12740,N_8826,N_9871);
or U12741 (N_12741,N_10572,N_11879);
or U12742 (N_12742,N_9206,N_9027);
nand U12743 (N_12743,N_8659,N_10215);
nor U12744 (N_12744,N_9879,N_9751);
or U12745 (N_12745,N_11049,N_8779);
or U12746 (N_12746,N_9706,N_11294);
or U12747 (N_12747,N_9215,N_10369);
or U12748 (N_12748,N_9755,N_10267);
nor U12749 (N_12749,N_8281,N_10272);
nor U12750 (N_12750,N_10781,N_11486);
xor U12751 (N_12751,N_11815,N_8332);
or U12752 (N_12752,N_8992,N_11780);
nand U12753 (N_12753,N_8031,N_9111);
and U12754 (N_12754,N_10421,N_11810);
nor U12755 (N_12755,N_11339,N_10939);
nor U12756 (N_12756,N_10190,N_10002);
or U12757 (N_12757,N_8350,N_11518);
or U12758 (N_12758,N_10035,N_10284);
nor U12759 (N_12759,N_8863,N_8823);
nand U12760 (N_12760,N_8302,N_10808);
and U12761 (N_12761,N_11991,N_8477);
or U12762 (N_12762,N_8187,N_9968);
nor U12763 (N_12763,N_9411,N_8524);
nand U12764 (N_12764,N_11940,N_8167);
and U12765 (N_12765,N_11750,N_10955);
xnor U12766 (N_12766,N_11447,N_11036);
nor U12767 (N_12767,N_8362,N_8317);
or U12768 (N_12768,N_9460,N_11976);
nand U12769 (N_12769,N_10835,N_11675);
nand U12770 (N_12770,N_9686,N_11567);
and U12771 (N_12771,N_10510,N_8555);
nor U12772 (N_12772,N_9930,N_10608);
and U12773 (N_12773,N_11717,N_9826);
and U12774 (N_12774,N_8988,N_11513);
nand U12775 (N_12775,N_9259,N_8519);
nand U12776 (N_12776,N_9906,N_11018);
nand U12777 (N_12777,N_10217,N_9900);
nand U12778 (N_12778,N_10950,N_10540);
nor U12779 (N_12779,N_9656,N_9895);
nor U12780 (N_12780,N_9445,N_8784);
xnor U12781 (N_12781,N_11253,N_11273);
and U12782 (N_12782,N_8715,N_11920);
and U12783 (N_12783,N_11114,N_8821);
nand U12784 (N_12784,N_9684,N_10445);
or U12785 (N_12785,N_11287,N_9605);
and U12786 (N_12786,N_11657,N_8595);
xnor U12787 (N_12787,N_11267,N_10810);
or U12788 (N_12788,N_11903,N_11373);
nor U12789 (N_12789,N_10244,N_8435);
nor U12790 (N_12790,N_10457,N_11402);
nor U12791 (N_12791,N_9181,N_8920);
nand U12792 (N_12792,N_10387,N_11262);
or U12793 (N_12793,N_9012,N_9889);
or U12794 (N_12794,N_9332,N_8954);
nand U12795 (N_12795,N_9718,N_9387);
and U12796 (N_12796,N_10032,N_9414);
nor U12797 (N_12797,N_9928,N_11136);
nand U12798 (N_12798,N_9479,N_11056);
and U12799 (N_12799,N_10152,N_10007);
xnor U12800 (N_12800,N_10418,N_10753);
nand U12801 (N_12801,N_11352,N_11683);
nor U12802 (N_12802,N_9149,N_10591);
or U12803 (N_12803,N_11208,N_10072);
xor U12804 (N_12804,N_11409,N_8717);
or U12805 (N_12805,N_10736,N_10161);
nor U12806 (N_12806,N_9824,N_11504);
nand U12807 (N_12807,N_10641,N_8218);
or U12808 (N_12808,N_11361,N_10459);
or U12809 (N_12809,N_11747,N_11231);
or U12810 (N_12810,N_9158,N_8093);
and U12811 (N_12811,N_9037,N_8207);
and U12812 (N_12812,N_11826,N_10930);
nand U12813 (N_12813,N_11201,N_9722);
xnor U12814 (N_12814,N_10611,N_10339);
nand U12815 (N_12815,N_10849,N_9349);
and U12816 (N_12816,N_9539,N_10512);
or U12817 (N_12817,N_9806,N_10336);
and U12818 (N_12818,N_11595,N_9601);
nand U12819 (N_12819,N_10499,N_11943);
nor U12820 (N_12820,N_8044,N_8325);
nor U12821 (N_12821,N_9178,N_11552);
nand U12822 (N_12822,N_10288,N_10871);
nor U12823 (N_12823,N_11605,N_8744);
nand U12824 (N_12824,N_8743,N_8520);
nor U12825 (N_12825,N_11620,N_9582);
or U12826 (N_12826,N_9659,N_11588);
or U12827 (N_12827,N_8705,N_11458);
or U12828 (N_12828,N_9191,N_11526);
or U12829 (N_12829,N_8179,N_9915);
or U12830 (N_12830,N_8989,N_10066);
nand U12831 (N_12831,N_9485,N_11374);
nor U12832 (N_12832,N_11300,N_8629);
nand U12833 (N_12833,N_11901,N_8567);
nand U12834 (N_12834,N_11851,N_9839);
nand U12835 (N_12835,N_10483,N_8513);
or U12836 (N_12836,N_10165,N_10841);
and U12837 (N_12837,N_8957,N_11237);
nand U12838 (N_12838,N_11260,N_10024);
or U12839 (N_12839,N_10974,N_8233);
nor U12840 (N_12840,N_11665,N_11692);
or U12841 (N_12841,N_10064,N_9959);
and U12842 (N_12842,N_8891,N_11837);
nand U12843 (N_12843,N_9966,N_9724);
and U12844 (N_12844,N_10163,N_8649);
and U12845 (N_12845,N_9204,N_8103);
or U12846 (N_12846,N_9557,N_10567);
or U12847 (N_12847,N_8033,N_9115);
nand U12848 (N_12848,N_11133,N_9698);
nand U12849 (N_12849,N_8574,N_8156);
nand U12850 (N_12850,N_11465,N_11410);
and U12851 (N_12851,N_11227,N_10179);
and U12852 (N_12852,N_9154,N_10056);
nand U12853 (N_12853,N_11910,N_9497);
nor U12854 (N_12854,N_9009,N_8636);
and U12855 (N_12855,N_10390,N_11650);
nand U12856 (N_12856,N_10571,N_10033);
and U12857 (N_12857,N_10710,N_9520);
and U12858 (N_12858,N_9421,N_11779);
or U12859 (N_12859,N_9787,N_9988);
and U12860 (N_12860,N_8105,N_10729);
nand U12861 (N_12861,N_10261,N_10771);
nand U12862 (N_12862,N_9584,N_9662);
nor U12863 (N_12863,N_11353,N_8124);
or U12864 (N_12864,N_8443,N_8188);
nand U12865 (N_12865,N_8929,N_10516);
or U12866 (N_12866,N_10916,N_11796);
and U12867 (N_12867,N_11633,N_10568);
nand U12868 (N_12868,N_10671,N_9780);
nand U12869 (N_12869,N_9252,N_9655);
or U12870 (N_12870,N_11557,N_10529);
or U12871 (N_12871,N_9950,N_8702);
nor U12872 (N_12872,N_11019,N_10093);
and U12873 (N_12873,N_9246,N_11964);
and U12874 (N_12874,N_11364,N_8253);
nor U12875 (N_12875,N_9955,N_11440);
or U12876 (N_12876,N_10245,N_10590);
or U12877 (N_12877,N_8095,N_11708);
nand U12878 (N_12878,N_9324,N_8382);
xnor U12879 (N_12879,N_11188,N_11739);
and U12880 (N_12880,N_11535,N_8333);
and U12881 (N_12881,N_10114,N_10170);
nand U12882 (N_12882,N_8533,N_11004);
nand U12883 (N_12883,N_10917,N_10147);
nor U12884 (N_12884,N_10081,N_10850);
or U12885 (N_12885,N_10305,N_8195);
nand U12886 (N_12886,N_9155,N_10242);
and U12887 (N_12887,N_8568,N_11957);
and U12888 (N_12888,N_10634,N_9961);
nand U12889 (N_12889,N_11550,N_9716);
nor U12890 (N_12890,N_11529,N_10680);
and U12891 (N_12891,N_11714,N_9808);
or U12892 (N_12892,N_8754,N_8750);
xor U12893 (N_12893,N_9249,N_8724);
or U12894 (N_12894,N_8385,N_10887);
or U12895 (N_12895,N_11947,N_8656);
nor U12896 (N_12896,N_11911,N_8800);
and U12897 (N_12897,N_11177,N_11659);
nand U12898 (N_12898,N_8374,N_10299);
and U12899 (N_12899,N_10905,N_8406);
nand U12900 (N_12900,N_8753,N_11742);
and U12901 (N_12901,N_11320,N_10229);
nor U12902 (N_12902,N_11768,N_11435);
nand U12903 (N_12903,N_8219,N_9058);
nor U12904 (N_12904,N_11653,N_11475);
nand U12905 (N_12905,N_8343,N_10107);
xnor U12906 (N_12906,N_8709,N_8151);
or U12907 (N_12907,N_11616,N_11344);
nor U12908 (N_12908,N_10670,N_10600);
nand U12909 (N_12909,N_11280,N_11250);
and U12910 (N_12910,N_9006,N_9025);
xor U12911 (N_12911,N_10405,N_8155);
nor U12912 (N_12912,N_9075,N_11422);
or U12913 (N_12913,N_8370,N_9878);
xnor U12914 (N_12914,N_11912,N_10739);
and U12915 (N_12915,N_9214,N_9603);
or U12916 (N_12916,N_11174,N_11450);
nor U12917 (N_12917,N_11008,N_10012);
or U12918 (N_12918,N_10260,N_8114);
nor U12919 (N_12919,N_8633,N_8969);
xor U12920 (N_12920,N_10490,N_10398);
and U12921 (N_12921,N_11163,N_10291);
and U12922 (N_12922,N_9733,N_9011);
nor U12923 (N_12923,N_11198,N_10845);
nand U12924 (N_12924,N_10154,N_11123);
and U12925 (N_12925,N_9053,N_10025);
nor U12926 (N_12926,N_10914,N_8273);
or U12927 (N_12927,N_8553,N_8146);
or U12928 (N_12928,N_11511,N_11809);
nor U12929 (N_12929,N_9869,N_8241);
or U12930 (N_12930,N_11579,N_8796);
and U12931 (N_12931,N_10796,N_9483);
or U12932 (N_12932,N_11871,N_10216);
nor U12933 (N_12933,N_10174,N_8592);
or U12934 (N_12934,N_10470,N_10598);
nand U12935 (N_12935,N_11926,N_8531);
or U12936 (N_12936,N_9844,N_8793);
and U12937 (N_12937,N_8359,N_10068);
and U12938 (N_12938,N_8181,N_10171);
xnor U12939 (N_12939,N_8682,N_9142);
nand U12940 (N_12940,N_9088,N_8389);
nand U12941 (N_12941,N_10100,N_9136);
nand U12942 (N_12942,N_11439,N_10896);
and U12943 (N_12943,N_10449,N_11669);
xnor U12944 (N_12944,N_8026,N_8890);
nor U12945 (N_12945,N_10737,N_9301);
and U12946 (N_12946,N_8379,N_8272);
and U12947 (N_12947,N_8417,N_8861);
or U12948 (N_12948,N_10181,N_11735);
nand U12949 (N_12949,N_10029,N_10430);
nor U12950 (N_12950,N_11642,N_11013);
nand U12951 (N_12951,N_8593,N_8720);
nor U12952 (N_12952,N_10996,N_11314);
and U12953 (N_12953,N_8538,N_11551);
nand U12954 (N_12954,N_10132,N_10902);
nor U12955 (N_12955,N_8078,N_9715);
xor U12956 (N_12956,N_8008,N_8675);
and U12957 (N_12957,N_9907,N_11003);
or U12958 (N_12958,N_9985,N_8689);
xor U12959 (N_12959,N_8104,N_11674);
and U12960 (N_12960,N_8150,N_9286);
or U12961 (N_12961,N_9472,N_11556);
or U12962 (N_12962,N_11494,N_11481);
nor U12963 (N_12963,N_11233,N_11492);
nor U12964 (N_12964,N_8203,N_8730);
nand U12965 (N_12965,N_8432,N_8526);
nor U12966 (N_12966,N_8622,N_11463);
and U12967 (N_12967,N_11351,N_11053);
nor U12968 (N_12968,N_8243,N_11379);
nor U12969 (N_12969,N_10791,N_10617);
nor U12970 (N_12970,N_9951,N_9979);
nand U12971 (N_12971,N_8549,N_8630);
or U12972 (N_12972,N_9296,N_9200);
nor U12973 (N_12973,N_11207,N_8597);
and U12974 (N_12974,N_10042,N_8699);
and U12975 (N_12975,N_11560,N_8316);
or U12976 (N_12976,N_8980,N_11047);
xnor U12977 (N_12977,N_9076,N_10899);
nand U12978 (N_12978,N_10840,N_8815);
xnor U12979 (N_12979,N_8372,N_11075);
and U12980 (N_12980,N_10432,N_9457);
nand U12981 (N_12981,N_10859,N_10117);
and U12982 (N_12982,N_10994,N_8216);
nand U12983 (N_12983,N_11581,N_11094);
nand U12984 (N_12984,N_9920,N_11433);
nand U12985 (N_12985,N_10069,N_8979);
or U12986 (N_12986,N_11236,N_8247);
or U12987 (N_12987,N_10844,N_11073);
and U12988 (N_12988,N_10797,N_9078);
nand U12989 (N_12989,N_10599,N_9303);
and U12990 (N_12990,N_8398,N_9014);
and U12991 (N_12991,N_11350,N_11323);
nand U12992 (N_12992,N_8006,N_11480);
or U12993 (N_12993,N_9224,N_10932);
and U12994 (N_12994,N_10662,N_10233);
or U12995 (N_12995,N_9008,N_8425);
or U12996 (N_12996,N_10468,N_10995);
or U12997 (N_12997,N_10391,N_8767);
nand U12998 (N_12998,N_10484,N_10433);
or U12999 (N_12999,N_11057,N_9810);
nor U13000 (N_13000,N_8559,N_8386);
and U13001 (N_13001,N_9954,N_10789);
and U13002 (N_13002,N_9148,N_9356);
nand U13003 (N_13003,N_8001,N_8326);
nand U13004 (N_13004,N_10225,N_9366);
nor U13005 (N_13005,N_11799,N_9566);
nor U13006 (N_13006,N_8964,N_8289);
nand U13007 (N_13007,N_10461,N_9967);
nor U13008 (N_13008,N_8859,N_8079);
and U13009 (N_13009,N_10362,N_11798);
nand U13010 (N_13010,N_8589,N_9408);
and U13011 (N_13011,N_11831,N_10864);
nor U13012 (N_13012,N_8982,N_9989);
nor U13013 (N_13013,N_9223,N_8698);
nor U13014 (N_13014,N_8183,N_10946);
or U13015 (N_13015,N_10506,N_8582);
nand U13016 (N_13016,N_10503,N_10554);
xor U13017 (N_13017,N_10981,N_10361);
and U13018 (N_13018,N_10800,N_8908);
nand U13019 (N_13019,N_9736,N_9661);
nand U13020 (N_13020,N_9300,N_9725);
nor U13021 (N_13021,N_8324,N_9370);
or U13022 (N_13022,N_9443,N_9653);
and U13023 (N_13023,N_11460,N_10765);
nand U13024 (N_13024,N_10296,N_11456);
nor U13025 (N_13025,N_8223,N_8413);
and U13026 (N_13026,N_8178,N_9717);
or U13027 (N_13027,N_10560,N_10558);
nand U13028 (N_13028,N_8941,N_11428);
nor U13029 (N_13029,N_8213,N_11835);
nor U13030 (N_13030,N_11376,N_8020);
or U13031 (N_13031,N_9935,N_10351);
xor U13032 (N_13032,N_11962,N_11935);
or U13033 (N_13033,N_9865,N_11590);
nor U13034 (N_13034,N_8190,N_9491);
or U13035 (N_13035,N_10919,N_11014);
and U13036 (N_13036,N_10980,N_9466);
and U13037 (N_13037,N_11689,N_10304);
and U13038 (N_13038,N_8614,N_9102);
or U13039 (N_13039,N_8356,N_8327);
xnor U13040 (N_13040,N_10967,N_9727);
xnor U13041 (N_13041,N_10984,N_8285);
nand U13042 (N_13042,N_9202,N_8928);
nor U13043 (N_13043,N_9641,N_9434);
nor U13044 (N_13044,N_11699,N_9852);
nor U13045 (N_13045,N_9433,N_9304);
and U13046 (N_13046,N_8246,N_10997);
nand U13047 (N_13047,N_10164,N_11519);
nand U13048 (N_13048,N_8923,N_9147);
and U13049 (N_13049,N_9328,N_11369);
nor U13050 (N_13050,N_11712,N_10123);
or U13051 (N_13051,N_10125,N_9226);
nand U13052 (N_13052,N_11454,N_9898);
nor U13053 (N_13053,N_10537,N_11175);
and U13054 (N_13054,N_8392,N_9763);
or U13055 (N_13055,N_11833,N_10214);
nor U13056 (N_13056,N_9099,N_10952);
nor U13057 (N_13057,N_11961,N_9146);
xnor U13058 (N_13058,N_8512,N_9875);
and U13059 (N_13059,N_10648,N_9110);
nand U13060 (N_13060,N_9323,N_11510);
nand U13061 (N_13061,N_9542,N_9822);
and U13062 (N_13062,N_10700,N_9729);
or U13063 (N_13063,N_9376,N_9140);
nor U13064 (N_13064,N_9337,N_9789);
or U13065 (N_13065,N_8718,N_11731);
nand U13066 (N_13066,N_10196,N_10793);
and U13067 (N_13067,N_8561,N_8950);
or U13068 (N_13068,N_8960,N_11938);
nor U13069 (N_13069,N_8532,N_10721);
nand U13070 (N_13070,N_9798,N_10809);
xor U13071 (N_13071,N_11525,N_11362);
and U13072 (N_13072,N_10776,N_10838);
or U13073 (N_13073,N_10718,N_8134);
nand U13074 (N_13074,N_10092,N_11263);
nor U13075 (N_13075,N_10811,N_9231);
and U13076 (N_13076,N_9219,N_11777);
xnor U13077 (N_13077,N_10237,N_8436);
or U13078 (N_13078,N_11989,N_9019);
or U13079 (N_13079,N_10236,N_11719);
nor U13080 (N_13080,N_10538,N_8639);
nand U13081 (N_13081,N_9043,N_9234);
nand U13082 (N_13082,N_10712,N_8113);
or U13083 (N_13083,N_9553,N_11576);
nor U13084 (N_13084,N_11375,N_9167);
and U13085 (N_13085,N_8983,N_11408);
and U13086 (N_13086,N_10119,N_9829);
xor U13087 (N_13087,N_8189,N_10609);
nand U13088 (N_13088,N_9685,N_10624);
and U13089 (N_13089,N_8300,N_8795);
nor U13090 (N_13090,N_9274,N_10592);
xor U13091 (N_13091,N_11682,N_8082);
or U13092 (N_13092,N_8323,N_9454);
xnor U13093 (N_13093,N_8161,N_11909);
and U13094 (N_13094,N_11459,N_9854);
nor U13095 (N_13095,N_11058,N_11257);
nor U13096 (N_13096,N_11660,N_10124);
or U13097 (N_13097,N_9294,N_9237);
or U13098 (N_13098,N_9644,N_8397);
xor U13099 (N_13099,N_8403,N_8500);
nor U13100 (N_13100,N_8118,N_9339);
nand U13101 (N_13101,N_9795,N_10248);
nand U13102 (N_13102,N_8766,N_9580);
nand U13103 (N_13103,N_9643,N_11649);
and U13104 (N_13104,N_10755,N_8147);
nand U13105 (N_13105,N_10894,N_11157);
or U13106 (N_13106,N_9343,N_10690);
nand U13107 (N_13107,N_8918,N_8405);
or U13108 (N_13108,N_10397,N_10706);
nor U13109 (N_13109,N_11593,N_10983);
or U13110 (N_13110,N_10866,N_11035);
and U13111 (N_13111,N_9257,N_9157);
nand U13112 (N_13112,N_8909,N_8335);
nor U13113 (N_13113,N_8723,N_11981);
or U13114 (N_13114,N_11523,N_11713);
nor U13115 (N_13115,N_8852,N_9511);
or U13116 (N_13116,N_11251,N_11986);
nor U13117 (N_13117,N_10717,N_8810);
nand U13118 (N_13118,N_11793,N_8635);
or U13119 (N_13119,N_8544,N_9045);
and U13120 (N_13120,N_9127,N_10672);
nand U13121 (N_13121,N_11246,N_8016);
or U13122 (N_13122,N_8427,N_8625);
or U13123 (N_13123,N_10373,N_8851);
or U13124 (N_13124,N_10322,N_8619);
or U13125 (N_13125,N_9123,N_11952);
nand U13126 (N_13126,N_9455,N_10115);
and U13127 (N_13127,N_8306,N_10686);
or U13128 (N_13128,N_9480,N_10273);
nand U13129 (N_13129,N_11611,N_10281);
nor U13130 (N_13130,N_11704,N_8516);
nand U13131 (N_13131,N_9284,N_10486);
or U13132 (N_13132,N_8937,N_8251);
nand U13133 (N_13133,N_8184,N_10818);
nand U13134 (N_13134,N_10316,N_9589);
nand U13135 (N_13135,N_9318,N_8539);
or U13136 (N_13136,N_11937,N_11496);
and U13137 (N_13137,N_8097,N_9606);
or U13138 (N_13138,N_9264,N_8211);
or U13139 (N_13139,N_10962,N_10222);
xor U13140 (N_13140,N_11543,N_11247);
nor U13141 (N_13141,N_9792,N_11854);
nand U13142 (N_13142,N_11270,N_10854);
nor U13143 (N_13143,N_9573,N_10434);
or U13144 (N_13144,N_8825,N_11178);
or U13145 (N_13145,N_8651,N_8706);
nor U13146 (N_13146,N_8904,N_9437);
nand U13147 (N_13147,N_11453,N_10455);
and U13148 (N_13148,N_10205,N_9484);
nor U13149 (N_13149,N_11801,N_10406);
nand U13150 (N_13150,N_8831,N_10404);
and U13151 (N_13151,N_8827,N_8011);
nand U13152 (N_13152,N_9315,N_11228);
and U13153 (N_13153,N_11933,N_10259);
nor U13154 (N_13154,N_8910,N_10454);
and U13155 (N_13155,N_10213,N_10942);
xor U13156 (N_13156,N_8140,N_8664);
nand U13157 (N_13157,N_11972,N_10723);
or U13158 (N_13158,N_11755,N_9791);
nand U13159 (N_13159,N_9797,N_9095);
nor U13160 (N_13160,N_9936,N_8172);
and U13161 (N_13161,N_11502,N_11062);
or U13162 (N_13162,N_11664,N_11030);
and U13163 (N_13163,N_10085,N_8734);
nor U13164 (N_13164,N_8358,N_10488);
nand U13165 (N_13165,N_11860,N_8077);
nor U13166 (N_13166,N_10286,N_10697);
nand U13167 (N_13167,N_11738,N_11960);
nand U13168 (N_13168,N_8423,N_9186);
nand U13169 (N_13169,N_10341,N_10988);
nor U13170 (N_13170,N_11830,N_9543);
or U13171 (N_13171,N_11121,N_10788);
xnor U13172 (N_13172,N_10178,N_10744);
nor U13173 (N_13173,N_9276,N_9198);
nand U13174 (N_13174,N_11873,N_10372);
nor U13175 (N_13175,N_8353,N_9105);
or U13176 (N_13176,N_9035,N_10965);
nand U13177 (N_13177,N_10113,N_9463);
and U13178 (N_13178,N_10986,N_10083);
xor U13179 (N_13179,N_11721,N_10740);
or U13180 (N_13180,N_9382,N_10497);
nor U13181 (N_13181,N_9531,N_10646);
or U13182 (N_13182,N_10713,N_10644);
and U13183 (N_13183,N_10619,N_8790);
or U13184 (N_13184,N_10757,N_10004);
nor U13185 (N_13185,N_9866,N_11726);
and U13186 (N_13186,N_8469,N_8946);
nand U13187 (N_13187,N_11627,N_11182);
and U13188 (N_13188,N_10556,N_10521);
and U13189 (N_13189,N_11023,N_8684);
and U13190 (N_13190,N_8643,N_8418);
or U13191 (N_13191,N_9769,N_11729);
nand U13192 (N_13192,N_9392,N_8004);
or U13193 (N_13193,N_9170,N_11108);
and U13194 (N_13194,N_9031,N_10500);
nand U13195 (N_13195,N_11417,N_11606);
nand U13196 (N_13196,N_8747,N_9447);
xnor U13197 (N_13197,N_8853,N_10565);
and U13198 (N_13198,N_10783,N_9925);
or U13199 (N_13199,N_9713,N_9578);
or U13200 (N_13200,N_11824,N_10110);
nand U13201 (N_13201,N_8284,N_11778);
nor U13202 (N_13202,N_10698,N_10356);
and U13203 (N_13203,N_10677,N_11096);
nor U13204 (N_13204,N_9404,N_8673);
nand U13205 (N_13205,N_8080,N_10999);
nand U13206 (N_13206,N_11391,N_8369);
nand U13207 (N_13207,N_9996,N_11148);
nor U13208 (N_13208,N_8509,N_9030);
nand U13209 (N_13209,N_11308,N_10943);
nand U13210 (N_13210,N_10386,N_10732);
nand U13211 (N_13211,N_10182,N_8906);
and U13212 (N_13212,N_8895,N_8741);
xor U13213 (N_13213,N_8974,N_10155);
nand U13214 (N_13214,N_11039,N_9974);
nor U13215 (N_13215,N_8975,N_9886);
nor U13216 (N_13216,N_10116,N_11400);
nand U13217 (N_13217,N_9492,N_10858);
or U13218 (N_13218,N_8613,N_8967);
nor U13219 (N_13219,N_11995,N_9770);
xor U13220 (N_13220,N_10954,N_9732);
nor U13221 (N_13221,N_9538,N_8953);
or U13222 (N_13222,N_9026,N_10071);
and U13223 (N_13223,N_8641,N_11691);
or U13224 (N_13224,N_8685,N_9080);
or U13225 (N_13225,N_11199,N_11420);
nand U13226 (N_13226,N_9040,N_10324);
and U13227 (N_13227,N_9481,N_10347);
nand U13228 (N_13228,N_10562,N_8377);
nand U13229 (N_13229,N_9034,N_11261);
nor U13230 (N_13230,N_9700,N_10875);
and U13231 (N_13231,N_9600,N_11340);
and U13232 (N_13232,N_11318,N_9720);
nor U13233 (N_13233,N_10275,N_8206);
and U13234 (N_13234,N_10293,N_10491);
nor U13235 (N_13235,N_11329,N_11325);
nor U13236 (N_13236,N_10923,N_8845);
nand U13237 (N_13237,N_8563,N_9583);
and U13238 (N_13238,N_8973,N_11490);
or U13239 (N_13239,N_9843,N_10173);
nand U13240 (N_13240,N_8071,N_8204);
and U13241 (N_13241,N_8157,N_11661);
or U13242 (N_13242,N_10920,N_8523);
or U13243 (N_13243,N_9061,N_10833);
or U13244 (N_13244,N_10446,N_8873);
and U13245 (N_13245,N_9239,N_8384);
nand U13246 (N_13246,N_11897,N_10956);
or U13247 (N_13247,N_10023,N_11844);
nor U13248 (N_13248,N_8084,N_11558);
xnor U13249 (N_13249,N_8412,N_8091);
or U13250 (N_13250,N_11538,N_8310);
or U13251 (N_13251,N_8367,N_9949);
or U13252 (N_13252,N_9125,N_11701);
and U13253 (N_13253,N_9507,N_10768);
nor U13254 (N_13254,N_9002,N_8931);
and U13255 (N_13255,N_9709,N_11599);
xnor U13256 (N_13256,N_10570,N_8771);
and U13257 (N_13257,N_9562,N_11264);
nand U13258 (N_13258,N_9338,N_9418);
nor U13259 (N_13259,N_8465,N_8822);
and U13260 (N_13260,N_8758,N_11338);
nor U13261 (N_13261,N_8751,N_8462);
xnor U13262 (N_13262,N_9310,N_8811);
nand U13263 (N_13263,N_10803,N_9650);
nand U13264 (N_13264,N_8978,N_9498);
or U13265 (N_13265,N_11936,N_8290);
or U13266 (N_13266,N_9948,N_11840);
or U13267 (N_13267,N_11055,N_11819);
and U13268 (N_13268,N_10684,N_11891);
nand U13269 (N_13269,N_10907,N_11469);
or U13270 (N_13270,N_8329,N_9381);
or U13271 (N_13271,N_11594,N_9518);
or U13272 (N_13272,N_10873,N_8607);
xor U13273 (N_13273,N_9073,N_10728);
and U13274 (N_13274,N_9326,N_10856);
and U13275 (N_13275,N_8015,N_8308);
or U13276 (N_13276,N_9398,N_10805);
nand U13277 (N_13277,N_11847,N_9163);
nor U13278 (N_13278,N_9477,N_8286);
nand U13279 (N_13279,N_8393,N_9063);
xor U13280 (N_13280,N_9490,N_8144);
and U13281 (N_13281,N_11274,N_10396);
and U13282 (N_13282,N_10922,N_9884);
and U13283 (N_13283,N_8828,N_10533);
nor U13284 (N_13284,N_11306,N_10828);
or U13285 (N_13285,N_8074,N_11955);
and U13286 (N_13286,N_11043,N_8070);
and U13287 (N_13287,N_11472,N_11794);
or U13288 (N_13288,N_10088,N_8609);
nor U13289 (N_13289,N_9976,N_9227);
or U13290 (N_13290,N_10579,N_9814);
nand U13291 (N_13291,N_11539,N_8439);
or U13292 (N_13292,N_9374,N_8455);
xor U13293 (N_13293,N_9532,N_11279);
nor U13294 (N_13294,N_8429,N_11766);
nand U13295 (N_13295,N_10798,N_8507);
and U13296 (N_13296,N_9919,N_9218);
nor U13297 (N_13297,N_10883,N_10059);
nand U13298 (N_13298,N_11678,N_11887);
xor U13299 (N_13299,N_8676,N_9731);
nand U13300 (N_13300,N_9660,N_8240);
nand U13301 (N_13301,N_8966,N_11992);
nand U13302 (N_13302,N_9793,N_11849);
nand U13303 (N_13303,N_10447,N_11283);
xnor U13304 (N_13304,N_10725,N_11209);
xnor U13305 (N_13305,N_9609,N_9593);
nand U13306 (N_13306,N_11613,N_8680);
or U13307 (N_13307,N_11152,N_8554);
or U13308 (N_13308,N_8208,N_8043);
or U13309 (N_13309,N_9835,N_11032);
nor U13310 (N_13310,N_8603,N_9238);
nand U13311 (N_13311,N_11821,N_8319);
nor U13312 (N_13312,N_9588,N_10605);
and U13313 (N_13313,N_8558,N_11679);
and U13314 (N_13314,N_9613,N_10062);
nor U13315 (N_13315,N_9171,N_9856);
nor U13316 (N_13316,N_11290,N_11067);
nor U13317 (N_13317,N_10441,N_9629);
nor U13318 (N_13318,N_11667,N_9807);
nand U13319 (N_13319,N_11737,N_10464);
nor U13320 (N_13320,N_10210,N_10743);
or U13321 (N_13321,N_10542,N_10971);
nor U13322 (N_13322,N_11761,N_11643);
and U13323 (N_13323,N_9947,N_10465);
nand U13324 (N_13324,N_8867,N_9697);
or U13325 (N_13325,N_8594,N_9396);
and U13326 (N_13326,N_9817,N_11956);
or U13327 (N_13327,N_10254,N_9737);
and U13328 (N_13328,N_10652,N_8305);
nor U13329 (N_13329,N_8850,N_9848);
nand U13330 (N_13330,N_8672,N_11064);
and U13331 (N_13331,N_9901,N_8100);
and U13332 (N_13332,N_11212,N_8576);
nor U13333 (N_13333,N_11522,N_9348);
and U13334 (N_13334,N_11345,N_9241);
nand U13335 (N_13335,N_8115,N_9280);
nor U13336 (N_13336,N_11559,N_11549);
nor U13337 (N_13337,N_11730,N_8088);
and U13338 (N_13338,N_11916,N_10440);
nor U13339 (N_13339,N_8126,N_11672);
and U13340 (N_13340,N_8722,N_11770);
or U13341 (N_13341,N_10526,N_11173);
and U13342 (N_13342,N_9909,N_9081);
and U13343 (N_13343,N_11010,N_11843);
and U13344 (N_13344,N_11452,N_11997);
nand U13345 (N_13345,N_8236,N_8746);
xnor U13346 (N_13346,N_8056,N_10750);
nor U13347 (N_13347,N_10596,N_8678);
nor U13348 (N_13348,N_11406,N_8467);
and U13349 (N_13349,N_11303,N_9614);
nand U13350 (N_13350,N_8764,N_11138);
nor U13351 (N_13351,N_10812,N_9939);
nor U13352 (N_13352,N_9311,N_11694);
and U13353 (N_13353,N_8089,N_10492);
xnor U13354 (N_13354,N_8288,N_10306);
and U13355 (N_13355,N_11240,N_8171);
nand U13356 (N_13356,N_10416,N_9041);
nand U13357 (N_13357,N_9997,N_9386);
nand U13358 (N_13358,N_9395,N_8271);
and U13359 (N_13359,N_9577,N_10436);
and U13360 (N_13360,N_11584,N_9714);
and U13361 (N_13361,N_8832,N_9288);
nor U13362 (N_13362,N_8951,N_9813);
nor U13363 (N_13363,N_8858,N_10987);
nor U13364 (N_13364,N_9818,N_8454);
nor U13365 (N_13365,N_11725,N_11902);
and U13366 (N_13366,N_11630,N_8719);
nor U13367 (N_13367,N_11656,N_11354);
nor U13368 (N_13368,N_9409,N_11982);
and U13369 (N_13369,N_11925,N_9621);
or U13370 (N_13370,N_10877,N_11707);
nor U13371 (N_13371,N_8017,N_11470);
nor U13372 (N_13372,N_10346,N_10295);
nor U13373 (N_13373,N_10511,N_10014);
nor U13374 (N_13374,N_11016,N_10087);
nor U13375 (N_13375,N_8296,N_11932);
and U13376 (N_13376,N_11127,N_9891);
nor U13377 (N_13377,N_9999,N_10280);
nor U13378 (N_13378,N_8259,N_9331);
or U13379 (N_13379,N_8338,N_11987);
nand U13380 (N_13380,N_10329,N_10209);
and U13381 (N_13381,N_8905,N_9216);
and U13382 (N_13382,N_8601,N_8903);
and U13383 (N_13383,N_10013,N_10442);
nor U13384 (N_13384,N_8882,N_11705);
or U13385 (N_13385,N_11528,N_10865);
nor U13386 (N_13386,N_8266,N_9500);
nor U13387 (N_13387,N_8578,N_11382);
nor U13388 (N_13388,N_9189,N_11413);
nand U13389 (N_13389,N_10427,N_8224);
or U13390 (N_13390,N_8158,N_9622);
nor U13391 (N_13391,N_9010,N_11533);
or U13392 (N_13392,N_8808,N_9765);
and U13393 (N_13393,N_10419,N_11524);
or U13394 (N_13394,N_11405,N_9334);
or U13395 (N_13395,N_8616,N_8035);
or U13396 (N_13396,N_8857,N_10402);
and U13397 (N_13397,N_11757,N_8239);
or U13398 (N_13398,N_8442,N_9728);
nor U13399 (N_13399,N_9921,N_10136);
and U13400 (N_13400,N_9636,N_11380);
nor U13401 (N_13401,N_9036,N_9849);
and U13402 (N_13402,N_11038,N_9341);
and U13403 (N_13403,N_8460,N_10420);
nor U13404 (N_13404,N_11996,N_11771);
nor U13405 (N_13405,N_10552,N_9565);
xor U13406 (N_13406,N_11154,N_10429);
or U13407 (N_13407,N_11746,N_9464);
nand U13408 (N_13408,N_11497,N_8484);
nand U13409 (N_13409,N_9422,N_11786);
nand U13410 (N_13410,N_11360,N_11811);
nor U13411 (N_13411,N_10985,N_10638);
and U13412 (N_13412,N_8585,N_8215);
nand U13413 (N_13413,N_11980,N_8990);
nor U13414 (N_13414,N_11272,N_9428);
or U13415 (N_13415,N_8037,N_9897);
xnor U13416 (N_13416,N_8802,N_8440);
or U13417 (N_13417,N_8529,N_9000);
and U13418 (N_13418,N_8865,N_9851);
nand U13419 (N_13419,N_11122,N_10911);
and U13420 (N_13420,N_11312,N_9602);
or U13421 (N_13421,N_10587,N_11241);
nor U13422 (N_13422,N_8291,N_9904);
xnor U13423 (N_13423,N_8939,N_10846);
nor U13424 (N_13424,N_8892,N_10872);
nand U13425 (N_13425,N_8263,N_10008);
nor U13426 (N_13426,N_10204,N_8160);
nor U13427 (N_13427,N_10921,N_8886);
and U13428 (N_13428,N_11244,N_9796);
nor U13429 (N_13429,N_8782,N_9689);
nand U13430 (N_13430,N_9265,N_8217);
nor U13431 (N_13431,N_9258,N_11769);
or U13432 (N_13432,N_9225,N_8655);
or U13433 (N_13433,N_10695,N_9007);
nor U13434 (N_13434,N_8174,N_10976);
or U13435 (N_13435,N_8848,N_10076);
nor U13436 (N_13436,N_10625,N_9646);
or U13437 (N_13437,N_10438,N_11950);
nor U13438 (N_13438,N_10368,N_8486);
or U13439 (N_13439,N_9320,N_9782);
and U13440 (N_13440,N_9269,N_8797);
and U13441 (N_13441,N_8488,N_9911);
and U13442 (N_13442,N_10159,N_8428);
and U13443 (N_13443,N_8772,N_11676);
or U13444 (N_13444,N_10603,N_9118);
or U13445 (N_13445,N_10101,N_11332);
or U13446 (N_13446,N_10536,N_11618);
and U13447 (N_13447,N_10664,N_9991);
nor U13448 (N_13448,N_8515,N_10103);
nor U13449 (N_13449,N_11304,N_8330);
and U13450 (N_13450,N_10169,N_10337);
nand U13451 (N_13451,N_9093,N_11820);
or U13452 (N_13452,N_10657,N_11946);
nor U13453 (N_13453,N_10935,N_9874);
nor U13454 (N_13454,N_10642,N_10451);
and U13455 (N_13455,N_9129,N_11693);
nor U13456 (N_13456,N_8152,N_8021);
nand U13457 (N_13457,N_11146,N_10018);
nand U13458 (N_13458,N_10198,N_11751);
and U13459 (N_13459,N_11900,N_8101);
nor U13460 (N_13460,N_9859,N_8770);
or U13461 (N_13461,N_9347,N_8788);
nor U13462 (N_13462,N_9302,N_10460);
xor U13463 (N_13463,N_9564,N_10041);
or U13464 (N_13464,N_10234,N_8242);
nand U13465 (N_13465,N_9091,N_10344);
nand U13466 (N_13466,N_11215,N_9322);
nor U13467 (N_13467,N_11563,N_9740);
and U13468 (N_13468,N_9821,N_10153);
or U13469 (N_13469,N_8839,N_10231);
nand U13470 (N_13470,N_9021,N_9179);
and U13471 (N_13471,N_8943,N_10297);
nor U13472 (N_13472,N_11160,N_10722);
nor U13473 (N_13473,N_9205,N_8809);
nand U13474 (N_13474,N_11917,N_9530);
nor U13475 (N_13475,N_8637,N_11773);
and U13476 (N_13476,N_8805,N_9262);
and U13477 (N_13477,N_11425,N_9047);
and U13478 (N_13478,N_11505,N_10960);
and U13479 (N_13479,N_9072,N_8650);
or U13480 (N_13480,N_11077,N_10477);
or U13481 (N_13481,N_8945,N_9594);
or U13482 (N_13482,N_8781,N_11206);
nand U13483 (N_13483,N_8842,N_11269);
and U13484 (N_13484,N_10474,N_9828);
nand U13485 (N_13485,N_9383,N_11461);
and U13486 (N_13486,N_10959,N_8055);
nor U13487 (N_13487,N_10250,N_11890);
nor U13488 (N_13488,N_9248,N_8426);
nand U13489 (N_13489,N_9176,N_10314);
nor U13490 (N_13490,N_8360,N_8458);
or U13491 (N_13491,N_8474,N_11765);
or U13492 (N_13492,N_10957,N_8461);
and U13493 (N_13493,N_8012,N_8463);
and U13494 (N_13494,N_8687,N_8628);
and U13495 (N_13495,N_8944,N_8841);
nand U13496 (N_13496,N_8282,N_11403);
xor U13497 (N_13497,N_11670,N_8491);
and U13498 (N_13498,N_8225,N_8408);
and U13499 (N_13499,N_8876,N_11908);
nor U13500 (N_13500,N_9971,N_9523);
and U13501 (N_13501,N_11884,N_8395);
nand U13502 (N_13502,N_10520,N_9607);
nand U13503 (N_13503,N_11575,N_10472);
and U13504 (N_13504,N_8054,N_9357);
nand U13505 (N_13505,N_8120,N_11754);
nor U13506 (N_13506,N_10593,N_9285);
nand U13507 (N_13507,N_11586,N_8688);
nor U13508 (N_13508,N_9313,N_10094);
nor U13509 (N_13509,N_10135,N_8818);
nand U13510 (N_13510,N_11690,N_11158);
and U13511 (N_13511,N_9213,N_8612);
nor U13512 (N_13512,N_8487,N_10912);
xor U13513 (N_13513,N_9293,N_8166);
and U13514 (N_13514,N_11234,N_10061);
and U13515 (N_13515,N_10604,N_8446);
and U13516 (N_13516,N_10843,N_9902);
xnor U13517 (N_13517,N_10650,N_10065);
nand U13518 (N_13518,N_9462,N_8366);
nand U13519 (N_13519,N_8856,N_9540);
xor U13520 (N_13520,N_11165,N_9352);
and U13521 (N_13521,N_9024,N_9667);
nor U13522 (N_13522,N_8404,N_8430);
nand U13523 (N_13523,N_8424,N_10370);
nand U13524 (N_13524,N_10431,N_10063);
nor U13525 (N_13525,N_8318,N_9228);
or U13526 (N_13526,N_11284,N_10048);
nor U13527 (N_13527,N_9106,N_10848);
xnor U13528 (N_13528,N_9128,N_11527);
and U13529 (N_13529,N_11203,N_9587);
xnor U13530 (N_13530,N_11416,N_10513);
and U13531 (N_13531,N_9013,N_9762);
and U13532 (N_13532,N_9781,N_8663);
or U13533 (N_13533,N_11088,N_10927);
or U13534 (N_13534,N_11196,N_10127);
nor U13535 (N_13535,N_11367,N_11867);
and U13536 (N_13536,N_8961,N_11885);
nand U13537 (N_13537,N_9756,N_10655);
and U13538 (N_13538,N_9627,N_10645);
and U13539 (N_13539,N_9482,N_10735);
and U13540 (N_13540,N_9282,N_10105);
nand U13541 (N_13541,N_9380,N_11602);
and U13542 (N_13542,N_10498,N_9640);
or U13543 (N_13543,N_11889,N_11386);
and U13544 (N_13544,N_9222,N_10830);
nand U13545 (N_13545,N_11072,N_9166);
or U13546 (N_13546,N_11859,N_11945);
nor U13547 (N_13547,N_11109,N_10352);
and U13548 (N_13548,N_10218,N_8378);
nand U13549 (N_13549,N_11009,N_10383);
nand U13550 (N_13550,N_9083,N_9647);
and U13551 (N_13551,N_10388,N_9747);
or U13552 (N_13552,N_11192,N_11104);
nor U13553 (N_13553,N_9777,N_8262);
or U13554 (N_13554,N_10212,N_8737);
nand U13555 (N_13555,N_11651,N_10444);
nor U13556 (N_13556,N_11046,N_11311);
and U13557 (N_13557,N_8714,N_11791);
nor U13558 (N_13558,N_8557,N_11219);
nor U13559 (N_13559,N_8170,N_10479);
nor U13560 (N_13560,N_9772,N_11256);
and U13561 (N_13561,N_9555,N_9893);
nor U13562 (N_13562,N_11363,N_8611);
nand U13563 (N_13563,N_8131,N_10759);
or U13564 (N_13564,N_10417,N_11697);
nor U13565 (N_13565,N_10885,N_11501);
or U13566 (N_13566,N_10016,N_11886);
nor U13567 (N_13567,N_10508,N_8700);
and U13568 (N_13568,N_11321,N_8222);
nand U13569 (N_13569,N_10711,N_8748);
nor U13570 (N_13570,N_10167,N_8668);
nor U13571 (N_13571,N_8792,N_9018);
and U13572 (N_13572,N_11442,N_10659);
or U13573 (N_13573,N_11479,N_10709);
or U13574 (N_13574,N_8030,N_11495);
or U13575 (N_13575,N_11578,N_11698);
nor U13576 (N_13576,N_11979,N_10891);
or U13577 (N_13577,N_11953,N_10379);
or U13578 (N_13578,N_9151,N_10614);
nor U13579 (N_13579,N_11948,N_11652);
nor U13580 (N_13580,N_9065,N_11614);
and U13581 (N_13581,N_8407,N_8059);
xor U13582 (N_13582,N_10067,N_9657);
and U13583 (N_13583,N_11482,N_9752);
or U13584 (N_13584,N_8163,N_9255);
and U13585 (N_13585,N_9084,N_11623);
xnor U13586 (N_13586,N_10819,N_11033);
xnor U13587 (N_13587,N_8387,N_9503);
nand U13588 (N_13588,N_11069,N_8061);
nand U13589 (N_13589,N_9273,N_8599);
and U13590 (N_13590,N_10948,N_8665);
or U13591 (N_13591,N_8736,N_11568);
or U13592 (N_13592,N_8762,N_9193);
nand U13593 (N_13593,N_10084,N_8738);
nor U13594 (N_13594,N_10232,N_11313);
xnor U13595 (N_13595,N_9232,N_9953);
and U13596 (N_13596,N_9612,N_8735);
or U13597 (N_13597,N_11564,N_10251);
and U13598 (N_13598,N_11282,N_9165);
nand U13599 (N_13599,N_11059,N_9858);
or U13600 (N_13600,N_10633,N_9703);
nor U13601 (N_13601,N_11415,N_10790);
xor U13602 (N_13602,N_8249,N_10668);
and U13603 (N_13603,N_11213,N_11733);
and U13604 (N_13604,N_9423,N_9055);
or U13605 (N_13605,N_9678,N_11965);
and U13606 (N_13606,N_9610,N_11102);
xnor U13607 (N_13607,N_10595,N_8476);
nand U13608 (N_13608,N_11190,N_10531);
and U13609 (N_13609,N_10331,N_10111);
and U13610 (N_13610,N_8855,N_10039);
nor U13611 (N_13611,N_10279,N_9495);
nor U13612 (N_13612,N_10343,N_11636);
and U13613 (N_13613,N_10785,N_11390);
or U13614 (N_13614,N_11343,N_11774);
nand U13615 (N_13615,N_11927,N_8036);
and U13616 (N_13616,N_9620,N_8315);
or U13617 (N_13617,N_9056,N_9778);
or U13618 (N_13618,N_11107,N_8139);
or U13619 (N_13619,N_11825,N_11226);
or U13620 (N_13620,N_11585,N_8598);
xnor U13621 (N_13621,N_11342,N_8022);
nand U13622 (N_13622,N_10597,N_8039);
xor U13623 (N_13623,N_9367,N_9033);
and U13624 (N_13624,N_9820,N_8527);
xor U13625 (N_13625,N_8708,N_10335);
nand U13626 (N_13626,N_11162,N_9268);
or U13627 (N_13627,N_9299,N_10158);
nand U13628 (N_13628,N_8548,N_10422);
and U13629 (N_13629,N_9668,N_11772);
or U13630 (N_13630,N_11005,N_11532);
nand U13631 (N_13631,N_9256,N_11185);
nand U13632 (N_13632,N_10961,N_9094);
or U13633 (N_13633,N_8749,N_9363);
nand U13634 (N_13634,N_9883,N_9336);
or U13635 (N_13635,N_11716,N_9090);
nor U13636 (N_13636,N_11464,N_8504);
nor U13637 (N_13637,N_10448,N_9312);
xor U13638 (N_13638,N_8420,N_11530);
or U13639 (N_13639,N_10658,N_10349);
and U13640 (N_13640,N_8731,N_11348);
and U13641 (N_13641,N_9441,N_8034);
and U13642 (N_13642,N_11517,N_8879);
and U13643 (N_13643,N_9645,N_8165);
nand U13644 (N_13644,N_11597,N_8887);
nor U13645 (N_13645,N_10495,N_10992);
xor U13646 (N_13646,N_9250,N_11068);
and U13647 (N_13647,N_10834,N_9918);
or U13648 (N_13648,N_8000,N_9670);
nand U13649 (N_13649,N_11852,N_8701);
nand U13650 (N_13650,N_9863,N_10055);
or U13651 (N_13651,N_10036,N_8297);
nor U13652 (N_13652,N_11983,N_10940);
or U13653 (N_13653,N_8368,N_11278);
or U13654 (N_13654,N_8063,N_8410);
or U13655 (N_13655,N_11128,N_9314);
or U13656 (N_13656,N_10494,N_11872);
nor U13657 (N_13657,N_8506,N_9924);
nand U13658 (N_13658,N_8588,N_11736);
xor U13659 (N_13659,N_11120,N_8314);
nand U13660 (N_13660,N_8846,N_8414);
xor U13661 (N_13661,N_9682,N_9537);
xor U13662 (N_13662,N_8185,N_10200);
or U13663 (N_13663,N_9220,N_10576);
and U13664 (N_13664,N_8502,N_9699);
and U13665 (N_13665,N_9192,N_9413);
or U13666 (N_13666,N_8072,N_9360);
or U13667 (N_13667,N_10632,N_8227);
xor U13668 (N_13668,N_8295,N_11431);
and U13669 (N_13669,N_9122,N_8106);
nand U13670 (N_13670,N_8993,N_11668);
xor U13671 (N_13671,N_11346,N_11135);
nand U13672 (N_13672,N_10636,N_8373);
nor U13673 (N_13673,N_9251,N_8336);
nand U13674 (N_13674,N_9899,N_8494);
nand U13675 (N_13675,N_8198,N_10199);
nor U13676 (N_13676,N_9240,N_10889);
nand U13677 (N_13677,N_11205,N_8501);
and U13678 (N_13678,N_11812,N_10365);
or U13679 (N_13679,N_9022,N_10450);
xor U13680 (N_13680,N_9235,N_11268);
xnor U13681 (N_13681,N_10890,N_9598);
or U13682 (N_13682,N_9705,N_9766);
nor U13683 (N_13683,N_8889,N_8182);
and U13684 (N_13684,N_10128,N_9425);
nor U13685 (N_13685,N_10020,N_9145);
or U13686 (N_13686,N_11646,N_11822);
or U13687 (N_13687,N_10574,N_11319);
or U13688 (N_13688,N_9847,N_8441);
nor U13689 (N_13689,N_8257,N_10108);
nand U13690 (N_13690,N_8566,N_9864);
or U13691 (N_13691,N_8900,N_10481);
and U13692 (N_13692,N_10239,N_8230);
and U13693 (N_13693,N_9695,N_9872);
nor U13694 (N_13694,N_9704,N_11954);
or U13695 (N_13695,N_11720,N_8051);
and U13696 (N_13696,N_10937,N_8837);
and U13697 (N_13697,N_9934,N_11455);
and U13698 (N_13698,N_9120,N_11193);
nor U13699 (N_13699,N_8396,N_9107);
nor U13700 (N_13700,N_11404,N_10086);
or U13701 (N_13701,N_8138,N_10364);
or U13702 (N_13702,N_9438,N_11371);
or U13703 (N_13703,N_10553,N_11006);
or U13704 (N_13704,N_8789,N_8466);
and U13705 (N_13705,N_8173,N_10660);
xor U13706 (N_13706,N_9458,N_11930);
and U13707 (N_13707,N_10471,N_11655);
nand U13708 (N_13708,N_8644,N_8337);
nor U13709 (N_13709,N_11507,N_11700);
xor U13710 (N_13710,N_10944,N_10045);
and U13711 (N_13711,N_9585,N_10366);
nor U13712 (N_13712,N_9963,N_11474);
nor U13713 (N_13713,N_9297,N_11150);
and U13714 (N_13714,N_11628,N_10030);
or U13715 (N_13715,N_8877,N_8304);
or U13716 (N_13716,N_9675,N_8234);
nor U13717 (N_13717,N_11087,N_10563);
and U13718 (N_13718,N_10371,N_10052);
or U13719 (N_13719,N_10639,N_11218);
and U13720 (N_13720,N_9152,N_8602);
or U13721 (N_13721,N_8298,N_11141);
or U13722 (N_13722,N_9742,N_8028);
or U13723 (N_13723,N_8935,N_10102);
or U13724 (N_13724,N_10452,N_9470);
nor U13725 (N_13725,N_9410,N_10327);
or U13726 (N_13726,N_10924,N_9776);
and U13727 (N_13727,N_10775,N_10006);
or U13728 (N_13728,N_11923,N_8984);
or U13729 (N_13729,N_9201,N_10881);
nand U13730 (N_13730,N_11905,N_9794);
nor U13731 (N_13731,N_11813,N_9440);
and U13732 (N_13732,N_11868,N_8897);
or U13733 (N_13733,N_10400,N_9242);
nor U13734 (N_13734,N_8018,N_9514);
nand U13735 (N_13735,N_8874,N_9506);
and U13736 (N_13736,N_9144,N_10047);
or U13737 (N_13737,N_8168,N_9444);
or U13738 (N_13738,N_9502,N_11204);
nand U13739 (N_13739,N_9604,N_11230);
or U13740 (N_13740,N_8009,N_9654);
nor U13741 (N_13741,N_10392,N_8075);
nor U13742 (N_13742,N_10411,N_8096);
or U13743 (N_13743,N_11292,N_11249);
nor U13744 (N_13744,N_10469,N_11856);
and U13745 (N_13745,N_10382,N_8040);
or U13746 (N_13746,N_10815,N_9245);
and U13747 (N_13747,N_11727,N_8679);
or U13748 (N_13748,N_8763,N_8361);
and U13749 (N_13749,N_8268,N_11149);
nor U13750 (N_13750,N_10389,N_8948);
nand U13751 (N_13751,N_8274,N_8053);
nor U13752 (N_13752,N_11118,N_10578);
or U13753 (N_13753,N_8838,N_9429);
or U13754 (N_13754,N_11336,N_8076);
or U13755 (N_13755,N_10929,N_9890);
nor U13756 (N_13756,N_11722,N_11115);
and U13757 (N_13757,N_9407,N_9023);
xnor U13758 (N_13758,N_11512,N_11572);
nand U13759 (N_13759,N_8193,N_10860);
or U13760 (N_13760,N_8775,N_8894);
xor U13761 (N_13761,N_11949,N_8200);
or U13762 (N_13762,N_8547,N_11444);
or U13763 (N_13763,N_8683,N_9066);
or U13764 (N_13764,N_10635,N_9384);
nand U13765 (N_13765,N_8307,N_11169);
and U13766 (N_13766,N_11569,N_9512);
nand U13767 (N_13767,N_11028,N_8732);
and U13768 (N_13768,N_9746,N_11368);
nand U13769 (N_13769,N_10375,N_10769);
nor U13770 (N_13770,N_8985,N_8162);
nand U13771 (N_13771,N_11070,N_9333);
nand U13772 (N_13772,N_9723,N_11629);
and U13773 (N_13773,N_8196,N_8798);
or U13774 (N_13774,N_10359,N_8854);
nand U13775 (N_13775,N_9937,N_9908);
nor U13776 (N_13776,N_10649,N_8005);
nand U13777 (N_13777,N_8791,N_8560);
and U13778 (N_13778,N_11436,N_9116);
and U13779 (N_13779,N_8482,N_10269);
nand U13780 (N_13780,N_10780,N_8902);
and U13781 (N_13781,N_11462,N_10131);
nor U13782 (N_13782,N_8914,N_8536);
nand U13783 (N_13783,N_11159,N_11776);
xor U13784 (N_13784,N_9028,N_9559);
nor U13785 (N_13785,N_10773,N_11427);
xor U13786 (N_13786,N_8872,N_11951);
nor U13787 (N_13787,N_11998,N_9734);
or U13788 (N_13788,N_10817,N_10489);
or U13789 (N_13789,N_10283,N_9571);
nor U13790 (N_13790,N_8065,N_9749);
and U13791 (N_13791,N_8804,N_10751);
or U13792 (N_13792,N_11787,N_11647);
nand U13793 (N_13793,N_9544,N_8955);
and U13794 (N_13794,N_11827,N_8128);
or U13795 (N_13795,N_9279,N_9133);
xor U13796 (N_13796,N_8580,N_9628);
or U13797 (N_13797,N_8958,N_11334);
xor U13798 (N_13798,N_10909,N_8380);
and U13799 (N_13799,N_11894,N_8710);
and U13800 (N_13800,N_10423,N_9253);
nand U13801 (N_13801,N_8600,N_10353);
and U13802 (N_13802,N_8777,N_10748);
and U13803 (N_13803,N_11814,N_8551);
or U13804 (N_13804,N_10300,N_8485);
nor U13805 (N_13805,N_10699,N_10746);
or U13806 (N_13806,N_10188,N_11969);
nand U13807 (N_13807,N_8492,N_8721);
and U13808 (N_13808,N_8674,N_10953);
or U13809 (N_13809,N_11634,N_11580);
nand U13810 (N_13810,N_8489,N_8543);
nand U13811 (N_13811,N_11467,N_9270);
and U13812 (N_13812,N_8087,N_11101);
or U13813 (N_13813,N_8057,N_11508);
nand U13814 (N_13814,N_11398,N_11658);
nor U13815 (N_13815,N_10070,N_8756);
nand U13816 (N_13816,N_8959,N_11223);
nand U13817 (N_13817,N_8479,N_10276);
nand U13818 (N_13818,N_9576,N_9468);
nor U13819 (N_13819,N_8617,N_10509);
and U13820 (N_13820,N_8459,N_9278);
or U13821 (N_13821,N_10874,N_11220);
nor U13822 (N_13822,N_9478,N_10058);
nand U13823 (N_13823,N_9946,N_8840);
nor U13824 (N_13824,N_11044,N_9412);
or U13825 (N_13825,N_9726,N_9138);
nand U13826 (N_13826,N_10726,N_9003);
or U13827 (N_13827,N_11281,N_10289);
and U13828 (N_13828,N_10345,N_11327);
xnor U13829 (N_13829,N_10144,N_11243);
nand U13830 (N_13830,N_8250,N_9819);
and U13831 (N_13831,N_10129,N_11106);
nor U13832 (N_13832,N_11002,N_9972);
nor U13833 (N_13833,N_11387,N_10975);
nand U13834 (N_13834,N_8901,N_9476);
or U13835 (N_13835,N_10137,N_9790);
nand U13836 (N_13836,N_11011,N_11012);
nor U13837 (N_13837,N_8919,N_9390);
nor U13838 (N_13838,N_10149,N_10807);
nor U13839 (N_13839,N_10716,N_10982);
nor U13840 (N_13840,N_11566,N_10168);
nand U13841 (N_13841,N_11471,N_10148);
and U13842 (N_13842,N_11414,N_9735);
nor U13843 (N_13843,N_10394,N_11328);
xnor U13844 (N_13844,N_10532,N_9748);
and U13845 (N_13845,N_10977,N_11052);
or U13846 (N_13846,N_9712,N_11200);
and U13847 (N_13847,N_11166,N_11711);
nor U13848 (N_13848,N_9388,N_8169);
nor U13849 (N_13849,N_10832,N_10317);
nand U13850 (N_13850,N_11895,N_10177);
or U13851 (N_13851,N_11555,N_10795);
nand U13852 (N_13852,N_10640,N_9554);
or U13853 (N_13853,N_8869,N_9786);
and U13854 (N_13854,N_9674,N_8354);
nor U13855 (N_13855,N_11275,N_10691);
nand U13856 (N_13856,N_10320,N_9281);
nand U13857 (N_13857,N_11000,N_9112);
nand U13858 (N_13858,N_9489,N_8029);
nor U13859 (N_13859,N_10517,N_11876);
or U13860 (N_13860,N_10878,N_10415);
and U13861 (N_13861,N_10947,N_11536);
nor U13862 (N_13862,N_8864,N_9721);
nand U13863 (N_13863,N_8704,N_8880);
xnor U13864 (N_13864,N_11931,N_11258);
and U13865 (N_13865,N_11994,N_11448);
nor U13866 (N_13866,N_11238,N_11695);
and U13867 (N_13867,N_9291,N_9521);
or U13868 (N_13868,N_10900,N_8888);
xor U13869 (N_13869,N_8276,N_8261);
nand U13870 (N_13870,N_8586,N_8445);
xor U13871 (N_13871,N_9940,N_11116);
nand U13872 (N_13872,N_8669,N_11309);
nor U13873 (N_13873,N_9126,N_9210);
nand U13874 (N_13874,N_10895,N_8917);
nand U13875 (N_13875,N_10203,N_10456);
nand U13876 (N_13876,N_10017,N_9956);
xnor U13877 (N_13877,N_9533,N_10575);
nor U13878 (N_13878,N_11839,N_8136);
and U13879 (N_13879,N_11624,N_8691);
or U13880 (N_13880,N_8448,N_8671);
and U13881 (N_13881,N_9071,N_10146);
nand U13882 (N_13882,N_8666,N_10719);
nor U13883 (N_13883,N_10767,N_10673);
nor U13884 (N_13884,N_10949,N_10226);
nor U13885 (N_13885,N_10588,N_11978);
xnor U13886 (N_13886,N_10355,N_10208);
or U13887 (N_13887,N_8214,N_11789);
nand U13888 (N_13888,N_9887,N_8422);
nor U13889 (N_13889,N_11803,N_10266);
nor U13890 (N_13890,N_10246,N_8108);
or U13891 (N_13891,N_8390,N_10731);
nand U13892 (N_13892,N_9221,N_11846);
nand U13893 (N_13893,N_11210,N_10577);
nand U13894 (N_13894,N_11050,N_10688);
and U13895 (N_13895,N_9941,N_10968);
nand U13896 (N_13896,N_9517,N_11582);
and U13897 (N_13897,N_8062,N_9345);
nand U13898 (N_13898,N_10302,N_10139);
and U13899 (N_13899,N_9527,N_8472);
and U13900 (N_13900,N_10820,N_11310);
and U13901 (N_13901,N_8972,N_11248);
nor U13902 (N_13902,N_8618,N_11603);
nand U13903 (N_13903,N_8450,N_8596);
nor U13904 (N_13904,N_11027,N_9141);
nor U13905 (N_13905,N_10219,N_8416);
and U13906 (N_13906,N_9079,N_8829);
xnor U13907 (N_13907,N_11571,N_9855);
nor U13908 (N_13908,N_8081,N_9568);
nand U13909 (N_13909,N_9130,N_9450);
or U13910 (N_13910,N_11184,N_9524);
and U13911 (N_13911,N_8623,N_11143);
nor U13912 (N_13912,N_11266,N_10779);
nand U13913 (N_13913,N_10934,N_10010);
xor U13914 (N_13914,N_9070,N_11899);
nor U13915 (N_13915,N_9156,N_11988);
or U13916 (N_13916,N_11491,N_9952);
and U13917 (N_13917,N_9342,N_9119);
and U13918 (N_13918,N_10863,N_10407);
nor U13919 (N_13919,N_9362,N_8927);
or U13920 (N_13920,N_9833,N_10142);
or U13921 (N_13921,N_10904,N_10701);
and U13922 (N_13922,N_11806,N_9880);
and U13923 (N_13923,N_8066,N_8457);
and U13924 (N_13924,N_11942,N_9267);
nand U13925 (N_13925,N_9321,N_8522);
or U13926 (N_13926,N_10522,N_11790);
xnor U13927 (N_13927,N_11478,N_8510);
nand U13928 (N_13928,N_10363,N_11758);
and U13929 (N_13929,N_10134,N_11644);
nor U13930 (N_13930,N_11869,N_10665);
nor U13931 (N_13931,N_10312,N_8924);
and U13932 (N_13932,N_8907,N_9960);
nand U13933 (N_13933,N_11322,N_11299);
nor U13934 (N_13934,N_10886,N_8610);
and U13935 (N_13935,N_9399,N_11706);
or U13936 (N_13936,N_9877,N_9870);
or U13937 (N_13937,N_8452,N_11688);
or U13938 (N_13938,N_8645,N_9677);
nand U13939 (N_13939,N_8473,N_11029);
and U13940 (N_13940,N_10462,N_11333);
and U13941 (N_13941,N_9671,N_9832);
nor U13942 (N_13942,N_8164,N_9190);
or U13943 (N_13943,N_9113,N_9400);
nand U13944 (N_13944,N_8401,N_10410);
nand U13945 (N_13945,N_9174,N_8962);
or U13946 (N_13946,N_9836,N_10193);
xor U13947 (N_13947,N_9137,N_8447);
nand U13948 (N_13948,N_8711,N_8344);
nor U13949 (N_13949,N_8313,N_10867);
nor U13950 (N_13950,N_9254,N_10908);
and U13951 (N_13951,N_9042,N_8112);
nand U13952 (N_13952,N_9335,N_10328);
nand U13953 (N_13953,N_11671,N_8349);
xnor U13954 (N_13954,N_11684,N_10034);
xnor U13955 (N_13955,N_8328,N_8768);
and U13956 (N_13956,N_8994,N_9516);
or U13957 (N_13957,N_9316,N_11145);
nand U13958 (N_13958,N_8534,N_11648);
nor U13959 (N_13959,N_11298,N_8123);
nand U13960 (N_13960,N_9207,N_9465);
xnor U13961 (N_13961,N_9229,N_8528);
nor U13962 (N_13962,N_11378,N_8019);
and U13963 (N_13963,N_8686,N_11080);
and U13964 (N_13964,N_9649,N_11326);
or U13965 (N_13965,N_10515,N_9917);
nor U13966 (N_13966,N_8229,N_10493);
and U13967 (N_13967,N_11760,N_9044);
xor U13968 (N_13968,N_9804,N_10252);
and U13969 (N_13969,N_8449,N_10079);
and U13970 (N_13970,N_9309,N_9658);
nor U13971 (N_13971,N_10897,N_8099);
nand U13972 (N_13972,N_10584,N_8444);
or U13973 (N_13973,N_11477,N_10211);
or U13974 (N_13974,N_8774,N_11763);
or U13975 (N_13975,N_8654,N_10015);
nor U13976 (N_13976,N_9702,N_9087);
nand U13977 (N_13977,N_10308,N_8232);
or U13978 (N_13978,N_10774,N_11040);
nor U13979 (N_13979,N_11276,N_8550);
and U13980 (N_13980,N_11394,N_11437);
nand U13981 (N_13981,N_8987,N_11443);
or U13982 (N_13982,N_10782,N_10741);
nor U13983 (N_13983,N_8341,N_8086);
or U13984 (N_13984,N_11105,N_11171);
and U13985 (N_13985,N_10263,N_8922);
or U13986 (N_13986,N_8109,N_10357);
nand U13987 (N_13987,N_10651,N_10936);
or U13988 (N_13988,N_10623,N_10191);
nand U13989 (N_13989,N_9180,N_10189);
nand U13990 (N_13990,N_11703,N_8415);
and U13991 (N_13991,N_11749,N_11500);
and U13992 (N_13992,N_8835,N_10292);
and U13993 (N_13993,N_8434,N_8755);
xor U13994 (N_13994,N_9745,N_9525);
nor U13995 (N_13995,N_11305,N_11609);
nor U13996 (N_13996,N_8545,N_8052);
or U13997 (N_13997,N_9632,N_10766);
and U13998 (N_13998,N_10548,N_11401);
or U13999 (N_13999,N_9551,N_11095);
and U14000 (N_14000,N_9864,N_8422);
or U14001 (N_14001,N_11400,N_9490);
or U14002 (N_14002,N_10433,N_11407);
and U14003 (N_14003,N_10458,N_11404);
nand U14004 (N_14004,N_10547,N_8389);
or U14005 (N_14005,N_9924,N_8322);
and U14006 (N_14006,N_10352,N_10374);
nor U14007 (N_14007,N_10805,N_9659);
xnor U14008 (N_14008,N_9707,N_10226);
nand U14009 (N_14009,N_11906,N_9013);
and U14010 (N_14010,N_10060,N_8940);
and U14011 (N_14011,N_8132,N_11504);
and U14012 (N_14012,N_9076,N_10743);
nand U14013 (N_14013,N_11792,N_9038);
nand U14014 (N_14014,N_9548,N_8282);
nand U14015 (N_14015,N_9855,N_9040);
or U14016 (N_14016,N_9624,N_9947);
nor U14017 (N_14017,N_8201,N_8591);
xnor U14018 (N_14018,N_9917,N_10206);
xor U14019 (N_14019,N_10063,N_8226);
and U14020 (N_14020,N_9196,N_9120);
xor U14021 (N_14021,N_9827,N_11406);
and U14022 (N_14022,N_11037,N_11692);
and U14023 (N_14023,N_10786,N_11337);
nor U14024 (N_14024,N_11239,N_9262);
nand U14025 (N_14025,N_11149,N_8168);
and U14026 (N_14026,N_11263,N_10892);
nor U14027 (N_14027,N_9783,N_11594);
and U14028 (N_14028,N_9820,N_11846);
nand U14029 (N_14029,N_11396,N_9051);
xnor U14030 (N_14030,N_9694,N_10836);
xnor U14031 (N_14031,N_8007,N_9378);
nand U14032 (N_14032,N_8511,N_9460);
or U14033 (N_14033,N_8049,N_10251);
nor U14034 (N_14034,N_10791,N_8865);
xnor U14035 (N_14035,N_11763,N_10947);
or U14036 (N_14036,N_9777,N_10112);
or U14037 (N_14037,N_9477,N_9552);
and U14038 (N_14038,N_11825,N_9593);
xor U14039 (N_14039,N_8311,N_10923);
nand U14040 (N_14040,N_11669,N_8147);
and U14041 (N_14041,N_8943,N_11249);
nand U14042 (N_14042,N_8982,N_10981);
xnor U14043 (N_14043,N_11554,N_8451);
nor U14044 (N_14044,N_10072,N_10031);
xor U14045 (N_14045,N_8549,N_10552);
nand U14046 (N_14046,N_9087,N_10976);
nor U14047 (N_14047,N_9532,N_9089);
nand U14048 (N_14048,N_8603,N_8847);
nor U14049 (N_14049,N_11833,N_11534);
and U14050 (N_14050,N_9568,N_11101);
or U14051 (N_14051,N_11141,N_8312);
and U14052 (N_14052,N_8634,N_8718);
and U14053 (N_14053,N_9278,N_8221);
or U14054 (N_14054,N_11332,N_11725);
and U14055 (N_14055,N_10268,N_11509);
nor U14056 (N_14056,N_9591,N_9619);
or U14057 (N_14057,N_9544,N_9087);
nand U14058 (N_14058,N_11347,N_11051);
nand U14059 (N_14059,N_11237,N_10018);
and U14060 (N_14060,N_10132,N_9636);
or U14061 (N_14061,N_10610,N_10076);
nor U14062 (N_14062,N_11422,N_10887);
xnor U14063 (N_14063,N_10205,N_11683);
and U14064 (N_14064,N_11343,N_10908);
or U14065 (N_14065,N_9691,N_11620);
nand U14066 (N_14066,N_8078,N_10335);
and U14067 (N_14067,N_11591,N_8666);
nor U14068 (N_14068,N_9925,N_9526);
or U14069 (N_14069,N_9872,N_9618);
nand U14070 (N_14070,N_10662,N_8808);
or U14071 (N_14071,N_8778,N_11231);
xor U14072 (N_14072,N_9408,N_9833);
nor U14073 (N_14073,N_8304,N_9346);
nor U14074 (N_14074,N_8962,N_11466);
nor U14075 (N_14075,N_8339,N_9230);
xnor U14076 (N_14076,N_8368,N_10735);
or U14077 (N_14077,N_8712,N_11290);
and U14078 (N_14078,N_9744,N_8415);
nand U14079 (N_14079,N_11710,N_8251);
nand U14080 (N_14080,N_8703,N_9806);
or U14081 (N_14081,N_9960,N_9566);
or U14082 (N_14082,N_10105,N_11193);
or U14083 (N_14083,N_8839,N_9330);
or U14084 (N_14084,N_10732,N_9336);
or U14085 (N_14085,N_10875,N_10724);
or U14086 (N_14086,N_11283,N_9204);
and U14087 (N_14087,N_8058,N_9549);
nand U14088 (N_14088,N_9104,N_8142);
nand U14089 (N_14089,N_9121,N_10661);
nor U14090 (N_14090,N_11411,N_10880);
and U14091 (N_14091,N_9314,N_8835);
nor U14092 (N_14092,N_11439,N_11596);
or U14093 (N_14093,N_9901,N_8901);
or U14094 (N_14094,N_8319,N_9904);
xnor U14095 (N_14095,N_11233,N_8078);
nor U14096 (N_14096,N_8385,N_8207);
nand U14097 (N_14097,N_9268,N_11219);
xnor U14098 (N_14098,N_9496,N_8297);
and U14099 (N_14099,N_11972,N_10202);
nand U14100 (N_14100,N_10760,N_11411);
nor U14101 (N_14101,N_11376,N_10399);
nand U14102 (N_14102,N_11789,N_9456);
or U14103 (N_14103,N_8830,N_9189);
nor U14104 (N_14104,N_9600,N_8397);
and U14105 (N_14105,N_10171,N_10687);
nand U14106 (N_14106,N_10177,N_11740);
xor U14107 (N_14107,N_11031,N_9297);
nand U14108 (N_14108,N_8209,N_11958);
or U14109 (N_14109,N_9698,N_8144);
nand U14110 (N_14110,N_8134,N_9665);
xnor U14111 (N_14111,N_11112,N_10765);
and U14112 (N_14112,N_11877,N_10169);
or U14113 (N_14113,N_8139,N_11269);
or U14114 (N_14114,N_8067,N_9191);
nand U14115 (N_14115,N_11979,N_11579);
and U14116 (N_14116,N_11470,N_8157);
nand U14117 (N_14117,N_8984,N_9703);
nor U14118 (N_14118,N_11140,N_9645);
or U14119 (N_14119,N_11352,N_9744);
and U14120 (N_14120,N_10111,N_8834);
xnor U14121 (N_14121,N_10512,N_10552);
nand U14122 (N_14122,N_9840,N_8331);
and U14123 (N_14123,N_9528,N_10099);
nand U14124 (N_14124,N_10581,N_9296);
or U14125 (N_14125,N_11174,N_10423);
or U14126 (N_14126,N_10743,N_8242);
or U14127 (N_14127,N_8651,N_8508);
and U14128 (N_14128,N_11916,N_9919);
xor U14129 (N_14129,N_8458,N_9456);
and U14130 (N_14130,N_11267,N_9898);
nor U14131 (N_14131,N_9788,N_9646);
and U14132 (N_14132,N_11748,N_8526);
nand U14133 (N_14133,N_11140,N_8478);
or U14134 (N_14134,N_9998,N_8160);
nor U14135 (N_14135,N_9245,N_10603);
or U14136 (N_14136,N_8555,N_9136);
nand U14137 (N_14137,N_10829,N_9631);
nor U14138 (N_14138,N_9357,N_10869);
nand U14139 (N_14139,N_9670,N_9154);
and U14140 (N_14140,N_10588,N_11931);
nand U14141 (N_14141,N_9282,N_10234);
and U14142 (N_14142,N_10966,N_11114);
nor U14143 (N_14143,N_10869,N_8429);
or U14144 (N_14144,N_10234,N_9319);
nand U14145 (N_14145,N_9157,N_8369);
or U14146 (N_14146,N_10243,N_8394);
nand U14147 (N_14147,N_8438,N_10832);
or U14148 (N_14148,N_9007,N_9388);
and U14149 (N_14149,N_8536,N_10104);
or U14150 (N_14150,N_9356,N_10443);
and U14151 (N_14151,N_8403,N_8054);
and U14152 (N_14152,N_8787,N_11131);
nand U14153 (N_14153,N_10963,N_9751);
nand U14154 (N_14154,N_9130,N_11342);
or U14155 (N_14155,N_11179,N_10791);
and U14156 (N_14156,N_11702,N_11593);
nand U14157 (N_14157,N_8473,N_11633);
or U14158 (N_14158,N_10935,N_10330);
or U14159 (N_14159,N_9376,N_9910);
nor U14160 (N_14160,N_11070,N_9417);
xnor U14161 (N_14161,N_8981,N_9004);
nand U14162 (N_14162,N_8461,N_9601);
nand U14163 (N_14163,N_10874,N_9005);
or U14164 (N_14164,N_9579,N_8365);
nand U14165 (N_14165,N_9741,N_11899);
and U14166 (N_14166,N_9083,N_9175);
and U14167 (N_14167,N_9888,N_10652);
or U14168 (N_14168,N_9568,N_9901);
and U14169 (N_14169,N_11317,N_8299);
nor U14170 (N_14170,N_11613,N_10296);
or U14171 (N_14171,N_11529,N_8580);
nand U14172 (N_14172,N_11636,N_8157);
nand U14173 (N_14173,N_9538,N_11576);
or U14174 (N_14174,N_11739,N_11199);
and U14175 (N_14175,N_9774,N_10021);
xor U14176 (N_14176,N_8613,N_9322);
or U14177 (N_14177,N_10413,N_10221);
nor U14178 (N_14178,N_10234,N_10975);
xnor U14179 (N_14179,N_8002,N_9959);
nand U14180 (N_14180,N_8897,N_9671);
nor U14181 (N_14181,N_8561,N_10720);
and U14182 (N_14182,N_9721,N_11366);
nand U14183 (N_14183,N_8113,N_8551);
or U14184 (N_14184,N_11767,N_8663);
nand U14185 (N_14185,N_11636,N_11009);
nor U14186 (N_14186,N_10335,N_8472);
nand U14187 (N_14187,N_9306,N_8168);
xor U14188 (N_14188,N_11358,N_11299);
and U14189 (N_14189,N_11137,N_8427);
nor U14190 (N_14190,N_8768,N_11663);
and U14191 (N_14191,N_8921,N_9111);
nor U14192 (N_14192,N_9476,N_9329);
nor U14193 (N_14193,N_10244,N_9290);
or U14194 (N_14194,N_10047,N_11987);
nand U14195 (N_14195,N_8181,N_9483);
and U14196 (N_14196,N_9196,N_11093);
or U14197 (N_14197,N_9018,N_8623);
or U14198 (N_14198,N_10693,N_9047);
or U14199 (N_14199,N_9383,N_10561);
xor U14200 (N_14200,N_9129,N_9446);
nor U14201 (N_14201,N_11734,N_8200);
nor U14202 (N_14202,N_10158,N_10125);
xnor U14203 (N_14203,N_10786,N_10123);
nand U14204 (N_14204,N_9461,N_8683);
or U14205 (N_14205,N_9697,N_10151);
nand U14206 (N_14206,N_9556,N_11718);
and U14207 (N_14207,N_9021,N_10550);
and U14208 (N_14208,N_11217,N_11124);
nand U14209 (N_14209,N_9538,N_10451);
nand U14210 (N_14210,N_8655,N_9194);
nor U14211 (N_14211,N_9415,N_10402);
xnor U14212 (N_14212,N_11695,N_11030);
nand U14213 (N_14213,N_10087,N_11591);
and U14214 (N_14214,N_9735,N_11309);
or U14215 (N_14215,N_8279,N_10207);
or U14216 (N_14216,N_10237,N_10752);
and U14217 (N_14217,N_8444,N_8180);
or U14218 (N_14218,N_11696,N_11190);
nor U14219 (N_14219,N_9233,N_8421);
or U14220 (N_14220,N_9708,N_11564);
or U14221 (N_14221,N_8511,N_9220);
xor U14222 (N_14222,N_8052,N_8344);
and U14223 (N_14223,N_11166,N_11287);
nand U14224 (N_14224,N_8325,N_11135);
xnor U14225 (N_14225,N_9916,N_10798);
nand U14226 (N_14226,N_9276,N_8570);
nor U14227 (N_14227,N_8345,N_11333);
nor U14228 (N_14228,N_9589,N_9435);
xor U14229 (N_14229,N_9846,N_9628);
and U14230 (N_14230,N_11672,N_10489);
nand U14231 (N_14231,N_9564,N_11825);
or U14232 (N_14232,N_9061,N_11703);
nand U14233 (N_14233,N_9691,N_8261);
nor U14234 (N_14234,N_8026,N_10607);
nand U14235 (N_14235,N_8315,N_8497);
nand U14236 (N_14236,N_8445,N_10176);
nand U14237 (N_14237,N_9167,N_10000);
nor U14238 (N_14238,N_8724,N_8245);
or U14239 (N_14239,N_11276,N_8979);
xnor U14240 (N_14240,N_9446,N_9849);
xnor U14241 (N_14241,N_11920,N_10834);
or U14242 (N_14242,N_8634,N_11063);
nand U14243 (N_14243,N_9335,N_10496);
nor U14244 (N_14244,N_8896,N_8180);
or U14245 (N_14245,N_10878,N_8230);
nor U14246 (N_14246,N_10398,N_8820);
xor U14247 (N_14247,N_11544,N_8855);
nor U14248 (N_14248,N_11524,N_9976);
or U14249 (N_14249,N_9635,N_10542);
nand U14250 (N_14250,N_9966,N_8663);
nand U14251 (N_14251,N_9496,N_9329);
xnor U14252 (N_14252,N_11068,N_9393);
nand U14253 (N_14253,N_10093,N_8830);
xnor U14254 (N_14254,N_8723,N_8983);
and U14255 (N_14255,N_9357,N_11376);
or U14256 (N_14256,N_8480,N_10887);
and U14257 (N_14257,N_8322,N_11254);
xnor U14258 (N_14258,N_11054,N_9579);
nand U14259 (N_14259,N_9591,N_11557);
or U14260 (N_14260,N_10856,N_10900);
and U14261 (N_14261,N_8730,N_10201);
nand U14262 (N_14262,N_8382,N_8262);
nor U14263 (N_14263,N_11555,N_11260);
nor U14264 (N_14264,N_11640,N_10852);
nor U14265 (N_14265,N_10011,N_10496);
or U14266 (N_14266,N_8244,N_11515);
nand U14267 (N_14267,N_8318,N_10117);
or U14268 (N_14268,N_11703,N_9741);
nor U14269 (N_14269,N_8074,N_11934);
nand U14270 (N_14270,N_8912,N_8201);
nand U14271 (N_14271,N_11610,N_8138);
nor U14272 (N_14272,N_8717,N_8933);
and U14273 (N_14273,N_10174,N_10145);
nor U14274 (N_14274,N_9038,N_11581);
nand U14275 (N_14275,N_10793,N_8703);
nor U14276 (N_14276,N_10213,N_11330);
nand U14277 (N_14277,N_11705,N_10288);
or U14278 (N_14278,N_11792,N_9691);
nand U14279 (N_14279,N_9558,N_10251);
xor U14280 (N_14280,N_8504,N_8297);
nor U14281 (N_14281,N_8272,N_9663);
or U14282 (N_14282,N_9069,N_9117);
nor U14283 (N_14283,N_8910,N_10187);
or U14284 (N_14284,N_11730,N_9103);
nand U14285 (N_14285,N_10020,N_10744);
xnor U14286 (N_14286,N_8623,N_11538);
or U14287 (N_14287,N_11727,N_8946);
or U14288 (N_14288,N_11949,N_9866);
and U14289 (N_14289,N_10995,N_8294);
xor U14290 (N_14290,N_9849,N_10531);
nor U14291 (N_14291,N_11088,N_8207);
nand U14292 (N_14292,N_8351,N_9661);
nor U14293 (N_14293,N_9736,N_8249);
or U14294 (N_14294,N_11827,N_11217);
nor U14295 (N_14295,N_11028,N_9537);
and U14296 (N_14296,N_9279,N_8371);
nor U14297 (N_14297,N_9193,N_8281);
or U14298 (N_14298,N_8173,N_9321);
nand U14299 (N_14299,N_9156,N_9502);
xnor U14300 (N_14300,N_10472,N_10998);
nand U14301 (N_14301,N_8537,N_10701);
or U14302 (N_14302,N_10972,N_10931);
or U14303 (N_14303,N_8120,N_11608);
or U14304 (N_14304,N_10699,N_9046);
nor U14305 (N_14305,N_9878,N_10699);
xnor U14306 (N_14306,N_8118,N_8529);
nand U14307 (N_14307,N_10952,N_9019);
xor U14308 (N_14308,N_8468,N_10532);
xor U14309 (N_14309,N_10426,N_9622);
xor U14310 (N_14310,N_8656,N_11385);
or U14311 (N_14311,N_10102,N_10543);
xnor U14312 (N_14312,N_10377,N_9540);
or U14313 (N_14313,N_9944,N_11433);
nand U14314 (N_14314,N_11643,N_11033);
nand U14315 (N_14315,N_9228,N_11733);
or U14316 (N_14316,N_9984,N_10563);
nand U14317 (N_14317,N_9832,N_11763);
nor U14318 (N_14318,N_9754,N_10265);
nand U14319 (N_14319,N_11942,N_10632);
nand U14320 (N_14320,N_10545,N_8236);
nand U14321 (N_14321,N_9938,N_10981);
nor U14322 (N_14322,N_11729,N_11248);
nor U14323 (N_14323,N_9088,N_9157);
and U14324 (N_14324,N_8896,N_9857);
or U14325 (N_14325,N_11126,N_9459);
and U14326 (N_14326,N_9278,N_9859);
nor U14327 (N_14327,N_11028,N_10316);
xnor U14328 (N_14328,N_10525,N_11901);
nand U14329 (N_14329,N_11332,N_10209);
nand U14330 (N_14330,N_11878,N_9629);
nor U14331 (N_14331,N_8846,N_11621);
xnor U14332 (N_14332,N_8093,N_10201);
and U14333 (N_14333,N_9968,N_10192);
or U14334 (N_14334,N_11001,N_8667);
nor U14335 (N_14335,N_10053,N_11868);
xnor U14336 (N_14336,N_11275,N_8459);
or U14337 (N_14337,N_8052,N_9776);
nor U14338 (N_14338,N_10277,N_8057);
nor U14339 (N_14339,N_9043,N_9659);
or U14340 (N_14340,N_8190,N_8948);
nor U14341 (N_14341,N_8443,N_9972);
and U14342 (N_14342,N_8178,N_11664);
xnor U14343 (N_14343,N_10474,N_8446);
nor U14344 (N_14344,N_10704,N_11297);
xor U14345 (N_14345,N_9475,N_9299);
nor U14346 (N_14346,N_8295,N_10857);
nand U14347 (N_14347,N_10403,N_8631);
and U14348 (N_14348,N_8745,N_10242);
nand U14349 (N_14349,N_8467,N_11139);
nor U14350 (N_14350,N_11566,N_11188);
and U14351 (N_14351,N_8703,N_8433);
nor U14352 (N_14352,N_8704,N_11597);
or U14353 (N_14353,N_10932,N_8780);
or U14354 (N_14354,N_11767,N_9378);
nor U14355 (N_14355,N_10192,N_10225);
nor U14356 (N_14356,N_10839,N_8150);
nor U14357 (N_14357,N_11474,N_10703);
xnor U14358 (N_14358,N_11020,N_8494);
nand U14359 (N_14359,N_11855,N_10589);
xnor U14360 (N_14360,N_9477,N_11111);
and U14361 (N_14361,N_10572,N_8066);
nor U14362 (N_14362,N_9573,N_8879);
xnor U14363 (N_14363,N_8701,N_10412);
nand U14364 (N_14364,N_8443,N_8813);
or U14365 (N_14365,N_9698,N_11285);
nor U14366 (N_14366,N_10205,N_11083);
nor U14367 (N_14367,N_9564,N_10131);
nand U14368 (N_14368,N_8009,N_10213);
nor U14369 (N_14369,N_10439,N_10113);
and U14370 (N_14370,N_10686,N_8513);
xnor U14371 (N_14371,N_8149,N_8385);
nand U14372 (N_14372,N_10686,N_10283);
nor U14373 (N_14373,N_8764,N_8768);
or U14374 (N_14374,N_10185,N_8856);
xnor U14375 (N_14375,N_10180,N_11851);
nor U14376 (N_14376,N_11310,N_8715);
or U14377 (N_14377,N_9479,N_11438);
nor U14378 (N_14378,N_10868,N_8503);
or U14379 (N_14379,N_10669,N_8398);
or U14380 (N_14380,N_11400,N_9551);
and U14381 (N_14381,N_11921,N_10617);
nor U14382 (N_14382,N_8699,N_10768);
nand U14383 (N_14383,N_8137,N_10625);
nand U14384 (N_14384,N_9901,N_10970);
or U14385 (N_14385,N_9917,N_11277);
or U14386 (N_14386,N_10100,N_10255);
xnor U14387 (N_14387,N_11076,N_9321);
and U14388 (N_14388,N_9357,N_11354);
and U14389 (N_14389,N_11531,N_11194);
nor U14390 (N_14390,N_9826,N_9132);
nand U14391 (N_14391,N_8313,N_10535);
nor U14392 (N_14392,N_9630,N_8464);
and U14393 (N_14393,N_8304,N_9712);
or U14394 (N_14394,N_9367,N_9364);
nand U14395 (N_14395,N_10745,N_8746);
or U14396 (N_14396,N_10070,N_8799);
nor U14397 (N_14397,N_10847,N_8841);
and U14398 (N_14398,N_10252,N_10233);
and U14399 (N_14399,N_9034,N_10012);
or U14400 (N_14400,N_8375,N_9742);
nand U14401 (N_14401,N_8178,N_9648);
nor U14402 (N_14402,N_9635,N_9429);
nand U14403 (N_14403,N_11760,N_8502);
and U14404 (N_14404,N_9316,N_11978);
nor U14405 (N_14405,N_8175,N_9895);
xnor U14406 (N_14406,N_10374,N_8190);
nand U14407 (N_14407,N_11518,N_11969);
or U14408 (N_14408,N_11522,N_9614);
or U14409 (N_14409,N_8861,N_11947);
nand U14410 (N_14410,N_10121,N_10093);
nor U14411 (N_14411,N_8243,N_10073);
xor U14412 (N_14412,N_8316,N_9081);
nand U14413 (N_14413,N_10621,N_10442);
or U14414 (N_14414,N_11844,N_10733);
nand U14415 (N_14415,N_11603,N_8169);
or U14416 (N_14416,N_9821,N_8517);
nand U14417 (N_14417,N_11087,N_8201);
nand U14418 (N_14418,N_10093,N_8086);
nor U14419 (N_14419,N_10847,N_10392);
nand U14420 (N_14420,N_11015,N_9944);
or U14421 (N_14421,N_11071,N_8760);
and U14422 (N_14422,N_10263,N_9734);
or U14423 (N_14423,N_9183,N_8433);
or U14424 (N_14424,N_9686,N_10392);
nor U14425 (N_14425,N_11419,N_8154);
or U14426 (N_14426,N_9434,N_9606);
nand U14427 (N_14427,N_8638,N_11968);
nor U14428 (N_14428,N_10373,N_9120);
nor U14429 (N_14429,N_8075,N_10817);
xor U14430 (N_14430,N_8928,N_9397);
and U14431 (N_14431,N_11039,N_10145);
or U14432 (N_14432,N_8153,N_9699);
nand U14433 (N_14433,N_10265,N_9837);
and U14434 (N_14434,N_9716,N_9007);
nor U14435 (N_14435,N_8979,N_9850);
and U14436 (N_14436,N_8006,N_8411);
and U14437 (N_14437,N_11673,N_9389);
and U14438 (N_14438,N_9911,N_8994);
nor U14439 (N_14439,N_10581,N_10935);
nand U14440 (N_14440,N_10869,N_9670);
nor U14441 (N_14441,N_10125,N_9218);
nand U14442 (N_14442,N_10298,N_9118);
nand U14443 (N_14443,N_8268,N_8892);
xor U14444 (N_14444,N_8845,N_10843);
nand U14445 (N_14445,N_10026,N_11752);
or U14446 (N_14446,N_8341,N_10295);
or U14447 (N_14447,N_8960,N_8376);
and U14448 (N_14448,N_10195,N_8163);
nor U14449 (N_14449,N_9926,N_11493);
or U14450 (N_14450,N_9572,N_9734);
nor U14451 (N_14451,N_9304,N_10408);
nand U14452 (N_14452,N_8562,N_10566);
or U14453 (N_14453,N_10246,N_10450);
nor U14454 (N_14454,N_11669,N_9235);
and U14455 (N_14455,N_8247,N_11752);
or U14456 (N_14456,N_8494,N_11812);
or U14457 (N_14457,N_10196,N_11512);
and U14458 (N_14458,N_10630,N_10622);
or U14459 (N_14459,N_10780,N_10844);
or U14460 (N_14460,N_11595,N_11693);
nand U14461 (N_14461,N_8969,N_10034);
nand U14462 (N_14462,N_8357,N_11498);
nor U14463 (N_14463,N_9354,N_9900);
nor U14464 (N_14464,N_9541,N_11952);
nand U14465 (N_14465,N_10818,N_10680);
or U14466 (N_14466,N_11265,N_11910);
nand U14467 (N_14467,N_8259,N_9846);
nor U14468 (N_14468,N_11734,N_11000);
nor U14469 (N_14469,N_8945,N_9647);
and U14470 (N_14470,N_8442,N_11867);
nand U14471 (N_14471,N_8358,N_8692);
xor U14472 (N_14472,N_8864,N_10821);
nor U14473 (N_14473,N_10340,N_9016);
nor U14474 (N_14474,N_8777,N_10716);
or U14475 (N_14475,N_9733,N_11144);
nor U14476 (N_14476,N_8854,N_9037);
xor U14477 (N_14477,N_11213,N_8940);
nor U14478 (N_14478,N_8583,N_8833);
xnor U14479 (N_14479,N_10152,N_9895);
xnor U14480 (N_14480,N_8811,N_8325);
nor U14481 (N_14481,N_10199,N_8293);
nand U14482 (N_14482,N_10398,N_10353);
nand U14483 (N_14483,N_10277,N_9513);
nor U14484 (N_14484,N_9074,N_9765);
nand U14485 (N_14485,N_10151,N_8505);
xor U14486 (N_14486,N_11834,N_9540);
nor U14487 (N_14487,N_8510,N_9689);
xor U14488 (N_14488,N_8022,N_10695);
nand U14489 (N_14489,N_9410,N_11951);
or U14490 (N_14490,N_10815,N_9599);
xnor U14491 (N_14491,N_8678,N_10019);
nor U14492 (N_14492,N_10862,N_10475);
nor U14493 (N_14493,N_10449,N_9723);
or U14494 (N_14494,N_8932,N_10938);
and U14495 (N_14495,N_11692,N_11318);
xor U14496 (N_14496,N_10415,N_9509);
nand U14497 (N_14497,N_9498,N_9214);
and U14498 (N_14498,N_10886,N_8871);
and U14499 (N_14499,N_11173,N_9519);
and U14500 (N_14500,N_10996,N_9310);
nor U14501 (N_14501,N_11433,N_11064);
or U14502 (N_14502,N_10923,N_9041);
nand U14503 (N_14503,N_10948,N_10546);
nor U14504 (N_14504,N_8084,N_8746);
or U14505 (N_14505,N_9008,N_10332);
nor U14506 (N_14506,N_9473,N_8989);
nor U14507 (N_14507,N_9301,N_10547);
xnor U14508 (N_14508,N_10740,N_9876);
xor U14509 (N_14509,N_8315,N_10758);
or U14510 (N_14510,N_8309,N_10508);
nor U14511 (N_14511,N_10962,N_10880);
nand U14512 (N_14512,N_10018,N_11074);
or U14513 (N_14513,N_9312,N_11196);
or U14514 (N_14514,N_8827,N_8989);
or U14515 (N_14515,N_11165,N_11881);
or U14516 (N_14516,N_9422,N_10223);
nor U14517 (N_14517,N_11098,N_11831);
nor U14518 (N_14518,N_10688,N_9622);
nor U14519 (N_14519,N_10246,N_10975);
nor U14520 (N_14520,N_11146,N_9215);
and U14521 (N_14521,N_10673,N_8882);
nand U14522 (N_14522,N_9197,N_10258);
or U14523 (N_14523,N_8684,N_8591);
nor U14524 (N_14524,N_9039,N_11325);
and U14525 (N_14525,N_8634,N_10820);
nand U14526 (N_14526,N_8416,N_9930);
nand U14527 (N_14527,N_9645,N_8351);
or U14528 (N_14528,N_9731,N_8825);
and U14529 (N_14529,N_9791,N_10318);
and U14530 (N_14530,N_10779,N_8172);
or U14531 (N_14531,N_11196,N_10500);
nor U14532 (N_14532,N_10533,N_8991);
and U14533 (N_14533,N_8821,N_10746);
or U14534 (N_14534,N_10418,N_10823);
nor U14535 (N_14535,N_8096,N_11627);
or U14536 (N_14536,N_9549,N_10957);
or U14537 (N_14537,N_11913,N_11189);
xor U14538 (N_14538,N_8607,N_10429);
nor U14539 (N_14539,N_10992,N_8180);
nor U14540 (N_14540,N_11748,N_10211);
or U14541 (N_14541,N_8815,N_11221);
nor U14542 (N_14542,N_11223,N_8590);
nor U14543 (N_14543,N_10411,N_8785);
nor U14544 (N_14544,N_10853,N_8251);
or U14545 (N_14545,N_11597,N_8632);
nand U14546 (N_14546,N_9082,N_9650);
nand U14547 (N_14547,N_8461,N_9173);
nor U14548 (N_14548,N_11813,N_9152);
and U14549 (N_14549,N_11765,N_9562);
and U14550 (N_14550,N_9640,N_9619);
and U14551 (N_14551,N_9201,N_10139);
nand U14552 (N_14552,N_9086,N_9106);
and U14553 (N_14553,N_9414,N_11057);
or U14554 (N_14554,N_11732,N_11638);
nand U14555 (N_14555,N_11862,N_9886);
or U14556 (N_14556,N_8646,N_11526);
and U14557 (N_14557,N_8827,N_8727);
nor U14558 (N_14558,N_8847,N_10579);
or U14559 (N_14559,N_10813,N_11020);
or U14560 (N_14560,N_11605,N_11502);
nand U14561 (N_14561,N_8271,N_11722);
or U14562 (N_14562,N_9469,N_11649);
nor U14563 (N_14563,N_9222,N_9862);
nand U14564 (N_14564,N_11418,N_11138);
nor U14565 (N_14565,N_10010,N_11873);
nor U14566 (N_14566,N_11971,N_10315);
nand U14567 (N_14567,N_8070,N_11407);
nand U14568 (N_14568,N_11610,N_10027);
nand U14569 (N_14569,N_9566,N_9217);
or U14570 (N_14570,N_9403,N_10806);
nor U14571 (N_14571,N_8946,N_10176);
nand U14572 (N_14572,N_10159,N_11086);
nor U14573 (N_14573,N_10590,N_10952);
and U14574 (N_14574,N_10244,N_11419);
nor U14575 (N_14575,N_10140,N_8760);
and U14576 (N_14576,N_9941,N_11379);
and U14577 (N_14577,N_9068,N_11937);
nor U14578 (N_14578,N_10637,N_10649);
nor U14579 (N_14579,N_11175,N_8688);
and U14580 (N_14580,N_11018,N_11669);
nand U14581 (N_14581,N_9926,N_11342);
nor U14582 (N_14582,N_11882,N_9575);
nor U14583 (N_14583,N_8905,N_8640);
and U14584 (N_14584,N_10103,N_9648);
and U14585 (N_14585,N_8579,N_8238);
and U14586 (N_14586,N_8320,N_8524);
nand U14587 (N_14587,N_10774,N_8366);
nor U14588 (N_14588,N_8196,N_8537);
nor U14589 (N_14589,N_9020,N_9297);
or U14590 (N_14590,N_8870,N_8771);
or U14591 (N_14591,N_8271,N_9636);
nand U14592 (N_14592,N_11345,N_8216);
or U14593 (N_14593,N_9248,N_9049);
and U14594 (N_14594,N_10848,N_8386);
and U14595 (N_14595,N_10557,N_10901);
xnor U14596 (N_14596,N_8443,N_9147);
or U14597 (N_14597,N_8463,N_8474);
and U14598 (N_14598,N_10322,N_8616);
xor U14599 (N_14599,N_10411,N_10742);
or U14600 (N_14600,N_8708,N_11098);
or U14601 (N_14601,N_11824,N_9301);
nand U14602 (N_14602,N_9332,N_8014);
and U14603 (N_14603,N_10754,N_9607);
nand U14604 (N_14604,N_11496,N_10376);
nor U14605 (N_14605,N_8332,N_11599);
nor U14606 (N_14606,N_11579,N_10496);
nor U14607 (N_14607,N_11436,N_9045);
nor U14608 (N_14608,N_11994,N_10910);
or U14609 (N_14609,N_9639,N_10847);
or U14610 (N_14610,N_9108,N_10792);
or U14611 (N_14611,N_10352,N_11392);
and U14612 (N_14612,N_11079,N_8914);
xnor U14613 (N_14613,N_10892,N_8807);
or U14614 (N_14614,N_11140,N_8503);
nor U14615 (N_14615,N_11934,N_10581);
and U14616 (N_14616,N_10927,N_9779);
nand U14617 (N_14617,N_8800,N_11006);
nand U14618 (N_14618,N_9443,N_10244);
nor U14619 (N_14619,N_11617,N_8120);
nor U14620 (N_14620,N_10677,N_8155);
or U14621 (N_14621,N_11810,N_11037);
or U14622 (N_14622,N_11002,N_8584);
or U14623 (N_14623,N_9735,N_9012);
nand U14624 (N_14624,N_8916,N_8133);
or U14625 (N_14625,N_10814,N_10916);
nand U14626 (N_14626,N_9084,N_9948);
or U14627 (N_14627,N_9543,N_9238);
and U14628 (N_14628,N_8953,N_10002);
nor U14629 (N_14629,N_8260,N_11723);
nor U14630 (N_14630,N_11453,N_8826);
or U14631 (N_14631,N_10800,N_9897);
nand U14632 (N_14632,N_8106,N_11828);
or U14633 (N_14633,N_8907,N_11367);
nor U14634 (N_14634,N_10015,N_11571);
or U14635 (N_14635,N_10825,N_10886);
and U14636 (N_14636,N_9519,N_8225);
or U14637 (N_14637,N_9343,N_10357);
xnor U14638 (N_14638,N_11921,N_11619);
or U14639 (N_14639,N_10882,N_9243);
nand U14640 (N_14640,N_9337,N_8574);
nand U14641 (N_14641,N_11659,N_9279);
or U14642 (N_14642,N_10146,N_10728);
nand U14643 (N_14643,N_8347,N_8365);
nand U14644 (N_14644,N_11857,N_10258);
nand U14645 (N_14645,N_8340,N_10573);
nor U14646 (N_14646,N_10402,N_9965);
nor U14647 (N_14647,N_8852,N_9757);
xor U14648 (N_14648,N_11274,N_8690);
nor U14649 (N_14649,N_11277,N_10664);
nor U14650 (N_14650,N_11225,N_9864);
or U14651 (N_14651,N_9366,N_9841);
nand U14652 (N_14652,N_10003,N_9879);
or U14653 (N_14653,N_10798,N_8721);
nand U14654 (N_14654,N_8017,N_11775);
nor U14655 (N_14655,N_8554,N_10511);
nor U14656 (N_14656,N_8529,N_8731);
and U14657 (N_14657,N_10160,N_9243);
or U14658 (N_14658,N_10985,N_10904);
or U14659 (N_14659,N_9323,N_8286);
nor U14660 (N_14660,N_9592,N_9488);
nor U14661 (N_14661,N_8679,N_11181);
or U14662 (N_14662,N_9709,N_8164);
xnor U14663 (N_14663,N_9617,N_10077);
xor U14664 (N_14664,N_11062,N_8400);
or U14665 (N_14665,N_11553,N_11827);
and U14666 (N_14666,N_9643,N_9967);
and U14667 (N_14667,N_8216,N_8946);
nor U14668 (N_14668,N_10087,N_8164);
and U14669 (N_14669,N_9935,N_10162);
nor U14670 (N_14670,N_8643,N_11695);
and U14671 (N_14671,N_8935,N_11484);
nor U14672 (N_14672,N_8788,N_9745);
nand U14673 (N_14673,N_8763,N_9939);
nand U14674 (N_14674,N_8110,N_9871);
or U14675 (N_14675,N_9242,N_8044);
nor U14676 (N_14676,N_10515,N_8076);
nand U14677 (N_14677,N_9461,N_11637);
or U14678 (N_14678,N_8668,N_10526);
or U14679 (N_14679,N_9409,N_11293);
nand U14680 (N_14680,N_10696,N_11950);
and U14681 (N_14681,N_11340,N_11049);
xnor U14682 (N_14682,N_9763,N_10651);
nand U14683 (N_14683,N_11327,N_10262);
or U14684 (N_14684,N_8327,N_8169);
nand U14685 (N_14685,N_10214,N_9578);
nor U14686 (N_14686,N_10240,N_11115);
xor U14687 (N_14687,N_8075,N_10581);
nand U14688 (N_14688,N_8538,N_9328);
nor U14689 (N_14689,N_8762,N_9213);
nor U14690 (N_14690,N_8791,N_10617);
or U14691 (N_14691,N_11783,N_9872);
nand U14692 (N_14692,N_9472,N_11205);
xor U14693 (N_14693,N_11745,N_8225);
and U14694 (N_14694,N_11916,N_8177);
nor U14695 (N_14695,N_10595,N_10394);
nand U14696 (N_14696,N_10110,N_9820);
nand U14697 (N_14697,N_10453,N_11267);
nand U14698 (N_14698,N_11116,N_9172);
and U14699 (N_14699,N_11217,N_9161);
and U14700 (N_14700,N_10136,N_8995);
and U14701 (N_14701,N_10675,N_11948);
nor U14702 (N_14702,N_10299,N_9170);
and U14703 (N_14703,N_9662,N_9448);
nor U14704 (N_14704,N_9740,N_11605);
or U14705 (N_14705,N_11990,N_8341);
or U14706 (N_14706,N_9765,N_8573);
nor U14707 (N_14707,N_10110,N_9602);
and U14708 (N_14708,N_11449,N_11512);
xnor U14709 (N_14709,N_10047,N_8530);
or U14710 (N_14710,N_10569,N_9542);
and U14711 (N_14711,N_11860,N_9522);
nor U14712 (N_14712,N_9297,N_8604);
xnor U14713 (N_14713,N_10273,N_11711);
or U14714 (N_14714,N_10938,N_10266);
and U14715 (N_14715,N_10023,N_8896);
nor U14716 (N_14716,N_11264,N_8580);
nand U14717 (N_14717,N_10275,N_10650);
or U14718 (N_14718,N_9380,N_10052);
or U14719 (N_14719,N_11183,N_10056);
nor U14720 (N_14720,N_11990,N_9097);
or U14721 (N_14721,N_10186,N_11208);
nor U14722 (N_14722,N_9501,N_9240);
or U14723 (N_14723,N_8055,N_11813);
nor U14724 (N_14724,N_11990,N_11644);
and U14725 (N_14725,N_11647,N_9596);
nand U14726 (N_14726,N_9706,N_8937);
and U14727 (N_14727,N_10824,N_9519);
or U14728 (N_14728,N_11107,N_8157);
xor U14729 (N_14729,N_8935,N_9086);
or U14730 (N_14730,N_10309,N_10466);
or U14731 (N_14731,N_9512,N_9665);
xnor U14732 (N_14732,N_10557,N_11134);
or U14733 (N_14733,N_9376,N_11024);
xnor U14734 (N_14734,N_9115,N_10168);
and U14735 (N_14735,N_10520,N_9143);
nand U14736 (N_14736,N_8876,N_8934);
xor U14737 (N_14737,N_10208,N_9327);
xor U14738 (N_14738,N_8443,N_10538);
and U14739 (N_14739,N_9497,N_11443);
or U14740 (N_14740,N_10980,N_10960);
or U14741 (N_14741,N_11982,N_9105);
or U14742 (N_14742,N_9152,N_11434);
nand U14743 (N_14743,N_11004,N_10118);
nor U14744 (N_14744,N_10590,N_9644);
xnor U14745 (N_14745,N_10283,N_11019);
xnor U14746 (N_14746,N_10516,N_8087);
or U14747 (N_14747,N_11585,N_8133);
or U14748 (N_14748,N_11045,N_8112);
or U14749 (N_14749,N_10515,N_11702);
xnor U14750 (N_14750,N_8286,N_8692);
nor U14751 (N_14751,N_8127,N_10402);
nor U14752 (N_14752,N_10255,N_9117);
and U14753 (N_14753,N_10929,N_8114);
nor U14754 (N_14754,N_8036,N_9389);
nor U14755 (N_14755,N_10117,N_10420);
nand U14756 (N_14756,N_10357,N_8319);
nand U14757 (N_14757,N_9150,N_8774);
nand U14758 (N_14758,N_10816,N_11188);
nor U14759 (N_14759,N_8552,N_9428);
nor U14760 (N_14760,N_8635,N_10833);
or U14761 (N_14761,N_8134,N_10163);
nor U14762 (N_14762,N_9087,N_9539);
nor U14763 (N_14763,N_10104,N_9795);
nand U14764 (N_14764,N_11292,N_9246);
and U14765 (N_14765,N_9259,N_11016);
nor U14766 (N_14766,N_10971,N_9579);
nand U14767 (N_14767,N_11088,N_10549);
nand U14768 (N_14768,N_10291,N_9240);
or U14769 (N_14769,N_11203,N_8236);
nor U14770 (N_14770,N_11782,N_11473);
nor U14771 (N_14771,N_10848,N_9707);
and U14772 (N_14772,N_8605,N_10115);
nand U14773 (N_14773,N_9835,N_11648);
nor U14774 (N_14774,N_11938,N_8049);
and U14775 (N_14775,N_11393,N_11221);
or U14776 (N_14776,N_9759,N_11984);
and U14777 (N_14777,N_10729,N_10152);
and U14778 (N_14778,N_9069,N_8478);
nor U14779 (N_14779,N_11188,N_10000);
or U14780 (N_14780,N_10716,N_10782);
nor U14781 (N_14781,N_11331,N_9727);
nor U14782 (N_14782,N_10361,N_10585);
nand U14783 (N_14783,N_9990,N_9890);
nand U14784 (N_14784,N_10908,N_10839);
nor U14785 (N_14785,N_8616,N_8421);
nor U14786 (N_14786,N_8242,N_8770);
and U14787 (N_14787,N_10812,N_11409);
nor U14788 (N_14788,N_8359,N_10709);
and U14789 (N_14789,N_8459,N_8355);
nand U14790 (N_14790,N_11809,N_11958);
nor U14791 (N_14791,N_11068,N_9145);
nand U14792 (N_14792,N_9224,N_9024);
or U14793 (N_14793,N_9666,N_9692);
nor U14794 (N_14794,N_8905,N_11212);
and U14795 (N_14795,N_8676,N_11223);
or U14796 (N_14796,N_9171,N_10614);
nor U14797 (N_14797,N_8972,N_10108);
or U14798 (N_14798,N_11139,N_9312);
xor U14799 (N_14799,N_11912,N_9866);
nand U14800 (N_14800,N_9357,N_11339);
nor U14801 (N_14801,N_10444,N_9805);
nor U14802 (N_14802,N_8229,N_8638);
and U14803 (N_14803,N_11258,N_9449);
nand U14804 (N_14804,N_10578,N_8675);
and U14805 (N_14805,N_8413,N_8584);
and U14806 (N_14806,N_8729,N_9583);
or U14807 (N_14807,N_11448,N_9437);
nand U14808 (N_14808,N_11840,N_9668);
nand U14809 (N_14809,N_10228,N_11187);
or U14810 (N_14810,N_10004,N_8544);
or U14811 (N_14811,N_11526,N_11773);
and U14812 (N_14812,N_11881,N_8609);
or U14813 (N_14813,N_10110,N_10930);
xnor U14814 (N_14814,N_9353,N_9427);
nor U14815 (N_14815,N_11914,N_8958);
nor U14816 (N_14816,N_9942,N_9496);
nor U14817 (N_14817,N_9993,N_8550);
and U14818 (N_14818,N_8737,N_10850);
and U14819 (N_14819,N_8913,N_9699);
nor U14820 (N_14820,N_9881,N_11746);
and U14821 (N_14821,N_9683,N_9315);
nor U14822 (N_14822,N_11358,N_10357);
nor U14823 (N_14823,N_9290,N_8663);
or U14824 (N_14824,N_8042,N_10910);
and U14825 (N_14825,N_10249,N_10522);
or U14826 (N_14826,N_9988,N_8783);
nor U14827 (N_14827,N_10757,N_9908);
or U14828 (N_14828,N_9260,N_8860);
nand U14829 (N_14829,N_8341,N_8664);
or U14830 (N_14830,N_9910,N_10016);
and U14831 (N_14831,N_11479,N_8423);
or U14832 (N_14832,N_11974,N_8077);
and U14833 (N_14833,N_10874,N_11048);
nand U14834 (N_14834,N_10661,N_10293);
and U14835 (N_14835,N_10721,N_9986);
nand U14836 (N_14836,N_8397,N_9670);
nand U14837 (N_14837,N_10626,N_11175);
nand U14838 (N_14838,N_8912,N_9621);
nor U14839 (N_14839,N_11328,N_9324);
nor U14840 (N_14840,N_11005,N_10821);
or U14841 (N_14841,N_8424,N_9434);
and U14842 (N_14842,N_8760,N_10843);
and U14843 (N_14843,N_11992,N_9264);
nor U14844 (N_14844,N_11213,N_9524);
nor U14845 (N_14845,N_8746,N_11051);
nand U14846 (N_14846,N_9637,N_8543);
and U14847 (N_14847,N_9849,N_11504);
nand U14848 (N_14848,N_11948,N_11213);
nor U14849 (N_14849,N_9698,N_8160);
or U14850 (N_14850,N_10793,N_8073);
nand U14851 (N_14851,N_8015,N_10719);
or U14852 (N_14852,N_10030,N_9361);
xnor U14853 (N_14853,N_9696,N_9970);
nand U14854 (N_14854,N_11951,N_9331);
and U14855 (N_14855,N_10272,N_9980);
or U14856 (N_14856,N_11644,N_10124);
and U14857 (N_14857,N_9623,N_8265);
or U14858 (N_14858,N_11157,N_8154);
or U14859 (N_14859,N_11965,N_8059);
nand U14860 (N_14860,N_8009,N_9558);
nand U14861 (N_14861,N_11269,N_10822);
xor U14862 (N_14862,N_9913,N_9506);
nor U14863 (N_14863,N_10661,N_11396);
and U14864 (N_14864,N_9586,N_10015);
and U14865 (N_14865,N_10290,N_9437);
nand U14866 (N_14866,N_11705,N_9857);
and U14867 (N_14867,N_9701,N_10496);
nand U14868 (N_14868,N_10688,N_9581);
or U14869 (N_14869,N_10897,N_8140);
or U14870 (N_14870,N_8667,N_10057);
or U14871 (N_14871,N_10794,N_9420);
and U14872 (N_14872,N_10900,N_11266);
or U14873 (N_14873,N_10394,N_9503);
or U14874 (N_14874,N_8778,N_9471);
nor U14875 (N_14875,N_10298,N_9548);
or U14876 (N_14876,N_9720,N_8827);
nor U14877 (N_14877,N_11616,N_9155);
nor U14878 (N_14878,N_10561,N_11967);
or U14879 (N_14879,N_8520,N_11838);
or U14880 (N_14880,N_8266,N_9477);
nand U14881 (N_14881,N_11053,N_9036);
or U14882 (N_14882,N_11847,N_10970);
nand U14883 (N_14883,N_8302,N_9400);
nor U14884 (N_14884,N_9601,N_9319);
and U14885 (N_14885,N_10265,N_11389);
nand U14886 (N_14886,N_11302,N_10034);
and U14887 (N_14887,N_10081,N_11822);
nor U14888 (N_14888,N_9413,N_8804);
and U14889 (N_14889,N_11189,N_10049);
nor U14890 (N_14890,N_10609,N_8905);
nor U14891 (N_14891,N_10588,N_8515);
xnor U14892 (N_14892,N_9337,N_9205);
and U14893 (N_14893,N_11828,N_10718);
and U14894 (N_14894,N_10749,N_9592);
or U14895 (N_14895,N_10237,N_11702);
or U14896 (N_14896,N_11805,N_9796);
and U14897 (N_14897,N_9562,N_9290);
nand U14898 (N_14898,N_8262,N_11209);
or U14899 (N_14899,N_11433,N_9437);
and U14900 (N_14900,N_8138,N_8626);
nand U14901 (N_14901,N_9313,N_11032);
or U14902 (N_14902,N_10427,N_9748);
or U14903 (N_14903,N_8164,N_10858);
nor U14904 (N_14904,N_11437,N_10917);
or U14905 (N_14905,N_11685,N_9477);
nand U14906 (N_14906,N_8919,N_8871);
nand U14907 (N_14907,N_9207,N_9320);
and U14908 (N_14908,N_11600,N_10044);
and U14909 (N_14909,N_10034,N_10064);
and U14910 (N_14910,N_8086,N_11036);
nand U14911 (N_14911,N_9070,N_9706);
and U14912 (N_14912,N_11455,N_11688);
nand U14913 (N_14913,N_8494,N_8929);
nor U14914 (N_14914,N_10357,N_10736);
or U14915 (N_14915,N_10294,N_9589);
or U14916 (N_14916,N_11013,N_8108);
and U14917 (N_14917,N_8876,N_11553);
nor U14918 (N_14918,N_9468,N_10362);
nor U14919 (N_14919,N_10112,N_8524);
nand U14920 (N_14920,N_8901,N_9762);
xor U14921 (N_14921,N_10794,N_11934);
or U14922 (N_14922,N_9146,N_9321);
nor U14923 (N_14923,N_10935,N_10344);
or U14924 (N_14924,N_8394,N_11593);
nor U14925 (N_14925,N_9745,N_9143);
nor U14926 (N_14926,N_10942,N_11374);
or U14927 (N_14927,N_9330,N_9959);
nand U14928 (N_14928,N_11681,N_9937);
and U14929 (N_14929,N_9472,N_11657);
and U14930 (N_14930,N_8808,N_9176);
or U14931 (N_14931,N_9420,N_11773);
or U14932 (N_14932,N_10847,N_8711);
and U14933 (N_14933,N_10039,N_9784);
xnor U14934 (N_14934,N_10548,N_11874);
xor U14935 (N_14935,N_8569,N_10022);
nor U14936 (N_14936,N_8103,N_10427);
nor U14937 (N_14937,N_10474,N_10538);
or U14938 (N_14938,N_8250,N_10792);
nand U14939 (N_14939,N_9007,N_10095);
nor U14940 (N_14940,N_10529,N_9239);
nor U14941 (N_14941,N_11057,N_11358);
and U14942 (N_14942,N_8574,N_8232);
xnor U14943 (N_14943,N_11589,N_11381);
nor U14944 (N_14944,N_9346,N_8227);
nor U14945 (N_14945,N_10653,N_11610);
and U14946 (N_14946,N_9832,N_10388);
or U14947 (N_14947,N_11106,N_10391);
and U14948 (N_14948,N_11985,N_9122);
nand U14949 (N_14949,N_8114,N_10558);
and U14950 (N_14950,N_11171,N_9822);
nor U14951 (N_14951,N_9178,N_11387);
nand U14952 (N_14952,N_9355,N_9916);
xor U14953 (N_14953,N_11067,N_8975);
nand U14954 (N_14954,N_9479,N_9550);
and U14955 (N_14955,N_9973,N_9704);
nand U14956 (N_14956,N_9443,N_9788);
nand U14957 (N_14957,N_10621,N_8205);
nor U14958 (N_14958,N_10673,N_11354);
and U14959 (N_14959,N_11193,N_11554);
nor U14960 (N_14960,N_10257,N_8149);
or U14961 (N_14961,N_8930,N_8475);
nand U14962 (N_14962,N_10342,N_10299);
nand U14963 (N_14963,N_8369,N_11076);
nor U14964 (N_14964,N_10850,N_8960);
or U14965 (N_14965,N_9795,N_10215);
and U14966 (N_14966,N_9433,N_11577);
and U14967 (N_14967,N_11835,N_11485);
nand U14968 (N_14968,N_11200,N_11030);
nor U14969 (N_14969,N_10225,N_9798);
nand U14970 (N_14970,N_10892,N_11497);
nand U14971 (N_14971,N_9602,N_9079);
nor U14972 (N_14972,N_10023,N_8206);
nand U14973 (N_14973,N_11959,N_10582);
nand U14974 (N_14974,N_8228,N_11653);
xnor U14975 (N_14975,N_11789,N_11010);
nand U14976 (N_14976,N_11184,N_8509);
and U14977 (N_14977,N_10069,N_9484);
or U14978 (N_14978,N_11060,N_10949);
and U14979 (N_14979,N_11170,N_11645);
and U14980 (N_14980,N_11568,N_8170);
and U14981 (N_14981,N_9319,N_11498);
nand U14982 (N_14982,N_8366,N_9973);
nor U14983 (N_14983,N_8054,N_9712);
and U14984 (N_14984,N_11010,N_10474);
nor U14985 (N_14985,N_11210,N_11230);
nand U14986 (N_14986,N_9594,N_8882);
or U14987 (N_14987,N_8532,N_11814);
nand U14988 (N_14988,N_11284,N_8297);
nand U14989 (N_14989,N_10891,N_10722);
nand U14990 (N_14990,N_10376,N_8734);
and U14991 (N_14991,N_9053,N_9598);
or U14992 (N_14992,N_11916,N_10336);
or U14993 (N_14993,N_10690,N_9104);
and U14994 (N_14994,N_10136,N_11409);
xnor U14995 (N_14995,N_11734,N_10318);
xnor U14996 (N_14996,N_10927,N_8784);
and U14997 (N_14997,N_8090,N_9070);
or U14998 (N_14998,N_9957,N_11890);
nand U14999 (N_14999,N_8084,N_8043);
and U15000 (N_15000,N_9656,N_11344);
nor U15001 (N_15001,N_8342,N_9223);
xnor U15002 (N_15002,N_10679,N_9767);
or U15003 (N_15003,N_10749,N_8839);
or U15004 (N_15004,N_8199,N_11104);
nand U15005 (N_15005,N_11386,N_8307);
nand U15006 (N_15006,N_9919,N_11781);
and U15007 (N_15007,N_9573,N_9754);
nand U15008 (N_15008,N_10899,N_11923);
nand U15009 (N_15009,N_8371,N_8064);
nand U15010 (N_15010,N_8447,N_9054);
or U15011 (N_15011,N_8813,N_11550);
nor U15012 (N_15012,N_11836,N_9452);
xor U15013 (N_15013,N_11491,N_8672);
and U15014 (N_15014,N_9705,N_10713);
nand U15015 (N_15015,N_11524,N_8448);
nor U15016 (N_15016,N_8545,N_10377);
nand U15017 (N_15017,N_9541,N_9332);
and U15018 (N_15018,N_9176,N_11771);
xor U15019 (N_15019,N_11764,N_10397);
nand U15020 (N_15020,N_10792,N_9081);
or U15021 (N_15021,N_11273,N_10250);
xor U15022 (N_15022,N_9999,N_11403);
nor U15023 (N_15023,N_8216,N_10180);
xnor U15024 (N_15024,N_11120,N_8466);
and U15025 (N_15025,N_8524,N_11548);
or U15026 (N_15026,N_10442,N_8643);
and U15027 (N_15027,N_11681,N_8474);
and U15028 (N_15028,N_8482,N_8120);
nand U15029 (N_15029,N_9418,N_11840);
nand U15030 (N_15030,N_10498,N_9454);
nor U15031 (N_15031,N_11039,N_11280);
nor U15032 (N_15032,N_8489,N_8394);
nand U15033 (N_15033,N_10705,N_8451);
and U15034 (N_15034,N_9996,N_9581);
and U15035 (N_15035,N_8785,N_11516);
nand U15036 (N_15036,N_8138,N_11416);
nand U15037 (N_15037,N_11752,N_8521);
xor U15038 (N_15038,N_8232,N_10871);
nor U15039 (N_15039,N_10961,N_10282);
nand U15040 (N_15040,N_9635,N_8100);
and U15041 (N_15041,N_10078,N_9244);
or U15042 (N_15042,N_10998,N_11240);
nor U15043 (N_15043,N_11343,N_10620);
and U15044 (N_15044,N_10607,N_9226);
nor U15045 (N_15045,N_11973,N_8292);
or U15046 (N_15046,N_11605,N_8143);
or U15047 (N_15047,N_11723,N_11434);
nand U15048 (N_15048,N_10643,N_11834);
or U15049 (N_15049,N_10367,N_10204);
and U15050 (N_15050,N_8216,N_11949);
and U15051 (N_15051,N_8448,N_9464);
nor U15052 (N_15052,N_11167,N_10651);
and U15053 (N_15053,N_10415,N_11700);
and U15054 (N_15054,N_9850,N_10514);
xnor U15055 (N_15055,N_11085,N_9748);
or U15056 (N_15056,N_8060,N_8655);
or U15057 (N_15057,N_9211,N_8068);
nand U15058 (N_15058,N_8339,N_10545);
and U15059 (N_15059,N_8283,N_9683);
or U15060 (N_15060,N_11201,N_11229);
nor U15061 (N_15061,N_9907,N_10763);
and U15062 (N_15062,N_11627,N_11775);
and U15063 (N_15063,N_8188,N_8945);
or U15064 (N_15064,N_11480,N_11250);
and U15065 (N_15065,N_8231,N_9955);
or U15066 (N_15066,N_11792,N_8479);
nand U15067 (N_15067,N_9898,N_11935);
nand U15068 (N_15068,N_11059,N_10145);
and U15069 (N_15069,N_10550,N_9858);
and U15070 (N_15070,N_9024,N_10449);
or U15071 (N_15071,N_9255,N_10139);
nand U15072 (N_15072,N_10122,N_8069);
xor U15073 (N_15073,N_11233,N_9429);
nor U15074 (N_15074,N_10833,N_11797);
nor U15075 (N_15075,N_10019,N_8186);
nand U15076 (N_15076,N_10338,N_11040);
nor U15077 (N_15077,N_10617,N_9710);
or U15078 (N_15078,N_11987,N_9227);
nand U15079 (N_15079,N_11904,N_10849);
xor U15080 (N_15080,N_9840,N_8401);
or U15081 (N_15081,N_11214,N_8306);
nor U15082 (N_15082,N_10987,N_11575);
or U15083 (N_15083,N_9592,N_10108);
or U15084 (N_15084,N_11291,N_9328);
nand U15085 (N_15085,N_9373,N_11453);
or U15086 (N_15086,N_9245,N_10226);
or U15087 (N_15087,N_9279,N_9972);
or U15088 (N_15088,N_10059,N_9873);
or U15089 (N_15089,N_9345,N_9777);
nor U15090 (N_15090,N_11808,N_8884);
nor U15091 (N_15091,N_11615,N_8490);
and U15092 (N_15092,N_11793,N_11329);
and U15093 (N_15093,N_10824,N_9983);
and U15094 (N_15094,N_10954,N_10226);
nor U15095 (N_15095,N_11462,N_11762);
or U15096 (N_15096,N_11278,N_9284);
and U15097 (N_15097,N_11615,N_9730);
or U15098 (N_15098,N_9859,N_9119);
or U15099 (N_15099,N_9467,N_10242);
or U15100 (N_15100,N_10183,N_11529);
nand U15101 (N_15101,N_10562,N_11099);
nand U15102 (N_15102,N_11640,N_9284);
and U15103 (N_15103,N_8044,N_10496);
nand U15104 (N_15104,N_9874,N_9625);
nand U15105 (N_15105,N_8752,N_11527);
xor U15106 (N_15106,N_8710,N_10059);
or U15107 (N_15107,N_11817,N_11977);
nor U15108 (N_15108,N_8575,N_10346);
nand U15109 (N_15109,N_9910,N_11945);
or U15110 (N_15110,N_8056,N_11689);
xor U15111 (N_15111,N_8725,N_10931);
xor U15112 (N_15112,N_10153,N_11643);
xor U15113 (N_15113,N_11176,N_10192);
xnor U15114 (N_15114,N_9265,N_8354);
and U15115 (N_15115,N_9713,N_10404);
nor U15116 (N_15116,N_10700,N_8058);
nand U15117 (N_15117,N_9878,N_11349);
and U15118 (N_15118,N_9186,N_11981);
nor U15119 (N_15119,N_10140,N_11405);
and U15120 (N_15120,N_8995,N_9571);
nor U15121 (N_15121,N_9143,N_8614);
and U15122 (N_15122,N_10262,N_8305);
and U15123 (N_15123,N_8345,N_10109);
or U15124 (N_15124,N_9854,N_11348);
or U15125 (N_15125,N_9674,N_9682);
nor U15126 (N_15126,N_8695,N_11422);
nor U15127 (N_15127,N_11478,N_11210);
nand U15128 (N_15128,N_9458,N_11438);
and U15129 (N_15129,N_9451,N_9731);
or U15130 (N_15130,N_11064,N_8171);
nand U15131 (N_15131,N_8633,N_10950);
nand U15132 (N_15132,N_9582,N_10496);
or U15133 (N_15133,N_8782,N_9864);
or U15134 (N_15134,N_9027,N_10779);
nand U15135 (N_15135,N_8423,N_10967);
nor U15136 (N_15136,N_8799,N_9477);
nor U15137 (N_15137,N_10063,N_8762);
nor U15138 (N_15138,N_8435,N_9634);
nand U15139 (N_15139,N_9091,N_10909);
xor U15140 (N_15140,N_11689,N_9701);
and U15141 (N_15141,N_9343,N_10731);
or U15142 (N_15142,N_11324,N_10033);
or U15143 (N_15143,N_8511,N_10170);
nand U15144 (N_15144,N_9136,N_8509);
xnor U15145 (N_15145,N_9590,N_9346);
nor U15146 (N_15146,N_9516,N_9575);
and U15147 (N_15147,N_10902,N_8780);
xor U15148 (N_15148,N_9181,N_10616);
or U15149 (N_15149,N_11818,N_10224);
nand U15150 (N_15150,N_10550,N_11779);
and U15151 (N_15151,N_8327,N_9086);
nor U15152 (N_15152,N_9714,N_10762);
nor U15153 (N_15153,N_8499,N_8731);
nand U15154 (N_15154,N_11805,N_10243);
or U15155 (N_15155,N_9952,N_9252);
nor U15156 (N_15156,N_8256,N_9582);
and U15157 (N_15157,N_11281,N_10854);
or U15158 (N_15158,N_8344,N_11989);
xor U15159 (N_15159,N_9114,N_10979);
nor U15160 (N_15160,N_11686,N_10255);
xor U15161 (N_15161,N_9404,N_8268);
nor U15162 (N_15162,N_9044,N_10227);
nor U15163 (N_15163,N_10284,N_10269);
nor U15164 (N_15164,N_8597,N_10475);
nor U15165 (N_15165,N_10000,N_11962);
and U15166 (N_15166,N_10180,N_8412);
nand U15167 (N_15167,N_10284,N_9262);
and U15168 (N_15168,N_11427,N_9647);
nand U15169 (N_15169,N_11697,N_9299);
nor U15170 (N_15170,N_8979,N_9788);
nor U15171 (N_15171,N_8785,N_9016);
nand U15172 (N_15172,N_8559,N_8152);
nand U15173 (N_15173,N_10342,N_11623);
or U15174 (N_15174,N_10116,N_10861);
and U15175 (N_15175,N_9046,N_8782);
nand U15176 (N_15176,N_10229,N_8076);
or U15177 (N_15177,N_9719,N_11464);
xor U15178 (N_15178,N_8206,N_11115);
nor U15179 (N_15179,N_11151,N_11899);
nand U15180 (N_15180,N_11576,N_11915);
nand U15181 (N_15181,N_9249,N_11000);
nand U15182 (N_15182,N_8687,N_10586);
or U15183 (N_15183,N_10685,N_9397);
nand U15184 (N_15184,N_8516,N_9876);
and U15185 (N_15185,N_11693,N_11800);
nor U15186 (N_15186,N_10851,N_8037);
nor U15187 (N_15187,N_10775,N_9318);
or U15188 (N_15188,N_9927,N_10634);
or U15189 (N_15189,N_11007,N_8909);
nand U15190 (N_15190,N_10758,N_11321);
nand U15191 (N_15191,N_8710,N_9202);
or U15192 (N_15192,N_10749,N_9486);
and U15193 (N_15193,N_9344,N_8297);
xnor U15194 (N_15194,N_8158,N_10228);
or U15195 (N_15195,N_9649,N_9289);
or U15196 (N_15196,N_10637,N_10315);
or U15197 (N_15197,N_11394,N_9919);
nand U15198 (N_15198,N_8732,N_8572);
or U15199 (N_15199,N_11285,N_9322);
nand U15200 (N_15200,N_8443,N_11044);
and U15201 (N_15201,N_9113,N_9728);
nand U15202 (N_15202,N_11872,N_9561);
nor U15203 (N_15203,N_10364,N_8770);
and U15204 (N_15204,N_10121,N_8646);
nor U15205 (N_15205,N_9978,N_10096);
nand U15206 (N_15206,N_9458,N_8635);
and U15207 (N_15207,N_10843,N_9133);
or U15208 (N_15208,N_9190,N_8249);
nor U15209 (N_15209,N_8903,N_9496);
xnor U15210 (N_15210,N_8032,N_10955);
xnor U15211 (N_15211,N_8742,N_10754);
xor U15212 (N_15212,N_8204,N_8009);
nand U15213 (N_15213,N_9574,N_8604);
xnor U15214 (N_15214,N_10331,N_8281);
and U15215 (N_15215,N_11345,N_9373);
and U15216 (N_15216,N_9181,N_8779);
nor U15217 (N_15217,N_8890,N_8992);
and U15218 (N_15218,N_8323,N_10868);
nand U15219 (N_15219,N_11501,N_9394);
xnor U15220 (N_15220,N_9809,N_9482);
nand U15221 (N_15221,N_8613,N_8222);
nor U15222 (N_15222,N_10437,N_10463);
nand U15223 (N_15223,N_11724,N_11160);
nor U15224 (N_15224,N_9961,N_8254);
nand U15225 (N_15225,N_9337,N_11534);
and U15226 (N_15226,N_11376,N_9184);
nor U15227 (N_15227,N_8694,N_10586);
nand U15228 (N_15228,N_8148,N_10802);
and U15229 (N_15229,N_10811,N_8152);
nand U15230 (N_15230,N_9034,N_8222);
nor U15231 (N_15231,N_11031,N_10150);
nor U15232 (N_15232,N_8288,N_9006);
nor U15233 (N_15233,N_10858,N_10158);
or U15234 (N_15234,N_8144,N_11566);
and U15235 (N_15235,N_9978,N_11092);
xor U15236 (N_15236,N_10033,N_10885);
xor U15237 (N_15237,N_8516,N_9346);
or U15238 (N_15238,N_11608,N_8108);
or U15239 (N_15239,N_9899,N_11270);
nor U15240 (N_15240,N_9580,N_11644);
nand U15241 (N_15241,N_9535,N_9252);
and U15242 (N_15242,N_10357,N_9137);
and U15243 (N_15243,N_9330,N_9338);
and U15244 (N_15244,N_8030,N_9887);
and U15245 (N_15245,N_9491,N_11216);
nand U15246 (N_15246,N_10823,N_10453);
nand U15247 (N_15247,N_8079,N_11601);
nor U15248 (N_15248,N_11457,N_10270);
xnor U15249 (N_15249,N_9821,N_9075);
nor U15250 (N_15250,N_11370,N_10968);
nor U15251 (N_15251,N_10645,N_11546);
xnor U15252 (N_15252,N_11508,N_10479);
or U15253 (N_15253,N_10475,N_8668);
and U15254 (N_15254,N_10682,N_9364);
or U15255 (N_15255,N_10191,N_8561);
nor U15256 (N_15256,N_10593,N_11473);
or U15257 (N_15257,N_10328,N_10662);
or U15258 (N_15258,N_8589,N_10969);
and U15259 (N_15259,N_10298,N_11689);
and U15260 (N_15260,N_10281,N_9548);
or U15261 (N_15261,N_8149,N_8448);
or U15262 (N_15262,N_10144,N_10891);
or U15263 (N_15263,N_8175,N_8993);
nand U15264 (N_15264,N_9095,N_9560);
or U15265 (N_15265,N_9552,N_8965);
and U15266 (N_15266,N_10759,N_8167);
and U15267 (N_15267,N_11761,N_11916);
nand U15268 (N_15268,N_9264,N_11066);
nor U15269 (N_15269,N_8695,N_10859);
nor U15270 (N_15270,N_9503,N_8334);
and U15271 (N_15271,N_8960,N_8480);
and U15272 (N_15272,N_10991,N_10164);
xnor U15273 (N_15273,N_8287,N_9599);
nand U15274 (N_15274,N_9191,N_11681);
nor U15275 (N_15275,N_10842,N_11388);
xnor U15276 (N_15276,N_10237,N_8486);
or U15277 (N_15277,N_9145,N_8261);
nor U15278 (N_15278,N_10666,N_9219);
or U15279 (N_15279,N_10479,N_10383);
xnor U15280 (N_15280,N_11547,N_10019);
or U15281 (N_15281,N_10819,N_8096);
and U15282 (N_15282,N_11447,N_9959);
and U15283 (N_15283,N_11448,N_8666);
and U15284 (N_15284,N_9865,N_10417);
xor U15285 (N_15285,N_11906,N_8138);
or U15286 (N_15286,N_10375,N_8967);
xnor U15287 (N_15287,N_10106,N_9214);
xor U15288 (N_15288,N_10227,N_8974);
and U15289 (N_15289,N_10651,N_9416);
xor U15290 (N_15290,N_8705,N_8611);
nor U15291 (N_15291,N_8548,N_11683);
nand U15292 (N_15292,N_9525,N_10800);
or U15293 (N_15293,N_8081,N_9053);
nand U15294 (N_15294,N_11908,N_11427);
xnor U15295 (N_15295,N_8589,N_8432);
nor U15296 (N_15296,N_10140,N_11568);
nor U15297 (N_15297,N_8828,N_8258);
nor U15298 (N_15298,N_8805,N_10398);
xnor U15299 (N_15299,N_11523,N_11879);
or U15300 (N_15300,N_9856,N_10964);
nand U15301 (N_15301,N_8507,N_10994);
or U15302 (N_15302,N_11893,N_10887);
and U15303 (N_15303,N_10168,N_11552);
nor U15304 (N_15304,N_8403,N_9586);
and U15305 (N_15305,N_9119,N_9792);
or U15306 (N_15306,N_11742,N_10292);
nand U15307 (N_15307,N_11726,N_11148);
or U15308 (N_15308,N_8478,N_9972);
nand U15309 (N_15309,N_8839,N_11091);
or U15310 (N_15310,N_10985,N_9997);
or U15311 (N_15311,N_8567,N_10556);
nor U15312 (N_15312,N_10311,N_9170);
xnor U15313 (N_15313,N_8949,N_8314);
nand U15314 (N_15314,N_9427,N_9298);
or U15315 (N_15315,N_9989,N_11965);
and U15316 (N_15316,N_10942,N_11356);
xnor U15317 (N_15317,N_11759,N_8670);
nor U15318 (N_15318,N_10033,N_9131);
and U15319 (N_15319,N_10315,N_9259);
nor U15320 (N_15320,N_10427,N_11618);
nor U15321 (N_15321,N_8527,N_9782);
and U15322 (N_15322,N_8070,N_8947);
nor U15323 (N_15323,N_10381,N_10955);
and U15324 (N_15324,N_9727,N_9819);
and U15325 (N_15325,N_9896,N_11042);
or U15326 (N_15326,N_9653,N_11804);
and U15327 (N_15327,N_9024,N_10939);
xor U15328 (N_15328,N_10567,N_10445);
nand U15329 (N_15329,N_10029,N_8510);
and U15330 (N_15330,N_8358,N_9097);
or U15331 (N_15331,N_8498,N_8386);
nand U15332 (N_15332,N_9060,N_10042);
and U15333 (N_15333,N_11305,N_9089);
or U15334 (N_15334,N_11857,N_11024);
xor U15335 (N_15335,N_11224,N_10441);
or U15336 (N_15336,N_8048,N_10347);
nand U15337 (N_15337,N_8330,N_11272);
or U15338 (N_15338,N_8616,N_9308);
or U15339 (N_15339,N_10144,N_9814);
or U15340 (N_15340,N_8437,N_9527);
nor U15341 (N_15341,N_11201,N_8811);
nor U15342 (N_15342,N_8886,N_9172);
or U15343 (N_15343,N_11986,N_8356);
nand U15344 (N_15344,N_11259,N_9916);
nand U15345 (N_15345,N_9825,N_10360);
or U15346 (N_15346,N_10379,N_11180);
nor U15347 (N_15347,N_10580,N_11707);
xor U15348 (N_15348,N_10709,N_9000);
nor U15349 (N_15349,N_8182,N_11730);
xnor U15350 (N_15350,N_10900,N_8663);
or U15351 (N_15351,N_10446,N_9328);
xor U15352 (N_15352,N_10383,N_8354);
xnor U15353 (N_15353,N_8839,N_8172);
or U15354 (N_15354,N_11826,N_11997);
nand U15355 (N_15355,N_8317,N_10427);
xor U15356 (N_15356,N_11270,N_11800);
nand U15357 (N_15357,N_10350,N_10220);
or U15358 (N_15358,N_8527,N_11481);
nor U15359 (N_15359,N_9651,N_9660);
nand U15360 (N_15360,N_8413,N_10028);
nand U15361 (N_15361,N_10254,N_8463);
nor U15362 (N_15362,N_8231,N_10131);
nor U15363 (N_15363,N_11735,N_11670);
nor U15364 (N_15364,N_11708,N_11514);
nor U15365 (N_15365,N_8599,N_11656);
nor U15366 (N_15366,N_11720,N_11295);
and U15367 (N_15367,N_9619,N_11556);
or U15368 (N_15368,N_9075,N_11873);
nand U15369 (N_15369,N_8308,N_9656);
or U15370 (N_15370,N_9032,N_11978);
and U15371 (N_15371,N_11884,N_10451);
nor U15372 (N_15372,N_8684,N_10681);
xnor U15373 (N_15373,N_11713,N_10362);
nor U15374 (N_15374,N_8319,N_8809);
nor U15375 (N_15375,N_9320,N_8148);
and U15376 (N_15376,N_10764,N_8901);
and U15377 (N_15377,N_11641,N_10838);
or U15378 (N_15378,N_11280,N_8503);
or U15379 (N_15379,N_11287,N_11971);
xnor U15380 (N_15380,N_11811,N_9206);
and U15381 (N_15381,N_9454,N_10338);
or U15382 (N_15382,N_11569,N_10033);
nand U15383 (N_15383,N_10606,N_8627);
or U15384 (N_15384,N_11487,N_9146);
nor U15385 (N_15385,N_8715,N_9424);
xnor U15386 (N_15386,N_8004,N_9006);
and U15387 (N_15387,N_11555,N_11587);
nand U15388 (N_15388,N_9059,N_11534);
nand U15389 (N_15389,N_10030,N_10036);
or U15390 (N_15390,N_11835,N_8464);
or U15391 (N_15391,N_9088,N_8357);
and U15392 (N_15392,N_8189,N_11634);
or U15393 (N_15393,N_9821,N_9123);
nor U15394 (N_15394,N_11726,N_11785);
and U15395 (N_15395,N_10347,N_8686);
nand U15396 (N_15396,N_8728,N_9398);
and U15397 (N_15397,N_10490,N_9743);
and U15398 (N_15398,N_10265,N_8180);
and U15399 (N_15399,N_9271,N_10445);
nand U15400 (N_15400,N_9313,N_8870);
and U15401 (N_15401,N_11122,N_8732);
or U15402 (N_15402,N_11763,N_10724);
nand U15403 (N_15403,N_10497,N_9804);
xnor U15404 (N_15404,N_11571,N_9286);
nor U15405 (N_15405,N_10323,N_10736);
nand U15406 (N_15406,N_10758,N_8066);
or U15407 (N_15407,N_9542,N_10179);
and U15408 (N_15408,N_9393,N_9475);
or U15409 (N_15409,N_11709,N_11459);
nand U15410 (N_15410,N_11708,N_9460);
nand U15411 (N_15411,N_11906,N_10316);
xor U15412 (N_15412,N_8132,N_10090);
nor U15413 (N_15413,N_9201,N_10376);
nor U15414 (N_15414,N_9499,N_11974);
or U15415 (N_15415,N_11880,N_8969);
or U15416 (N_15416,N_11843,N_8805);
or U15417 (N_15417,N_8447,N_9076);
and U15418 (N_15418,N_9863,N_11489);
nor U15419 (N_15419,N_8407,N_9963);
nor U15420 (N_15420,N_10069,N_8871);
and U15421 (N_15421,N_10632,N_9876);
or U15422 (N_15422,N_11728,N_11619);
xnor U15423 (N_15423,N_11467,N_11293);
xor U15424 (N_15424,N_11965,N_9350);
nor U15425 (N_15425,N_10874,N_8525);
nand U15426 (N_15426,N_11327,N_9462);
nand U15427 (N_15427,N_10748,N_9304);
and U15428 (N_15428,N_8455,N_11017);
xnor U15429 (N_15429,N_11242,N_10488);
nand U15430 (N_15430,N_9975,N_8708);
and U15431 (N_15431,N_11532,N_9605);
nor U15432 (N_15432,N_9851,N_9222);
nor U15433 (N_15433,N_9578,N_11979);
nand U15434 (N_15434,N_9118,N_10952);
nor U15435 (N_15435,N_8855,N_9567);
nand U15436 (N_15436,N_8640,N_11591);
xnor U15437 (N_15437,N_9293,N_9068);
and U15438 (N_15438,N_10021,N_10573);
and U15439 (N_15439,N_10428,N_9702);
or U15440 (N_15440,N_11782,N_10522);
nand U15441 (N_15441,N_11001,N_11411);
and U15442 (N_15442,N_9533,N_10755);
nand U15443 (N_15443,N_9648,N_9537);
xor U15444 (N_15444,N_8375,N_9588);
nand U15445 (N_15445,N_9900,N_8503);
nand U15446 (N_15446,N_10210,N_8212);
nand U15447 (N_15447,N_9878,N_9702);
nor U15448 (N_15448,N_9109,N_11956);
nand U15449 (N_15449,N_10895,N_8306);
or U15450 (N_15450,N_8397,N_10382);
xnor U15451 (N_15451,N_10858,N_10307);
xnor U15452 (N_15452,N_10251,N_11448);
nor U15453 (N_15453,N_10378,N_9255);
and U15454 (N_15454,N_11793,N_8630);
nor U15455 (N_15455,N_11232,N_11646);
and U15456 (N_15456,N_9344,N_11130);
or U15457 (N_15457,N_9425,N_10726);
xor U15458 (N_15458,N_10202,N_10485);
xnor U15459 (N_15459,N_9725,N_11914);
and U15460 (N_15460,N_9029,N_10077);
and U15461 (N_15461,N_8234,N_9138);
or U15462 (N_15462,N_9061,N_10147);
nor U15463 (N_15463,N_9700,N_9466);
nand U15464 (N_15464,N_10271,N_8868);
nor U15465 (N_15465,N_9075,N_8408);
or U15466 (N_15466,N_11446,N_8167);
or U15467 (N_15467,N_10529,N_8190);
nand U15468 (N_15468,N_8191,N_9060);
and U15469 (N_15469,N_10836,N_9852);
and U15470 (N_15470,N_11192,N_11921);
nor U15471 (N_15471,N_11641,N_9514);
and U15472 (N_15472,N_8907,N_9719);
nor U15473 (N_15473,N_10865,N_11014);
xor U15474 (N_15474,N_9612,N_8102);
or U15475 (N_15475,N_10823,N_9664);
or U15476 (N_15476,N_9530,N_11650);
and U15477 (N_15477,N_8623,N_9156);
nor U15478 (N_15478,N_11765,N_10582);
nor U15479 (N_15479,N_8684,N_9647);
or U15480 (N_15480,N_8472,N_10374);
and U15481 (N_15481,N_8189,N_10024);
xnor U15482 (N_15482,N_10203,N_8011);
nand U15483 (N_15483,N_10343,N_9153);
nand U15484 (N_15484,N_8296,N_8783);
nor U15485 (N_15485,N_10865,N_11918);
nor U15486 (N_15486,N_8911,N_9786);
nor U15487 (N_15487,N_11084,N_8396);
or U15488 (N_15488,N_11717,N_8748);
and U15489 (N_15489,N_11867,N_11813);
nand U15490 (N_15490,N_8395,N_10117);
or U15491 (N_15491,N_9444,N_9855);
and U15492 (N_15492,N_10940,N_11676);
nor U15493 (N_15493,N_10603,N_11814);
xor U15494 (N_15494,N_9782,N_9228);
nor U15495 (N_15495,N_9212,N_9941);
nand U15496 (N_15496,N_8658,N_8022);
nor U15497 (N_15497,N_11082,N_11857);
and U15498 (N_15498,N_9484,N_8030);
nor U15499 (N_15499,N_11143,N_11230);
or U15500 (N_15500,N_9862,N_9307);
and U15501 (N_15501,N_10966,N_10290);
or U15502 (N_15502,N_11040,N_11436);
nor U15503 (N_15503,N_10571,N_9690);
nand U15504 (N_15504,N_11427,N_8346);
nor U15505 (N_15505,N_9260,N_9898);
nand U15506 (N_15506,N_8070,N_8014);
nand U15507 (N_15507,N_11090,N_8896);
and U15508 (N_15508,N_8314,N_10923);
nor U15509 (N_15509,N_8194,N_9225);
or U15510 (N_15510,N_8534,N_9908);
or U15511 (N_15511,N_8495,N_11439);
nand U15512 (N_15512,N_10570,N_11305);
and U15513 (N_15513,N_9343,N_11681);
or U15514 (N_15514,N_9518,N_10786);
nor U15515 (N_15515,N_8331,N_11638);
nand U15516 (N_15516,N_8735,N_9359);
nor U15517 (N_15517,N_10829,N_10621);
and U15518 (N_15518,N_10549,N_10297);
xor U15519 (N_15519,N_10674,N_10041);
nand U15520 (N_15520,N_11432,N_9869);
and U15521 (N_15521,N_11930,N_10740);
xnor U15522 (N_15522,N_9154,N_8555);
nor U15523 (N_15523,N_8275,N_8566);
or U15524 (N_15524,N_8090,N_9743);
xor U15525 (N_15525,N_8474,N_8716);
nor U15526 (N_15526,N_8456,N_8588);
nor U15527 (N_15527,N_9738,N_11397);
nor U15528 (N_15528,N_10502,N_9474);
xnor U15529 (N_15529,N_9222,N_8251);
or U15530 (N_15530,N_9110,N_9298);
xor U15531 (N_15531,N_9313,N_10599);
nand U15532 (N_15532,N_8298,N_9361);
nor U15533 (N_15533,N_10064,N_10794);
or U15534 (N_15534,N_8997,N_11087);
nor U15535 (N_15535,N_11230,N_9469);
nor U15536 (N_15536,N_11397,N_9563);
nor U15537 (N_15537,N_8900,N_11860);
or U15538 (N_15538,N_10913,N_9960);
nor U15539 (N_15539,N_11567,N_8948);
and U15540 (N_15540,N_10751,N_11623);
nor U15541 (N_15541,N_10926,N_9015);
or U15542 (N_15542,N_11313,N_9516);
nand U15543 (N_15543,N_10786,N_9388);
nor U15544 (N_15544,N_11722,N_10816);
nor U15545 (N_15545,N_9914,N_9864);
or U15546 (N_15546,N_8313,N_11060);
and U15547 (N_15547,N_10399,N_11498);
xor U15548 (N_15548,N_11388,N_9169);
and U15549 (N_15549,N_9034,N_8200);
or U15550 (N_15550,N_8253,N_10759);
nand U15551 (N_15551,N_8730,N_11730);
xnor U15552 (N_15552,N_10022,N_11802);
nor U15553 (N_15553,N_10192,N_10914);
nand U15554 (N_15554,N_11494,N_9429);
xnor U15555 (N_15555,N_8748,N_11813);
nor U15556 (N_15556,N_8113,N_8579);
nand U15557 (N_15557,N_9917,N_8617);
nor U15558 (N_15558,N_9652,N_9998);
or U15559 (N_15559,N_8572,N_10537);
xor U15560 (N_15560,N_10539,N_9746);
nor U15561 (N_15561,N_11769,N_11922);
and U15562 (N_15562,N_10116,N_9579);
and U15563 (N_15563,N_10971,N_8027);
nand U15564 (N_15564,N_11354,N_9480);
or U15565 (N_15565,N_8205,N_8896);
nor U15566 (N_15566,N_11099,N_9193);
nand U15567 (N_15567,N_8113,N_9087);
xnor U15568 (N_15568,N_10519,N_10371);
and U15569 (N_15569,N_11498,N_11733);
and U15570 (N_15570,N_8631,N_9066);
nor U15571 (N_15571,N_9565,N_8634);
and U15572 (N_15572,N_10903,N_11227);
xnor U15573 (N_15573,N_8594,N_11861);
nand U15574 (N_15574,N_11825,N_10085);
and U15575 (N_15575,N_10093,N_8350);
and U15576 (N_15576,N_10750,N_11707);
nand U15577 (N_15577,N_11907,N_10400);
nor U15578 (N_15578,N_11730,N_9951);
xor U15579 (N_15579,N_10929,N_10741);
nand U15580 (N_15580,N_8859,N_8642);
or U15581 (N_15581,N_10916,N_8425);
and U15582 (N_15582,N_9864,N_11598);
nor U15583 (N_15583,N_8807,N_9978);
nand U15584 (N_15584,N_8272,N_10685);
nand U15585 (N_15585,N_9782,N_8365);
nor U15586 (N_15586,N_11727,N_10786);
and U15587 (N_15587,N_8815,N_9118);
and U15588 (N_15588,N_11885,N_10924);
or U15589 (N_15589,N_8108,N_9276);
nor U15590 (N_15590,N_10323,N_10876);
nand U15591 (N_15591,N_10391,N_11676);
or U15592 (N_15592,N_11147,N_10021);
and U15593 (N_15593,N_11739,N_8290);
or U15594 (N_15594,N_8108,N_10835);
xor U15595 (N_15595,N_10704,N_9605);
nor U15596 (N_15596,N_9065,N_9663);
nand U15597 (N_15597,N_10599,N_10905);
nor U15598 (N_15598,N_11746,N_9869);
nor U15599 (N_15599,N_8656,N_8746);
and U15600 (N_15600,N_9000,N_8740);
and U15601 (N_15601,N_11253,N_8871);
and U15602 (N_15602,N_11279,N_8728);
xnor U15603 (N_15603,N_9083,N_11118);
xnor U15604 (N_15604,N_11691,N_10971);
or U15605 (N_15605,N_8456,N_11266);
nor U15606 (N_15606,N_9727,N_10594);
and U15607 (N_15607,N_11218,N_10017);
and U15608 (N_15608,N_10242,N_10512);
nor U15609 (N_15609,N_9456,N_11621);
or U15610 (N_15610,N_9503,N_8528);
or U15611 (N_15611,N_11535,N_8784);
and U15612 (N_15612,N_10930,N_9827);
and U15613 (N_15613,N_8074,N_10893);
nor U15614 (N_15614,N_9582,N_11592);
nor U15615 (N_15615,N_9873,N_11032);
or U15616 (N_15616,N_11759,N_8414);
xor U15617 (N_15617,N_9890,N_9331);
nand U15618 (N_15618,N_11503,N_11609);
nor U15619 (N_15619,N_10450,N_10334);
and U15620 (N_15620,N_11042,N_8813);
xor U15621 (N_15621,N_8573,N_10190);
and U15622 (N_15622,N_11402,N_8485);
xnor U15623 (N_15623,N_9835,N_10222);
and U15624 (N_15624,N_10384,N_8140);
nand U15625 (N_15625,N_11574,N_8140);
nor U15626 (N_15626,N_11589,N_9883);
nand U15627 (N_15627,N_9000,N_10145);
and U15628 (N_15628,N_8882,N_9415);
nor U15629 (N_15629,N_8276,N_11174);
and U15630 (N_15630,N_8524,N_10328);
nand U15631 (N_15631,N_9760,N_9608);
or U15632 (N_15632,N_10046,N_10669);
xnor U15633 (N_15633,N_10925,N_8928);
and U15634 (N_15634,N_11393,N_11381);
or U15635 (N_15635,N_9678,N_10872);
nand U15636 (N_15636,N_10536,N_11436);
and U15637 (N_15637,N_10774,N_8945);
or U15638 (N_15638,N_10242,N_9486);
or U15639 (N_15639,N_9957,N_11969);
or U15640 (N_15640,N_8028,N_11243);
xnor U15641 (N_15641,N_9508,N_8059);
nand U15642 (N_15642,N_11309,N_11166);
nand U15643 (N_15643,N_9162,N_10129);
xor U15644 (N_15644,N_9572,N_8789);
nand U15645 (N_15645,N_8707,N_10543);
or U15646 (N_15646,N_8923,N_8461);
nand U15647 (N_15647,N_9045,N_10760);
nor U15648 (N_15648,N_8695,N_10415);
xor U15649 (N_15649,N_11146,N_10697);
or U15650 (N_15650,N_10536,N_8835);
nand U15651 (N_15651,N_9602,N_11196);
or U15652 (N_15652,N_11062,N_9133);
nand U15653 (N_15653,N_11835,N_9588);
xor U15654 (N_15654,N_11396,N_10481);
or U15655 (N_15655,N_8478,N_11228);
nand U15656 (N_15656,N_9779,N_8844);
and U15657 (N_15657,N_11176,N_10940);
or U15658 (N_15658,N_11838,N_9517);
and U15659 (N_15659,N_11757,N_11335);
nand U15660 (N_15660,N_9904,N_10185);
nand U15661 (N_15661,N_9724,N_10526);
or U15662 (N_15662,N_9447,N_10498);
or U15663 (N_15663,N_8966,N_11007);
nor U15664 (N_15664,N_8768,N_10225);
or U15665 (N_15665,N_11598,N_11313);
or U15666 (N_15666,N_10625,N_8145);
xnor U15667 (N_15667,N_11700,N_10860);
nor U15668 (N_15668,N_8108,N_8407);
or U15669 (N_15669,N_11326,N_11513);
or U15670 (N_15670,N_9908,N_10079);
xor U15671 (N_15671,N_11366,N_10061);
nor U15672 (N_15672,N_11391,N_10489);
and U15673 (N_15673,N_11287,N_11010);
nand U15674 (N_15674,N_10231,N_10118);
and U15675 (N_15675,N_8584,N_8033);
or U15676 (N_15676,N_10210,N_11540);
nand U15677 (N_15677,N_9063,N_10934);
nand U15678 (N_15678,N_8258,N_9584);
or U15679 (N_15679,N_11441,N_9867);
xnor U15680 (N_15680,N_9708,N_11344);
nor U15681 (N_15681,N_10465,N_8439);
nor U15682 (N_15682,N_11376,N_11851);
nor U15683 (N_15683,N_11940,N_10378);
nand U15684 (N_15684,N_11325,N_11431);
nand U15685 (N_15685,N_11896,N_11682);
nor U15686 (N_15686,N_11466,N_8862);
or U15687 (N_15687,N_10203,N_9698);
nand U15688 (N_15688,N_9936,N_9823);
and U15689 (N_15689,N_10669,N_10159);
or U15690 (N_15690,N_8906,N_8370);
nand U15691 (N_15691,N_9021,N_8330);
nor U15692 (N_15692,N_8691,N_9832);
nand U15693 (N_15693,N_11315,N_9839);
or U15694 (N_15694,N_9712,N_8173);
or U15695 (N_15695,N_8409,N_9176);
or U15696 (N_15696,N_9199,N_8203);
or U15697 (N_15697,N_10911,N_11974);
or U15698 (N_15698,N_10646,N_8001);
and U15699 (N_15699,N_11874,N_11722);
and U15700 (N_15700,N_10506,N_9392);
nand U15701 (N_15701,N_8115,N_10707);
and U15702 (N_15702,N_11660,N_8781);
or U15703 (N_15703,N_11888,N_10501);
xnor U15704 (N_15704,N_10941,N_8090);
nor U15705 (N_15705,N_8471,N_8219);
and U15706 (N_15706,N_9097,N_11182);
or U15707 (N_15707,N_9022,N_9735);
and U15708 (N_15708,N_10918,N_10674);
or U15709 (N_15709,N_8311,N_8727);
nor U15710 (N_15710,N_8537,N_8138);
nor U15711 (N_15711,N_10286,N_8709);
nor U15712 (N_15712,N_9654,N_8802);
nor U15713 (N_15713,N_10333,N_10077);
and U15714 (N_15714,N_9349,N_11994);
and U15715 (N_15715,N_11395,N_10816);
nand U15716 (N_15716,N_9222,N_10400);
or U15717 (N_15717,N_8132,N_8738);
nor U15718 (N_15718,N_9019,N_11719);
nor U15719 (N_15719,N_10805,N_9320);
nor U15720 (N_15720,N_8330,N_10809);
nor U15721 (N_15721,N_8325,N_10145);
nand U15722 (N_15722,N_9486,N_8803);
and U15723 (N_15723,N_9126,N_9872);
nor U15724 (N_15724,N_9432,N_9869);
and U15725 (N_15725,N_11790,N_10546);
and U15726 (N_15726,N_11798,N_10850);
nand U15727 (N_15727,N_9333,N_11952);
or U15728 (N_15728,N_8263,N_9341);
xor U15729 (N_15729,N_11738,N_8345);
or U15730 (N_15730,N_11323,N_9823);
and U15731 (N_15731,N_10169,N_9905);
or U15732 (N_15732,N_8679,N_11627);
nor U15733 (N_15733,N_9736,N_9597);
nor U15734 (N_15734,N_11052,N_10886);
nand U15735 (N_15735,N_9904,N_10740);
or U15736 (N_15736,N_11463,N_10909);
or U15737 (N_15737,N_9726,N_8521);
or U15738 (N_15738,N_8213,N_11009);
nand U15739 (N_15739,N_8590,N_8815);
nor U15740 (N_15740,N_9907,N_10349);
nand U15741 (N_15741,N_9647,N_10948);
and U15742 (N_15742,N_9046,N_9700);
nand U15743 (N_15743,N_10622,N_11376);
nor U15744 (N_15744,N_10948,N_10236);
xor U15745 (N_15745,N_8636,N_11087);
nand U15746 (N_15746,N_8770,N_11799);
nand U15747 (N_15747,N_8710,N_10163);
nand U15748 (N_15748,N_9311,N_8917);
xor U15749 (N_15749,N_11624,N_9415);
and U15750 (N_15750,N_8502,N_10357);
or U15751 (N_15751,N_9316,N_8566);
nand U15752 (N_15752,N_10715,N_8892);
nor U15753 (N_15753,N_9583,N_11830);
nor U15754 (N_15754,N_9896,N_10533);
nor U15755 (N_15755,N_9107,N_10732);
nand U15756 (N_15756,N_9653,N_8785);
xnor U15757 (N_15757,N_8893,N_11292);
nor U15758 (N_15758,N_10532,N_8144);
or U15759 (N_15759,N_8862,N_10089);
nand U15760 (N_15760,N_8527,N_10181);
and U15761 (N_15761,N_9551,N_8318);
nand U15762 (N_15762,N_11702,N_10446);
nand U15763 (N_15763,N_8109,N_8084);
nand U15764 (N_15764,N_8544,N_8822);
or U15765 (N_15765,N_11895,N_8783);
nand U15766 (N_15766,N_10516,N_8214);
and U15767 (N_15767,N_10796,N_9756);
or U15768 (N_15768,N_11616,N_10003);
nor U15769 (N_15769,N_11419,N_9499);
nor U15770 (N_15770,N_9708,N_8946);
nand U15771 (N_15771,N_9556,N_9506);
and U15772 (N_15772,N_9125,N_11284);
or U15773 (N_15773,N_11676,N_8981);
and U15774 (N_15774,N_8250,N_9154);
nand U15775 (N_15775,N_8986,N_9180);
or U15776 (N_15776,N_9867,N_11263);
and U15777 (N_15777,N_11683,N_10585);
nand U15778 (N_15778,N_8558,N_8603);
nor U15779 (N_15779,N_11583,N_11546);
nand U15780 (N_15780,N_9870,N_10173);
nand U15781 (N_15781,N_10212,N_10600);
or U15782 (N_15782,N_8125,N_11542);
nor U15783 (N_15783,N_9167,N_8336);
xnor U15784 (N_15784,N_8795,N_11161);
and U15785 (N_15785,N_8673,N_9252);
nor U15786 (N_15786,N_9570,N_10003);
nor U15787 (N_15787,N_11827,N_9066);
or U15788 (N_15788,N_8793,N_8996);
nor U15789 (N_15789,N_9263,N_10474);
nor U15790 (N_15790,N_9049,N_10577);
nor U15791 (N_15791,N_8791,N_9664);
or U15792 (N_15792,N_11261,N_11064);
nor U15793 (N_15793,N_11172,N_9901);
nor U15794 (N_15794,N_11832,N_8791);
and U15795 (N_15795,N_9950,N_8909);
nor U15796 (N_15796,N_9378,N_11909);
nand U15797 (N_15797,N_10542,N_10011);
or U15798 (N_15798,N_10393,N_8556);
nand U15799 (N_15799,N_11147,N_9335);
or U15800 (N_15800,N_11051,N_10186);
nor U15801 (N_15801,N_8332,N_10283);
or U15802 (N_15802,N_8359,N_9617);
nor U15803 (N_15803,N_10604,N_10248);
or U15804 (N_15804,N_10524,N_11384);
and U15805 (N_15805,N_11887,N_8597);
or U15806 (N_15806,N_8196,N_8749);
and U15807 (N_15807,N_9070,N_8855);
nor U15808 (N_15808,N_9747,N_11611);
xor U15809 (N_15809,N_10984,N_8966);
or U15810 (N_15810,N_10433,N_10197);
nand U15811 (N_15811,N_8856,N_11949);
xnor U15812 (N_15812,N_11071,N_8828);
nand U15813 (N_15813,N_10657,N_11494);
and U15814 (N_15814,N_9563,N_9179);
and U15815 (N_15815,N_9819,N_9394);
nand U15816 (N_15816,N_10332,N_11655);
or U15817 (N_15817,N_8813,N_11251);
nand U15818 (N_15818,N_11466,N_11622);
and U15819 (N_15819,N_10632,N_9777);
nand U15820 (N_15820,N_9605,N_8452);
or U15821 (N_15821,N_10632,N_10427);
or U15822 (N_15822,N_8658,N_9383);
nor U15823 (N_15823,N_8172,N_10711);
nor U15824 (N_15824,N_11197,N_11728);
or U15825 (N_15825,N_10280,N_9495);
or U15826 (N_15826,N_9313,N_8744);
or U15827 (N_15827,N_9884,N_11888);
nor U15828 (N_15828,N_9146,N_10133);
and U15829 (N_15829,N_10045,N_9986);
nand U15830 (N_15830,N_9381,N_8800);
or U15831 (N_15831,N_11025,N_11105);
nor U15832 (N_15832,N_9567,N_11480);
and U15833 (N_15833,N_9404,N_11349);
xor U15834 (N_15834,N_8496,N_9883);
or U15835 (N_15835,N_10104,N_8982);
and U15836 (N_15836,N_11675,N_10793);
nand U15837 (N_15837,N_9750,N_9814);
nor U15838 (N_15838,N_9565,N_10145);
nor U15839 (N_15839,N_9847,N_8517);
or U15840 (N_15840,N_11270,N_10483);
or U15841 (N_15841,N_9465,N_9824);
xor U15842 (N_15842,N_9655,N_11670);
xor U15843 (N_15843,N_9814,N_10201);
or U15844 (N_15844,N_11174,N_8462);
xnor U15845 (N_15845,N_8205,N_11101);
nand U15846 (N_15846,N_11238,N_9233);
or U15847 (N_15847,N_11818,N_10135);
or U15848 (N_15848,N_11010,N_10728);
nor U15849 (N_15849,N_11483,N_11283);
or U15850 (N_15850,N_8343,N_9213);
xor U15851 (N_15851,N_8690,N_11208);
and U15852 (N_15852,N_8239,N_9125);
and U15853 (N_15853,N_11529,N_10083);
nor U15854 (N_15854,N_11751,N_9650);
nor U15855 (N_15855,N_8762,N_11427);
nor U15856 (N_15856,N_11844,N_8365);
xnor U15857 (N_15857,N_10552,N_9593);
nand U15858 (N_15858,N_11959,N_10885);
or U15859 (N_15859,N_11602,N_9982);
or U15860 (N_15860,N_10344,N_8446);
and U15861 (N_15861,N_11167,N_10380);
and U15862 (N_15862,N_11048,N_10990);
or U15863 (N_15863,N_9956,N_11822);
or U15864 (N_15864,N_8855,N_11694);
nor U15865 (N_15865,N_10567,N_10127);
nand U15866 (N_15866,N_10325,N_9252);
and U15867 (N_15867,N_9686,N_8681);
or U15868 (N_15868,N_10129,N_9765);
nand U15869 (N_15869,N_9138,N_9862);
nand U15870 (N_15870,N_11645,N_11866);
or U15871 (N_15871,N_11017,N_9314);
and U15872 (N_15872,N_11637,N_11706);
or U15873 (N_15873,N_9096,N_8497);
or U15874 (N_15874,N_10819,N_9480);
and U15875 (N_15875,N_10763,N_8429);
or U15876 (N_15876,N_8979,N_8546);
nor U15877 (N_15877,N_10849,N_9770);
nor U15878 (N_15878,N_10464,N_10216);
nand U15879 (N_15879,N_10617,N_10186);
nor U15880 (N_15880,N_11761,N_9810);
xnor U15881 (N_15881,N_9290,N_9399);
and U15882 (N_15882,N_11071,N_11159);
nor U15883 (N_15883,N_10861,N_9503);
nor U15884 (N_15884,N_11392,N_8289);
nor U15885 (N_15885,N_8370,N_9219);
nand U15886 (N_15886,N_11205,N_8652);
and U15887 (N_15887,N_9105,N_8283);
or U15888 (N_15888,N_11832,N_8739);
nand U15889 (N_15889,N_11579,N_8930);
nand U15890 (N_15890,N_10922,N_8525);
and U15891 (N_15891,N_8151,N_10687);
or U15892 (N_15892,N_8414,N_8793);
and U15893 (N_15893,N_11633,N_9792);
and U15894 (N_15894,N_10509,N_8920);
and U15895 (N_15895,N_9515,N_11099);
nand U15896 (N_15896,N_9720,N_9678);
nor U15897 (N_15897,N_8099,N_9910);
or U15898 (N_15898,N_9775,N_9164);
nor U15899 (N_15899,N_9474,N_9302);
or U15900 (N_15900,N_10431,N_10024);
or U15901 (N_15901,N_8976,N_9273);
or U15902 (N_15902,N_10255,N_9319);
nand U15903 (N_15903,N_8158,N_8726);
nand U15904 (N_15904,N_9829,N_8311);
and U15905 (N_15905,N_11489,N_8152);
and U15906 (N_15906,N_8795,N_8692);
nand U15907 (N_15907,N_8116,N_8392);
or U15908 (N_15908,N_11384,N_9112);
nor U15909 (N_15909,N_10828,N_11160);
xor U15910 (N_15910,N_11596,N_8842);
or U15911 (N_15911,N_8955,N_8368);
xor U15912 (N_15912,N_10063,N_9341);
and U15913 (N_15913,N_9297,N_9559);
nor U15914 (N_15914,N_10324,N_10382);
or U15915 (N_15915,N_10328,N_8361);
nor U15916 (N_15916,N_10303,N_8333);
or U15917 (N_15917,N_10583,N_10440);
or U15918 (N_15918,N_11810,N_8364);
and U15919 (N_15919,N_8268,N_10712);
nor U15920 (N_15920,N_8629,N_8378);
or U15921 (N_15921,N_10417,N_8198);
xnor U15922 (N_15922,N_11983,N_10115);
or U15923 (N_15923,N_8853,N_11316);
or U15924 (N_15924,N_10456,N_8283);
nand U15925 (N_15925,N_10024,N_8380);
nor U15926 (N_15926,N_11015,N_11991);
or U15927 (N_15927,N_11856,N_8469);
nand U15928 (N_15928,N_11260,N_8404);
nand U15929 (N_15929,N_11141,N_8758);
nor U15930 (N_15930,N_9840,N_9739);
and U15931 (N_15931,N_11725,N_9324);
nor U15932 (N_15932,N_9049,N_10771);
nand U15933 (N_15933,N_10930,N_10802);
or U15934 (N_15934,N_8723,N_8621);
nand U15935 (N_15935,N_8978,N_9416);
nand U15936 (N_15936,N_10711,N_11524);
nand U15937 (N_15937,N_9430,N_11745);
nor U15938 (N_15938,N_8955,N_8222);
nand U15939 (N_15939,N_9212,N_9804);
nand U15940 (N_15940,N_8864,N_10795);
and U15941 (N_15941,N_10532,N_11752);
or U15942 (N_15942,N_9683,N_10674);
and U15943 (N_15943,N_10770,N_9059);
nand U15944 (N_15944,N_10208,N_9587);
nor U15945 (N_15945,N_11584,N_11967);
nand U15946 (N_15946,N_11900,N_8521);
or U15947 (N_15947,N_11835,N_9698);
and U15948 (N_15948,N_9364,N_8819);
nor U15949 (N_15949,N_11842,N_11293);
and U15950 (N_15950,N_8352,N_11990);
or U15951 (N_15951,N_9473,N_9052);
nor U15952 (N_15952,N_8807,N_8307);
nand U15953 (N_15953,N_11963,N_9976);
or U15954 (N_15954,N_9957,N_9755);
or U15955 (N_15955,N_9248,N_11818);
and U15956 (N_15956,N_9696,N_11964);
nor U15957 (N_15957,N_11556,N_9931);
and U15958 (N_15958,N_11332,N_11869);
nor U15959 (N_15959,N_10858,N_8657);
nor U15960 (N_15960,N_9725,N_8471);
and U15961 (N_15961,N_9847,N_8356);
nand U15962 (N_15962,N_9288,N_8632);
nand U15963 (N_15963,N_11000,N_8394);
and U15964 (N_15964,N_9154,N_9203);
nor U15965 (N_15965,N_8191,N_10999);
xnor U15966 (N_15966,N_11718,N_8961);
or U15967 (N_15967,N_9246,N_9173);
and U15968 (N_15968,N_10902,N_8382);
or U15969 (N_15969,N_8494,N_10384);
or U15970 (N_15970,N_10478,N_10921);
xor U15971 (N_15971,N_9080,N_9136);
nor U15972 (N_15972,N_11700,N_8408);
and U15973 (N_15973,N_8159,N_8352);
and U15974 (N_15974,N_10106,N_8036);
nor U15975 (N_15975,N_10773,N_11436);
xor U15976 (N_15976,N_11370,N_8893);
nand U15977 (N_15977,N_9673,N_9701);
and U15978 (N_15978,N_8403,N_11291);
and U15979 (N_15979,N_8356,N_10006);
or U15980 (N_15980,N_10926,N_9457);
nand U15981 (N_15981,N_8344,N_8296);
nor U15982 (N_15982,N_8553,N_10925);
or U15983 (N_15983,N_10424,N_10953);
nor U15984 (N_15984,N_10548,N_8362);
nand U15985 (N_15985,N_10120,N_10608);
nand U15986 (N_15986,N_11446,N_11959);
or U15987 (N_15987,N_9847,N_8855);
nor U15988 (N_15988,N_11106,N_9199);
or U15989 (N_15989,N_10878,N_8431);
xor U15990 (N_15990,N_8481,N_8986);
nor U15991 (N_15991,N_9495,N_9536);
and U15992 (N_15992,N_8785,N_8533);
and U15993 (N_15993,N_11895,N_11724);
nand U15994 (N_15994,N_9315,N_9273);
nor U15995 (N_15995,N_11336,N_10785);
nor U15996 (N_15996,N_10550,N_8462);
and U15997 (N_15997,N_9106,N_9009);
or U15998 (N_15998,N_9776,N_8624);
or U15999 (N_15999,N_8161,N_8165);
or U16000 (N_16000,N_15338,N_15422);
nand U16001 (N_16001,N_15109,N_14595);
nor U16002 (N_16002,N_14330,N_13017);
nand U16003 (N_16003,N_12006,N_12743);
nor U16004 (N_16004,N_15264,N_15611);
nor U16005 (N_16005,N_14229,N_13454);
nor U16006 (N_16006,N_13163,N_15220);
nand U16007 (N_16007,N_14814,N_14018);
nand U16008 (N_16008,N_14806,N_12486);
and U16009 (N_16009,N_15533,N_15067);
nand U16010 (N_16010,N_14833,N_14775);
or U16011 (N_16011,N_14510,N_14299);
and U16012 (N_16012,N_13652,N_14365);
nand U16013 (N_16013,N_13190,N_15224);
nor U16014 (N_16014,N_15580,N_14934);
and U16015 (N_16015,N_14070,N_15794);
nand U16016 (N_16016,N_15496,N_14618);
xnor U16017 (N_16017,N_14863,N_15071);
xnor U16018 (N_16018,N_14946,N_12101);
xor U16019 (N_16019,N_12253,N_13626);
and U16020 (N_16020,N_12352,N_12891);
or U16021 (N_16021,N_14243,N_13380);
or U16022 (N_16022,N_13110,N_12808);
or U16023 (N_16023,N_12497,N_13134);
or U16024 (N_16024,N_13693,N_14706);
xor U16025 (N_16025,N_13650,N_14060);
nand U16026 (N_16026,N_14849,N_15810);
nand U16027 (N_16027,N_15487,N_14826);
or U16028 (N_16028,N_15500,N_15107);
or U16029 (N_16029,N_14388,N_12385);
or U16030 (N_16030,N_13765,N_12334);
and U16031 (N_16031,N_13420,N_12060);
nand U16032 (N_16032,N_14281,N_12027);
nand U16033 (N_16033,N_15767,N_12750);
xor U16034 (N_16034,N_14100,N_14959);
nor U16035 (N_16035,N_15193,N_14000);
and U16036 (N_16036,N_13256,N_13273);
xor U16037 (N_16037,N_12045,N_12211);
and U16038 (N_16038,N_15662,N_13522);
or U16039 (N_16039,N_14160,N_12168);
or U16040 (N_16040,N_14976,N_12143);
or U16041 (N_16041,N_13629,N_13744);
nand U16042 (N_16042,N_12389,N_14444);
nor U16043 (N_16043,N_14542,N_13912);
and U16044 (N_16044,N_14106,N_14237);
or U16045 (N_16045,N_12462,N_12179);
nor U16046 (N_16046,N_15212,N_13392);
and U16047 (N_16047,N_12766,N_14025);
and U16048 (N_16048,N_15238,N_14024);
nor U16049 (N_16049,N_13731,N_14581);
nand U16050 (N_16050,N_13569,N_14817);
nor U16051 (N_16051,N_14749,N_12569);
nand U16052 (N_16052,N_14065,N_12853);
or U16053 (N_16053,N_14726,N_15476);
and U16054 (N_16054,N_12991,N_14327);
and U16055 (N_16055,N_14439,N_12845);
nor U16056 (N_16056,N_13007,N_12167);
nand U16057 (N_16057,N_14906,N_13348);
nand U16058 (N_16058,N_15166,N_12559);
nor U16059 (N_16059,N_12841,N_13145);
nand U16060 (N_16060,N_15684,N_15352);
and U16061 (N_16061,N_14443,N_15625);
and U16062 (N_16062,N_15255,N_14851);
or U16063 (N_16063,N_12884,N_12321);
and U16064 (N_16064,N_12964,N_13700);
and U16065 (N_16065,N_13516,N_12860);
xor U16066 (N_16066,N_15572,N_12127);
xor U16067 (N_16067,N_15630,N_15734);
and U16068 (N_16068,N_13992,N_13651);
xnor U16069 (N_16069,N_12344,N_15041);
nor U16070 (N_16070,N_15294,N_13265);
and U16071 (N_16071,N_13571,N_15874);
nor U16072 (N_16072,N_15781,N_15965);
and U16073 (N_16073,N_13597,N_14297);
nor U16074 (N_16074,N_12975,N_13185);
or U16075 (N_16075,N_15601,N_14455);
and U16076 (N_16076,N_15498,N_15334);
and U16077 (N_16077,N_14489,N_13328);
nor U16078 (N_16078,N_13258,N_13051);
or U16079 (N_16079,N_14614,N_12191);
or U16080 (N_16080,N_15010,N_13404);
nand U16081 (N_16081,N_13409,N_13010);
nor U16082 (N_16082,N_13451,N_13029);
and U16083 (N_16083,N_14175,N_15455);
and U16084 (N_16084,N_15605,N_12839);
and U16085 (N_16085,N_14720,N_13077);
nor U16086 (N_16086,N_13776,N_13524);
and U16087 (N_16087,N_15800,N_13779);
nor U16088 (N_16088,N_13786,N_12250);
and U16089 (N_16089,N_13669,N_14232);
nor U16090 (N_16090,N_14421,N_13115);
nor U16091 (N_16091,N_14820,N_15353);
and U16092 (N_16092,N_15447,N_15218);
nor U16093 (N_16093,N_15236,N_14370);
xnor U16094 (N_16094,N_14066,N_13961);
and U16095 (N_16095,N_13488,N_14957);
or U16096 (N_16096,N_15813,N_13839);
nand U16097 (N_16097,N_15252,N_13216);
and U16098 (N_16098,N_14326,N_13820);
and U16099 (N_16099,N_15749,N_13098);
or U16100 (N_16100,N_12647,N_14710);
and U16101 (N_16101,N_14046,N_13493);
and U16102 (N_16102,N_13337,N_15791);
nand U16103 (N_16103,N_14801,N_15714);
nor U16104 (N_16104,N_14717,N_12069);
and U16105 (N_16105,N_13986,N_15648);
nor U16106 (N_16106,N_13898,N_14225);
and U16107 (N_16107,N_12986,N_14042);
and U16108 (N_16108,N_14377,N_13095);
or U16109 (N_16109,N_13641,N_12171);
xor U16110 (N_16110,N_13170,N_12567);
nor U16111 (N_16111,N_15708,N_15124);
or U16112 (N_16112,N_14150,N_13906);
nand U16113 (N_16113,N_14051,N_14883);
nand U16114 (N_16114,N_12402,N_15511);
nor U16115 (N_16115,N_14955,N_12077);
or U16116 (N_16116,N_13657,N_12166);
or U16117 (N_16117,N_15545,N_14763);
or U16118 (N_16118,N_12008,N_15406);
xor U16119 (N_16119,N_15310,N_13993);
xor U16120 (N_16120,N_13772,N_12652);
xnor U16121 (N_16121,N_13654,N_14908);
and U16122 (N_16122,N_15509,N_14875);
or U16123 (N_16123,N_14156,N_13477);
nor U16124 (N_16124,N_12565,N_15348);
and U16125 (N_16125,N_14292,N_14916);
and U16126 (N_16126,N_12675,N_13585);
xor U16127 (N_16127,N_14651,N_12295);
or U16128 (N_16128,N_14274,N_13685);
nor U16129 (N_16129,N_15633,N_12798);
nor U16130 (N_16130,N_12679,N_13479);
xor U16131 (N_16131,N_15504,N_14559);
or U16132 (N_16132,N_12862,N_12815);
nand U16133 (N_16133,N_14534,N_14166);
and U16134 (N_16134,N_15642,N_12310);
or U16135 (N_16135,N_14850,N_14802);
nand U16136 (N_16136,N_14333,N_15996);
or U16137 (N_16137,N_15553,N_13630);
and U16138 (N_16138,N_13468,N_15741);
nand U16139 (N_16139,N_12709,N_15631);
and U16140 (N_16140,N_12837,N_14563);
and U16141 (N_16141,N_13034,N_15022);
nand U16142 (N_16142,N_14668,N_12151);
and U16143 (N_16143,N_14502,N_15102);
and U16144 (N_16144,N_13166,N_12056);
nor U16145 (N_16145,N_15106,N_15740);
xnor U16146 (N_16146,N_12973,N_12135);
or U16147 (N_16147,N_14901,N_14712);
xnor U16148 (N_16148,N_12463,N_13842);
and U16149 (N_16149,N_12552,N_13949);
nand U16150 (N_16150,N_13633,N_15766);
nand U16151 (N_16151,N_15940,N_14480);
and U16152 (N_16152,N_12036,N_15024);
and U16153 (N_16153,N_13833,N_14625);
nand U16154 (N_16154,N_14186,N_15594);
or U16155 (N_16155,N_14585,N_14354);
and U16156 (N_16156,N_15974,N_15614);
and U16157 (N_16157,N_12443,N_15443);
nor U16158 (N_16158,N_13778,N_12020);
or U16159 (N_16159,N_14089,N_12011);
or U16160 (N_16160,N_13092,N_12941);
nand U16161 (N_16161,N_13297,N_14499);
or U16162 (N_16162,N_14990,N_13997);
nor U16163 (N_16163,N_14022,N_14484);
and U16164 (N_16164,N_13545,N_12067);
nor U16165 (N_16165,N_14218,N_15247);
nor U16166 (N_16166,N_13774,N_13557);
nor U16167 (N_16167,N_15566,N_13313);
xnor U16168 (N_16168,N_13040,N_13807);
nand U16169 (N_16169,N_14291,N_13818);
nand U16170 (N_16170,N_13977,N_14117);
and U16171 (N_16171,N_12693,N_14570);
or U16172 (N_16172,N_12180,N_15925);
and U16173 (N_16173,N_13677,N_13976);
nor U16174 (N_16174,N_12984,N_14895);
xor U16175 (N_16175,N_14538,N_12651);
nor U16176 (N_16176,N_12384,N_14135);
or U16177 (N_16177,N_14234,N_14647);
nor U16178 (N_16178,N_14737,N_14188);
or U16179 (N_16179,N_12142,N_12208);
nand U16180 (N_16180,N_14164,N_14304);
and U16181 (N_16181,N_15692,N_12949);
and U16182 (N_16182,N_15482,N_12790);
nor U16183 (N_16183,N_13223,N_12734);
nand U16184 (N_16184,N_13277,N_13823);
xor U16185 (N_16185,N_12013,N_12787);
xnor U16186 (N_16186,N_14986,N_14242);
nor U16187 (N_16187,N_15872,N_12404);
or U16188 (N_16188,N_13683,N_13427);
or U16189 (N_16189,N_13103,N_14578);
nor U16190 (N_16190,N_14399,N_15429);
or U16191 (N_16191,N_14357,N_14606);
and U16192 (N_16192,N_15340,N_12394);
nand U16193 (N_16193,N_14886,N_15196);
and U16194 (N_16194,N_12585,N_14645);
nor U16195 (N_16195,N_14925,N_15211);
nor U16196 (N_16196,N_13220,N_12538);
nand U16197 (N_16197,N_12773,N_13863);
and U16198 (N_16198,N_13725,N_15761);
nand U16199 (N_16199,N_15574,N_15694);
nand U16200 (N_16200,N_14283,N_15624);
or U16201 (N_16201,N_12943,N_12413);
or U16202 (N_16202,N_13219,N_13125);
and U16203 (N_16203,N_14011,N_14743);
xnor U16204 (N_16204,N_15062,N_12562);
and U16205 (N_16205,N_13728,N_14674);
nor U16206 (N_16206,N_14180,N_15955);
nand U16207 (N_16207,N_13004,N_13504);
or U16208 (N_16208,N_12279,N_15672);
xor U16209 (N_16209,N_13470,N_12451);
nor U16210 (N_16210,N_13987,N_15819);
and U16211 (N_16211,N_15315,N_15650);
xnor U16212 (N_16212,N_13999,N_13866);
nand U16213 (N_16213,N_14879,N_14996);
and U16214 (N_16214,N_15277,N_12681);
and U16215 (N_16215,N_15359,N_14069);
nor U16216 (N_16216,N_12627,N_13503);
and U16217 (N_16217,N_14336,N_13974);
nor U16218 (N_16218,N_13696,N_13081);
nor U16219 (N_16219,N_14653,N_15537);
and U16220 (N_16220,N_14192,N_14193);
or U16221 (N_16221,N_14536,N_14398);
nand U16222 (N_16222,N_13023,N_14579);
or U16223 (N_16223,N_12178,N_15042);
and U16224 (N_16224,N_14774,N_14861);
or U16225 (N_16225,N_15226,N_12418);
or U16226 (N_16226,N_12115,N_14389);
or U16227 (N_16227,N_13925,N_15462);
nand U16228 (N_16228,N_12969,N_15367);
nand U16229 (N_16229,N_12267,N_15478);
or U16230 (N_16230,N_12610,N_13330);
and U16231 (N_16231,N_12905,N_14437);
and U16232 (N_16232,N_14257,N_12556);
nand U16233 (N_16233,N_13604,N_14496);
xnor U16234 (N_16234,N_13798,N_13981);
nand U16235 (N_16235,N_14482,N_13784);
nor U16236 (N_16236,N_15680,N_15835);
or U16237 (N_16237,N_15322,N_12296);
xnor U16238 (N_16238,N_14224,N_14251);
nor U16239 (N_16239,N_14719,N_15050);
nand U16240 (N_16240,N_13106,N_14063);
or U16241 (N_16241,N_14555,N_12085);
xor U16242 (N_16242,N_15671,N_15936);
or U16243 (N_16243,N_13858,N_14786);
nand U16244 (N_16244,N_12993,N_15239);
and U16245 (N_16245,N_13064,N_13593);
or U16246 (N_16246,N_13462,N_15863);
nor U16247 (N_16247,N_12868,N_12123);
and U16248 (N_16248,N_13116,N_13591);
nor U16249 (N_16249,N_12770,N_13229);
nand U16250 (N_16250,N_14639,N_13411);
nor U16251 (N_16251,N_14129,N_12519);
or U16252 (N_16252,N_15139,N_12201);
xor U16253 (N_16253,N_12932,N_15030);
nand U16254 (N_16254,N_14074,N_15779);
or U16255 (N_16255,N_12602,N_14753);
xnor U16256 (N_16256,N_13336,N_12529);
or U16257 (N_16257,N_15341,N_13038);
or U16258 (N_16258,N_14738,N_14628);
nand U16259 (N_16259,N_15829,N_13162);
nor U16260 (N_16260,N_12325,N_12138);
xor U16261 (N_16261,N_13828,N_12924);
nand U16262 (N_16262,N_15091,N_15728);
or U16263 (N_16263,N_15392,N_12909);
and U16264 (N_16264,N_15303,N_12098);
and U16265 (N_16265,N_12769,N_14321);
nand U16266 (N_16266,N_14605,N_12611);
nor U16267 (N_16267,N_13235,N_13300);
nor U16268 (N_16268,N_12458,N_15858);
or U16269 (N_16269,N_15964,N_13400);
nor U16270 (N_16270,N_14580,N_14664);
nor U16271 (N_16271,N_15824,N_14880);
nor U16272 (N_16272,N_15944,N_15745);
or U16273 (N_16273,N_13737,N_12748);
nor U16274 (N_16274,N_14638,N_13595);
or U16275 (N_16275,N_15421,N_15691);
or U16276 (N_16276,N_14268,N_13046);
or U16277 (N_16277,N_15817,N_13027);
nor U16278 (N_16278,N_13837,N_12664);
nor U16279 (N_16279,N_12614,N_12412);
or U16280 (N_16280,N_15904,N_15921);
xor U16281 (N_16281,N_15233,N_14222);
xnor U16282 (N_16282,N_13446,N_13936);
or U16283 (N_16283,N_14495,N_13838);
and U16284 (N_16284,N_14187,N_13009);
and U16285 (N_16285,N_14921,N_12516);
nand U16286 (N_16286,N_14865,N_15929);
or U16287 (N_16287,N_14620,N_14467);
and U16288 (N_16288,N_13801,N_15470);
nor U16289 (N_16289,N_14815,N_15544);
nand U16290 (N_16290,N_13016,N_13035);
or U16291 (N_16291,N_15870,N_15908);
nor U16292 (N_16292,N_13721,N_14953);
or U16293 (N_16293,N_13485,N_15616);
and U16294 (N_16294,N_12351,N_12161);
nor U16295 (N_16295,N_15197,N_15815);
or U16296 (N_16296,N_15901,N_13291);
and U16297 (N_16297,N_12236,N_15877);
xnor U16298 (N_16298,N_15612,N_12820);
or U16299 (N_16299,N_14407,N_14692);
and U16300 (N_16300,N_15147,N_13590);
and U16301 (N_16301,N_15201,N_15770);
and U16302 (N_16302,N_15841,N_13849);
nor U16303 (N_16303,N_15349,N_13024);
and U16304 (N_16304,N_14746,N_12136);
nor U16305 (N_16305,N_15912,N_12999);
nand U16306 (N_16306,N_15049,N_12873);
and U16307 (N_16307,N_12582,N_13180);
and U16308 (N_16308,N_13860,N_14572);
or U16309 (N_16309,N_12335,N_15913);
nand U16310 (N_16310,N_15926,N_14183);
and U16311 (N_16311,N_12324,N_14394);
xnor U16312 (N_16312,N_13391,N_14617);
xor U16313 (N_16313,N_13295,N_15737);
nand U16314 (N_16314,N_12882,N_12465);
nor U16315 (N_16315,N_13740,N_13289);
and U16316 (N_16316,N_13169,N_15419);
nor U16317 (N_16317,N_13568,N_12239);
or U16318 (N_16318,N_14823,N_13979);
nand U16319 (N_16319,N_12205,N_12946);
nor U16320 (N_16320,N_13803,N_14083);
and U16321 (N_16321,N_15618,N_15599);
nor U16322 (N_16322,N_13260,N_15727);
and U16323 (N_16323,N_12896,N_15356);
and U16324 (N_16324,N_13781,N_15095);
nand U16325 (N_16325,N_13543,N_12812);
and U16326 (N_16326,N_15405,N_13674);
or U16327 (N_16327,N_15742,N_14830);
nand U16328 (N_16328,N_13698,N_13745);
or U16329 (N_16329,N_15526,N_14152);
or U16330 (N_16330,N_15444,N_15715);
or U16331 (N_16331,N_13676,N_13533);
nand U16332 (N_16332,N_15654,N_14470);
nor U16333 (N_16333,N_12517,N_13018);
nand U16334 (N_16334,N_13114,N_15307);
or U16335 (N_16335,N_13492,N_15845);
or U16336 (N_16336,N_15804,N_14624);
and U16337 (N_16337,N_15304,N_12217);
nand U16338 (N_16338,N_14217,N_12106);
nor U16339 (N_16339,N_12926,N_15079);
nor U16340 (N_16340,N_13775,N_14386);
or U16341 (N_16341,N_12545,N_12978);
or U16342 (N_16342,N_14667,N_15070);
nor U16343 (N_16343,N_15257,N_12717);
xnor U16344 (N_16344,N_15665,N_12739);
nand U16345 (N_16345,N_12423,N_13567);
and U16346 (N_16346,N_12019,N_12426);
nand U16347 (N_16347,N_13773,N_15129);
or U16348 (N_16348,N_14363,N_15373);
and U16349 (N_16349,N_14825,N_12885);
and U16350 (N_16350,N_14026,N_14887);
or U16351 (N_16351,N_12212,N_14529);
and U16352 (N_16352,N_12714,N_15222);
and U16353 (N_16353,N_14867,N_14813);
and U16354 (N_16354,N_13443,N_13250);
and U16355 (N_16355,N_13717,N_12015);
and U16356 (N_16356,N_12230,N_12219);
or U16357 (N_16357,N_12190,N_13965);
xor U16358 (N_16358,N_15923,N_12775);
nand U16359 (N_16359,N_12245,N_13448);
nand U16360 (N_16360,N_14805,N_15646);
nor U16361 (N_16361,N_15882,N_14781);
nor U16362 (N_16362,N_13201,N_14372);
nand U16363 (N_16363,N_15871,N_14423);
or U16364 (N_16364,N_12796,N_15632);
nor U16365 (N_16365,N_13234,N_13850);
or U16366 (N_16366,N_15426,N_12030);
nand U16367 (N_16367,N_14369,N_12738);
nor U16368 (N_16368,N_12476,N_15418);
xnor U16369 (N_16369,N_15298,N_13157);
nor U16370 (N_16370,N_15903,N_13130);
nor U16371 (N_16371,N_13613,N_13834);
and U16372 (N_16372,N_12540,N_14951);
or U16373 (N_16373,N_14009,N_12009);
or U16374 (N_16374,N_12629,N_14432);
nand U16375 (N_16375,N_15404,N_15021);
and U16376 (N_16376,N_13791,N_12176);
nor U16377 (N_16377,N_15973,N_15583);
xnor U16378 (N_16378,N_15792,N_13374);
and U16379 (N_16379,N_12512,N_14872);
nand U16380 (N_16380,N_15358,N_15957);
or U16381 (N_16381,N_15271,N_15951);
or U16382 (N_16382,N_15494,N_15560);
and U16383 (N_16383,N_12125,N_13598);
or U16384 (N_16384,N_14045,N_12827);
nor U16385 (N_16385,N_12718,N_14505);
nor U16386 (N_16386,N_13200,N_15150);
nor U16387 (N_16387,N_14923,N_12410);
or U16388 (N_16388,N_15155,N_12081);
nand U16389 (N_16389,N_12297,N_12712);
or U16390 (N_16390,N_15688,N_13099);
nor U16391 (N_16391,N_13228,N_13347);
and U16392 (N_16392,N_12348,N_12415);
nor U16393 (N_16393,N_12831,N_13396);
nor U16394 (N_16394,N_15488,N_15347);
or U16395 (N_16395,N_15245,N_14235);
xnor U16396 (N_16396,N_12648,N_15956);
nand U16397 (N_16397,N_14793,N_13878);
and U16398 (N_16398,N_15036,N_12972);
nand U16399 (N_16399,N_12243,N_12071);
or U16400 (N_16400,N_12114,N_15126);
nand U16401 (N_16401,N_12357,N_12273);
nor U16402 (N_16402,N_13455,N_15812);
or U16403 (N_16403,N_14465,N_12522);
xor U16404 (N_16404,N_14163,N_14039);
nor U16405 (N_16405,N_14558,N_15600);
and U16406 (N_16406,N_12526,N_15939);
and U16407 (N_16407,N_12560,N_12803);
nor U16408 (N_16408,N_13910,N_15012);
nand U16409 (N_16409,N_12643,N_12899);
or U16410 (N_16410,N_13857,N_13713);
nand U16411 (N_16411,N_13436,N_15753);
nand U16412 (N_16412,N_15472,N_12988);
nor U16413 (N_16413,N_14684,N_12042);
nand U16414 (N_16414,N_12680,N_12425);
nand U16415 (N_16415,N_12164,N_13565);
and U16416 (N_16416,N_13527,N_15213);
nand U16417 (N_16417,N_14642,N_14450);
or U16418 (N_16418,N_13546,N_15552);
xnor U16419 (N_16419,N_13671,N_14704);
or U16420 (N_16420,N_13108,N_12515);
nand U16421 (N_16421,N_12441,N_12968);
and U16422 (N_16422,N_14528,N_15777);
or U16423 (N_16423,N_14006,N_15256);
and U16424 (N_16424,N_14461,N_15788);
or U16425 (N_16425,N_12473,N_14409);
and U16426 (N_16426,N_13580,N_15515);
or U16427 (N_16427,N_14691,N_15948);
and U16428 (N_16428,N_14412,N_14378);
nand U16429 (N_16429,N_15620,N_14782);
and U16430 (N_16430,N_15011,N_14991);
nor U16431 (N_16431,N_15698,N_12655);
nand U16432 (N_16432,N_13406,N_15640);
nand U16433 (N_16433,N_15941,N_14967);
nand U16434 (N_16434,N_13517,N_14107);
nand U16435 (N_16435,N_15342,N_13579);
and U16436 (N_16436,N_14195,N_14052);
and U16437 (N_16437,N_14085,N_12628);
and U16438 (N_16438,N_12049,N_14189);
nor U16439 (N_16439,N_12086,N_13702);
and U16440 (N_16440,N_13670,N_12343);
or U16441 (N_16441,N_12504,N_13296);
or U16442 (N_16442,N_12755,N_14522);
nor U16443 (N_16443,N_13605,N_15313);
nand U16444 (N_16444,N_15730,N_12752);
and U16445 (N_16445,N_13014,N_15602);
nand U16446 (N_16446,N_12293,N_14114);
or U16447 (N_16447,N_15549,N_14239);
nor U16448 (N_16448,N_12810,N_15289);
or U16449 (N_16449,N_12925,N_14860);
nor U16450 (N_16450,N_13188,N_13309);
xnor U16451 (N_16451,N_12158,N_12501);
or U16452 (N_16452,N_15953,N_13394);
nor U16453 (N_16453,N_12104,N_15986);
nand U16454 (N_16454,N_12005,N_15412);
or U16455 (N_16455,N_12814,N_14891);
nand U16456 (N_16456,N_12215,N_14448);
nand U16457 (N_16457,N_14105,N_15805);
and U16458 (N_16458,N_14290,N_14263);
nand U16459 (N_16459,N_12561,N_13008);
nor U16460 (N_16460,N_14462,N_12888);
or U16461 (N_16461,N_15541,N_14220);
xor U16462 (N_16462,N_12468,N_14788);
or U16463 (N_16463,N_13854,N_13730);
nand U16464 (N_16464,N_14745,N_15834);
or U16465 (N_16465,N_15732,N_15410);
or U16466 (N_16466,N_13464,N_12740);
nand U16467 (N_16467,N_14172,N_13375);
and U16468 (N_16468,N_14862,N_13418);
nand U16469 (N_16469,N_13830,N_14727);
or U16470 (N_16470,N_15591,N_12280);
nand U16471 (N_16471,N_15004,N_15171);
or U16472 (N_16472,N_13520,N_14077);
nor U16473 (N_16473,N_13782,N_15435);
nand U16474 (N_16474,N_13043,N_14596);
xor U16475 (N_16475,N_12350,N_12674);
and U16476 (N_16476,N_14834,N_12301);
or U16477 (N_16477,N_15157,N_12877);
xor U16478 (N_16478,N_13761,N_12626);
nor U16479 (N_16479,N_14751,N_13584);
nor U16480 (N_16480,N_14611,N_13015);
or U16481 (N_16481,N_15508,N_14115);
nor U16482 (N_16482,N_13069,N_14776);
or U16483 (N_16483,N_12154,N_13031);
or U16484 (N_16484,N_15626,N_12040);
and U16485 (N_16485,N_14707,N_14512);
or U16486 (N_16486,N_15408,N_13575);
or U16487 (N_16487,N_14718,N_14371);
and U16488 (N_16488,N_15507,N_15219);
nor U16489 (N_16489,N_13748,N_13746);
and U16490 (N_16490,N_15199,N_14373);
nand U16491 (N_16491,N_15638,N_13658);
nor U16492 (N_16492,N_15275,N_15263);
and U16493 (N_16493,N_13563,N_12874);
and U16494 (N_16494,N_14509,N_13708);
xnor U16495 (N_16495,N_14714,N_12194);
or U16496 (N_16496,N_12435,N_12121);
nand U16497 (N_16497,N_14173,N_14413);
nand U16498 (N_16498,N_13882,N_13777);
nor U16499 (N_16499,N_12923,N_15718);
and U16500 (N_16500,N_12883,N_14593);
nor U16501 (N_16501,N_12240,N_12861);
or U16502 (N_16502,N_14869,N_12469);
and U16503 (N_16503,N_13689,N_15786);
and U16504 (N_16504,N_14178,N_14629);
and U16505 (N_16505,N_15297,N_15176);
nand U16506 (N_16506,N_12128,N_12900);
or U16507 (N_16507,N_15311,N_13012);
or U16508 (N_16508,N_15585,N_13254);
and U16509 (N_16509,N_13891,N_12959);
nor U16510 (N_16510,N_12252,N_15182);
nor U16511 (N_16511,N_13224,N_12044);
or U16512 (N_16512,N_12307,N_15883);
and U16513 (N_16513,N_14138,N_14963);
nor U16514 (N_16514,N_14007,N_14313);
xnor U16515 (N_16515,N_12759,N_12726);
nor U16516 (N_16516,N_15325,N_15430);
nor U16517 (N_16517,N_13824,N_15505);
nand U16518 (N_16518,N_14770,N_13528);
nor U16519 (N_16519,N_12854,N_13919);
nand U16520 (N_16520,N_13926,N_12231);
or U16521 (N_16521,N_12095,N_13970);
nand U16522 (N_16522,N_15007,N_14108);
and U16523 (N_16523,N_15649,N_14610);
nand U16524 (N_16524,N_12365,N_14553);
nand U16525 (N_16525,N_15584,N_12510);
nor U16526 (N_16526,N_12131,N_14562);
and U16527 (N_16527,N_12035,N_13371);
or U16528 (N_16528,N_13867,N_15937);
and U16529 (N_16529,N_15615,N_13549);
and U16530 (N_16530,N_15032,N_14278);
nor U16531 (N_16531,N_13226,N_13975);
nor U16532 (N_16532,N_14672,N_14168);
and U16533 (N_16533,N_12588,N_13495);
and U16534 (N_16534,N_15374,N_15980);
nand U16535 (N_16535,N_13726,N_12054);
or U16536 (N_16536,N_14944,N_12150);
or U16537 (N_16537,N_13639,N_12604);
or U16538 (N_16538,N_15628,N_12671);
nor U16539 (N_16539,N_13570,N_12915);
and U16540 (N_16540,N_13124,N_12401);
and U16541 (N_16541,N_14504,N_13682);
and U16542 (N_16542,N_12043,N_14084);
nand U16543 (N_16543,N_13075,N_13734);
nor U16544 (N_16544,N_15202,N_12590);
or U16545 (N_16545,N_15380,N_14109);
xnor U16546 (N_16546,N_13982,N_15158);
and U16547 (N_16547,N_14660,N_12615);
nand U16548 (N_16548,N_12491,N_12314);
nand U16549 (N_16549,N_15997,N_15945);
nor U16550 (N_16550,N_14530,N_15866);
nor U16551 (N_16551,N_12672,N_13073);
nor U16552 (N_16552,N_15441,N_13877);
xor U16553 (N_16553,N_14004,N_12551);
nor U16554 (N_16554,N_12945,N_14984);
or U16555 (N_16555,N_15604,N_15296);
nand U16556 (N_16556,N_13489,N_13117);
nand U16557 (N_16557,N_14387,N_15034);
nor U16558 (N_16558,N_13532,N_13832);
nand U16559 (N_16559,N_14974,N_12890);
nand U16560 (N_16560,N_14344,N_12898);
and U16561 (N_16561,N_13876,N_15383);
nand U16562 (N_16562,N_15899,N_15907);
or U16563 (N_16563,N_12857,N_14909);
nor U16564 (N_16564,N_12741,N_12508);
nor U16565 (N_16565,N_12448,N_13422);
and U16566 (N_16566,N_14818,N_12341);
or U16567 (N_16567,N_15009,N_12185);
nand U16568 (N_16568,N_12704,N_12794);
or U16569 (N_16569,N_15711,N_13059);
xor U16570 (N_16570,N_13601,N_12699);
nand U16571 (N_16571,N_14125,N_13251);
xnor U16572 (N_16572,N_13353,N_13230);
xnor U16573 (N_16573,N_13263,N_13884);
and U16574 (N_16574,N_14789,N_13026);
nor U16575 (N_16575,N_12395,N_14141);
and U16576 (N_16576,N_15471,N_13240);
nand U16577 (N_16577,N_14174,N_13183);
nand U16578 (N_16578,N_12537,N_14131);
nor U16579 (N_16579,N_12482,N_12112);
and U16580 (N_16580,N_12791,N_14328);
or U16581 (N_16581,N_15606,N_15789);
nor U16582 (N_16582,N_12836,N_13189);
and U16583 (N_16583,N_15832,N_14343);
and U16584 (N_16584,N_15658,N_12918);
nand U16585 (N_16585,N_12713,N_13937);
nor U16586 (N_16586,N_12875,N_12916);
and U16587 (N_16587,N_12484,N_14641);
nor U16588 (N_16588,N_13354,N_12264);
nor U16589 (N_16589,N_12288,N_13452);
nor U16590 (N_16590,N_15363,N_13617);
nand U16591 (N_16591,N_14739,N_13127);
and U16592 (N_16592,N_13271,N_13541);
and U16593 (N_16593,N_15379,N_13988);
nand U16594 (N_16594,N_15878,N_15397);
nand U16595 (N_16595,N_15796,N_12485);
or U16596 (N_16596,N_15163,N_14898);
or U16597 (N_16597,N_13290,N_13624);
nand U16598 (N_16598,N_14408,N_14663);
nor U16599 (N_16599,N_12971,N_14212);
nand U16600 (N_16600,N_14419,N_15860);
or U16601 (N_16601,N_13054,N_14016);
xor U16602 (N_16602,N_13768,N_15439);
or U16603 (N_16603,N_13523,N_15133);
nand U16604 (N_16604,N_14116,N_13608);
nor U16605 (N_16605,N_15733,N_13248);
and U16606 (N_16606,N_15525,N_15249);
and U16607 (N_16607,N_15229,N_14569);
or U16608 (N_16608,N_14184,N_14029);
nand U16609 (N_16609,N_15806,N_13921);
or U16610 (N_16610,N_15667,N_13058);
and U16611 (N_16611,N_12456,N_15780);
nor U16612 (N_16612,N_14282,N_12603);
or U16613 (N_16613,N_13764,N_12257);
nand U16614 (N_16614,N_12302,N_15634);
nor U16615 (N_16615,N_13453,N_12368);
xor U16616 (N_16616,N_14418,N_12823);
nand U16617 (N_16617,N_14907,N_14310);
nand U16618 (N_16618,N_15803,N_15474);
nand U16619 (N_16619,N_15044,N_13221);
nor U16620 (N_16620,N_13151,N_14219);
xnor U16621 (N_16621,N_12886,N_15485);
and U16622 (N_16622,N_14474,N_14079);
nor U16623 (N_16623,N_15331,N_15750);
nand U16624 (N_16624,N_12105,N_13582);
and U16625 (N_16625,N_15040,N_15959);
and U16626 (N_16626,N_14970,N_14431);
nor U16627 (N_16627,N_12763,N_14159);
nand U16628 (N_16628,N_13193,N_13105);
nand U16629 (N_16629,N_12102,N_12129);
and U16630 (N_16630,N_13853,N_15453);
and U16631 (N_16631,N_14521,N_15273);
nand U16632 (N_16632,N_12170,N_14347);
and U16633 (N_16633,N_12229,N_12711);
and U16634 (N_16634,N_13795,N_15895);
or U16635 (N_16635,N_15861,N_12303);
xnor U16636 (N_16636,N_15451,N_13471);
nor U16637 (N_16637,N_13197,N_14197);
and U16638 (N_16638,N_15849,N_14736);
nor U16639 (N_16639,N_15595,N_14403);
or U16640 (N_16640,N_15530,N_12683);
nor U16641 (N_16641,N_14803,N_12571);
nor U16642 (N_16642,N_13028,N_15890);
or U16643 (N_16643,N_13377,N_15712);
and U16644 (N_16644,N_15014,N_13021);
nand U16645 (N_16645,N_12144,N_12625);
nand U16646 (N_16646,N_14767,N_12471);
or U16647 (N_16647,N_14368,N_14937);
or U16648 (N_16648,N_12851,N_12092);
or U16649 (N_16649,N_15954,N_12554);
and U16650 (N_16650,N_15394,N_13177);
nand U16651 (N_16651,N_15846,N_12779);
nor U16652 (N_16652,N_13126,N_14837);
or U16653 (N_16653,N_15920,N_12998);
xor U16654 (N_16654,N_14250,N_13720);
nand U16655 (N_16655,N_14659,N_13886);
or U16656 (N_16656,N_13344,N_14279);
or U16657 (N_16657,N_15240,N_12119);
and U16658 (N_16658,N_12479,N_14678);
nand U16659 (N_16659,N_14238,N_12367);
nor U16660 (N_16660,N_13173,N_12237);
and U16661 (N_16661,N_15839,N_12459);
nor U16662 (N_16662,N_14557,N_12449);
and U16663 (N_16663,N_12431,N_12157);
or U16664 (N_16664,N_13953,N_13205);
or U16665 (N_16665,N_14027,N_15837);
nand U16666 (N_16666,N_14203,N_13331);
or U16667 (N_16667,N_13955,N_14646);
and U16668 (N_16668,N_13316,N_12361);
or U16669 (N_16669,N_15077,N_14201);
or U16670 (N_16670,N_14043,N_13080);
or U16671 (N_16671,N_13252,N_14685);
nor U16672 (N_16672,N_14381,N_15057);
xnor U16673 (N_16673,N_12342,N_14656);
or U16674 (N_16674,N_14098,N_15862);
and U16675 (N_16675,N_13431,N_12970);
nor U16676 (N_16676,N_15230,N_13540);
and U16677 (N_16677,N_12624,N_12710);
nand U16678 (N_16678,N_14270,N_15413);
nor U16679 (N_16679,N_12742,N_15932);
nor U16680 (N_16680,N_13680,N_15563);
and U16681 (N_16681,N_14795,N_13628);
and U16682 (N_16682,N_15719,N_14846);
and U16683 (N_16683,N_14082,N_13065);
nor U16684 (N_16684,N_12091,N_15069);
and U16685 (N_16685,N_14366,N_12446);
nand U16686 (N_16686,N_15529,N_14400);
nand U16687 (N_16687,N_12028,N_15270);
xor U16688 (N_16688,N_12226,N_14227);
nand U16689 (N_16689,N_12023,N_15274);
xor U16690 (N_16690,N_14999,N_13753);
or U16691 (N_16691,N_15651,N_12152);
nor U16692 (N_16692,N_13822,N_12963);
nor U16693 (N_16693,N_15177,N_14648);
xnor U16694 (N_16694,N_12631,N_14878);
nand U16695 (N_16695,N_14936,N_12047);
and U16696 (N_16696,N_15204,N_14005);
nor U16697 (N_16697,N_12399,N_12246);
xor U16698 (N_16698,N_12130,N_12041);
or U16699 (N_16699,N_14417,N_14631);
nand U16700 (N_16700,N_15195,N_13661);
nor U16701 (N_16701,N_13929,N_15116);
nor U16702 (N_16702,N_12606,N_13583);
or U16703 (N_16703,N_12544,N_14729);
or U16704 (N_16704,N_12878,N_13036);
and U16705 (N_16705,N_13738,N_14713);
or U16706 (N_16706,N_14332,N_14881);
nor U16707 (N_16707,N_14314,N_14915);
and U16708 (N_16708,N_12109,N_12444);
or U16709 (N_16709,N_15607,N_13287);
nor U16710 (N_16710,N_15776,N_14273);
xor U16711 (N_16711,N_15723,N_13686);
nor U16712 (N_16712,N_14787,N_14513);
nand U16713 (N_16713,N_13805,N_13141);
or U16714 (N_16714,N_12665,N_12558);
nand U16715 (N_16715,N_12965,N_12908);
or U16716 (N_16716,N_13140,N_15169);
nand U16717 (N_16717,N_12535,N_13766);
nor U16718 (N_16718,N_14154,N_15251);
and U16719 (N_16719,N_14799,N_14700);
nand U16720 (N_16720,N_15016,N_15039);
nor U16721 (N_16721,N_12824,N_15360);
xor U16722 (N_16722,N_15382,N_12427);
nor U16723 (N_16723,N_13282,N_13596);
and U16724 (N_16724,N_13610,N_14603);
nor U16725 (N_16725,N_15952,N_15637);
nor U16726 (N_16726,N_15389,N_12962);
nor U16727 (N_16727,N_12645,N_14933);
or U16728 (N_16728,N_15966,N_13736);
xor U16729 (N_16729,N_12424,N_14240);
or U16730 (N_16730,N_15434,N_12780);
or U16731 (N_16731,N_15596,N_14223);
or U16732 (N_16732,N_13142,N_14140);
or U16733 (N_16733,N_12619,N_12518);
nor U16734 (N_16734,N_14829,N_13351);
and U16735 (N_16735,N_14938,N_14733);
and U16736 (N_16736,N_15339,N_14599);
or U16737 (N_16737,N_12145,N_15317);
or U16738 (N_16738,N_12224,N_13061);
nor U16739 (N_16739,N_14615,N_15143);
nand U16740 (N_16740,N_14272,N_15464);
nor U16741 (N_16741,N_15868,N_15217);
nor U16742 (N_16742,N_14958,N_15610);
nor U16743 (N_16743,N_13994,N_12701);
nor U16744 (N_16744,N_12079,N_12548);
nor U16745 (N_16745,N_15048,N_13278);
nand U16746 (N_16746,N_12733,N_12189);
or U16747 (N_16747,N_12686,N_12646);
xnor U16748 (N_16748,N_15663,N_15205);
or U16749 (N_16749,N_15666,N_14101);
nor U16750 (N_16750,N_15087,N_14401);
nor U16751 (N_16751,N_12724,N_14893);
nor U16752 (N_16752,N_15765,N_12284);
nand U16753 (N_16753,N_14627,N_13547);
nor U16754 (N_16754,N_12578,N_12137);
or U16755 (N_16755,N_14324,N_12193);
or U16756 (N_16756,N_15838,N_15532);
or U16757 (N_16757,N_15122,N_15467);
and U16758 (N_16758,N_14228,N_15055);
nand U16759 (N_16759,N_14705,N_14030);
nor U16760 (N_16760,N_14864,N_12593);
nor U16761 (N_16761,N_12934,N_13892);
nand U16762 (N_16762,N_15971,N_12002);
xor U16763 (N_16763,N_13956,N_15915);
nand U16764 (N_16764,N_15922,N_14438);
and U16765 (N_16765,N_15085,N_14634);
nor U16766 (N_16766,N_13437,N_14650);
nand U16767 (N_16767,N_13681,N_14723);
and U16768 (N_16768,N_12966,N_14785);
or U16769 (N_16769,N_14167,N_12829);
or U16770 (N_16770,N_15958,N_15884);
and U16771 (N_16771,N_15551,N_12880);
or U16772 (N_16772,N_13222,N_13856);
xor U16773 (N_16773,N_14346,N_15627);
or U16774 (N_16774,N_15621,N_14554);
nor U16775 (N_16775,N_12347,N_14068);
nand U16776 (N_16776,N_13249,N_13701);
nor U16777 (N_16777,N_12363,N_15774);
or U16778 (N_16778,N_12388,N_12498);
or U16779 (N_16779,N_14551,N_12326);
nand U16780 (N_16780,N_13447,N_14300);
nand U16781 (N_16781,N_13942,N_13370);
xnor U16782 (N_16782,N_13088,N_15043);
xnor U16783 (N_16783,N_13047,N_13817);
nor U16784 (N_16784,N_12360,N_14930);
and U16785 (N_16785,N_14658,N_15465);
or U16786 (N_16786,N_12055,N_13074);
and U16787 (N_16787,N_14335,N_12272);
or U16788 (N_16788,N_14670,N_13544);
and U16789 (N_16789,N_15301,N_12269);
and U16790 (N_16790,N_13553,N_12802);
nand U16791 (N_16791,N_13358,N_13338);
xnor U16792 (N_16792,N_14067,N_13078);
or U16793 (N_16793,N_13413,N_12223);
nand U16794 (N_16794,N_15608,N_12894);
nand U16795 (N_16795,N_13405,N_15402);
nand U16796 (N_16796,N_13440,N_13855);
nand U16797 (N_16797,N_12196,N_13259);
nand U16798 (N_16798,N_14110,N_15635);
and U16799 (N_16799,N_13368,N_12074);
nand U16800 (N_16800,N_14750,N_14036);
or U16801 (N_16801,N_15244,N_13294);
nor U16802 (N_16802,N_14725,N_13561);
or U16803 (N_16803,N_12525,N_15019);
or U16804 (N_16804,N_13362,N_14613);
or U16805 (N_16805,N_15370,N_12657);
and U16806 (N_16806,N_12202,N_12238);
nor U16807 (N_16807,N_12902,N_15081);
or U16808 (N_16808,N_12383,N_14014);
nand U16809 (N_16809,N_15454,N_13401);
or U16810 (N_16810,N_14076,N_14758);
nor U16811 (N_16811,N_13460,N_13924);
nor U16812 (N_16812,N_12799,N_15440);
nor U16813 (N_16813,N_14385,N_14920);
xor U16814 (N_16814,N_12113,N_15653);
nor U16815 (N_16815,N_15558,N_13484);
nand U16816 (N_16816,N_12440,N_14561);
nand U16817 (N_16817,N_12141,N_14422);
nand U16818 (N_16818,N_15536,N_13962);
and U16819 (N_16819,N_13410,N_13432);
or U16820 (N_16820,N_13957,N_14609);
nand U16821 (N_16821,N_12706,N_13762);
nand U16822 (N_16822,N_13900,N_13231);
nand U16823 (N_16823,N_12566,N_12678);
nor U16824 (N_16824,N_15025,N_12608);
nand U16825 (N_16825,N_13308,N_13048);
nor U16826 (N_16826,N_15198,N_12457);
nor U16827 (N_16827,N_12450,N_14289);
nand U16828 (N_16828,N_13558,N_12495);
nor U16829 (N_16829,N_15499,N_14755);
and U16830 (N_16830,N_15578,N_12420);
nand U16831 (N_16831,N_12957,N_12481);
nor U16832 (N_16832,N_12004,N_15105);
or U16833 (N_16833,N_13888,N_13444);
nor U16834 (N_16834,N_14402,N_15333);
and U16835 (N_16835,N_13373,N_13668);
nand U16836 (N_16836,N_15816,N_13551);
nor U16837 (N_16837,N_15047,N_14340);
nand U16838 (N_16838,N_13699,N_13894);
nor U16839 (N_16839,N_12828,N_15556);
nand U16840 (N_16840,N_14679,N_13952);
and U16841 (N_16841,N_13577,N_13243);
and U16842 (N_16842,N_14929,N_14322);
xnor U16843 (N_16843,N_15232,N_15372);
nand U16844 (N_16844,N_15335,N_14541);
xor U16845 (N_16845,N_12801,N_15989);
or U16846 (N_16846,N_13320,N_14093);
xor U16847 (N_16847,N_13237,N_12550);
and U16848 (N_16848,N_15473,N_14452);
and U16849 (N_16849,N_15265,N_15768);
nor U16850 (N_16850,N_15506,N_12433);
and U16851 (N_16851,N_14583,N_15366);
and U16852 (N_16852,N_14094,N_14157);
nand U16853 (N_16853,N_13171,N_15655);
nor U16854 (N_16854,N_13643,N_15286);
xor U16855 (N_16855,N_15994,N_13100);
nor U16856 (N_16856,N_13213,N_14962);
or U16857 (N_16857,N_14454,N_13182);
nor U16858 (N_16858,N_12345,N_12702);
nor U16859 (N_16859,N_13918,N_14249);
and U16860 (N_16860,N_13324,N_14731);
nand U16861 (N_16861,N_15074,N_15864);
or U16862 (N_16862,N_13743,N_14473);
nand U16863 (N_16863,N_15354,N_12833);
and U16864 (N_16864,N_15486,N_14506);
nor U16865 (N_16865,N_15111,N_15854);
or U16866 (N_16866,N_15378,N_13827);
nand U16867 (N_16867,N_14533,N_14960);
nor U16868 (N_16868,N_14034,N_15278);
nand U16869 (N_16869,N_15652,N_13242);
and U16870 (N_16870,N_15351,N_15764);
or U16871 (N_16871,N_15151,N_13076);
and U16872 (N_16872,N_12800,N_13562);
nor U16873 (N_16873,N_13637,N_12445);
and U16874 (N_16874,N_13767,N_13967);
xor U16875 (N_16875,N_13262,N_13480);
nor U16876 (N_16876,N_14661,N_13463);
nand U16877 (N_16877,N_14426,N_13215);
nand U16878 (N_16878,N_12850,N_14525);
nand U16879 (N_16879,N_15098,N_12181);
nor U16880 (N_16880,N_13102,N_13366);
or U16881 (N_16881,N_12870,N_12089);
or U16882 (N_16882,N_15246,N_13502);
and U16883 (N_16883,N_14306,N_15448);
nand U16884 (N_16884,N_13360,N_15362);
or U16885 (N_16885,N_15721,N_15174);
nor U16886 (N_16886,N_15407,N_12511);
nor U16887 (N_16887,N_12847,N_15970);
nand U16888 (N_16888,N_12454,N_15117);
nor U16889 (N_16889,N_15592,N_15054);
nor U16890 (N_16890,N_13499,N_13174);
nor U16891 (N_16891,N_13616,N_15720);
nor U16892 (N_16892,N_13889,N_15258);
nor U16893 (N_16893,N_15279,N_15947);
xnor U16894 (N_16894,N_12464,N_14698);
nor U16895 (N_16895,N_14015,N_14630);
and U16896 (N_16896,N_12403,N_12398);
nand U16897 (N_16897,N_15534,N_14772);
nor U16898 (N_16898,N_15942,N_13361);
and U16899 (N_16899,N_14345,N_12982);
nor U16900 (N_16900,N_14112,N_14768);
nor U16901 (N_16901,N_12822,N_13403);
and U16902 (N_16902,N_15173,N_13812);
nand U16903 (N_16903,N_13176,N_12442);
or U16904 (N_16904,N_13049,N_13896);
and U16905 (N_16905,N_13983,N_13678);
or U16906 (N_16906,N_13346,N_15066);
nor U16907 (N_16907,N_12872,N_12634);
nor U16908 (N_16908,N_12249,N_13461);
nand U16909 (N_16909,N_15822,N_13032);
nand U16910 (N_16910,N_12955,N_15709);
nor U16911 (N_16911,N_13625,N_13359);
nor U16912 (N_16912,N_15976,N_12466);
nand U16913 (N_16913,N_13425,N_14560);
nand U16914 (N_16914,N_12477,N_15597);
nand U16915 (N_16915,N_15262,N_14155);
or U16916 (N_16916,N_15415,N_14924);
nand U16917 (N_16917,N_14702,N_14831);
nor U16918 (N_16918,N_12613,N_14978);
or U16919 (N_16919,N_13241,N_12084);
or U16920 (N_16920,N_13372,N_15518);
nor U16921 (N_16921,N_15364,N_15140);
nor U16922 (N_16922,N_12177,N_14144);
nor U16923 (N_16923,N_14118,N_13559);
and U16924 (N_16924,N_15194,N_12553);
nor U16925 (N_16925,N_13872,N_15754);
and U16926 (N_16926,N_15752,N_13835);
nand U16927 (N_16927,N_15928,N_13433);
nor U16928 (N_16928,N_13530,N_12555);
nand U16929 (N_16929,N_13672,N_15857);
nand U16930 (N_16930,N_14972,N_13632);
nor U16931 (N_16931,N_13663,N_12981);
xnor U16932 (N_16932,N_13950,N_12271);
nand U16933 (N_16933,N_15847,N_14680);
and U16934 (N_16934,N_15769,N_14293);
nand U16935 (N_16935,N_12953,N_13587);
nand U16936 (N_16936,N_14191,N_12897);
nand U16937 (N_16937,N_15183,N_13573);
or U16938 (N_16938,N_14383,N_13187);
xnor U16939 (N_16939,N_14190,N_15013);
or U16940 (N_16940,N_14932,N_14230);
nand U16941 (N_16941,N_14688,N_14643);
nand U16942 (N_16942,N_15458,N_14842);
nand U16943 (N_16943,N_15830,N_12386);
nor U16944 (N_16944,N_12199,N_14549);
or U16945 (N_16945,N_14367,N_13357);
nand U16946 (N_16946,N_15573,N_12031);
nor U16947 (N_16947,N_13703,N_13931);
or U16948 (N_16948,N_14226,N_15587);
or U16949 (N_16949,N_13206,N_15979);
or U16950 (N_16950,N_14493,N_13497);
or U16951 (N_16951,N_12989,N_12636);
or U16952 (N_16952,N_12090,N_15782);
nand U16953 (N_16953,N_14675,N_14910);
or U16954 (N_16954,N_15759,N_14545);
nand U16955 (N_16955,N_14500,N_14577);
nand U16956 (N_16956,N_12786,N_12018);
or U16957 (N_16957,N_13156,N_15384);
or U16958 (N_16958,N_15679,N_12703);
or U16959 (N_16959,N_14102,N_15420);
and U16960 (N_16960,N_15988,N_15477);
nand U16961 (N_16961,N_12947,N_12422);
or U16962 (N_16962,N_13914,N_12220);
xnor U16963 (N_16963,N_14427,N_12317);
nand U16964 (N_16964,N_15035,N_12600);
or U16965 (N_16965,N_15990,N_15452);
nand U16966 (N_16966,N_14845,N_12134);
nor U16967 (N_16967,N_13194,N_14078);
or U16968 (N_16968,N_12000,N_12830);
nand U16969 (N_16969,N_14205,N_13714);
or U16970 (N_16970,N_12842,N_14012);
or U16971 (N_16971,N_15254,N_15726);
and U16972 (N_16972,N_13508,N_15227);
and U16973 (N_16973,N_15540,N_15668);
nand U16974 (N_16974,N_15755,N_12782);
or U16975 (N_16975,N_14134,N_15268);
or U16976 (N_16976,N_13233,N_13272);
and U16977 (N_16977,N_15216,N_15983);
nand U16978 (N_16978,N_12234,N_13618);
or U16979 (N_16979,N_13211,N_15097);
and U16980 (N_16980,N_13649,N_15215);
nand U16981 (N_16981,N_14149,N_14721);
xor U16982 (N_16982,N_12735,N_12889);
or U16983 (N_16983,N_15425,N_15542);
or U16984 (N_16984,N_13172,N_14356);
nand U16985 (N_16985,N_15909,N_13275);
and U16986 (N_16986,N_13846,N_14436);
and U16987 (N_16987,N_12387,N_12174);
or U16988 (N_16988,N_13192,N_15906);
or U16989 (N_16989,N_15590,N_14103);
or U16990 (N_16990,N_13227,N_14361);
nor U16991 (N_16991,N_15881,N_15411);
nand U16992 (N_16992,N_14295,N_12865);
or U16993 (N_16993,N_14416,N_15501);
or U16994 (N_16994,N_14086,N_12904);
nand U16995 (N_16995,N_13066,N_14797);
or U16996 (N_16996,N_14351,N_14342);
nand U16997 (N_16997,N_15623,N_14247);
and U16998 (N_16998,N_14153,N_15490);
nand U16999 (N_16999,N_13128,N_14632);
xor U17000 (N_17000,N_12370,N_14683);
nor U17001 (N_17001,N_14756,N_15466);
nor U17002 (N_17002,N_14543,N_12140);
nand U17003 (N_17003,N_13381,N_14050);
nand U17004 (N_17004,N_15214,N_14002);
and U17005 (N_17005,N_13474,N_12720);
xor U17006 (N_17006,N_12961,N_12381);
nand U17007 (N_17007,N_13416,N_12784);
and U17008 (N_17008,N_14884,N_14088);
nor U17009 (N_17009,N_14892,N_14734);
xor U17010 (N_17010,N_14137,N_15704);
and U17011 (N_17011,N_13286,N_13387);
or U17012 (N_17012,N_15266,N_13780);
or U17013 (N_17013,N_13627,N_13688);
or U17014 (N_17014,N_13288,N_15059);
and U17015 (N_17015,N_15241,N_12952);
nor U17016 (N_17016,N_13450,N_12110);
and U17017 (N_17017,N_12514,N_15493);
or U17018 (N_17018,N_15189,N_12694);
and U17019 (N_17019,N_13865,N_13239);
nor U17020 (N_17020,N_15018,N_15345);
nor U17021 (N_17021,N_15609,N_13323);
nand U17022 (N_17022,N_12494,N_15814);
or U17023 (N_17023,N_15368,N_14919);
xor U17024 (N_17024,N_14374,N_14676);
and U17025 (N_17025,N_12292,N_12819);
or U17026 (N_17026,N_14132,N_14406);
nor U17027 (N_17027,N_14927,N_14928);
nor U17028 (N_17028,N_15292,N_14148);
xnor U17029 (N_17029,N_14253,N_15369);
nor U17030 (N_17030,N_14586,N_15023);
nand U17031 (N_17031,N_12990,N_14453);
or U17032 (N_17032,N_12620,N_15221);
xor U17033 (N_17033,N_14301,N_12059);
nand U17034 (N_17034,N_14576,N_12439);
or U17035 (N_17035,N_13096,N_15569);
nand U17036 (N_17036,N_14515,N_12316);
nor U17037 (N_17037,N_15589,N_14547);
or U17038 (N_17038,N_14591,N_13101);
nor U17039 (N_17039,N_14215,N_12783);
nor U17040 (N_17040,N_12543,N_14914);
or U17041 (N_17041,N_12058,N_15121);
and U17042 (N_17042,N_15283,N_13383);
nand U17043 (N_17043,N_12736,N_15641);
nand U17044 (N_17044,N_15869,N_12268);
and U17045 (N_17045,N_13915,N_13135);
or U17046 (N_17046,N_13318,N_13640);
nand U17047 (N_17047,N_15503,N_12762);
xnor U17048 (N_17048,N_13788,N_12806);
nand U17049 (N_17049,N_12116,N_13070);
nand U17050 (N_17050,N_15459,N_15399);
nor U17051 (N_17051,N_13666,N_12323);
or U17052 (N_17052,N_14550,N_13885);
or U17053 (N_17053,N_15557,N_14821);
nor U17054 (N_17054,N_14854,N_15784);
and U17055 (N_17055,N_12729,N_15190);
nor U17056 (N_17056,N_13184,N_15701);
or U17057 (N_17057,N_12282,N_15778);
xnor U17058 (N_17058,N_12397,N_15843);
nand U17059 (N_17059,N_14994,N_13244);
and U17060 (N_17060,N_13167,N_15629);
nor U17061 (N_17061,N_13269,N_13526);
or U17062 (N_17062,N_13566,N_14699);
nand U17063 (N_17063,N_14548,N_15450);
nand U17064 (N_17064,N_14451,N_15853);
or U17065 (N_17065,N_12705,N_12907);
xnor U17066 (N_17066,N_13638,N_12751);
nor U17067 (N_17067,N_15479,N_15280);
or U17068 (N_17068,N_14181,N_12195);
nor U17069 (N_17069,N_12183,N_12318);
nand U17070 (N_17070,N_12737,N_13507);
and U17071 (N_17071,N_15992,N_13903);
nand U17072 (N_17072,N_12073,N_12232);
and U17073 (N_17073,N_13810,N_12642);
nor U17074 (N_17074,N_14017,N_15387);
nand U17075 (N_17075,N_15180,N_12320);
or U17076 (N_17076,N_15876,N_13747);
nand U17077 (N_17077,N_12843,N_15125);
nand U17078 (N_17078,N_12339,N_13715);
nor U17079 (N_17079,N_15053,N_13367);
nand U17080 (N_17080,N_13345,N_12568);
and U17081 (N_17081,N_15725,N_13491);
or U17082 (N_17082,N_15005,N_14507);
nor U17083 (N_17083,N_15891,N_13852);
nor U17084 (N_17084,N_13376,N_14151);
and U17085 (N_17085,N_13576,N_15206);
and U17086 (N_17086,N_12840,N_12478);
nor U17087 (N_17087,N_12583,N_15328);
or U17088 (N_17088,N_13398,N_15586);
xor U17089 (N_17089,N_15078,N_12520);
nand U17090 (N_17090,N_14246,N_15000);
nor U17091 (N_17091,N_12744,N_15645);
and U17092 (N_17092,N_15787,N_13945);
and U17093 (N_17093,N_15388,N_13139);
xor U17094 (N_17094,N_14589,N_13136);
or U17095 (N_17095,N_14490,N_13843);
nor U17096 (N_17096,N_14352,N_15337);
or U17097 (N_17097,N_15261,N_14487);
or U17098 (N_17098,N_15702,N_14859);
and U17099 (N_17099,N_14935,N_12596);
and U17100 (N_17100,N_12541,N_15132);
nor U17101 (N_17101,N_14911,N_15825);
nor U17102 (N_17102,N_13989,N_13264);
or U17103 (N_17103,N_14655,N_15661);
and U17104 (N_17104,N_15187,N_13705);
nor U17105 (N_17105,N_12500,N_14415);
and U17106 (N_17106,N_14690,N_12623);
and U17107 (N_17107,N_13572,N_14001);
or U17108 (N_17108,N_12380,N_14165);
nand U17109 (N_17109,N_15826,N_14626);
nand U17110 (N_17110,N_13386,N_15414);
or U17111 (N_17111,N_14280,N_14973);
or U17112 (N_17112,N_13861,N_12879);
or U17113 (N_17113,N_12983,N_12929);
nor U17114 (N_17114,N_14382,N_14031);
nor U17115 (N_17115,N_13208,N_15210);
nor U17116 (N_17116,N_15910,N_15203);
or U17117 (N_17117,N_14457,N_12480);
nor U17118 (N_17118,N_12447,N_13168);
nand U17119 (N_17119,N_13487,N_13694);
nor U17120 (N_17120,N_15927,N_13057);
or U17121 (N_17121,N_12754,N_13449);
and U17122 (N_17122,N_15999,N_15100);
nand U17123 (N_17123,N_15880,N_14244);
nand U17124 (N_17124,N_13041,N_15695);
and U17125 (N_17125,N_13901,N_12745);
nor U17126 (N_17126,N_14716,N_15031);
nand U17127 (N_17127,N_15075,N_14985);
nor U17128 (N_17128,N_12414,N_12032);
nor U17129 (N_17129,N_13506,N_15700);
nor U17130 (N_17130,N_15659,N_12460);
or U17131 (N_17131,N_13928,N_14701);
and U17132 (N_17132,N_13611,N_14003);
nor U17133 (N_17133,N_15527,N_14694);
nand U17134 (N_17134,N_14392,N_13122);
or U17135 (N_17135,N_15156,N_13179);
or U17136 (N_17136,N_15886,N_15568);
and U17137 (N_17137,N_13763,N_14968);
nor U17138 (N_17138,N_13787,N_13232);
and U17139 (N_17139,N_12658,N_13586);
or U17140 (N_17140,N_13390,N_15706);
nor U17141 (N_17141,N_13349,N_15060);
and U17142 (N_17142,N_12187,N_13195);
nand U17143 (N_17143,N_14206,N_14904);
or U17144 (N_17144,N_15456,N_13954);
or U17145 (N_17145,N_14091,N_12669);
or U17146 (N_17146,N_13321,N_13606);
xor U17147 (N_17147,N_13556,N_12346);
and U17148 (N_17148,N_13724,N_13093);
and U17149 (N_17149,N_15089,N_14468);
and U17150 (N_17150,N_14302,N_14520);
nor U17151 (N_17151,N_14844,N_13793);
and U17152 (N_17152,N_14337,N_12490);
and U17153 (N_17153,N_14669,N_12235);
and U17154 (N_17154,N_13644,N_15131);
nand U17155 (N_17155,N_13301,N_12954);
or U17156 (N_17156,N_12980,N_13402);
nand U17157 (N_17157,N_13144,N_12995);
nand U17158 (N_17158,N_14566,N_13332);
or U17159 (N_17159,N_13315,N_12364);
and U17160 (N_17160,N_14633,N_13435);
nor U17161 (N_17161,N_13087,N_15038);
xnor U17162 (N_17162,N_14023,N_14355);
and U17163 (N_17163,N_15138,N_14485);
nand U17164 (N_17164,N_14265,N_14979);
and U17165 (N_17165,N_13684,N_15427);
nand U17166 (N_17166,N_15531,N_14104);
and U17167 (N_17167,N_14564,N_13094);
and U17168 (N_17168,N_15949,N_13339);
nand U17169 (N_17169,N_15168,N_14428);
and U17170 (N_17170,N_15562,N_14133);
nor U17171 (N_17171,N_12372,N_13466);
nor U17172 (N_17172,N_15757,N_14722);
nor U17173 (N_17173,N_12016,N_13958);
and U17174 (N_17174,N_13963,N_14761);
nor U17175 (N_17175,N_12075,N_14565);
nor U17176 (N_17176,N_13948,N_13030);
and U17177 (N_17177,N_12375,N_13690);
and U17178 (N_17178,N_13304,N_14982);
nor U17179 (N_17179,N_15678,N_12083);
nor U17180 (N_17180,N_13467,N_13588);
nand U17181 (N_17181,N_13389,N_15329);
nor U17182 (N_17182,N_12467,N_13478);
and U17183 (N_17183,N_12117,N_13712);
and U17184 (N_17184,N_15346,N_12809);
or U17185 (N_17185,N_14211,N_15020);
nand U17186 (N_17186,N_12241,N_12730);
nor U17187 (N_17187,N_14208,N_14130);
and U17188 (N_17188,N_14592,N_12871);
nor U17189 (N_17189,N_12635,N_13851);
nor U17190 (N_17190,N_12169,N_12684);
nand U17191 (N_17191,N_13274,N_12148);
nand U17192 (N_17192,N_13960,N_12688);
nor U17193 (N_17193,N_12940,N_12175);
or U17194 (N_17194,N_15773,N_12996);
and U17195 (N_17195,N_12563,N_13426);
nand U17196 (N_17196,N_15001,N_13535);
and U17197 (N_17197,N_14338,N_15713);
and U17198 (N_17198,N_14621,N_13175);
xnor U17199 (N_17199,N_13119,N_12753);
xnor U17200 (N_17200,N_13317,N_15083);
nor U17201 (N_17201,N_13341,N_13796);
nor U17202 (N_17202,N_13729,N_12663);
nand U17203 (N_17203,N_14075,N_13916);
nand U17204 (N_17204,N_15188,N_13472);
or U17205 (N_17205,N_13514,N_13247);
or U17206 (N_17206,N_12797,N_13006);
and U17207 (N_17207,N_12793,N_14841);
and U17208 (N_17208,N_15318,N_14980);
or U17209 (N_17209,N_13564,N_15893);
and U17210 (N_17210,N_12777,N_12197);
or U17211 (N_17211,N_12542,N_14594);
and U17212 (N_17212,N_15463,N_15480);
nand U17213 (N_17213,N_13927,N_14233);
nor U17214 (N_17214,N_12419,N_14926);
and U17215 (N_17215,N_15887,N_12254);
nor U17216 (N_17216,N_13123,N_14194);
nor U17217 (N_17217,N_15523,N_15859);
and U17218 (N_17218,N_13864,N_12725);
xor U17219 (N_17219,N_14899,N_15225);
nand U17220 (N_17220,N_14424,N_13365);
and U17221 (N_17221,N_13783,N_12922);
or U17222 (N_17222,N_15554,N_12052);
and U17223 (N_17223,N_13723,N_13521);
nand U17224 (N_17224,N_13922,N_13751);
xnor U17225 (N_17225,N_13133,N_14435);
and U17226 (N_17226,N_14516,N_12228);
nand U17227 (N_17227,N_13631,N_13369);
or U17228 (N_17228,N_14997,N_13311);
nor U17229 (N_17229,N_14478,N_12409);
nor U17230 (N_17230,N_13203,N_13340);
nor U17231 (N_17231,N_13749,N_12133);
or U17232 (N_17232,N_13067,N_13146);
or U17233 (N_17233,N_15738,N_13662);
xor U17234 (N_17234,N_15416,N_15739);
and U17235 (N_17235,N_12242,N_12708);
nor U17236 (N_17236,N_13515,N_15442);
and U17237 (N_17237,N_12103,N_13667);
and U17238 (N_17238,N_14248,N_12225);
nor U17239 (N_17239,N_15821,N_13181);
nor U17240 (N_17240,N_13679,N_14836);
and U17241 (N_17241,N_12691,N_12162);
xor U17242 (N_17242,N_12778,N_14459);
nor U17243 (N_17243,N_13257,N_14213);
or U17244 (N_17244,N_15686,N_13212);
or U17245 (N_17245,N_13414,N_12640);
nor U17246 (N_17246,N_13759,N_14792);
or U17247 (N_17247,N_14475,N_15101);
nand U17248 (N_17248,N_12338,N_12276);
and U17249 (N_17249,N_14730,N_13307);
or U17250 (N_17250,N_12406,N_13752);
nor U17251 (N_17251,N_14276,N_14329);
or U17252 (N_17252,N_14097,N_14696);
and U17253 (N_17253,N_12374,N_12263);
and U17254 (N_17254,N_13821,N_13552);
and U17255 (N_17255,N_14902,N_13056);
nor U17256 (N_17256,N_14057,N_14640);
and U17257 (N_17257,N_13594,N_13819);
and U17258 (N_17258,N_15856,N_13161);
or U17259 (N_17259,N_14939,N_15302);
nand U17260 (N_17260,N_14765,N_15660);
nor U17261 (N_17261,N_12987,N_13039);
and U17262 (N_17262,N_12760,N_14518);
or U17263 (N_17263,N_12920,N_14742);
nand U17264 (N_17264,N_15287,N_15284);
nor U17265 (N_17265,N_12416,N_15191);
xor U17266 (N_17266,N_14956,N_14198);
nor U17267 (N_17267,N_13923,N_15762);
and U17268 (N_17268,N_15468,N_12072);
or U17269 (N_17269,N_13408,N_14317);
nor U17270 (N_17270,N_12088,N_14430);
nor U17271 (N_17271,N_14095,N_12139);
and U17272 (N_17272,N_13966,N_15502);
and U17273 (N_17273,N_13695,N_12956);
and U17274 (N_17274,N_15390,N_14947);
nand U17275 (N_17275,N_12156,N_14777);
or U17276 (N_17276,N_14800,N_13636);
nor U17277 (N_17277,N_14619,N_12436);
nand U17278 (N_17278,N_13303,N_15795);
nor U17279 (N_17279,N_14665,N_15094);
or U17280 (N_17280,N_12256,N_14434);
nor U17281 (N_17281,N_14113,N_13326);
and U17282 (N_17282,N_15968,N_14481);
nand U17283 (N_17283,N_12093,N_13814);
nand U17284 (N_17284,N_12505,N_13306);
and U17285 (N_17285,N_15192,N_15306);
nand U17286 (N_17286,N_12534,N_12064);
nand U17287 (N_17287,N_12294,N_14810);
and U17288 (N_17288,N_12690,N_14913);
or U17289 (N_17289,N_12933,N_14759);
nor U17290 (N_17290,N_14359,N_13844);
and U17291 (N_17291,N_15961,N_12126);
and U17292 (N_17292,N_12666,N_12696);
xor U17293 (N_17293,N_14397,N_15120);
nor U17294 (N_17294,N_14827,N_12697);
xnor U17295 (N_17295,N_13537,N_14757);
or U17296 (N_17296,N_15546,N_15336);
or U17297 (N_17297,N_12182,N_14010);
nand U17298 (N_17298,N_15141,N_15052);
and U17299 (N_17299,N_14771,N_12728);
nand U17300 (N_17300,N_12287,N_13062);
and U17301 (N_17301,N_12094,N_13706);
nor U17302 (N_17302,N_13393,N_13458);
or U17303 (N_17303,N_12429,N_13281);
nand U17304 (N_17304,N_15178,N_12155);
or U17305 (N_17305,N_12483,N_12621);
and U17306 (N_17306,N_12428,N_14773);
and U17307 (N_17307,N_14210,N_15744);
xor U17308 (N_17308,N_12207,N_13019);
xnor U17309 (N_17309,N_15512,N_14271);
or U17310 (N_17310,N_13155,N_15361);
xor U17311 (N_17311,N_14393,N_13415);
xnor U17312 (N_17312,N_15428,N_12661);
and U17313 (N_17313,N_13742,N_13995);
or U17314 (N_17314,N_13808,N_12499);
nor U17315 (N_17315,N_13893,N_15998);
or U17316 (N_17316,N_14824,N_12107);
nor U17317 (N_17317,N_14391,N_13207);
nor U17318 (N_17318,N_13806,N_12532);
or U17319 (N_17319,N_15823,N_14087);
or U17320 (N_17320,N_12291,N_13947);
and U17321 (N_17321,N_14199,N_15731);
nand U17322 (N_17322,N_13459,N_15885);
nand U17323 (N_17323,N_15137,N_15371);
nand U17324 (N_17324,N_15931,N_14983);
nand U17325 (N_17325,N_15598,N_14170);
nand U17326 (N_17326,N_14760,N_14950);
nand U17327 (N_17327,N_14196,N_13279);
nor U17328 (N_17328,N_12682,N_14169);
and U17329 (N_17329,N_13946,N_13707);
nor U17330 (N_17330,N_12192,N_12931);
and U17331 (N_17331,N_12051,N_12976);
nand U17332 (N_17332,N_13111,N_15538);
nand U17333 (N_17333,N_14856,N_12785);
nand U17334 (N_17334,N_14588,N_13589);
nand U17335 (N_17335,N_13574,N_14472);
nor U17336 (N_17336,N_13457,N_12111);
and U17337 (N_17337,N_15705,N_13660);
nand U17338 (N_17338,N_15919,N_12618);
or U17339 (N_17339,N_12289,N_14894);
nor U17340 (N_17340,N_15905,N_15914);
nand U17341 (N_17341,N_12100,N_14081);
nand U17342 (N_17342,N_12673,N_15724);
nand U17343 (N_17343,N_15675,N_13873);
and U17344 (N_17344,N_14214,N_13068);
or U17345 (N_17345,N_13727,N_12392);
or U17346 (N_17346,N_12349,N_12721);
or U17347 (N_17347,N_14889,N_13935);
nand U17348 (N_17348,N_14896,N_12050);
xnor U17349 (N_17349,N_15084,N_14922);
nand U17350 (N_17350,N_12489,N_12698);
and U17351 (N_17351,N_12328,N_15167);
nor U17352 (N_17352,N_15894,N_12974);
nand U17353 (N_17353,N_13825,N_14843);
nand U17354 (N_17354,N_12676,N_12203);
and U17355 (N_17355,N_12146,N_13642);
or U17356 (N_17356,N_15930,N_15875);
or U17357 (N_17357,N_15267,N_12599);
and U17358 (N_17358,N_15555,N_15438);
and U17359 (N_17359,N_15223,N_12408);
nor U17360 (N_17360,N_13319,N_13655);
or U17361 (N_17361,N_12887,N_14852);
nand U17362 (N_17362,N_12186,N_14259);
nor U17363 (N_17363,N_12859,N_14590);
xor U17364 (N_17364,N_12632,N_14308);
nor U17365 (N_17365,N_12337,N_15559);
or U17366 (N_17366,N_15250,N_14790);
or U17367 (N_17367,N_15401,N_12265);
nand U17368 (N_17368,N_12816,N_14597);
or U17369 (N_17369,N_14202,N_12813);
nor U17370 (N_17370,N_13476,N_15088);
nand U17371 (N_17371,N_13800,N_13847);
nor U17372 (N_17372,N_13881,N_14987);
nor U17373 (N_17373,N_15736,N_13266);
nand U17374 (N_17374,N_13137,N_15403);
nand U17375 (N_17375,N_12805,N_15670);
or U17376 (N_17376,N_12977,N_14318);
or U17377 (N_17377,N_13980,N_12825);
or U17378 (N_17378,N_12209,N_12580);
nand U17379 (N_17379,N_14780,N_13534);
and U17380 (N_17380,N_14995,N_12881);
or U17381 (N_17381,N_14049,N_15417);
nand U17382 (N_17382,N_15879,N_13811);
and U17383 (N_17383,N_15299,N_13815);
nor U17384 (N_17384,N_12391,N_14546);
nand U17385 (N_17385,N_13158,N_12846);
nand U17386 (N_17386,N_14458,N_15581);
xnor U17387 (N_17387,N_15514,N_14486);
and U17388 (N_17388,N_12758,N_13011);
xor U17389 (N_17389,N_12617,N_14090);
and U17390 (N_17390,N_12014,N_13904);
xnor U17391 (N_17391,N_15991,N_14380);
nor U17392 (N_17392,N_14122,N_15343);
or U17393 (N_17393,N_12455,N_13869);
nand U17394 (N_17394,N_14981,N_14260);
and U17395 (N_17395,N_12080,N_12938);
and U17396 (N_17396,N_14405,N_14871);
or U17397 (N_17397,N_12792,N_12716);
or U17398 (N_17398,N_14334,N_13756);
nor U17399 (N_17399,N_13060,N_12589);
nand U17400 (N_17400,N_12376,N_12772);
and U17401 (N_17401,N_12507,N_14573);
or U17402 (N_17402,N_15916,N_14523);
or U17403 (N_17403,N_15051,N_13120);
nand U17404 (N_17404,N_12163,N_15685);
nor U17405 (N_17405,N_14816,N_15565);
nor U17406 (N_17406,N_15118,N_12099);
nor U17407 (N_17407,N_15185,N_12487);
nor U17408 (N_17408,N_14449,N_15099);
and U17409 (N_17409,N_13198,N_15689);
and U17410 (N_17410,N_15497,N_13165);
nand U17411 (N_17411,N_14703,N_12354);
nand U17412 (N_17412,N_14791,N_12506);
nor U17413 (N_17413,N_13612,N_12259);
nand U17414 (N_17414,N_13794,N_13789);
nor U17415 (N_17415,N_13645,N_15260);
and U17416 (N_17416,N_15130,N_14584);
or U17417 (N_17417,N_15295,N_14686);
nand U17418 (N_17418,N_14965,N_13809);
and U17419 (N_17419,N_15017,N_12811);
or U17420 (N_17420,N_15561,N_13969);
and U17421 (N_17421,N_15386,N_12218);
xor U17422 (N_17422,N_13692,N_13255);
nand U17423 (N_17423,N_12311,N_12573);
or U17424 (N_17424,N_13902,N_14019);
and U17425 (N_17425,N_14073,N_15687);
nand U17426 (N_17426,N_15798,N_13089);
nor U17427 (N_17427,N_13991,N_13711);
and U17428 (N_17428,N_14255,N_15644);
nand U17429 (N_17429,N_12612,N_14264);
nor U17430 (N_17430,N_13719,N_14917);
nand U17431 (N_17431,N_14779,N_12503);
nand U17432 (N_17432,N_12764,N_14649);
xor U17433 (N_17433,N_15850,N_14764);
nor U17434 (N_17434,N_15833,N_15082);
nand U17435 (N_17435,N_13880,N_14033);
nand U17436 (N_17436,N_14305,N_13829);
nand U17437 (N_17437,N_15135,N_12771);
and U17438 (N_17438,N_12153,N_12914);
nor U17439 (N_17439,N_15037,N_14096);
or U17440 (N_17440,N_13490,N_14677);
nand U17441 (N_17441,N_14526,N_13355);
nor U17442 (N_17442,N_14882,N_12944);
and U17443 (N_17443,N_12863,N_15716);
or U17444 (N_17444,N_14466,N_14028);
or U17445 (N_17445,N_15984,N_14209);
nand U17446 (N_17446,N_14977,N_15520);
nand U17447 (N_17447,N_12939,N_13675);
and U17448 (N_17448,N_13998,N_15237);
nor U17449 (N_17449,N_14544,N_13634);
or U17450 (N_17450,N_13908,N_13002);
or U17451 (N_17451,N_14671,N_13469);
xnor U17452 (N_17452,N_12281,N_12216);
nand U17453 (N_17453,N_14966,N_12147);
xor U17454 (N_17454,N_14769,N_14616);
nand U17455 (N_17455,N_13548,N_13104);
and U17456 (N_17456,N_13084,N_14766);
and U17457 (N_17457,N_13739,N_13430);
or U17458 (N_17458,N_13687,N_15751);
nand U17459 (N_17459,N_15090,N_13005);
xor U17460 (N_17460,N_15208,N_12306);
nand U17461 (N_17461,N_12315,N_15110);
xor U17462 (N_17462,N_14410,N_13599);
and U17463 (N_17463,N_13245,N_12576);
and U17464 (N_17464,N_12461,N_14812);
or U17465 (N_17465,N_15184,N_14540);
and U17466 (N_17466,N_12575,N_14058);
or U17467 (N_17467,N_13968,N_12967);
and U17468 (N_17468,N_13481,N_15186);
nor U17469 (N_17469,N_15181,N_13930);
or U17470 (N_17470,N_12244,N_15735);
and U17471 (N_17471,N_14949,N_14574);
and U17472 (N_17472,N_14539,N_12667);
xor U17473 (N_17473,N_12597,N_13868);
and U17474 (N_17474,N_13578,N_12333);
and U17475 (N_17475,N_12379,N_14162);
and U17476 (N_17476,N_12393,N_13542);
nor U17477 (N_17477,N_12855,N_12536);
or U17478 (N_17478,N_14657,N_14303);
and U17479 (N_17479,N_15029,N_14071);
nor U17480 (N_17480,N_12275,N_13770);
and U17481 (N_17481,N_13984,N_13388);
nand U17482 (N_17482,N_14940,N_14147);
nand U17483 (N_17483,N_12033,N_13943);
or U17484 (N_17484,N_12198,N_15312);
or U17485 (N_17485,N_14142,N_15513);
nand U17486 (N_17486,N_14492,N_15760);
nor U17487 (N_17487,N_12921,N_13118);
and U17488 (N_17488,N_12930,N_14873);
nand U17489 (N_17489,N_14582,N_13697);
and U17490 (N_17490,N_12835,N_12437);
and U17491 (N_17491,N_15033,N_13623);
nand U17492 (N_17492,N_12592,N_12649);
nor U17493 (N_17493,N_14460,N_15152);
or U17494 (N_17494,N_14477,N_14762);
nor U17495 (N_17495,N_15519,N_14552);
nand U17496 (N_17496,N_12757,N_14252);
nand U17497 (N_17497,N_14307,N_13132);
nor U17498 (N_17498,N_15086,N_12407);
nand U17499 (N_17499,N_12411,N_14556);
nor U17500 (N_17500,N_14612,N_14254);
nor U17501 (N_17501,N_14277,N_12332);
and U17502 (N_17502,N_14807,N_12012);
nor U17503 (N_17503,N_13933,N_14682);
nand U17504 (N_17504,N_12660,N_12788);
and U17505 (N_17505,N_14414,N_14689);
nand U17506 (N_17506,N_14853,N_14158);
xor U17507 (N_17507,N_15344,N_15924);
nand U17508 (N_17508,N_13342,N_13109);
nor U17509 (N_17509,N_14711,N_13138);
nor U17510 (N_17510,N_14176,N_12299);
and U17511 (N_17511,N_14360,N_14256);
nand U17512 (N_17512,N_13379,N_12747);
or U17513 (N_17513,N_15243,N_15457);
nand U17514 (N_17514,N_14471,N_15460);
nand U17515 (N_17515,N_14840,N_15064);
nor U17516 (N_17516,N_13268,N_15548);
nand U17517 (N_17517,N_15528,N_12159);
xnor U17518 (N_17518,N_15068,N_13831);
xor U17519 (N_17519,N_13920,N_15282);
and U17520 (N_17520,N_12029,N_13445);
nand U17521 (N_17521,N_12492,N_12656);
and U17522 (N_17522,N_13159,N_13217);
or U17523 (N_17523,N_13293,N_14236);
and U17524 (N_17524,N_15603,N_14441);
nand U17525 (N_17525,N_14445,N_15481);
or U17526 (N_17526,N_12723,N_15673);
nor U17527 (N_17527,N_12685,N_12985);
and U17528 (N_17528,N_14362,N_15865);
and U17529 (N_17529,N_12767,N_14784);
xor U17530 (N_17530,N_12960,N_14231);
and U17531 (N_17531,N_12378,N_15811);
nor U17532 (N_17532,N_15207,N_12390);
or U17533 (N_17533,N_14494,N_14503);
nor U17534 (N_17534,N_15003,N_14905);
nor U17535 (N_17535,N_13152,N_12807);
or U17536 (N_17536,N_15290,N_15797);
nor U17537 (N_17537,N_15818,N_12025);
nand U17538 (N_17538,N_15747,N_13531);
and U17539 (N_17539,N_13284,N_12521);
nand U17540 (N_17540,N_15484,N_14855);
or U17541 (N_17541,N_14952,N_15892);
nand U17542 (N_17542,N_15355,N_15142);
or U17543 (N_17543,N_13270,N_13053);
or U17544 (N_17544,N_13329,N_14080);
or U17545 (N_17545,N_12336,N_13310);
and U17546 (N_17546,N_12034,N_13550);
and U17547 (N_17547,N_15272,N_12421);
nand U17548 (N_17548,N_15492,N_14396);
or U17549 (N_17549,N_12173,N_15431);
nand U17550 (N_17550,N_12048,N_12818);
and U17551 (N_17551,N_14662,N_12472);
or U17552 (N_17552,N_15162,N_12858);
nor U17553 (N_17553,N_13673,N_13285);
nor U17554 (N_17554,N_14433,N_13238);
nand U17555 (N_17555,N_12149,N_12283);
nand U17556 (N_17556,N_12834,N_14600);
nor U17557 (N_17557,N_14128,N_14517);
xnor U17558 (N_17558,N_14358,N_12003);
nand U17559 (N_17559,N_12432,N_12547);
nand U17560 (N_17560,N_14037,N_14425);
nor U17561 (N_17561,N_13218,N_13292);
xor U17562 (N_17562,N_13600,N_13757);
nand U17563 (N_17563,N_12453,N_15808);
xnor U17564 (N_17564,N_12677,N_14267);
nand U17565 (N_17565,N_15575,N_14848);
xnor U17566 (N_17566,N_14989,N_12382);
nand U17567 (N_17567,N_12065,N_15112);
and U17568 (N_17568,N_14993,N_14744);
nor U17569 (N_17569,N_13150,N_14942);
nand U17570 (N_17570,N_14748,N_14866);
nor U17571 (N_17571,N_13072,N_15707);
and U17572 (N_17572,N_14783,N_13704);
or U17573 (N_17573,N_13439,N_15982);
or U17574 (N_17574,N_13407,N_14491);
or U17575 (N_17575,N_15722,N_13498);
or U17576 (N_17576,N_14404,N_15396);
or U17577 (N_17577,N_13973,N_13792);
or U17578 (N_17578,N_12659,N_14601);
and U17579 (N_17579,N_13653,N_12601);
or U17580 (N_17580,N_12662,N_13554);
and U17581 (N_17581,N_13862,N_12937);
or U17582 (N_17582,N_14054,N_12068);
and U17583 (N_17583,N_14945,N_15323);
or U17584 (N_17584,N_13750,N_14035);
or U17585 (N_17585,N_15449,N_13941);
and U17586 (N_17586,N_15179,N_13939);
or U17587 (N_17587,N_14008,N_15398);
and U17588 (N_17588,N_15867,N_15888);
and U17589 (N_17589,N_15436,N_13438);
xor U17590 (N_17590,N_13419,N_15900);
xor U17591 (N_17591,N_15775,N_15161);
nand U17592 (N_17592,N_14693,N_12452);
nand U17593 (N_17593,N_14136,N_15248);
or U17594 (N_17594,N_15228,N_14794);
nor U17595 (N_17595,N_12247,N_12210);
nor U17596 (N_17596,N_13505,N_14654);
nand U17597 (N_17597,N_12832,N_15381);
and U17598 (N_17598,N_15699,N_13305);
nand U17599 (N_17599,N_14587,N_12070);
nand U17600 (N_17600,N_13691,N_13442);
nor U17601 (N_17601,N_15104,N_14868);
nand U17602 (N_17602,N_12260,N_13607);
or U17603 (N_17603,N_13210,N_12727);
or U17604 (N_17604,N_13799,N_12255);
nand U17605 (N_17605,N_15898,N_12120);
xnor U17606 (N_17606,N_15073,N_12331);
xor U17607 (N_17607,N_13836,N_14064);
and U17608 (N_17608,N_15144,N_12638);
nand U17609 (N_17609,N_14429,N_15172);
nor U17610 (N_17610,N_12329,N_14145);
or U17611 (N_17611,N_12523,N_12893);
and U17612 (N_17612,N_15981,N_13536);
nor U17613 (N_17613,N_12700,N_12609);
nand U17614 (N_17614,N_15851,N_14835);
nor U17615 (N_17615,N_14740,N_14379);
nor U17616 (N_17616,N_13500,N_15588);
nand U17617 (N_17617,N_14442,N_12756);
and U17618 (N_17618,N_13003,N_12502);
or U17619 (N_17619,N_13875,N_13934);
xor U17620 (N_17620,N_12639,N_13399);
nor U17621 (N_17621,N_15682,N_13364);
nand U17622 (N_17622,N_13899,N_12046);
and U17623 (N_17623,N_14735,N_15946);
and U17624 (N_17624,N_13334,N_14221);
nand U17625 (N_17625,N_15076,N_15622);
nand U17626 (N_17626,N_15291,N_12901);
nand U17627 (N_17627,N_12261,N_12761);
nand U17628 (N_17628,N_13614,N_13592);
or U17629 (N_17629,N_13148,N_14179);
nor U17630 (N_17630,N_15145,N_12689);
nand U17631 (N_17631,N_14216,N_14602);
nor U17632 (N_17632,N_13424,N_15309);
nand U17633 (N_17633,N_14456,N_13001);
nor U17634 (N_17634,N_15165,N_14819);
nor U17635 (N_17635,N_14728,N_12670);
or U17636 (N_17636,N_12108,N_12958);
or U17637 (N_17637,N_12493,N_14954);
nand U17638 (N_17638,N_13804,N_12849);
or U17639 (N_17639,N_12731,N_13659);
or U17640 (N_17640,N_12574,N_14311);
xor U17641 (N_17641,N_12637,N_15028);
or U17642 (N_17642,N_12616,N_15092);
nand U17643 (N_17643,N_14126,N_14497);
or U17644 (N_17644,N_13760,N_13518);
nand U17645 (N_17645,N_14514,N_15423);
and U17646 (N_17646,N_14681,N_14635);
xnor U17647 (N_17647,N_15093,N_15080);
xnor U17648 (N_17648,N_14048,N_13160);
nor U17649 (N_17649,N_15950,N_15643);
or U17650 (N_17650,N_14508,N_14822);
and U17651 (N_17651,N_12715,N_15703);
or U17652 (N_17652,N_14204,N_13848);
and U17653 (N_17653,N_14839,N_13441);
nor U17654 (N_17654,N_12188,N_12057);
nor U17655 (N_17655,N_14511,N_15134);
or U17656 (N_17656,N_13236,N_14903);
nor U17657 (N_17657,N_15756,N_14666);
nor U17658 (N_17658,N_13153,N_14975);
nand U17659 (N_17659,N_15108,N_14575);
and U17660 (N_17660,N_14245,N_14524);
and U17661 (N_17661,N_14123,N_15567);
nor U17662 (N_17662,N_12838,N_15758);
nor U17663 (N_17663,N_12528,N_13917);
and U17664 (N_17664,N_13352,N_13052);
xnor U17665 (N_17665,N_12290,N_13519);
nor U17666 (N_17666,N_13343,N_14798);
or U17667 (N_17667,N_12184,N_12509);
nand U17668 (N_17668,N_15619,N_15376);
xnor U17669 (N_17669,N_15446,N_12286);
or U17670 (N_17670,N_12817,N_12362);
xnor U17671 (N_17671,N_14857,N_14608);
and U17672 (N_17672,N_14161,N_12438);
and U17673 (N_17673,N_13429,N_15269);
and U17674 (N_17674,N_12749,N_12062);
nor U17675 (N_17675,N_13090,N_15276);
nor U17676 (N_17676,N_15063,N_12001);
or U17677 (N_17677,N_15852,N_14828);
or U17678 (N_17678,N_15170,N_15288);
nor U17679 (N_17679,N_13621,N_13509);
or U17680 (N_17680,N_14607,N_14858);
or U17681 (N_17681,N_15393,N_13870);
nand U17682 (N_17682,N_13907,N_12305);
xnor U17683 (N_17683,N_13143,N_15577);
and U17684 (N_17684,N_12586,N_13771);
nand U17685 (N_17685,N_13615,N_12768);
xnor U17686 (N_17686,N_15985,N_12906);
nor U17687 (N_17687,N_12319,N_15046);
nand U17688 (N_17688,N_15960,N_13434);
or U17689 (N_17689,N_14339,N_12488);
nand U17690 (N_17690,N_14262,N_13412);
nor U17691 (N_17691,N_12124,N_12204);
and U17692 (N_17692,N_12572,N_13718);
nor U17693 (N_17693,N_12010,N_14697);
or U17694 (N_17694,N_12251,N_14323);
and U17695 (N_17695,N_13990,N_12082);
nor U17696 (N_17696,N_15639,N_13178);
or U17697 (N_17697,N_13511,N_12266);
or U17698 (N_17698,N_15820,N_12598);
xor U17699 (N_17699,N_13428,N_12304);
nor U17700 (N_17700,N_15972,N_13191);
or U17701 (N_17701,N_14943,N_12911);
and U17702 (N_17702,N_12496,N_15332);
nand U17703 (N_17703,N_15933,N_15807);
nand U17704 (N_17704,N_15570,N_15424);
nor U17705 (N_17705,N_15136,N_14636);
or U17706 (N_17706,N_15934,N_15783);
xnor U17707 (N_17707,N_14838,N_13813);
xor U17708 (N_17708,N_15969,N_12912);
or U17709 (N_17709,N_13620,N_14948);
or U17710 (N_17710,N_13513,N_12172);
nor U17711 (N_17711,N_14532,N_13897);
nor U17712 (N_17712,N_14119,N_15491);
or U17713 (N_17713,N_13196,N_12895);
and U17714 (N_17714,N_15710,N_14146);
nand U17715 (N_17715,N_14623,N_13665);
nand U17716 (N_17716,N_13648,N_12577);
nor U17717 (N_17717,N_14013,N_15461);
nand U17718 (N_17718,N_12248,N_14885);
and U17719 (N_17719,N_14747,N_15963);
or U17720 (N_17720,N_14870,N_14124);
and U17721 (N_17721,N_12024,N_15831);
and U17722 (N_17722,N_13735,N_13841);
nand U17723 (N_17723,N_13482,N_14376);
and U17724 (N_17724,N_13496,N_12668);
nand U17725 (N_17725,N_13085,N_14567);
nand U17726 (N_17726,N_15377,N_13149);
nand U17727 (N_17727,N_14375,N_13826);
or U17728 (N_17728,N_14673,N_12910);
and U17729 (N_17729,N_12221,N_15072);
nand U17730 (N_17730,N_15571,N_15873);
and U17731 (N_17731,N_15917,N_15350);
nand U17732 (N_17732,N_13722,N_13246);
or U17733 (N_17733,N_15281,N_15801);
or U17734 (N_17734,N_12309,N_13529);
nor U17735 (N_17735,N_12581,N_12867);
and U17736 (N_17736,N_14637,N_14463);
nand U17737 (N_17737,N_12579,N_14320);
or U17738 (N_17738,N_14294,N_15433);
and U17739 (N_17739,N_15576,N_14501);
nand U17740 (N_17740,N_15676,N_14832);
and U17741 (N_17741,N_13785,N_12353);
nor U17742 (N_17742,N_12206,N_12285);
or U17743 (N_17743,N_15889,N_12570);
or U17744 (N_17744,N_15259,N_12038);
and U17745 (N_17745,N_13395,N_12848);
or U17746 (N_17746,N_15746,N_12591);
nor U17747 (N_17747,N_12017,N_12687);
or U17748 (N_17748,N_12653,N_15400);
nand U17749 (N_17749,N_15008,N_13091);
nor U17750 (N_17750,N_15827,N_15128);
nand U17751 (N_17751,N_12359,N_12417);
nand U17752 (N_17752,N_15235,N_13710);
or U17753 (N_17753,N_15967,N_15327);
or U17754 (N_17754,N_12948,N_12061);
and U17755 (N_17755,N_15896,N_12270);
and U17756 (N_17756,N_14464,N_13603);
and U17757 (N_17757,N_14900,N_12524);
nor U17758 (N_17758,N_15664,N_15242);
nand U17759 (N_17759,N_12527,N_14808);
or U17760 (N_17760,N_14182,N_15149);
nand U17761 (N_17761,N_12076,N_15771);
xor U17762 (N_17762,N_14469,N_13214);
nand U17763 (N_17763,N_13267,N_12327);
and U17764 (N_17764,N_15844,N_14062);
nand U17765 (N_17765,N_15326,N_14316);
or U17766 (N_17766,N_13261,N_15975);
or U17767 (N_17767,N_12200,N_12405);
xor U17768 (N_17768,N_12078,N_14804);
nand U17769 (N_17769,N_13486,N_13050);
xnor U17770 (N_17770,N_15683,N_14258);
or U17771 (N_17771,N_13475,N_14143);
nor U17772 (N_17772,N_14811,N_15935);
nand U17773 (N_17773,N_13186,N_15061);
nor U17774 (N_17774,N_12233,N_14121);
or U17775 (N_17775,N_15717,N_13314);
and U17776 (N_17776,N_13964,N_13911);
or U17777 (N_17777,N_13560,N_15593);
and U17778 (N_17778,N_15160,N_13581);
or U17779 (N_17779,N_14341,N_13602);
nor U17780 (N_17780,N_12022,N_14177);
and U17781 (N_17781,N_14040,N_12531);
nand U17782 (N_17782,N_13741,N_14604);
nand U17783 (N_17783,N_13147,N_12869);
nand U17784 (N_17784,N_12278,N_14298);
nor U17785 (N_17785,N_12549,N_15799);
and U17786 (N_17786,N_14890,N_15522);
nor U17787 (N_17787,N_12096,N_15127);
nand U17788 (N_17788,N_14809,N_12605);
or U17789 (N_17789,N_14309,N_14527);
nand U17790 (N_17790,N_13020,N_13758);
and U17791 (N_17791,N_15096,N_15978);
or U17792 (N_17792,N_14897,N_14440);
xor U17793 (N_17793,N_13845,N_13253);
nor U17794 (N_17794,N_13938,N_12722);
nor U17795 (N_17795,N_15164,N_14998);
nor U17796 (N_17796,N_13732,N_13647);
nand U17797 (N_17797,N_13209,N_13932);
nor U17798 (N_17798,N_15897,N_15316);
or U17799 (N_17799,N_14171,N_15617);
nor U17800 (N_17800,N_14476,N_14053);
nor U17801 (N_17801,N_12607,N_14732);
nor U17802 (N_17802,N_12355,N_12533);
nor U17803 (N_17803,N_14488,N_15234);
nor U17804 (N_17804,N_12118,N_13335);
or U17805 (N_17805,N_12732,N_12160);
or U17806 (N_17806,N_14319,N_14111);
nor U17807 (N_17807,N_12928,N_12530);
or U17808 (N_17808,N_13204,N_15006);
and U17809 (N_17809,N_15321,N_15677);
and U17810 (N_17810,N_15432,N_15495);
nand U17811 (N_17811,N_15840,N_14061);
or U17812 (N_17812,N_15681,N_13350);
xnor U17813 (N_17813,N_12313,N_14072);
nand U17814 (N_17814,N_12584,N_15743);
or U17815 (N_17815,N_13874,N_14752);
nand U17816 (N_17816,N_12430,N_13656);
and U17817 (N_17817,N_15365,N_12546);
or U17818 (N_17818,N_12695,N_13619);
and U17819 (N_17819,N_13733,N_12122);
or U17820 (N_17820,N_15539,N_14446);
and U17821 (N_17821,N_13384,N_14537);
and U17822 (N_17822,N_14888,N_12707);
nor U17823 (N_17823,N_12795,N_14200);
nand U17824 (N_17824,N_12856,N_12371);
or U17825 (N_17825,N_12935,N_14874);
and U17826 (N_17826,N_13769,N_14568);
or U17827 (N_17827,N_14964,N_13276);
and U17828 (N_17828,N_14325,N_14353);
or U17829 (N_17829,N_12165,N_15836);
xnor U17830 (N_17830,N_15231,N_12633);
or U17831 (N_17831,N_12844,N_14687);
and U17832 (N_17832,N_14941,N_13079);
nor U17833 (N_17833,N_14315,N_13840);
and U17834 (N_17834,N_12951,N_13996);
and U17835 (N_17835,N_12340,N_15918);
xnor U17836 (N_17836,N_13754,N_12650);
or U17837 (N_17837,N_15308,N_15785);
and U17838 (N_17838,N_15209,N_13302);
or U17839 (N_17839,N_15395,N_13283);
or U17840 (N_17840,N_14185,N_15790);
or U17841 (N_17841,N_14535,N_15647);
or U17842 (N_17842,N_13790,N_15564);
nand U17843 (N_17843,N_13512,N_12312);
and U17844 (N_17844,N_14056,N_12513);
or U17845 (N_17845,N_13322,N_15314);
nor U17846 (N_17846,N_15391,N_13909);
or U17847 (N_17847,N_14877,N_13971);
or U17848 (N_17848,N_15324,N_13086);
and U17849 (N_17849,N_14287,N_14207);
nor U17850 (N_17850,N_12434,N_12222);
nor U17851 (N_17851,N_13063,N_13483);
nor U17852 (N_17852,N_15305,N_12630);
xnor U17853 (N_17853,N_13333,N_13883);
nor U17854 (N_17854,N_15483,N_13312);
nand U17855 (N_17855,N_12936,N_13013);
and U17856 (N_17856,N_14912,N_14531);
nand U17857 (N_17857,N_14261,N_13539);
or U17858 (N_17858,N_13417,N_15995);
nor U17859 (N_17859,N_13473,N_15656);
nor U17860 (N_17860,N_14021,N_12821);
and U17861 (N_17861,N_12308,N_14644);
xnor U17862 (N_17862,N_13113,N_13944);
and U17863 (N_17863,N_14038,N_15200);
xor U17864 (N_17864,N_14971,N_13664);
or U17865 (N_17865,N_13378,N_13042);
or U17866 (N_17866,N_12776,N_13709);
and U17867 (N_17867,N_14695,N_14754);
nor U17868 (N_17868,N_12852,N_14988);
or U17869 (N_17869,N_13555,N_13421);
nand U17870 (N_17870,N_15550,N_14395);
xor U17871 (N_17871,N_15058,N_15469);
nand U17872 (N_17872,N_14044,N_13802);
nor U17873 (N_17873,N_15547,N_13797);
nand U17874 (N_17874,N_15114,N_12475);
nand U17875 (N_17875,N_13905,N_15330);
and U17876 (N_17876,N_15579,N_12213);
or U17877 (N_17877,N_15148,N_14992);
xor U17878 (N_17878,N_14847,N_14047);
and U17879 (N_17879,N_14796,N_13280);
nand U17880 (N_17880,N_13538,N_14709);
or U17881 (N_17881,N_15065,N_12330);
xor U17882 (N_17882,N_15119,N_12997);
xnor U17883 (N_17883,N_12026,N_15146);
nand U17884 (N_17884,N_14961,N_14288);
nor U17885 (N_17885,N_14622,N_15943);
nor U17886 (N_17886,N_15103,N_14384);
or U17887 (N_17887,N_12258,N_13097);
or U17888 (N_17888,N_15516,N_12654);
nand U17889 (N_17889,N_13044,N_15977);
nor U17890 (N_17890,N_15911,N_13465);
or U17891 (N_17891,N_12622,N_14479);
nor U17892 (N_17892,N_12087,N_15855);
or U17893 (N_17893,N_12356,N_13510);
and U17894 (N_17894,N_14286,N_13913);
xnor U17895 (N_17895,N_13755,N_12917);
or U17896 (N_17896,N_12919,N_15613);
or U17897 (N_17897,N_12876,N_14931);
xor U17898 (N_17898,N_13985,N_15793);
or U17899 (N_17899,N_15636,N_13879);
nor U17900 (N_17900,N_15517,N_14420);
nand U17901 (N_17901,N_12765,N_13622);
and U17902 (N_17902,N_13959,N_15693);
nand U17903 (N_17903,N_12927,N_15113);
nand U17904 (N_17904,N_13107,N_13083);
or U17905 (N_17905,N_12474,N_12781);
nand U17906 (N_17906,N_15375,N_12277);
nor U17907 (N_17907,N_15993,N_14331);
nor U17908 (N_17908,N_13385,N_14715);
nor U17909 (N_17909,N_13327,N_15437);
nand U17910 (N_17910,N_12007,N_14598);
and U17911 (N_17911,N_14348,N_15026);
and U17912 (N_17912,N_14483,N_13525);
and U17913 (N_17913,N_12377,N_12298);
or U17914 (N_17914,N_13037,N_15938);
nor U17915 (N_17915,N_12358,N_13887);
nand U17916 (N_17916,N_12369,N_13154);
nor U17917 (N_17917,N_13045,N_13972);
nand U17918 (N_17918,N_14312,N_12097);
xor U17919 (N_17919,N_12366,N_13022);
or U17920 (N_17920,N_14876,N_15285);
and U17921 (N_17921,N_14041,N_13299);
xnor U17922 (N_17922,N_12994,N_13071);
nor U17923 (N_17923,N_13609,N_14350);
nand U17924 (N_17924,N_12789,N_13716);
or U17925 (N_17925,N_12400,N_14390);
nand U17926 (N_17926,N_14296,N_15690);
and U17927 (N_17927,N_13951,N_13940);
xor U17928 (N_17928,N_12039,N_15015);
nand U17929 (N_17929,N_13131,N_15293);
xnor U17930 (N_17930,N_14918,N_13121);
nor U17931 (N_17931,N_15489,N_14411);
or U17932 (N_17932,N_14269,N_13025);
or U17933 (N_17933,N_12644,N_12214);
or U17934 (N_17934,N_13164,N_13423);
and U17935 (N_17935,N_12641,N_14284);
or U17936 (N_17936,N_14120,N_14364);
nand U17937 (N_17937,N_15842,N_12587);
or U17938 (N_17938,N_14059,N_15056);
xnor U17939 (N_17939,N_15357,N_15253);
or U17940 (N_17940,N_12227,N_15045);
nor U17941 (N_17941,N_13033,N_15475);
xnor U17942 (N_17942,N_13325,N_12373);
nand U17943 (N_17943,N_15657,N_13895);
nor U17944 (N_17944,N_15535,N_13082);
nand U17945 (N_17945,N_15697,N_14032);
and U17946 (N_17946,N_15510,N_12470);
or U17947 (N_17947,N_15772,N_12564);
xnor U17948 (N_17948,N_12746,N_15902);
nand U17949 (N_17949,N_15987,N_13225);
or U17950 (N_17950,N_12595,N_15962);
nand U17951 (N_17951,N_14275,N_12804);
and U17952 (N_17952,N_15300,N_14099);
nor U17953 (N_17953,N_13635,N_12950);
and U17954 (N_17954,N_14285,N_13055);
xnor U17955 (N_17955,N_14778,N_13129);
or U17956 (N_17956,N_12892,N_15543);
nand U17957 (N_17957,N_15319,N_14349);
and U17958 (N_17958,N_12021,N_15524);
nor U17959 (N_17959,N_12992,N_12274);
nand U17960 (N_17960,N_12719,N_15696);
nor U17961 (N_17961,N_13298,N_14969);
nand U17962 (N_17962,N_13890,N_12774);
nand U17963 (N_17963,N_15729,N_14241);
nand U17964 (N_17964,N_15582,N_15669);
xnor U17965 (N_17965,N_12300,N_13871);
and U17966 (N_17966,N_12942,N_15027);
and U17967 (N_17967,N_15154,N_15175);
or U17968 (N_17968,N_12539,N_12396);
nand U17969 (N_17969,N_15159,N_13199);
nor U17970 (N_17970,N_14092,N_14498);
or U17971 (N_17971,N_12913,N_15409);
and U17972 (N_17972,N_15809,N_12557);
nor U17973 (N_17973,N_13456,N_14020);
nor U17974 (N_17974,N_13382,N_15763);
nor U17975 (N_17975,N_12262,N_15674);
or U17976 (N_17976,N_12864,N_12322);
and U17977 (N_17977,N_13501,N_15320);
nor U17978 (N_17978,N_15002,N_14741);
nor U17979 (N_17979,N_12692,N_14519);
and U17980 (N_17980,N_14055,N_15385);
or U17981 (N_17981,N_15153,N_13112);
and U17982 (N_17982,N_13363,N_14139);
nor U17983 (N_17983,N_13202,N_14571);
xnor U17984 (N_17984,N_13646,N_14708);
nand U17985 (N_17985,N_12063,N_13859);
or U17986 (N_17986,N_15848,N_14652);
or U17987 (N_17987,N_14724,N_15828);
nand U17988 (N_17988,N_12866,N_15445);
nand U17989 (N_17989,N_15802,N_15748);
nand U17990 (N_17990,N_12903,N_12066);
and U17991 (N_17991,N_12053,N_14447);
or U17992 (N_17992,N_13356,N_15115);
nor U17993 (N_17993,N_13494,N_13816);
nand U17994 (N_17994,N_13978,N_12594);
nand U17995 (N_17995,N_14127,N_14266);
nand U17996 (N_17996,N_12826,N_15123);
nand U17997 (N_17997,N_13397,N_15521);
and U17998 (N_17998,N_12979,N_12037);
nand U17999 (N_17999,N_13000,N_12132);
nand U18000 (N_18000,N_15669,N_14877);
and U18001 (N_18001,N_12559,N_13265);
and U18002 (N_18002,N_15401,N_13440);
or U18003 (N_18003,N_12185,N_12926);
or U18004 (N_18004,N_15126,N_15954);
or U18005 (N_18005,N_14762,N_13489);
or U18006 (N_18006,N_13955,N_15360);
or U18007 (N_18007,N_15525,N_14309);
nor U18008 (N_18008,N_13258,N_13160);
and U18009 (N_18009,N_13560,N_12524);
nor U18010 (N_18010,N_15815,N_15808);
and U18011 (N_18011,N_12632,N_13360);
nand U18012 (N_18012,N_12340,N_12258);
and U18013 (N_18013,N_13072,N_14610);
nand U18014 (N_18014,N_12960,N_15906);
nand U18015 (N_18015,N_14930,N_15938);
nor U18016 (N_18016,N_15730,N_12382);
nand U18017 (N_18017,N_15545,N_12596);
and U18018 (N_18018,N_14321,N_15932);
nor U18019 (N_18019,N_12891,N_12465);
or U18020 (N_18020,N_13286,N_12025);
nand U18021 (N_18021,N_12971,N_15855);
and U18022 (N_18022,N_14456,N_15537);
nand U18023 (N_18023,N_15747,N_13798);
and U18024 (N_18024,N_12031,N_15886);
and U18025 (N_18025,N_14612,N_12618);
nor U18026 (N_18026,N_12612,N_14252);
nor U18027 (N_18027,N_15071,N_12685);
or U18028 (N_18028,N_12736,N_12408);
xor U18029 (N_18029,N_12430,N_15946);
or U18030 (N_18030,N_15871,N_15308);
nor U18031 (N_18031,N_13035,N_15568);
nor U18032 (N_18032,N_15523,N_12950);
nor U18033 (N_18033,N_15039,N_14571);
nor U18034 (N_18034,N_15772,N_14610);
xor U18035 (N_18035,N_13160,N_15719);
nor U18036 (N_18036,N_13499,N_15591);
nand U18037 (N_18037,N_12930,N_12629);
nor U18038 (N_18038,N_14524,N_15260);
xnor U18039 (N_18039,N_12253,N_12046);
and U18040 (N_18040,N_15408,N_12589);
nor U18041 (N_18041,N_12298,N_12055);
nand U18042 (N_18042,N_14068,N_15813);
nor U18043 (N_18043,N_12306,N_15239);
and U18044 (N_18044,N_15493,N_12844);
or U18045 (N_18045,N_15251,N_15609);
or U18046 (N_18046,N_13976,N_14139);
nand U18047 (N_18047,N_13323,N_12682);
or U18048 (N_18048,N_12645,N_15064);
xnor U18049 (N_18049,N_12601,N_12207);
nor U18050 (N_18050,N_13153,N_14022);
nand U18051 (N_18051,N_14607,N_12328);
or U18052 (N_18052,N_13840,N_13971);
or U18053 (N_18053,N_12063,N_12773);
nor U18054 (N_18054,N_13779,N_15232);
and U18055 (N_18055,N_13789,N_12888);
nand U18056 (N_18056,N_12434,N_12462);
nand U18057 (N_18057,N_14842,N_13483);
or U18058 (N_18058,N_14281,N_14568);
and U18059 (N_18059,N_13966,N_12074);
and U18060 (N_18060,N_13775,N_12665);
or U18061 (N_18061,N_12313,N_14388);
nor U18062 (N_18062,N_14985,N_14144);
nor U18063 (N_18063,N_12342,N_13759);
and U18064 (N_18064,N_14332,N_12567);
or U18065 (N_18065,N_13956,N_13545);
or U18066 (N_18066,N_13838,N_15601);
or U18067 (N_18067,N_14920,N_15109);
nor U18068 (N_18068,N_14589,N_14545);
xor U18069 (N_18069,N_14908,N_15050);
nor U18070 (N_18070,N_13467,N_14492);
and U18071 (N_18071,N_15852,N_13180);
xnor U18072 (N_18072,N_15590,N_14954);
or U18073 (N_18073,N_15649,N_14587);
and U18074 (N_18074,N_12470,N_14363);
and U18075 (N_18075,N_15316,N_15368);
nand U18076 (N_18076,N_12924,N_13049);
nand U18077 (N_18077,N_13846,N_14519);
nor U18078 (N_18078,N_15595,N_15440);
nand U18079 (N_18079,N_13474,N_14713);
nor U18080 (N_18080,N_12359,N_14002);
and U18081 (N_18081,N_13253,N_12263);
nor U18082 (N_18082,N_14245,N_14603);
xnor U18083 (N_18083,N_12733,N_15134);
nor U18084 (N_18084,N_15602,N_15017);
nor U18085 (N_18085,N_12690,N_13091);
or U18086 (N_18086,N_12201,N_13671);
and U18087 (N_18087,N_15087,N_14049);
or U18088 (N_18088,N_13134,N_12183);
and U18089 (N_18089,N_15147,N_12555);
or U18090 (N_18090,N_13045,N_14746);
nor U18091 (N_18091,N_12404,N_13199);
nand U18092 (N_18092,N_13602,N_13727);
nand U18093 (N_18093,N_13040,N_14526);
or U18094 (N_18094,N_14824,N_14648);
nand U18095 (N_18095,N_12628,N_12471);
xor U18096 (N_18096,N_12161,N_14052);
nor U18097 (N_18097,N_13260,N_12455);
nand U18098 (N_18098,N_12086,N_12699);
nand U18099 (N_18099,N_12808,N_13086);
or U18100 (N_18100,N_14847,N_12620);
and U18101 (N_18101,N_14505,N_12717);
nor U18102 (N_18102,N_14362,N_15366);
nor U18103 (N_18103,N_12210,N_13959);
and U18104 (N_18104,N_15766,N_12487);
or U18105 (N_18105,N_14654,N_15209);
and U18106 (N_18106,N_15519,N_13454);
or U18107 (N_18107,N_15443,N_12926);
nor U18108 (N_18108,N_15111,N_13553);
or U18109 (N_18109,N_14902,N_13023);
or U18110 (N_18110,N_12342,N_15808);
and U18111 (N_18111,N_15366,N_15990);
or U18112 (N_18112,N_12921,N_12382);
or U18113 (N_18113,N_14481,N_15348);
or U18114 (N_18114,N_14083,N_12552);
nor U18115 (N_18115,N_14987,N_13957);
nand U18116 (N_18116,N_14098,N_14859);
nor U18117 (N_18117,N_13621,N_15370);
nand U18118 (N_18118,N_14526,N_12788);
or U18119 (N_18119,N_12089,N_12759);
nor U18120 (N_18120,N_15334,N_14601);
nor U18121 (N_18121,N_12985,N_14342);
nand U18122 (N_18122,N_14153,N_12743);
xor U18123 (N_18123,N_13561,N_12489);
nand U18124 (N_18124,N_12162,N_13174);
nor U18125 (N_18125,N_13279,N_13562);
xor U18126 (N_18126,N_15620,N_13197);
nand U18127 (N_18127,N_12185,N_14893);
xor U18128 (N_18128,N_13582,N_14632);
and U18129 (N_18129,N_13234,N_14068);
and U18130 (N_18130,N_15644,N_13713);
and U18131 (N_18131,N_12644,N_12113);
or U18132 (N_18132,N_14033,N_14544);
nor U18133 (N_18133,N_13981,N_12565);
xnor U18134 (N_18134,N_15398,N_12476);
nand U18135 (N_18135,N_12777,N_14519);
xor U18136 (N_18136,N_14707,N_12970);
nor U18137 (N_18137,N_15814,N_12934);
nor U18138 (N_18138,N_13395,N_14142);
xor U18139 (N_18139,N_15249,N_14761);
or U18140 (N_18140,N_13509,N_12772);
or U18141 (N_18141,N_14293,N_14112);
and U18142 (N_18142,N_15781,N_14143);
nand U18143 (N_18143,N_14417,N_12605);
and U18144 (N_18144,N_13309,N_15760);
and U18145 (N_18145,N_14181,N_14898);
and U18146 (N_18146,N_13408,N_12595);
and U18147 (N_18147,N_12891,N_13798);
xor U18148 (N_18148,N_14891,N_13140);
nand U18149 (N_18149,N_13831,N_12962);
nor U18150 (N_18150,N_13415,N_15911);
and U18151 (N_18151,N_12822,N_13586);
or U18152 (N_18152,N_15542,N_15790);
nor U18153 (N_18153,N_14948,N_13693);
nand U18154 (N_18154,N_12415,N_14115);
or U18155 (N_18155,N_14796,N_13720);
and U18156 (N_18156,N_15850,N_15695);
or U18157 (N_18157,N_15227,N_15672);
and U18158 (N_18158,N_14864,N_12475);
nand U18159 (N_18159,N_12072,N_14597);
and U18160 (N_18160,N_14904,N_12001);
nand U18161 (N_18161,N_12290,N_13942);
and U18162 (N_18162,N_14266,N_12954);
nor U18163 (N_18163,N_13057,N_15881);
nand U18164 (N_18164,N_15797,N_12935);
and U18165 (N_18165,N_13206,N_13953);
nor U18166 (N_18166,N_12959,N_14620);
or U18167 (N_18167,N_14014,N_13766);
nand U18168 (N_18168,N_13094,N_12665);
or U18169 (N_18169,N_14952,N_12489);
and U18170 (N_18170,N_12721,N_12203);
and U18171 (N_18171,N_13821,N_14676);
and U18172 (N_18172,N_15013,N_13469);
nor U18173 (N_18173,N_14430,N_14387);
nand U18174 (N_18174,N_14966,N_14611);
nor U18175 (N_18175,N_15646,N_12358);
and U18176 (N_18176,N_12071,N_13518);
or U18177 (N_18177,N_14608,N_12108);
xor U18178 (N_18178,N_14508,N_13440);
or U18179 (N_18179,N_12339,N_12694);
or U18180 (N_18180,N_12610,N_14865);
xnor U18181 (N_18181,N_14095,N_15441);
or U18182 (N_18182,N_12027,N_15480);
or U18183 (N_18183,N_12624,N_12121);
nand U18184 (N_18184,N_14278,N_15882);
and U18185 (N_18185,N_12649,N_14072);
nor U18186 (N_18186,N_12007,N_15497);
xor U18187 (N_18187,N_14761,N_12104);
nor U18188 (N_18188,N_14607,N_13366);
nand U18189 (N_18189,N_14670,N_12783);
nand U18190 (N_18190,N_14427,N_14606);
and U18191 (N_18191,N_13970,N_12148);
nor U18192 (N_18192,N_12245,N_14052);
nand U18193 (N_18193,N_13784,N_12856);
nor U18194 (N_18194,N_13872,N_14536);
or U18195 (N_18195,N_12634,N_15854);
nand U18196 (N_18196,N_13083,N_13625);
nor U18197 (N_18197,N_12343,N_12187);
or U18198 (N_18198,N_15945,N_12075);
xor U18199 (N_18199,N_15067,N_13002);
and U18200 (N_18200,N_13489,N_15955);
or U18201 (N_18201,N_15287,N_14403);
xnor U18202 (N_18202,N_15165,N_12659);
and U18203 (N_18203,N_13617,N_14913);
xnor U18204 (N_18204,N_15891,N_12538);
nor U18205 (N_18205,N_14748,N_13938);
nand U18206 (N_18206,N_15497,N_15806);
or U18207 (N_18207,N_12304,N_12791);
xor U18208 (N_18208,N_15514,N_15008);
nor U18209 (N_18209,N_13108,N_15148);
nand U18210 (N_18210,N_12512,N_13471);
xnor U18211 (N_18211,N_14549,N_13561);
nand U18212 (N_18212,N_15316,N_13503);
nor U18213 (N_18213,N_14306,N_14789);
xor U18214 (N_18214,N_12522,N_15541);
and U18215 (N_18215,N_15613,N_12248);
nand U18216 (N_18216,N_15171,N_12165);
nor U18217 (N_18217,N_15112,N_14419);
nand U18218 (N_18218,N_15170,N_13520);
nor U18219 (N_18219,N_12323,N_14490);
nand U18220 (N_18220,N_14711,N_12316);
or U18221 (N_18221,N_14760,N_13892);
xor U18222 (N_18222,N_13847,N_14202);
nor U18223 (N_18223,N_13317,N_15796);
nand U18224 (N_18224,N_15860,N_15249);
nand U18225 (N_18225,N_14814,N_13841);
or U18226 (N_18226,N_14230,N_12561);
and U18227 (N_18227,N_12715,N_12282);
nand U18228 (N_18228,N_13119,N_12711);
nor U18229 (N_18229,N_12654,N_15719);
nor U18230 (N_18230,N_13148,N_14599);
or U18231 (N_18231,N_13672,N_15695);
or U18232 (N_18232,N_13434,N_13374);
nand U18233 (N_18233,N_14586,N_13247);
or U18234 (N_18234,N_15301,N_12094);
or U18235 (N_18235,N_13511,N_12666);
xor U18236 (N_18236,N_15789,N_13544);
nor U18237 (N_18237,N_14575,N_12284);
nand U18238 (N_18238,N_15731,N_13696);
and U18239 (N_18239,N_13732,N_12001);
and U18240 (N_18240,N_14131,N_14386);
and U18241 (N_18241,N_12419,N_14257);
nor U18242 (N_18242,N_14802,N_13508);
and U18243 (N_18243,N_12293,N_13986);
nand U18244 (N_18244,N_14757,N_15955);
xor U18245 (N_18245,N_12881,N_12407);
nand U18246 (N_18246,N_14939,N_13983);
and U18247 (N_18247,N_15241,N_15385);
and U18248 (N_18248,N_15526,N_14831);
or U18249 (N_18249,N_15419,N_13627);
nand U18250 (N_18250,N_13541,N_14533);
or U18251 (N_18251,N_15597,N_13429);
and U18252 (N_18252,N_15918,N_12566);
and U18253 (N_18253,N_15489,N_12681);
and U18254 (N_18254,N_12713,N_12146);
and U18255 (N_18255,N_14339,N_15808);
or U18256 (N_18256,N_15517,N_13041);
or U18257 (N_18257,N_14951,N_12968);
or U18258 (N_18258,N_14160,N_13728);
nand U18259 (N_18259,N_15253,N_13224);
and U18260 (N_18260,N_12806,N_12209);
nor U18261 (N_18261,N_14745,N_14596);
or U18262 (N_18262,N_12495,N_12778);
xnor U18263 (N_18263,N_14318,N_12812);
and U18264 (N_18264,N_15826,N_12803);
or U18265 (N_18265,N_12927,N_13284);
nor U18266 (N_18266,N_14072,N_12971);
nor U18267 (N_18267,N_15115,N_12537);
nor U18268 (N_18268,N_13727,N_15372);
and U18269 (N_18269,N_12801,N_15469);
nand U18270 (N_18270,N_15153,N_12716);
and U18271 (N_18271,N_12879,N_13433);
and U18272 (N_18272,N_13610,N_12192);
or U18273 (N_18273,N_14102,N_12709);
nand U18274 (N_18274,N_15024,N_12054);
nand U18275 (N_18275,N_13755,N_12494);
nand U18276 (N_18276,N_13914,N_12620);
nand U18277 (N_18277,N_13523,N_12381);
nor U18278 (N_18278,N_13316,N_12967);
nor U18279 (N_18279,N_13988,N_13558);
nand U18280 (N_18280,N_14476,N_14627);
and U18281 (N_18281,N_13677,N_14999);
nand U18282 (N_18282,N_14960,N_15519);
nor U18283 (N_18283,N_15478,N_12647);
nand U18284 (N_18284,N_13867,N_12298);
nand U18285 (N_18285,N_12183,N_14117);
and U18286 (N_18286,N_12399,N_12730);
and U18287 (N_18287,N_15869,N_15377);
and U18288 (N_18288,N_14322,N_14698);
nor U18289 (N_18289,N_13950,N_12292);
nor U18290 (N_18290,N_15763,N_13985);
and U18291 (N_18291,N_12921,N_13697);
and U18292 (N_18292,N_14417,N_12568);
nand U18293 (N_18293,N_12049,N_15836);
xnor U18294 (N_18294,N_14189,N_15747);
xnor U18295 (N_18295,N_13615,N_12860);
or U18296 (N_18296,N_15436,N_14063);
nor U18297 (N_18297,N_12910,N_15530);
and U18298 (N_18298,N_13868,N_13828);
or U18299 (N_18299,N_13640,N_12912);
nor U18300 (N_18300,N_12823,N_15443);
nor U18301 (N_18301,N_15356,N_14659);
xor U18302 (N_18302,N_12808,N_14685);
xnor U18303 (N_18303,N_13670,N_15753);
and U18304 (N_18304,N_14560,N_14237);
or U18305 (N_18305,N_14891,N_15025);
or U18306 (N_18306,N_14153,N_12286);
or U18307 (N_18307,N_14746,N_13314);
nor U18308 (N_18308,N_12212,N_14059);
and U18309 (N_18309,N_15951,N_15200);
nand U18310 (N_18310,N_12899,N_13037);
and U18311 (N_18311,N_13076,N_12560);
nor U18312 (N_18312,N_12444,N_15456);
nor U18313 (N_18313,N_14935,N_13983);
xor U18314 (N_18314,N_15806,N_14175);
or U18315 (N_18315,N_15911,N_14952);
and U18316 (N_18316,N_15891,N_12070);
or U18317 (N_18317,N_13270,N_15844);
xnor U18318 (N_18318,N_14434,N_12382);
nand U18319 (N_18319,N_13139,N_14598);
and U18320 (N_18320,N_14832,N_15950);
nand U18321 (N_18321,N_15447,N_13388);
or U18322 (N_18322,N_13622,N_14406);
nor U18323 (N_18323,N_14984,N_15959);
and U18324 (N_18324,N_12061,N_14863);
xnor U18325 (N_18325,N_15627,N_13107);
and U18326 (N_18326,N_13467,N_14096);
xnor U18327 (N_18327,N_13695,N_12660);
xor U18328 (N_18328,N_13250,N_12391);
nor U18329 (N_18329,N_14553,N_14371);
nand U18330 (N_18330,N_14641,N_15682);
xor U18331 (N_18331,N_15041,N_13515);
or U18332 (N_18332,N_15317,N_15726);
and U18333 (N_18333,N_15499,N_14193);
or U18334 (N_18334,N_15040,N_12591);
and U18335 (N_18335,N_12416,N_14263);
or U18336 (N_18336,N_14684,N_13191);
nor U18337 (N_18337,N_12119,N_13614);
or U18338 (N_18338,N_14903,N_15418);
nand U18339 (N_18339,N_15427,N_13839);
or U18340 (N_18340,N_12893,N_13879);
nand U18341 (N_18341,N_13402,N_13922);
and U18342 (N_18342,N_14217,N_14518);
nand U18343 (N_18343,N_15712,N_14288);
xnor U18344 (N_18344,N_14581,N_15494);
or U18345 (N_18345,N_13234,N_12264);
or U18346 (N_18346,N_12789,N_13803);
nand U18347 (N_18347,N_14554,N_14450);
nand U18348 (N_18348,N_14256,N_13213);
or U18349 (N_18349,N_12129,N_12957);
nor U18350 (N_18350,N_13397,N_12546);
nor U18351 (N_18351,N_12622,N_13357);
or U18352 (N_18352,N_14531,N_12875);
nand U18353 (N_18353,N_14768,N_13566);
nor U18354 (N_18354,N_13360,N_14803);
nor U18355 (N_18355,N_14032,N_15424);
and U18356 (N_18356,N_15198,N_15669);
or U18357 (N_18357,N_12401,N_12225);
and U18358 (N_18358,N_15122,N_13105);
nand U18359 (N_18359,N_14698,N_12957);
and U18360 (N_18360,N_12961,N_13693);
nand U18361 (N_18361,N_14356,N_12067);
xor U18362 (N_18362,N_15474,N_15910);
and U18363 (N_18363,N_15821,N_14281);
or U18364 (N_18364,N_12636,N_15746);
nand U18365 (N_18365,N_13390,N_12931);
and U18366 (N_18366,N_15840,N_14161);
and U18367 (N_18367,N_14792,N_13898);
or U18368 (N_18368,N_14538,N_14793);
nor U18369 (N_18369,N_15207,N_13775);
nor U18370 (N_18370,N_12680,N_12142);
nor U18371 (N_18371,N_15721,N_12845);
nor U18372 (N_18372,N_14123,N_15370);
xor U18373 (N_18373,N_12390,N_12655);
nor U18374 (N_18374,N_14419,N_14488);
nand U18375 (N_18375,N_14227,N_13123);
nor U18376 (N_18376,N_12261,N_13294);
xnor U18377 (N_18377,N_13924,N_15146);
and U18378 (N_18378,N_13306,N_14810);
or U18379 (N_18379,N_13023,N_14983);
and U18380 (N_18380,N_14265,N_15924);
xnor U18381 (N_18381,N_13379,N_12398);
nor U18382 (N_18382,N_15666,N_14547);
nor U18383 (N_18383,N_13075,N_15232);
xnor U18384 (N_18384,N_12358,N_14800);
nor U18385 (N_18385,N_12518,N_12999);
or U18386 (N_18386,N_14349,N_14814);
xnor U18387 (N_18387,N_12614,N_12625);
nor U18388 (N_18388,N_14316,N_14165);
and U18389 (N_18389,N_13306,N_14506);
or U18390 (N_18390,N_14542,N_14568);
or U18391 (N_18391,N_14870,N_12973);
and U18392 (N_18392,N_14716,N_14861);
nor U18393 (N_18393,N_15657,N_12000);
nor U18394 (N_18394,N_12653,N_12833);
nor U18395 (N_18395,N_14378,N_12827);
or U18396 (N_18396,N_13045,N_13393);
nand U18397 (N_18397,N_13129,N_14571);
nand U18398 (N_18398,N_13030,N_12743);
nand U18399 (N_18399,N_14359,N_13780);
and U18400 (N_18400,N_15032,N_15943);
nand U18401 (N_18401,N_12739,N_15086);
and U18402 (N_18402,N_13101,N_12446);
and U18403 (N_18403,N_12775,N_12783);
xnor U18404 (N_18404,N_13054,N_12880);
nand U18405 (N_18405,N_13133,N_12690);
or U18406 (N_18406,N_14966,N_15117);
and U18407 (N_18407,N_15367,N_14760);
nand U18408 (N_18408,N_12173,N_15773);
nor U18409 (N_18409,N_14491,N_13799);
nand U18410 (N_18410,N_12788,N_13047);
or U18411 (N_18411,N_12446,N_12287);
or U18412 (N_18412,N_12875,N_14110);
nor U18413 (N_18413,N_13299,N_13790);
and U18414 (N_18414,N_14731,N_15152);
or U18415 (N_18415,N_13953,N_14011);
nor U18416 (N_18416,N_12278,N_13093);
nand U18417 (N_18417,N_15125,N_14966);
and U18418 (N_18418,N_13647,N_15505);
and U18419 (N_18419,N_15623,N_14255);
or U18420 (N_18420,N_15045,N_12117);
nor U18421 (N_18421,N_14819,N_15997);
nor U18422 (N_18422,N_13998,N_13660);
nor U18423 (N_18423,N_14771,N_12362);
xor U18424 (N_18424,N_12086,N_15755);
and U18425 (N_18425,N_13807,N_15225);
and U18426 (N_18426,N_15271,N_12528);
nand U18427 (N_18427,N_12284,N_14302);
xor U18428 (N_18428,N_14856,N_12453);
or U18429 (N_18429,N_15277,N_15996);
or U18430 (N_18430,N_15703,N_15252);
or U18431 (N_18431,N_14659,N_12123);
or U18432 (N_18432,N_13327,N_14370);
and U18433 (N_18433,N_14520,N_15545);
nand U18434 (N_18434,N_14468,N_12506);
xnor U18435 (N_18435,N_15668,N_12349);
xor U18436 (N_18436,N_12026,N_12239);
or U18437 (N_18437,N_14113,N_14895);
or U18438 (N_18438,N_15975,N_14270);
nand U18439 (N_18439,N_12066,N_13613);
nor U18440 (N_18440,N_12118,N_15490);
xnor U18441 (N_18441,N_13191,N_14579);
and U18442 (N_18442,N_13210,N_12668);
and U18443 (N_18443,N_14194,N_14286);
and U18444 (N_18444,N_14514,N_15794);
and U18445 (N_18445,N_12353,N_13076);
nor U18446 (N_18446,N_14208,N_14168);
and U18447 (N_18447,N_15818,N_15444);
or U18448 (N_18448,N_13716,N_15212);
and U18449 (N_18449,N_14429,N_13255);
nor U18450 (N_18450,N_14719,N_14254);
or U18451 (N_18451,N_12747,N_14129);
nand U18452 (N_18452,N_15015,N_14249);
nor U18453 (N_18453,N_12291,N_13664);
and U18454 (N_18454,N_14957,N_12563);
nor U18455 (N_18455,N_14647,N_15134);
and U18456 (N_18456,N_12247,N_14639);
xnor U18457 (N_18457,N_14183,N_15505);
or U18458 (N_18458,N_15664,N_14715);
nor U18459 (N_18459,N_15203,N_13292);
and U18460 (N_18460,N_13181,N_15649);
nor U18461 (N_18461,N_13042,N_12929);
or U18462 (N_18462,N_14502,N_13457);
and U18463 (N_18463,N_15318,N_13658);
nor U18464 (N_18464,N_15526,N_12082);
and U18465 (N_18465,N_13018,N_14540);
nor U18466 (N_18466,N_14097,N_12041);
nand U18467 (N_18467,N_14074,N_12278);
and U18468 (N_18468,N_14024,N_13833);
nor U18469 (N_18469,N_15099,N_14349);
xor U18470 (N_18470,N_15882,N_15491);
or U18471 (N_18471,N_15172,N_14814);
or U18472 (N_18472,N_14392,N_13359);
nor U18473 (N_18473,N_15533,N_14244);
or U18474 (N_18474,N_14047,N_15456);
nor U18475 (N_18475,N_14232,N_14932);
nor U18476 (N_18476,N_13637,N_14693);
or U18477 (N_18477,N_15367,N_12380);
nor U18478 (N_18478,N_15020,N_13524);
and U18479 (N_18479,N_15524,N_12490);
and U18480 (N_18480,N_13972,N_12541);
nand U18481 (N_18481,N_15234,N_12380);
nor U18482 (N_18482,N_12212,N_12458);
or U18483 (N_18483,N_14169,N_14751);
nand U18484 (N_18484,N_15590,N_15056);
nor U18485 (N_18485,N_13114,N_15523);
nor U18486 (N_18486,N_13295,N_14410);
nor U18487 (N_18487,N_13299,N_15619);
nor U18488 (N_18488,N_12968,N_12289);
nor U18489 (N_18489,N_12781,N_12976);
or U18490 (N_18490,N_13436,N_12364);
nor U18491 (N_18491,N_15765,N_15614);
nand U18492 (N_18492,N_12356,N_12327);
nand U18493 (N_18493,N_14738,N_12063);
nand U18494 (N_18494,N_12168,N_12119);
nor U18495 (N_18495,N_14278,N_15265);
nand U18496 (N_18496,N_12561,N_13299);
and U18497 (N_18497,N_14285,N_14296);
and U18498 (N_18498,N_14397,N_13639);
and U18499 (N_18499,N_14250,N_14717);
or U18500 (N_18500,N_14755,N_15161);
or U18501 (N_18501,N_13717,N_15520);
nor U18502 (N_18502,N_14356,N_12715);
nor U18503 (N_18503,N_12327,N_12616);
and U18504 (N_18504,N_12153,N_15271);
nor U18505 (N_18505,N_15991,N_13699);
and U18506 (N_18506,N_15762,N_13794);
and U18507 (N_18507,N_14341,N_12972);
or U18508 (N_18508,N_13824,N_15388);
or U18509 (N_18509,N_12668,N_14736);
or U18510 (N_18510,N_13928,N_14141);
nand U18511 (N_18511,N_15248,N_15644);
and U18512 (N_18512,N_13381,N_14909);
and U18513 (N_18513,N_13182,N_12611);
or U18514 (N_18514,N_14467,N_14555);
nand U18515 (N_18515,N_13728,N_15594);
nor U18516 (N_18516,N_12670,N_13202);
nand U18517 (N_18517,N_13021,N_15282);
and U18518 (N_18518,N_15843,N_12494);
or U18519 (N_18519,N_13700,N_12320);
nand U18520 (N_18520,N_14727,N_13991);
nor U18521 (N_18521,N_15388,N_14856);
nor U18522 (N_18522,N_14650,N_12104);
and U18523 (N_18523,N_14723,N_14083);
nand U18524 (N_18524,N_12085,N_14170);
nor U18525 (N_18525,N_12158,N_13367);
nand U18526 (N_18526,N_12716,N_13774);
or U18527 (N_18527,N_13561,N_12781);
nand U18528 (N_18528,N_12794,N_14743);
nand U18529 (N_18529,N_13118,N_14412);
nand U18530 (N_18530,N_14761,N_14759);
and U18531 (N_18531,N_12712,N_14598);
xor U18532 (N_18532,N_14890,N_13659);
nor U18533 (N_18533,N_14726,N_12196);
and U18534 (N_18534,N_15352,N_15668);
nor U18535 (N_18535,N_15505,N_14307);
or U18536 (N_18536,N_13426,N_13277);
or U18537 (N_18537,N_14033,N_14419);
nand U18538 (N_18538,N_14610,N_13508);
nand U18539 (N_18539,N_15164,N_12571);
or U18540 (N_18540,N_12194,N_15608);
and U18541 (N_18541,N_14216,N_14899);
xor U18542 (N_18542,N_13497,N_14544);
or U18543 (N_18543,N_13179,N_14663);
nor U18544 (N_18544,N_15673,N_12032);
or U18545 (N_18545,N_12337,N_14678);
nand U18546 (N_18546,N_14404,N_15368);
or U18547 (N_18547,N_15441,N_15345);
nand U18548 (N_18548,N_13015,N_14873);
or U18549 (N_18549,N_15111,N_15443);
and U18550 (N_18550,N_12138,N_12406);
nand U18551 (N_18551,N_13601,N_14240);
nand U18552 (N_18552,N_15305,N_15910);
nor U18553 (N_18553,N_15288,N_15804);
nand U18554 (N_18554,N_14880,N_13753);
nor U18555 (N_18555,N_13159,N_12513);
or U18556 (N_18556,N_13189,N_12785);
and U18557 (N_18557,N_15870,N_13696);
nor U18558 (N_18558,N_13194,N_15952);
xor U18559 (N_18559,N_13066,N_15457);
nand U18560 (N_18560,N_15066,N_15621);
nor U18561 (N_18561,N_13393,N_12599);
and U18562 (N_18562,N_15790,N_13829);
and U18563 (N_18563,N_13771,N_13321);
or U18564 (N_18564,N_12644,N_12236);
or U18565 (N_18565,N_15064,N_12372);
and U18566 (N_18566,N_13272,N_15072);
nor U18567 (N_18567,N_13671,N_14909);
or U18568 (N_18568,N_15842,N_12652);
or U18569 (N_18569,N_13989,N_15553);
or U18570 (N_18570,N_13672,N_14149);
or U18571 (N_18571,N_15561,N_13607);
xor U18572 (N_18572,N_12870,N_15626);
and U18573 (N_18573,N_14000,N_13485);
nand U18574 (N_18574,N_12358,N_12447);
and U18575 (N_18575,N_15127,N_13945);
nand U18576 (N_18576,N_12749,N_12239);
or U18577 (N_18577,N_13325,N_14909);
and U18578 (N_18578,N_12379,N_14980);
nor U18579 (N_18579,N_15051,N_15069);
nand U18580 (N_18580,N_13237,N_14455);
and U18581 (N_18581,N_14878,N_13521);
or U18582 (N_18582,N_12926,N_12042);
nand U18583 (N_18583,N_14132,N_12914);
nand U18584 (N_18584,N_12604,N_14763);
xnor U18585 (N_18585,N_15507,N_14228);
and U18586 (N_18586,N_12359,N_14894);
and U18587 (N_18587,N_13796,N_13790);
nor U18588 (N_18588,N_12156,N_15393);
nor U18589 (N_18589,N_15459,N_15798);
and U18590 (N_18590,N_12595,N_14120);
nand U18591 (N_18591,N_12930,N_12975);
nand U18592 (N_18592,N_15646,N_15904);
nor U18593 (N_18593,N_15381,N_12064);
nand U18594 (N_18594,N_13231,N_15476);
nor U18595 (N_18595,N_15833,N_15984);
nor U18596 (N_18596,N_14747,N_14966);
and U18597 (N_18597,N_14139,N_15262);
and U18598 (N_18598,N_14017,N_13371);
xor U18599 (N_18599,N_13763,N_15677);
and U18600 (N_18600,N_14828,N_14878);
nand U18601 (N_18601,N_14890,N_15479);
nand U18602 (N_18602,N_12005,N_12961);
xnor U18603 (N_18603,N_12908,N_15379);
and U18604 (N_18604,N_12729,N_15026);
or U18605 (N_18605,N_14698,N_12144);
xor U18606 (N_18606,N_12644,N_14640);
and U18607 (N_18607,N_14226,N_14534);
nor U18608 (N_18608,N_12291,N_13960);
and U18609 (N_18609,N_13191,N_15225);
or U18610 (N_18610,N_12790,N_13865);
nand U18611 (N_18611,N_12312,N_13459);
or U18612 (N_18612,N_15280,N_14366);
nor U18613 (N_18613,N_14578,N_15502);
nand U18614 (N_18614,N_12267,N_15459);
and U18615 (N_18615,N_15068,N_13142);
or U18616 (N_18616,N_13508,N_14290);
and U18617 (N_18617,N_13253,N_14194);
and U18618 (N_18618,N_14526,N_15511);
nand U18619 (N_18619,N_12688,N_13586);
or U18620 (N_18620,N_15412,N_12436);
or U18621 (N_18621,N_14100,N_14439);
nand U18622 (N_18622,N_15798,N_13035);
and U18623 (N_18623,N_14867,N_15133);
or U18624 (N_18624,N_13694,N_15412);
and U18625 (N_18625,N_12038,N_14454);
xnor U18626 (N_18626,N_12793,N_12714);
and U18627 (N_18627,N_12791,N_15144);
or U18628 (N_18628,N_12612,N_14596);
and U18629 (N_18629,N_13717,N_14843);
xnor U18630 (N_18630,N_15946,N_13352);
or U18631 (N_18631,N_14258,N_12252);
or U18632 (N_18632,N_14933,N_14632);
and U18633 (N_18633,N_12072,N_15169);
nand U18634 (N_18634,N_14055,N_14792);
xnor U18635 (N_18635,N_15287,N_14008);
or U18636 (N_18636,N_12232,N_14834);
nand U18637 (N_18637,N_15191,N_15535);
and U18638 (N_18638,N_15542,N_14303);
and U18639 (N_18639,N_13757,N_15319);
nand U18640 (N_18640,N_15780,N_13112);
nor U18641 (N_18641,N_14865,N_12403);
xnor U18642 (N_18642,N_14971,N_15729);
nand U18643 (N_18643,N_12365,N_14161);
and U18644 (N_18644,N_12544,N_14667);
xnor U18645 (N_18645,N_13273,N_14793);
and U18646 (N_18646,N_13228,N_12249);
and U18647 (N_18647,N_13992,N_15044);
nor U18648 (N_18648,N_14353,N_12180);
nand U18649 (N_18649,N_13187,N_12133);
nand U18650 (N_18650,N_14876,N_15445);
nand U18651 (N_18651,N_15134,N_15466);
and U18652 (N_18652,N_15969,N_12767);
nand U18653 (N_18653,N_14977,N_12938);
nand U18654 (N_18654,N_12866,N_12862);
and U18655 (N_18655,N_15155,N_13740);
and U18656 (N_18656,N_14237,N_15950);
nor U18657 (N_18657,N_14276,N_15868);
xor U18658 (N_18658,N_13407,N_12876);
nor U18659 (N_18659,N_14075,N_14459);
nand U18660 (N_18660,N_14900,N_14521);
nor U18661 (N_18661,N_15944,N_12615);
xnor U18662 (N_18662,N_14577,N_13190);
nand U18663 (N_18663,N_14423,N_14550);
or U18664 (N_18664,N_15191,N_14886);
or U18665 (N_18665,N_14169,N_14584);
nor U18666 (N_18666,N_14879,N_14965);
nand U18667 (N_18667,N_13252,N_15799);
or U18668 (N_18668,N_15078,N_12548);
nor U18669 (N_18669,N_12773,N_14588);
nand U18670 (N_18670,N_15639,N_14064);
xor U18671 (N_18671,N_12407,N_12071);
or U18672 (N_18672,N_14139,N_14438);
and U18673 (N_18673,N_12466,N_14458);
nand U18674 (N_18674,N_12124,N_14157);
and U18675 (N_18675,N_15629,N_14037);
and U18676 (N_18676,N_15656,N_12158);
nor U18677 (N_18677,N_15750,N_15204);
or U18678 (N_18678,N_14254,N_12983);
nand U18679 (N_18679,N_12367,N_15727);
nor U18680 (N_18680,N_13302,N_12947);
or U18681 (N_18681,N_13730,N_12068);
nor U18682 (N_18682,N_15009,N_13845);
and U18683 (N_18683,N_15244,N_15556);
nor U18684 (N_18684,N_13450,N_13213);
or U18685 (N_18685,N_15050,N_15764);
or U18686 (N_18686,N_12898,N_13936);
xnor U18687 (N_18687,N_13928,N_12273);
or U18688 (N_18688,N_14009,N_13747);
or U18689 (N_18689,N_14294,N_13154);
nor U18690 (N_18690,N_13444,N_14328);
nor U18691 (N_18691,N_15077,N_14463);
and U18692 (N_18692,N_12901,N_12684);
nand U18693 (N_18693,N_15923,N_14040);
nand U18694 (N_18694,N_15478,N_14814);
or U18695 (N_18695,N_12517,N_15630);
nor U18696 (N_18696,N_13259,N_13104);
nand U18697 (N_18697,N_12388,N_15793);
nor U18698 (N_18698,N_15647,N_12763);
nand U18699 (N_18699,N_14613,N_15372);
nor U18700 (N_18700,N_13553,N_15642);
nand U18701 (N_18701,N_14400,N_15846);
nor U18702 (N_18702,N_13037,N_15937);
nor U18703 (N_18703,N_13493,N_14614);
or U18704 (N_18704,N_14848,N_15752);
xor U18705 (N_18705,N_15298,N_12385);
nand U18706 (N_18706,N_14019,N_13042);
and U18707 (N_18707,N_14402,N_13139);
nor U18708 (N_18708,N_12864,N_13914);
and U18709 (N_18709,N_12950,N_12954);
and U18710 (N_18710,N_13374,N_14048);
nor U18711 (N_18711,N_12583,N_13404);
nand U18712 (N_18712,N_13902,N_14327);
nor U18713 (N_18713,N_15890,N_14547);
or U18714 (N_18714,N_12352,N_13327);
and U18715 (N_18715,N_12652,N_12354);
nor U18716 (N_18716,N_13810,N_13046);
nand U18717 (N_18717,N_12551,N_15044);
nand U18718 (N_18718,N_14372,N_15402);
or U18719 (N_18719,N_15507,N_12757);
nor U18720 (N_18720,N_12017,N_15581);
nor U18721 (N_18721,N_12716,N_13843);
nor U18722 (N_18722,N_12163,N_13265);
nor U18723 (N_18723,N_13257,N_14103);
nand U18724 (N_18724,N_15560,N_15571);
nand U18725 (N_18725,N_14322,N_14185);
and U18726 (N_18726,N_14139,N_14768);
nor U18727 (N_18727,N_13849,N_15079);
nand U18728 (N_18728,N_14988,N_13198);
or U18729 (N_18729,N_12440,N_12854);
or U18730 (N_18730,N_13279,N_14082);
and U18731 (N_18731,N_15506,N_15793);
nor U18732 (N_18732,N_14599,N_14859);
nand U18733 (N_18733,N_14978,N_15439);
nor U18734 (N_18734,N_15766,N_12022);
nand U18735 (N_18735,N_14015,N_15113);
nand U18736 (N_18736,N_13344,N_14424);
or U18737 (N_18737,N_12509,N_15927);
nand U18738 (N_18738,N_14105,N_14319);
or U18739 (N_18739,N_14882,N_12434);
nand U18740 (N_18740,N_13588,N_13952);
nand U18741 (N_18741,N_14194,N_15006);
nor U18742 (N_18742,N_15122,N_15693);
or U18743 (N_18743,N_14278,N_13190);
and U18744 (N_18744,N_13008,N_14969);
nand U18745 (N_18745,N_15819,N_13399);
nand U18746 (N_18746,N_15611,N_15487);
xor U18747 (N_18747,N_14479,N_13022);
nor U18748 (N_18748,N_15501,N_15932);
or U18749 (N_18749,N_12333,N_12084);
and U18750 (N_18750,N_13549,N_15660);
and U18751 (N_18751,N_12340,N_14631);
nor U18752 (N_18752,N_13793,N_12859);
and U18753 (N_18753,N_13498,N_14108);
or U18754 (N_18754,N_13069,N_14844);
nand U18755 (N_18755,N_14601,N_13280);
nand U18756 (N_18756,N_15066,N_13429);
nand U18757 (N_18757,N_13801,N_13893);
nor U18758 (N_18758,N_15281,N_12877);
and U18759 (N_18759,N_13545,N_14100);
xnor U18760 (N_18760,N_14006,N_13225);
nand U18761 (N_18761,N_13085,N_15157);
nor U18762 (N_18762,N_15366,N_14340);
nor U18763 (N_18763,N_15175,N_13772);
or U18764 (N_18764,N_14930,N_12230);
nor U18765 (N_18765,N_13050,N_15522);
nor U18766 (N_18766,N_15417,N_14335);
and U18767 (N_18767,N_15682,N_13514);
xor U18768 (N_18768,N_13126,N_13268);
nor U18769 (N_18769,N_12531,N_12323);
or U18770 (N_18770,N_13213,N_15125);
nor U18771 (N_18771,N_12413,N_14483);
and U18772 (N_18772,N_12009,N_15183);
or U18773 (N_18773,N_15523,N_12927);
or U18774 (N_18774,N_14182,N_13032);
and U18775 (N_18775,N_15576,N_14084);
nand U18776 (N_18776,N_13939,N_13582);
nor U18777 (N_18777,N_12806,N_15554);
and U18778 (N_18778,N_14792,N_15745);
nor U18779 (N_18779,N_14726,N_15071);
and U18780 (N_18780,N_14173,N_13914);
and U18781 (N_18781,N_13409,N_14085);
nor U18782 (N_18782,N_12861,N_15201);
xnor U18783 (N_18783,N_14530,N_13732);
and U18784 (N_18784,N_15165,N_15753);
and U18785 (N_18785,N_13926,N_14568);
nor U18786 (N_18786,N_12407,N_15627);
or U18787 (N_18787,N_13179,N_12598);
and U18788 (N_18788,N_15430,N_12777);
and U18789 (N_18789,N_15470,N_13322);
and U18790 (N_18790,N_13549,N_13388);
or U18791 (N_18791,N_15596,N_12428);
and U18792 (N_18792,N_15217,N_15609);
nand U18793 (N_18793,N_12069,N_15451);
nor U18794 (N_18794,N_13155,N_13009);
nor U18795 (N_18795,N_14907,N_13352);
nor U18796 (N_18796,N_15807,N_14436);
and U18797 (N_18797,N_12357,N_13243);
and U18798 (N_18798,N_15890,N_12007);
or U18799 (N_18799,N_13737,N_12711);
or U18800 (N_18800,N_15745,N_15139);
and U18801 (N_18801,N_13220,N_13573);
and U18802 (N_18802,N_15947,N_15752);
nor U18803 (N_18803,N_15389,N_12580);
xor U18804 (N_18804,N_15866,N_12712);
xor U18805 (N_18805,N_15424,N_12653);
nand U18806 (N_18806,N_12259,N_12066);
nand U18807 (N_18807,N_12618,N_15808);
nand U18808 (N_18808,N_15389,N_14981);
and U18809 (N_18809,N_14731,N_13317);
xor U18810 (N_18810,N_15499,N_13859);
and U18811 (N_18811,N_12600,N_12579);
nor U18812 (N_18812,N_12582,N_15955);
nand U18813 (N_18813,N_13034,N_14763);
xor U18814 (N_18814,N_12658,N_13157);
and U18815 (N_18815,N_12405,N_12953);
nand U18816 (N_18816,N_13771,N_12689);
or U18817 (N_18817,N_14588,N_13751);
and U18818 (N_18818,N_14729,N_15954);
xnor U18819 (N_18819,N_15842,N_13407);
or U18820 (N_18820,N_14227,N_15796);
nand U18821 (N_18821,N_14090,N_14264);
nand U18822 (N_18822,N_12558,N_14610);
nor U18823 (N_18823,N_15877,N_13147);
and U18824 (N_18824,N_12555,N_14813);
and U18825 (N_18825,N_12976,N_13017);
nand U18826 (N_18826,N_15973,N_15136);
or U18827 (N_18827,N_12540,N_14034);
nand U18828 (N_18828,N_13556,N_15693);
or U18829 (N_18829,N_13887,N_13764);
nand U18830 (N_18830,N_14253,N_12976);
and U18831 (N_18831,N_14110,N_13262);
xnor U18832 (N_18832,N_13288,N_13453);
nand U18833 (N_18833,N_12607,N_12148);
xnor U18834 (N_18834,N_12564,N_12083);
nor U18835 (N_18835,N_14030,N_13732);
nor U18836 (N_18836,N_12035,N_14800);
nand U18837 (N_18837,N_13063,N_14129);
or U18838 (N_18838,N_13819,N_14517);
and U18839 (N_18839,N_13998,N_12197);
and U18840 (N_18840,N_15930,N_12409);
or U18841 (N_18841,N_13655,N_13134);
or U18842 (N_18842,N_12927,N_12586);
nand U18843 (N_18843,N_14750,N_15680);
or U18844 (N_18844,N_13396,N_13674);
and U18845 (N_18845,N_12524,N_12899);
and U18846 (N_18846,N_15494,N_12557);
or U18847 (N_18847,N_12828,N_13744);
xnor U18848 (N_18848,N_13537,N_13148);
or U18849 (N_18849,N_12561,N_15887);
and U18850 (N_18850,N_13392,N_15097);
nand U18851 (N_18851,N_14840,N_15872);
nor U18852 (N_18852,N_15506,N_13167);
xnor U18853 (N_18853,N_15500,N_15892);
nand U18854 (N_18854,N_12953,N_14482);
and U18855 (N_18855,N_14693,N_13310);
nor U18856 (N_18856,N_12944,N_15422);
or U18857 (N_18857,N_12453,N_15399);
or U18858 (N_18858,N_14546,N_14934);
nand U18859 (N_18859,N_13149,N_14001);
and U18860 (N_18860,N_12194,N_12851);
nor U18861 (N_18861,N_12045,N_13410);
and U18862 (N_18862,N_12018,N_12493);
nor U18863 (N_18863,N_15390,N_12318);
or U18864 (N_18864,N_14789,N_15652);
or U18865 (N_18865,N_13750,N_13560);
or U18866 (N_18866,N_15431,N_15778);
nand U18867 (N_18867,N_12766,N_13874);
nand U18868 (N_18868,N_15811,N_15025);
nor U18869 (N_18869,N_12541,N_15936);
or U18870 (N_18870,N_12030,N_12516);
nand U18871 (N_18871,N_15033,N_14023);
and U18872 (N_18872,N_12815,N_15994);
or U18873 (N_18873,N_14384,N_12688);
nand U18874 (N_18874,N_14478,N_14210);
nor U18875 (N_18875,N_12708,N_15704);
and U18876 (N_18876,N_15382,N_13944);
nor U18877 (N_18877,N_13128,N_14187);
or U18878 (N_18878,N_13955,N_14592);
and U18879 (N_18879,N_15975,N_15059);
or U18880 (N_18880,N_12291,N_14060);
xor U18881 (N_18881,N_13976,N_14998);
nand U18882 (N_18882,N_13396,N_12513);
nor U18883 (N_18883,N_15984,N_12898);
or U18884 (N_18884,N_12265,N_14112);
xnor U18885 (N_18885,N_12373,N_12892);
xor U18886 (N_18886,N_12434,N_12107);
or U18887 (N_18887,N_14065,N_13150);
and U18888 (N_18888,N_14952,N_12194);
and U18889 (N_18889,N_14215,N_12774);
and U18890 (N_18890,N_14978,N_15714);
nand U18891 (N_18891,N_15396,N_14309);
xor U18892 (N_18892,N_14068,N_14874);
nand U18893 (N_18893,N_14595,N_13974);
or U18894 (N_18894,N_13791,N_12974);
xnor U18895 (N_18895,N_13422,N_15270);
or U18896 (N_18896,N_15555,N_15497);
nand U18897 (N_18897,N_13924,N_14493);
nand U18898 (N_18898,N_12474,N_14260);
or U18899 (N_18899,N_13376,N_15807);
nand U18900 (N_18900,N_13698,N_13058);
nor U18901 (N_18901,N_15565,N_13311);
nor U18902 (N_18902,N_15736,N_13823);
or U18903 (N_18903,N_12346,N_13579);
and U18904 (N_18904,N_15792,N_12645);
or U18905 (N_18905,N_12602,N_13516);
or U18906 (N_18906,N_15178,N_12092);
nand U18907 (N_18907,N_12123,N_12335);
and U18908 (N_18908,N_12196,N_15186);
nor U18909 (N_18909,N_13265,N_12245);
or U18910 (N_18910,N_12811,N_15563);
and U18911 (N_18911,N_14949,N_14871);
nand U18912 (N_18912,N_14196,N_13872);
or U18913 (N_18913,N_12883,N_14545);
or U18914 (N_18914,N_15779,N_12697);
nand U18915 (N_18915,N_14441,N_15097);
nand U18916 (N_18916,N_12326,N_15571);
nand U18917 (N_18917,N_15921,N_12666);
xnor U18918 (N_18918,N_15624,N_15696);
nor U18919 (N_18919,N_14602,N_15149);
or U18920 (N_18920,N_13155,N_14304);
or U18921 (N_18921,N_12934,N_14929);
or U18922 (N_18922,N_15733,N_15056);
nand U18923 (N_18923,N_12378,N_12269);
nand U18924 (N_18924,N_15628,N_14990);
nor U18925 (N_18925,N_12143,N_12541);
nand U18926 (N_18926,N_12711,N_15539);
nor U18927 (N_18927,N_12205,N_14474);
or U18928 (N_18928,N_15594,N_13784);
xor U18929 (N_18929,N_14274,N_12410);
nor U18930 (N_18930,N_15782,N_12597);
or U18931 (N_18931,N_15901,N_13951);
nor U18932 (N_18932,N_14060,N_13997);
nand U18933 (N_18933,N_13663,N_13026);
nand U18934 (N_18934,N_15418,N_15538);
and U18935 (N_18935,N_12074,N_13851);
nor U18936 (N_18936,N_14648,N_12833);
and U18937 (N_18937,N_15830,N_15562);
nor U18938 (N_18938,N_12499,N_15369);
nand U18939 (N_18939,N_15396,N_15445);
nor U18940 (N_18940,N_12368,N_14529);
nor U18941 (N_18941,N_15500,N_12972);
xor U18942 (N_18942,N_14835,N_12356);
or U18943 (N_18943,N_12620,N_12566);
nand U18944 (N_18944,N_12411,N_13015);
nand U18945 (N_18945,N_12295,N_12383);
nor U18946 (N_18946,N_12346,N_12215);
nand U18947 (N_18947,N_15644,N_15825);
and U18948 (N_18948,N_12357,N_13615);
and U18949 (N_18949,N_14766,N_15203);
nand U18950 (N_18950,N_12699,N_12018);
xor U18951 (N_18951,N_14190,N_13720);
nor U18952 (N_18952,N_15426,N_14637);
or U18953 (N_18953,N_13266,N_15550);
xnor U18954 (N_18954,N_12554,N_12658);
xor U18955 (N_18955,N_15395,N_12250);
xor U18956 (N_18956,N_12101,N_14970);
nand U18957 (N_18957,N_13926,N_15428);
nor U18958 (N_18958,N_13513,N_15309);
nand U18959 (N_18959,N_13385,N_12867);
or U18960 (N_18960,N_14305,N_15842);
and U18961 (N_18961,N_12690,N_12535);
or U18962 (N_18962,N_13607,N_14109);
xor U18963 (N_18963,N_12198,N_15858);
or U18964 (N_18964,N_14777,N_15748);
and U18965 (N_18965,N_13978,N_14928);
nand U18966 (N_18966,N_14298,N_15227);
nor U18967 (N_18967,N_13683,N_15753);
nand U18968 (N_18968,N_14130,N_12700);
nand U18969 (N_18969,N_14612,N_13295);
or U18970 (N_18970,N_15126,N_15507);
xnor U18971 (N_18971,N_12947,N_12518);
nand U18972 (N_18972,N_15171,N_12894);
and U18973 (N_18973,N_14809,N_13325);
and U18974 (N_18974,N_12446,N_15774);
and U18975 (N_18975,N_13430,N_13484);
and U18976 (N_18976,N_14127,N_12133);
nand U18977 (N_18977,N_13463,N_15290);
nor U18978 (N_18978,N_12076,N_15882);
and U18979 (N_18979,N_15523,N_15623);
nand U18980 (N_18980,N_15895,N_12625);
and U18981 (N_18981,N_12857,N_12442);
and U18982 (N_18982,N_14184,N_13178);
nor U18983 (N_18983,N_13394,N_14573);
or U18984 (N_18984,N_13578,N_13142);
nand U18985 (N_18985,N_13037,N_14909);
nand U18986 (N_18986,N_13817,N_12024);
nor U18987 (N_18987,N_13073,N_14455);
or U18988 (N_18988,N_12175,N_12187);
nor U18989 (N_18989,N_15978,N_15461);
or U18990 (N_18990,N_14097,N_13966);
nand U18991 (N_18991,N_12361,N_15534);
or U18992 (N_18992,N_12223,N_12322);
nor U18993 (N_18993,N_13928,N_13139);
or U18994 (N_18994,N_15293,N_15980);
or U18995 (N_18995,N_12489,N_14402);
and U18996 (N_18996,N_13253,N_13918);
and U18997 (N_18997,N_14038,N_12680);
or U18998 (N_18998,N_14886,N_15322);
or U18999 (N_18999,N_12902,N_12321);
or U19000 (N_19000,N_14263,N_12003);
xnor U19001 (N_19001,N_12439,N_12012);
nor U19002 (N_19002,N_14423,N_14110);
nor U19003 (N_19003,N_14584,N_15630);
nor U19004 (N_19004,N_12833,N_15492);
and U19005 (N_19005,N_13606,N_13651);
or U19006 (N_19006,N_13214,N_12618);
nand U19007 (N_19007,N_12277,N_15317);
or U19008 (N_19008,N_13146,N_13838);
nand U19009 (N_19009,N_15066,N_12276);
nand U19010 (N_19010,N_13027,N_14562);
nor U19011 (N_19011,N_12058,N_13767);
nand U19012 (N_19012,N_12098,N_15212);
nor U19013 (N_19013,N_13027,N_14370);
and U19014 (N_19014,N_12950,N_14574);
and U19015 (N_19015,N_15112,N_14030);
nor U19016 (N_19016,N_15055,N_15038);
or U19017 (N_19017,N_15046,N_14670);
nor U19018 (N_19018,N_14514,N_14110);
nor U19019 (N_19019,N_12739,N_15585);
nor U19020 (N_19020,N_15255,N_14906);
or U19021 (N_19021,N_15194,N_15989);
nand U19022 (N_19022,N_13273,N_15798);
nor U19023 (N_19023,N_13046,N_14334);
and U19024 (N_19024,N_14947,N_12686);
nor U19025 (N_19025,N_12786,N_15950);
nand U19026 (N_19026,N_15891,N_14167);
or U19027 (N_19027,N_15400,N_14703);
and U19028 (N_19028,N_13050,N_13295);
and U19029 (N_19029,N_15087,N_12516);
and U19030 (N_19030,N_15229,N_13835);
nor U19031 (N_19031,N_14188,N_12348);
or U19032 (N_19032,N_14591,N_13488);
and U19033 (N_19033,N_15624,N_12210);
nor U19034 (N_19034,N_14920,N_13255);
or U19035 (N_19035,N_15060,N_12017);
nand U19036 (N_19036,N_12335,N_15936);
and U19037 (N_19037,N_15286,N_13275);
nor U19038 (N_19038,N_14042,N_15164);
nand U19039 (N_19039,N_13725,N_12572);
and U19040 (N_19040,N_12842,N_14894);
and U19041 (N_19041,N_14871,N_15558);
or U19042 (N_19042,N_13668,N_13004);
nand U19043 (N_19043,N_14896,N_14401);
and U19044 (N_19044,N_14871,N_13017);
and U19045 (N_19045,N_15310,N_12387);
nor U19046 (N_19046,N_14482,N_13723);
nor U19047 (N_19047,N_13635,N_14007);
nor U19048 (N_19048,N_13893,N_15536);
or U19049 (N_19049,N_15327,N_14808);
nand U19050 (N_19050,N_14453,N_12089);
nand U19051 (N_19051,N_15569,N_13302);
and U19052 (N_19052,N_13648,N_13711);
nor U19053 (N_19053,N_12926,N_13968);
and U19054 (N_19054,N_12872,N_13128);
nor U19055 (N_19055,N_13987,N_12988);
or U19056 (N_19056,N_14137,N_14123);
and U19057 (N_19057,N_12300,N_12942);
nand U19058 (N_19058,N_15162,N_13615);
nand U19059 (N_19059,N_12594,N_15505);
and U19060 (N_19060,N_15743,N_13535);
nand U19061 (N_19061,N_14236,N_13038);
or U19062 (N_19062,N_13555,N_13227);
nand U19063 (N_19063,N_12911,N_15873);
nand U19064 (N_19064,N_13761,N_12435);
or U19065 (N_19065,N_14710,N_12083);
nand U19066 (N_19066,N_14595,N_14101);
xnor U19067 (N_19067,N_14766,N_13823);
nor U19068 (N_19068,N_12009,N_14656);
and U19069 (N_19069,N_14921,N_15959);
or U19070 (N_19070,N_14786,N_14122);
or U19071 (N_19071,N_14675,N_15705);
xnor U19072 (N_19072,N_13648,N_13420);
nor U19073 (N_19073,N_14991,N_12033);
and U19074 (N_19074,N_15576,N_15053);
nand U19075 (N_19075,N_12526,N_14227);
and U19076 (N_19076,N_15414,N_15904);
nor U19077 (N_19077,N_12121,N_12128);
and U19078 (N_19078,N_15356,N_15274);
and U19079 (N_19079,N_14119,N_14932);
nor U19080 (N_19080,N_13814,N_12543);
or U19081 (N_19081,N_13331,N_13243);
nor U19082 (N_19082,N_15150,N_12538);
and U19083 (N_19083,N_14629,N_13324);
and U19084 (N_19084,N_12483,N_13108);
nor U19085 (N_19085,N_12292,N_14342);
nand U19086 (N_19086,N_12138,N_14326);
nand U19087 (N_19087,N_14129,N_13902);
xor U19088 (N_19088,N_15808,N_15337);
nand U19089 (N_19089,N_15705,N_12481);
and U19090 (N_19090,N_14180,N_13322);
nand U19091 (N_19091,N_15399,N_15238);
nor U19092 (N_19092,N_14767,N_12096);
nand U19093 (N_19093,N_12687,N_12837);
or U19094 (N_19094,N_14849,N_14670);
and U19095 (N_19095,N_13613,N_14432);
or U19096 (N_19096,N_14478,N_14998);
nand U19097 (N_19097,N_14731,N_13151);
or U19098 (N_19098,N_13027,N_12401);
and U19099 (N_19099,N_12397,N_12853);
nand U19100 (N_19100,N_12776,N_15426);
nand U19101 (N_19101,N_14294,N_14910);
nand U19102 (N_19102,N_12737,N_12823);
and U19103 (N_19103,N_15970,N_15602);
or U19104 (N_19104,N_12197,N_12715);
nor U19105 (N_19105,N_12085,N_13297);
nand U19106 (N_19106,N_13289,N_13535);
nand U19107 (N_19107,N_15051,N_15845);
or U19108 (N_19108,N_14901,N_15258);
or U19109 (N_19109,N_13711,N_14430);
and U19110 (N_19110,N_15021,N_12480);
nor U19111 (N_19111,N_12665,N_14546);
xnor U19112 (N_19112,N_13213,N_13507);
and U19113 (N_19113,N_15826,N_15439);
and U19114 (N_19114,N_12068,N_12880);
or U19115 (N_19115,N_12485,N_15048);
or U19116 (N_19116,N_12995,N_15547);
and U19117 (N_19117,N_14930,N_13434);
or U19118 (N_19118,N_13959,N_15256);
and U19119 (N_19119,N_13904,N_12914);
or U19120 (N_19120,N_14497,N_12678);
nor U19121 (N_19121,N_14704,N_13487);
nor U19122 (N_19122,N_14767,N_14662);
nand U19123 (N_19123,N_13791,N_12964);
nor U19124 (N_19124,N_15874,N_12942);
nand U19125 (N_19125,N_15613,N_13234);
or U19126 (N_19126,N_14224,N_12305);
nand U19127 (N_19127,N_14567,N_13274);
or U19128 (N_19128,N_13590,N_12878);
nand U19129 (N_19129,N_13059,N_14748);
or U19130 (N_19130,N_12797,N_13086);
nand U19131 (N_19131,N_13611,N_14789);
or U19132 (N_19132,N_14984,N_13212);
nor U19133 (N_19133,N_14653,N_15623);
xnor U19134 (N_19134,N_15845,N_13643);
or U19135 (N_19135,N_15543,N_12692);
nor U19136 (N_19136,N_12181,N_15147);
nand U19137 (N_19137,N_12316,N_13810);
or U19138 (N_19138,N_13025,N_14183);
nor U19139 (N_19139,N_15073,N_15775);
nand U19140 (N_19140,N_15992,N_14572);
nand U19141 (N_19141,N_13273,N_12691);
nand U19142 (N_19142,N_15480,N_15170);
and U19143 (N_19143,N_12299,N_15846);
nand U19144 (N_19144,N_14115,N_12963);
xnor U19145 (N_19145,N_12950,N_13742);
or U19146 (N_19146,N_14036,N_14038);
xnor U19147 (N_19147,N_15220,N_13908);
nand U19148 (N_19148,N_15589,N_12087);
xnor U19149 (N_19149,N_13191,N_13474);
or U19150 (N_19150,N_15035,N_14211);
and U19151 (N_19151,N_14245,N_13857);
and U19152 (N_19152,N_14790,N_14069);
nand U19153 (N_19153,N_14338,N_12985);
or U19154 (N_19154,N_13359,N_13955);
nand U19155 (N_19155,N_15174,N_12116);
and U19156 (N_19156,N_14285,N_15864);
xnor U19157 (N_19157,N_13953,N_12896);
nor U19158 (N_19158,N_12913,N_13968);
and U19159 (N_19159,N_14726,N_12670);
or U19160 (N_19160,N_15756,N_12062);
xor U19161 (N_19161,N_13683,N_14459);
and U19162 (N_19162,N_14551,N_12890);
and U19163 (N_19163,N_12442,N_14859);
nand U19164 (N_19164,N_14299,N_15894);
nor U19165 (N_19165,N_14483,N_15770);
nor U19166 (N_19166,N_12568,N_12240);
nand U19167 (N_19167,N_13252,N_13573);
and U19168 (N_19168,N_15141,N_13614);
or U19169 (N_19169,N_14554,N_13381);
nor U19170 (N_19170,N_13811,N_12932);
xor U19171 (N_19171,N_14097,N_14319);
and U19172 (N_19172,N_13496,N_12916);
nor U19173 (N_19173,N_13346,N_13897);
xnor U19174 (N_19174,N_12655,N_15699);
and U19175 (N_19175,N_12963,N_13418);
nand U19176 (N_19176,N_12216,N_14203);
nand U19177 (N_19177,N_13101,N_12341);
and U19178 (N_19178,N_14785,N_12725);
and U19179 (N_19179,N_14228,N_12401);
or U19180 (N_19180,N_14829,N_12460);
and U19181 (N_19181,N_14721,N_12759);
and U19182 (N_19182,N_12425,N_14065);
xnor U19183 (N_19183,N_12969,N_14900);
and U19184 (N_19184,N_13246,N_15555);
xor U19185 (N_19185,N_15067,N_13356);
nor U19186 (N_19186,N_12560,N_13131);
nand U19187 (N_19187,N_15727,N_13029);
nand U19188 (N_19188,N_13535,N_12325);
or U19189 (N_19189,N_12232,N_15682);
and U19190 (N_19190,N_13502,N_15553);
and U19191 (N_19191,N_15249,N_12654);
nor U19192 (N_19192,N_14168,N_15924);
or U19193 (N_19193,N_13256,N_13619);
nand U19194 (N_19194,N_14298,N_14840);
xnor U19195 (N_19195,N_12314,N_12290);
or U19196 (N_19196,N_14444,N_14947);
nor U19197 (N_19197,N_14896,N_13935);
nor U19198 (N_19198,N_15499,N_14238);
and U19199 (N_19199,N_14510,N_12880);
or U19200 (N_19200,N_15570,N_13221);
nand U19201 (N_19201,N_15068,N_13293);
xor U19202 (N_19202,N_15768,N_15678);
nor U19203 (N_19203,N_15095,N_14298);
or U19204 (N_19204,N_12235,N_13989);
and U19205 (N_19205,N_12380,N_15933);
and U19206 (N_19206,N_12817,N_15917);
or U19207 (N_19207,N_15443,N_13117);
nor U19208 (N_19208,N_13668,N_14819);
nor U19209 (N_19209,N_13264,N_14343);
nand U19210 (N_19210,N_13647,N_12121);
nor U19211 (N_19211,N_15519,N_14741);
and U19212 (N_19212,N_12120,N_12425);
nor U19213 (N_19213,N_14809,N_15921);
and U19214 (N_19214,N_13458,N_12422);
and U19215 (N_19215,N_15036,N_13043);
or U19216 (N_19216,N_12345,N_12304);
or U19217 (N_19217,N_13243,N_12679);
nand U19218 (N_19218,N_12345,N_13180);
xnor U19219 (N_19219,N_12074,N_15909);
nand U19220 (N_19220,N_15049,N_14797);
and U19221 (N_19221,N_13761,N_15898);
and U19222 (N_19222,N_14581,N_15915);
and U19223 (N_19223,N_14139,N_15678);
xnor U19224 (N_19224,N_12804,N_12916);
nor U19225 (N_19225,N_15871,N_12411);
xnor U19226 (N_19226,N_15545,N_12897);
xnor U19227 (N_19227,N_14486,N_15592);
and U19228 (N_19228,N_14178,N_14524);
and U19229 (N_19229,N_14270,N_15614);
nand U19230 (N_19230,N_15844,N_15805);
nand U19231 (N_19231,N_15961,N_15200);
nor U19232 (N_19232,N_12602,N_15065);
nor U19233 (N_19233,N_13996,N_15345);
nand U19234 (N_19234,N_12426,N_12092);
or U19235 (N_19235,N_13446,N_13839);
nor U19236 (N_19236,N_13070,N_13934);
nor U19237 (N_19237,N_13228,N_15849);
nand U19238 (N_19238,N_13156,N_13519);
nor U19239 (N_19239,N_12693,N_13554);
nand U19240 (N_19240,N_14902,N_13299);
and U19241 (N_19241,N_12353,N_13335);
or U19242 (N_19242,N_13408,N_12467);
nand U19243 (N_19243,N_15440,N_15163);
and U19244 (N_19244,N_13721,N_15018);
nor U19245 (N_19245,N_12572,N_12275);
and U19246 (N_19246,N_14845,N_14160);
nor U19247 (N_19247,N_15664,N_14689);
nor U19248 (N_19248,N_14113,N_13981);
or U19249 (N_19249,N_15710,N_14317);
nand U19250 (N_19250,N_13902,N_15525);
nor U19251 (N_19251,N_15894,N_14873);
nand U19252 (N_19252,N_13862,N_15285);
nand U19253 (N_19253,N_13244,N_13401);
and U19254 (N_19254,N_15280,N_13049);
and U19255 (N_19255,N_12343,N_14583);
or U19256 (N_19256,N_14426,N_13927);
xor U19257 (N_19257,N_14051,N_14156);
nand U19258 (N_19258,N_15170,N_15983);
or U19259 (N_19259,N_14479,N_15537);
and U19260 (N_19260,N_13909,N_14424);
and U19261 (N_19261,N_15567,N_14612);
or U19262 (N_19262,N_14170,N_13193);
nor U19263 (N_19263,N_15733,N_13565);
nor U19264 (N_19264,N_12779,N_15618);
xor U19265 (N_19265,N_13538,N_14119);
and U19266 (N_19266,N_14256,N_14282);
nor U19267 (N_19267,N_13055,N_13999);
and U19268 (N_19268,N_14030,N_15152);
or U19269 (N_19269,N_12449,N_12069);
nor U19270 (N_19270,N_14127,N_13451);
nand U19271 (N_19271,N_13273,N_14176);
nand U19272 (N_19272,N_14467,N_15650);
xor U19273 (N_19273,N_13873,N_12050);
xor U19274 (N_19274,N_15345,N_12144);
nor U19275 (N_19275,N_14089,N_12455);
nand U19276 (N_19276,N_14914,N_12876);
nand U19277 (N_19277,N_12845,N_13803);
nand U19278 (N_19278,N_15196,N_15237);
or U19279 (N_19279,N_13920,N_13359);
or U19280 (N_19280,N_13022,N_13093);
nor U19281 (N_19281,N_13502,N_14993);
nor U19282 (N_19282,N_13225,N_14258);
or U19283 (N_19283,N_14500,N_14891);
nor U19284 (N_19284,N_14144,N_13413);
or U19285 (N_19285,N_15253,N_14209);
and U19286 (N_19286,N_13291,N_12756);
and U19287 (N_19287,N_12389,N_12732);
or U19288 (N_19288,N_15590,N_14916);
or U19289 (N_19289,N_15629,N_14703);
nor U19290 (N_19290,N_14805,N_13708);
and U19291 (N_19291,N_12649,N_13155);
nor U19292 (N_19292,N_12218,N_12607);
nor U19293 (N_19293,N_13281,N_14498);
and U19294 (N_19294,N_13547,N_14456);
and U19295 (N_19295,N_12904,N_14666);
and U19296 (N_19296,N_15792,N_15224);
or U19297 (N_19297,N_13996,N_12030);
nor U19298 (N_19298,N_12548,N_14685);
and U19299 (N_19299,N_12029,N_15337);
and U19300 (N_19300,N_12956,N_15839);
nand U19301 (N_19301,N_12698,N_12704);
and U19302 (N_19302,N_12193,N_15716);
nor U19303 (N_19303,N_13948,N_15857);
nor U19304 (N_19304,N_15564,N_12831);
xnor U19305 (N_19305,N_15224,N_15773);
or U19306 (N_19306,N_12974,N_13324);
or U19307 (N_19307,N_15476,N_14366);
or U19308 (N_19308,N_14403,N_14652);
nand U19309 (N_19309,N_14878,N_14729);
and U19310 (N_19310,N_14923,N_13641);
or U19311 (N_19311,N_12788,N_13415);
or U19312 (N_19312,N_13957,N_13264);
and U19313 (N_19313,N_13977,N_12420);
or U19314 (N_19314,N_12272,N_12496);
nand U19315 (N_19315,N_14259,N_12587);
and U19316 (N_19316,N_14924,N_14682);
and U19317 (N_19317,N_13136,N_14729);
nor U19318 (N_19318,N_13845,N_14043);
and U19319 (N_19319,N_12880,N_15714);
and U19320 (N_19320,N_12445,N_14639);
xnor U19321 (N_19321,N_14962,N_14512);
or U19322 (N_19322,N_14224,N_15759);
nor U19323 (N_19323,N_12947,N_13996);
nor U19324 (N_19324,N_12859,N_12278);
and U19325 (N_19325,N_12680,N_13686);
nand U19326 (N_19326,N_13904,N_14784);
nand U19327 (N_19327,N_15607,N_14458);
nor U19328 (N_19328,N_13662,N_15012);
nand U19329 (N_19329,N_13492,N_15956);
and U19330 (N_19330,N_15075,N_12982);
nand U19331 (N_19331,N_13616,N_14385);
or U19332 (N_19332,N_12970,N_14498);
or U19333 (N_19333,N_14514,N_12853);
nor U19334 (N_19334,N_12938,N_13633);
nor U19335 (N_19335,N_14127,N_15151);
nor U19336 (N_19336,N_13062,N_14653);
nor U19337 (N_19337,N_15647,N_13029);
nor U19338 (N_19338,N_14469,N_15507);
nor U19339 (N_19339,N_15352,N_14121);
nor U19340 (N_19340,N_12365,N_15318);
nor U19341 (N_19341,N_14729,N_13767);
or U19342 (N_19342,N_12308,N_13357);
nand U19343 (N_19343,N_15922,N_14754);
nor U19344 (N_19344,N_13108,N_14537);
nor U19345 (N_19345,N_15980,N_13300);
and U19346 (N_19346,N_13216,N_13600);
nor U19347 (N_19347,N_12810,N_15144);
nor U19348 (N_19348,N_15680,N_13012);
nand U19349 (N_19349,N_15086,N_14791);
nor U19350 (N_19350,N_12094,N_15983);
nor U19351 (N_19351,N_12319,N_12642);
nand U19352 (N_19352,N_13081,N_14017);
nor U19353 (N_19353,N_12214,N_12889);
nor U19354 (N_19354,N_15485,N_15814);
nand U19355 (N_19355,N_14488,N_13228);
nor U19356 (N_19356,N_13451,N_13799);
or U19357 (N_19357,N_14150,N_13869);
and U19358 (N_19358,N_15676,N_13087);
nor U19359 (N_19359,N_12143,N_13828);
xnor U19360 (N_19360,N_14019,N_13746);
and U19361 (N_19361,N_14763,N_13415);
xor U19362 (N_19362,N_15372,N_15053);
and U19363 (N_19363,N_12790,N_13302);
or U19364 (N_19364,N_12627,N_15274);
nor U19365 (N_19365,N_12881,N_14522);
nor U19366 (N_19366,N_14112,N_15861);
and U19367 (N_19367,N_14557,N_15807);
nand U19368 (N_19368,N_15778,N_13283);
and U19369 (N_19369,N_14344,N_14465);
nand U19370 (N_19370,N_14996,N_15938);
xor U19371 (N_19371,N_14157,N_12913);
or U19372 (N_19372,N_14848,N_13921);
nor U19373 (N_19373,N_14251,N_14872);
nand U19374 (N_19374,N_15372,N_15593);
nand U19375 (N_19375,N_12283,N_15760);
or U19376 (N_19376,N_14755,N_15103);
or U19377 (N_19377,N_15061,N_12331);
nand U19378 (N_19378,N_12935,N_14602);
nand U19379 (N_19379,N_15364,N_13499);
nor U19380 (N_19380,N_15802,N_13526);
or U19381 (N_19381,N_15389,N_12470);
xor U19382 (N_19382,N_12123,N_12361);
or U19383 (N_19383,N_12441,N_12933);
or U19384 (N_19384,N_12957,N_15895);
nor U19385 (N_19385,N_12477,N_12828);
or U19386 (N_19386,N_12232,N_12446);
nor U19387 (N_19387,N_13943,N_15904);
xor U19388 (N_19388,N_15038,N_14760);
or U19389 (N_19389,N_12177,N_13402);
nor U19390 (N_19390,N_12854,N_13379);
nor U19391 (N_19391,N_12118,N_14362);
and U19392 (N_19392,N_15330,N_14635);
nand U19393 (N_19393,N_13227,N_13063);
and U19394 (N_19394,N_14511,N_14393);
and U19395 (N_19395,N_14004,N_12889);
and U19396 (N_19396,N_13266,N_13344);
and U19397 (N_19397,N_13992,N_15215);
xnor U19398 (N_19398,N_12293,N_12307);
or U19399 (N_19399,N_14134,N_14953);
nand U19400 (N_19400,N_12934,N_13385);
nand U19401 (N_19401,N_15309,N_14666);
xnor U19402 (N_19402,N_14211,N_12437);
or U19403 (N_19403,N_15846,N_13681);
or U19404 (N_19404,N_15793,N_14724);
nor U19405 (N_19405,N_13710,N_15050);
nand U19406 (N_19406,N_15314,N_14666);
nor U19407 (N_19407,N_12362,N_14787);
nor U19408 (N_19408,N_15360,N_13805);
or U19409 (N_19409,N_15403,N_13188);
nand U19410 (N_19410,N_14325,N_13164);
or U19411 (N_19411,N_13048,N_14632);
and U19412 (N_19412,N_14301,N_12986);
nor U19413 (N_19413,N_13324,N_12800);
nand U19414 (N_19414,N_14329,N_14437);
and U19415 (N_19415,N_14190,N_15495);
or U19416 (N_19416,N_12849,N_13956);
nor U19417 (N_19417,N_13355,N_13726);
nor U19418 (N_19418,N_15646,N_13133);
or U19419 (N_19419,N_14643,N_12223);
nand U19420 (N_19420,N_15317,N_13946);
nand U19421 (N_19421,N_15605,N_12366);
nor U19422 (N_19422,N_14784,N_13759);
and U19423 (N_19423,N_13339,N_14950);
or U19424 (N_19424,N_15325,N_13956);
and U19425 (N_19425,N_15611,N_14149);
nand U19426 (N_19426,N_13653,N_14002);
nand U19427 (N_19427,N_14166,N_13300);
and U19428 (N_19428,N_13297,N_14084);
nor U19429 (N_19429,N_14848,N_12090);
nor U19430 (N_19430,N_15062,N_14724);
or U19431 (N_19431,N_14019,N_14403);
or U19432 (N_19432,N_12060,N_13059);
and U19433 (N_19433,N_14420,N_13281);
nor U19434 (N_19434,N_13394,N_15841);
nor U19435 (N_19435,N_14180,N_13007);
or U19436 (N_19436,N_13000,N_15566);
nor U19437 (N_19437,N_13337,N_12697);
or U19438 (N_19438,N_13480,N_14418);
and U19439 (N_19439,N_13804,N_13648);
or U19440 (N_19440,N_13742,N_15920);
and U19441 (N_19441,N_15592,N_12070);
nand U19442 (N_19442,N_14089,N_14099);
or U19443 (N_19443,N_14483,N_13019);
and U19444 (N_19444,N_12931,N_12211);
xor U19445 (N_19445,N_12237,N_13038);
or U19446 (N_19446,N_14226,N_15202);
xnor U19447 (N_19447,N_12185,N_12565);
nor U19448 (N_19448,N_13296,N_13035);
or U19449 (N_19449,N_13211,N_12656);
xnor U19450 (N_19450,N_13605,N_15933);
nand U19451 (N_19451,N_12835,N_14017);
or U19452 (N_19452,N_15455,N_15433);
nand U19453 (N_19453,N_15711,N_15284);
and U19454 (N_19454,N_13615,N_15664);
nor U19455 (N_19455,N_14743,N_14856);
or U19456 (N_19456,N_15611,N_14495);
and U19457 (N_19457,N_15457,N_13884);
xnor U19458 (N_19458,N_15338,N_13737);
nor U19459 (N_19459,N_13779,N_14463);
and U19460 (N_19460,N_13979,N_14945);
or U19461 (N_19461,N_15374,N_14552);
and U19462 (N_19462,N_15858,N_15019);
nor U19463 (N_19463,N_12139,N_12089);
or U19464 (N_19464,N_13612,N_13240);
and U19465 (N_19465,N_13294,N_13180);
or U19466 (N_19466,N_14360,N_14363);
and U19467 (N_19467,N_12199,N_15887);
or U19468 (N_19468,N_15139,N_14919);
and U19469 (N_19469,N_15734,N_12597);
or U19470 (N_19470,N_12322,N_13704);
xnor U19471 (N_19471,N_12726,N_14851);
and U19472 (N_19472,N_14370,N_15522);
nor U19473 (N_19473,N_14450,N_14114);
or U19474 (N_19474,N_14514,N_14485);
nand U19475 (N_19475,N_15221,N_15768);
and U19476 (N_19476,N_13302,N_15272);
and U19477 (N_19477,N_12869,N_14163);
nand U19478 (N_19478,N_15673,N_14777);
or U19479 (N_19479,N_14703,N_14726);
nor U19480 (N_19480,N_13858,N_13895);
nor U19481 (N_19481,N_13519,N_12264);
nor U19482 (N_19482,N_12112,N_14929);
and U19483 (N_19483,N_13408,N_12735);
or U19484 (N_19484,N_14239,N_14468);
nor U19485 (N_19485,N_12544,N_14086);
nor U19486 (N_19486,N_15112,N_13582);
nand U19487 (N_19487,N_12006,N_15705);
nor U19488 (N_19488,N_15565,N_14316);
or U19489 (N_19489,N_13911,N_12570);
or U19490 (N_19490,N_12955,N_12193);
nor U19491 (N_19491,N_12713,N_14395);
and U19492 (N_19492,N_14241,N_15313);
nand U19493 (N_19493,N_15804,N_14678);
nor U19494 (N_19494,N_14928,N_12860);
nor U19495 (N_19495,N_15661,N_13138);
nor U19496 (N_19496,N_13576,N_13388);
nand U19497 (N_19497,N_14911,N_13126);
nand U19498 (N_19498,N_12513,N_13284);
nand U19499 (N_19499,N_14878,N_13192);
or U19500 (N_19500,N_13864,N_14571);
nand U19501 (N_19501,N_15274,N_15115);
nand U19502 (N_19502,N_15259,N_13269);
nor U19503 (N_19503,N_12611,N_15648);
nand U19504 (N_19504,N_12675,N_12740);
or U19505 (N_19505,N_12004,N_12843);
or U19506 (N_19506,N_12706,N_12339);
or U19507 (N_19507,N_13092,N_14965);
nor U19508 (N_19508,N_14716,N_15889);
or U19509 (N_19509,N_13320,N_14517);
nor U19510 (N_19510,N_14869,N_15029);
or U19511 (N_19511,N_14311,N_15263);
and U19512 (N_19512,N_12990,N_14190);
and U19513 (N_19513,N_13365,N_13456);
nand U19514 (N_19514,N_15382,N_13789);
nor U19515 (N_19515,N_14199,N_13931);
nand U19516 (N_19516,N_15840,N_14938);
and U19517 (N_19517,N_12448,N_14038);
nand U19518 (N_19518,N_12219,N_12809);
and U19519 (N_19519,N_13965,N_15961);
and U19520 (N_19520,N_15442,N_12293);
nand U19521 (N_19521,N_13384,N_13572);
nor U19522 (N_19522,N_13422,N_15659);
or U19523 (N_19523,N_12899,N_12254);
nand U19524 (N_19524,N_13571,N_13765);
or U19525 (N_19525,N_15102,N_15421);
and U19526 (N_19526,N_13947,N_13999);
and U19527 (N_19527,N_15646,N_15358);
nor U19528 (N_19528,N_15479,N_12183);
and U19529 (N_19529,N_15299,N_13294);
nor U19530 (N_19530,N_15967,N_15946);
or U19531 (N_19531,N_14777,N_15747);
nor U19532 (N_19532,N_15094,N_15734);
and U19533 (N_19533,N_13716,N_12382);
nor U19534 (N_19534,N_14745,N_15097);
or U19535 (N_19535,N_12359,N_14117);
xnor U19536 (N_19536,N_14086,N_12733);
nand U19537 (N_19537,N_15225,N_13442);
nor U19538 (N_19538,N_13654,N_13111);
or U19539 (N_19539,N_13223,N_14554);
nor U19540 (N_19540,N_12742,N_15471);
nor U19541 (N_19541,N_13335,N_12666);
xor U19542 (N_19542,N_15174,N_12899);
xor U19543 (N_19543,N_14495,N_14828);
nor U19544 (N_19544,N_14473,N_12618);
and U19545 (N_19545,N_14022,N_15089);
or U19546 (N_19546,N_15232,N_12528);
xor U19547 (N_19547,N_13407,N_12157);
nor U19548 (N_19548,N_14077,N_15380);
xor U19549 (N_19549,N_13684,N_14698);
nor U19550 (N_19550,N_13448,N_15062);
and U19551 (N_19551,N_15599,N_15626);
and U19552 (N_19552,N_12893,N_12129);
or U19553 (N_19553,N_12752,N_14304);
nand U19554 (N_19554,N_15362,N_14176);
nand U19555 (N_19555,N_15669,N_13672);
nand U19556 (N_19556,N_13283,N_14447);
and U19557 (N_19557,N_13279,N_14878);
nand U19558 (N_19558,N_14357,N_15528);
nor U19559 (N_19559,N_13159,N_15811);
or U19560 (N_19560,N_14098,N_13425);
xnor U19561 (N_19561,N_15065,N_14365);
and U19562 (N_19562,N_15202,N_13905);
nand U19563 (N_19563,N_14419,N_12058);
nand U19564 (N_19564,N_12450,N_13629);
and U19565 (N_19565,N_14324,N_15372);
nor U19566 (N_19566,N_13691,N_12032);
nor U19567 (N_19567,N_13724,N_14683);
xor U19568 (N_19568,N_14895,N_15274);
nand U19569 (N_19569,N_14277,N_13274);
nor U19570 (N_19570,N_14125,N_14583);
or U19571 (N_19571,N_12281,N_12978);
nor U19572 (N_19572,N_15352,N_13809);
nand U19573 (N_19573,N_14229,N_12641);
nand U19574 (N_19574,N_14050,N_15611);
and U19575 (N_19575,N_14270,N_13660);
and U19576 (N_19576,N_14573,N_14504);
nand U19577 (N_19577,N_13884,N_15430);
or U19578 (N_19578,N_15360,N_13845);
or U19579 (N_19579,N_13950,N_12113);
or U19580 (N_19580,N_13206,N_13483);
or U19581 (N_19581,N_12363,N_13717);
nor U19582 (N_19582,N_15559,N_13416);
nand U19583 (N_19583,N_15113,N_13236);
or U19584 (N_19584,N_14754,N_12963);
and U19585 (N_19585,N_15460,N_13364);
nor U19586 (N_19586,N_14021,N_12811);
nand U19587 (N_19587,N_13520,N_13845);
nand U19588 (N_19588,N_12727,N_12295);
or U19589 (N_19589,N_15322,N_15684);
or U19590 (N_19590,N_15474,N_15079);
nor U19591 (N_19591,N_13326,N_15562);
nor U19592 (N_19592,N_13716,N_15348);
xnor U19593 (N_19593,N_15690,N_13327);
nand U19594 (N_19594,N_14233,N_15543);
nand U19595 (N_19595,N_12087,N_15149);
nand U19596 (N_19596,N_13638,N_14040);
nor U19597 (N_19597,N_14276,N_15031);
or U19598 (N_19598,N_14449,N_15023);
nand U19599 (N_19599,N_14672,N_14489);
and U19600 (N_19600,N_14767,N_15103);
or U19601 (N_19601,N_14192,N_12211);
nor U19602 (N_19602,N_12071,N_15837);
and U19603 (N_19603,N_14140,N_13698);
or U19604 (N_19604,N_14334,N_13698);
and U19605 (N_19605,N_13895,N_15664);
or U19606 (N_19606,N_15237,N_12304);
nor U19607 (N_19607,N_13510,N_14195);
or U19608 (N_19608,N_12161,N_14416);
nor U19609 (N_19609,N_15201,N_14019);
nand U19610 (N_19610,N_13333,N_14352);
or U19611 (N_19611,N_15261,N_12272);
and U19612 (N_19612,N_14735,N_15796);
or U19613 (N_19613,N_12112,N_13046);
or U19614 (N_19614,N_12553,N_12557);
xnor U19615 (N_19615,N_13891,N_14961);
and U19616 (N_19616,N_12711,N_13901);
nor U19617 (N_19617,N_13938,N_15668);
and U19618 (N_19618,N_12356,N_15169);
nand U19619 (N_19619,N_14615,N_15598);
xor U19620 (N_19620,N_14443,N_13489);
nand U19621 (N_19621,N_15478,N_13728);
nand U19622 (N_19622,N_14287,N_13965);
xor U19623 (N_19623,N_14752,N_13202);
or U19624 (N_19624,N_15579,N_14527);
nand U19625 (N_19625,N_12056,N_12124);
nor U19626 (N_19626,N_14649,N_14751);
or U19627 (N_19627,N_15350,N_13388);
or U19628 (N_19628,N_12414,N_13333);
nor U19629 (N_19629,N_15576,N_14523);
or U19630 (N_19630,N_14360,N_14370);
xor U19631 (N_19631,N_15123,N_15763);
nand U19632 (N_19632,N_13469,N_13074);
or U19633 (N_19633,N_15368,N_14846);
and U19634 (N_19634,N_12034,N_14551);
nand U19635 (N_19635,N_14629,N_15938);
nand U19636 (N_19636,N_15848,N_12225);
nor U19637 (N_19637,N_14142,N_14483);
and U19638 (N_19638,N_15289,N_15767);
and U19639 (N_19639,N_13223,N_14221);
nand U19640 (N_19640,N_15830,N_13466);
nand U19641 (N_19641,N_15775,N_12875);
nand U19642 (N_19642,N_14808,N_12638);
nor U19643 (N_19643,N_13484,N_14238);
or U19644 (N_19644,N_12138,N_13263);
nand U19645 (N_19645,N_14587,N_14869);
nand U19646 (N_19646,N_15525,N_15653);
nor U19647 (N_19647,N_15604,N_13299);
or U19648 (N_19648,N_13519,N_12804);
nand U19649 (N_19649,N_13767,N_12710);
and U19650 (N_19650,N_15020,N_15082);
nor U19651 (N_19651,N_15303,N_12099);
or U19652 (N_19652,N_15484,N_15148);
or U19653 (N_19653,N_14399,N_15784);
and U19654 (N_19654,N_15847,N_12304);
nand U19655 (N_19655,N_13704,N_12620);
and U19656 (N_19656,N_12940,N_15393);
nor U19657 (N_19657,N_15049,N_12724);
and U19658 (N_19658,N_13819,N_15460);
and U19659 (N_19659,N_14498,N_14549);
and U19660 (N_19660,N_13443,N_15386);
and U19661 (N_19661,N_15971,N_12549);
nor U19662 (N_19662,N_13216,N_13368);
xor U19663 (N_19663,N_14339,N_15652);
and U19664 (N_19664,N_14206,N_12266);
or U19665 (N_19665,N_13895,N_12784);
and U19666 (N_19666,N_13531,N_15933);
nor U19667 (N_19667,N_12658,N_12532);
or U19668 (N_19668,N_13312,N_12737);
or U19669 (N_19669,N_12407,N_13814);
or U19670 (N_19670,N_12297,N_13235);
or U19671 (N_19671,N_15248,N_12284);
and U19672 (N_19672,N_13402,N_13778);
nand U19673 (N_19673,N_15380,N_12339);
or U19674 (N_19674,N_15878,N_15289);
and U19675 (N_19675,N_14310,N_14812);
xnor U19676 (N_19676,N_12826,N_12829);
and U19677 (N_19677,N_15000,N_15155);
and U19678 (N_19678,N_14142,N_13244);
and U19679 (N_19679,N_15527,N_12669);
nand U19680 (N_19680,N_14479,N_13974);
or U19681 (N_19681,N_12867,N_15516);
or U19682 (N_19682,N_12610,N_13313);
and U19683 (N_19683,N_14468,N_13058);
and U19684 (N_19684,N_14846,N_13753);
or U19685 (N_19685,N_14932,N_14662);
nand U19686 (N_19686,N_13092,N_15311);
nand U19687 (N_19687,N_14448,N_12653);
and U19688 (N_19688,N_12593,N_12799);
or U19689 (N_19689,N_14569,N_13226);
nand U19690 (N_19690,N_14833,N_13007);
nor U19691 (N_19691,N_14865,N_12576);
or U19692 (N_19692,N_13605,N_14752);
or U19693 (N_19693,N_15869,N_14663);
or U19694 (N_19694,N_14024,N_13975);
and U19695 (N_19695,N_12839,N_12721);
nor U19696 (N_19696,N_13208,N_13361);
and U19697 (N_19697,N_12586,N_12260);
nor U19698 (N_19698,N_15681,N_13764);
or U19699 (N_19699,N_15297,N_14345);
nor U19700 (N_19700,N_15666,N_12459);
nand U19701 (N_19701,N_13774,N_13599);
and U19702 (N_19702,N_12086,N_15797);
xor U19703 (N_19703,N_12785,N_12334);
and U19704 (N_19704,N_15539,N_12826);
nand U19705 (N_19705,N_13583,N_14140);
or U19706 (N_19706,N_14018,N_15522);
nand U19707 (N_19707,N_13332,N_15754);
xnor U19708 (N_19708,N_12681,N_15605);
or U19709 (N_19709,N_13110,N_15411);
nor U19710 (N_19710,N_13459,N_12699);
nand U19711 (N_19711,N_14216,N_12720);
nor U19712 (N_19712,N_15871,N_15207);
nand U19713 (N_19713,N_14333,N_13065);
xor U19714 (N_19714,N_12435,N_13467);
nor U19715 (N_19715,N_13111,N_15226);
nand U19716 (N_19716,N_14212,N_12847);
nand U19717 (N_19717,N_14262,N_14271);
and U19718 (N_19718,N_12222,N_15108);
nand U19719 (N_19719,N_15826,N_12888);
or U19720 (N_19720,N_14630,N_13148);
nor U19721 (N_19721,N_12857,N_15896);
xnor U19722 (N_19722,N_15952,N_15151);
nor U19723 (N_19723,N_15703,N_12359);
xor U19724 (N_19724,N_13032,N_15739);
xor U19725 (N_19725,N_12690,N_15993);
xnor U19726 (N_19726,N_12798,N_12118);
nand U19727 (N_19727,N_12513,N_14038);
nor U19728 (N_19728,N_14109,N_15424);
nor U19729 (N_19729,N_14131,N_13021);
nor U19730 (N_19730,N_15553,N_12978);
nor U19731 (N_19731,N_12660,N_13358);
xnor U19732 (N_19732,N_15870,N_14224);
and U19733 (N_19733,N_12993,N_14313);
xor U19734 (N_19734,N_12702,N_15192);
and U19735 (N_19735,N_12294,N_13250);
and U19736 (N_19736,N_13730,N_15207);
and U19737 (N_19737,N_14007,N_13359);
or U19738 (N_19738,N_12058,N_14124);
and U19739 (N_19739,N_13627,N_15483);
and U19740 (N_19740,N_12050,N_15464);
nand U19741 (N_19741,N_14945,N_14288);
or U19742 (N_19742,N_13264,N_13747);
nor U19743 (N_19743,N_15077,N_15832);
nand U19744 (N_19744,N_12571,N_15798);
nand U19745 (N_19745,N_13389,N_15108);
and U19746 (N_19746,N_13859,N_12633);
and U19747 (N_19747,N_14429,N_15219);
nand U19748 (N_19748,N_13828,N_14699);
nand U19749 (N_19749,N_13009,N_13575);
xor U19750 (N_19750,N_14099,N_13705);
nor U19751 (N_19751,N_12063,N_14926);
nor U19752 (N_19752,N_12564,N_15261);
or U19753 (N_19753,N_15045,N_13870);
or U19754 (N_19754,N_13337,N_12082);
nor U19755 (N_19755,N_13993,N_15558);
nor U19756 (N_19756,N_12399,N_12779);
and U19757 (N_19757,N_12853,N_15237);
nor U19758 (N_19758,N_15402,N_15677);
nor U19759 (N_19759,N_13232,N_12919);
or U19760 (N_19760,N_12487,N_13379);
and U19761 (N_19761,N_14343,N_15161);
nand U19762 (N_19762,N_13952,N_12841);
or U19763 (N_19763,N_14070,N_12244);
and U19764 (N_19764,N_12289,N_13629);
or U19765 (N_19765,N_15852,N_12625);
nor U19766 (N_19766,N_14417,N_13052);
nor U19767 (N_19767,N_15425,N_13985);
xor U19768 (N_19768,N_15294,N_15943);
or U19769 (N_19769,N_13525,N_14486);
and U19770 (N_19770,N_13671,N_15274);
and U19771 (N_19771,N_12282,N_14819);
nand U19772 (N_19772,N_14031,N_12286);
nand U19773 (N_19773,N_13544,N_15775);
nand U19774 (N_19774,N_13452,N_12005);
or U19775 (N_19775,N_14126,N_13173);
nand U19776 (N_19776,N_14581,N_14738);
and U19777 (N_19777,N_12943,N_15126);
nor U19778 (N_19778,N_15153,N_14232);
nor U19779 (N_19779,N_12470,N_13673);
and U19780 (N_19780,N_13755,N_14952);
or U19781 (N_19781,N_13165,N_12749);
xor U19782 (N_19782,N_15296,N_12508);
nor U19783 (N_19783,N_14983,N_13994);
or U19784 (N_19784,N_12503,N_13856);
or U19785 (N_19785,N_13503,N_13222);
or U19786 (N_19786,N_15765,N_12500);
xnor U19787 (N_19787,N_15082,N_12464);
nand U19788 (N_19788,N_13037,N_12800);
nor U19789 (N_19789,N_12306,N_15912);
xnor U19790 (N_19790,N_15206,N_15782);
or U19791 (N_19791,N_13337,N_12536);
xor U19792 (N_19792,N_15243,N_14888);
and U19793 (N_19793,N_14968,N_12513);
or U19794 (N_19794,N_14553,N_13419);
or U19795 (N_19795,N_15454,N_13297);
and U19796 (N_19796,N_15768,N_12725);
nand U19797 (N_19797,N_13674,N_12826);
nand U19798 (N_19798,N_12708,N_13893);
nand U19799 (N_19799,N_12190,N_12653);
nand U19800 (N_19800,N_12355,N_12668);
or U19801 (N_19801,N_12799,N_12035);
or U19802 (N_19802,N_15346,N_13502);
and U19803 (N_19803,N_14500,N_14246);
nand U19804 (N_19804,N_14457,N_12599);
nand U19805 (N_19805,N_12483,N_14154);
nand U19806 (N_19806,N_14910,N_15822);
and U19807 (N_19807,N_14105,N_14721);
nand U19808 (N_19808,N_13822,N_15461);
and U19809 (N_19809,N_14182,N_15353);
and U19810 (N_19810,N_14223,N_14387);
nor U19811 (N_19811,N_13572,N_13700);
nor U19812 (N_19812,N_15999,N_15799);
or U19813 (N_19813,N_12400,N_14778);
nor U19814 (N_19814,N_14327,N_15475);
or U19815 (N_19815,N_14079,N_13742);
and U19816 (N_19816,N_15399,N_12508);
nor U19817 (N_19817,N_15248,N_15753);
nor U19818 (N_19818,N_12118,N_15394);
and U19819 (N_19819,N_14143,N_14845);
nor U19820 (N_19820,N_12022,N_12850);
or U19821 (N_19821,N_12614,N_14065);
nand U19822 (N_19822,N_12694,N_13465);
xor U19823 (N_19823,N_12178,N_12735);
or U19824 (N_19824,N_15305,N_15581);
or U19825 (N_19825,N_15981,N_13354);
or U19826 (N_19826,N_12682,N_12195);
nor U19827 (N_19827,N_13942,N_15044);
nor U19828 (N_19828,N_14067,N_13252);
nand U19829 (N_19829,N_15106,N_13261);
or U19830 (N_19830,N_13623,N_14495);
and U19831 (N_19831,N_15735,N_12399);
or U19832 (N_19832,N_14569,N_14525);
nor U19833 (N_19833,N_12607,N_14536);
nand U19834 (N_19834,N_12934,N_13537);
and U19835 (N_19835,N_13397,N_12201);
or U19836 (N_19836,N_13992,N_15587);
and U19837 (N_19837,N_13307,N_13473);
or U19838 (N_19838,N_15280,N_13571);
and U19839 (N_19839,N_12111,N_14301);
or U19840 (N_19840,N_12366,N_15354);
and U19841 (N_19841,N_14464,N_15015);
or U19842 (N_19842,N_12981,N_12514);
and U19843 (N_19843,N_12083,N_14950);
nor U19844 (N_19844,N_13357,N_15673);
nor U19845 (N_19845,N_15370,N_14995);
nor U19846 (N_19846,N_13530,N_14119);
or U19847 (N_19847,N_13003,N_13774);
or U19848 (N_19848,N_14648,N_12126);
or U19849 (N_19849,N_15155,N_15272);
xor U19850 (N_19850,N_13680,N_12860);
nand U19851 (N_19851,N_13562,N_14049);
nor U19852 (N_19852,N_12810,N_12135);
or U19853 (N_19853,N_13608,N_14061);
xor U19854 (N_19854,N_15570,N_15422);
nor U19855 (N_19855,N_14793,N_15615);
nor U19856 (N_19856,N_13420,N_12158);
or U19857 (N_19857,N_15933,N_13767);
nor U19858 (N_19858,N_15943,N_14442);
or U19859 (N_19859,N_15001,N_13907);
nand U19860 (N_19860,N_13869,N_12156);
xor U19861 (N_19861,N_15771,N_13724);
nand U19862 (N_19862,N_14280,N_15411);
and U19863 (N_19863,N_12030,N_15280);
xor U19864 (N_19864,N_15770,N_15210);
nand U19865 (N_19865,N_15032,N_12240);
and U19866 (N_19866,N_15630,N_12331);
and U19867 (N_19867,N_14753,N_13674);
and U19868 (N_19868,N_13149,N_13627);
nand U19869 (N_19869,N_13250,N_13074);
nand U19870 (N_19870,N_15506,N_13125);
or U19871 (N_19871,N_14410,N_13806);
nor U19872 (N_19872,N_13680,N_12049);
nand U19873 (N_19873,N_14114,N_15216);
and U19874 (N_19874,N_15415,N_15099);
nand U19875 (N_19875,N_13416,N_14939);
xor U19876 (N_19876,N_13946,N_12263);
nand U19877 (N_19877,N_15558,N_12922);
or U19878 (N_19878,N_14510,N_14663);
or U19879 (N_19879,N_12326,N_14564);
nand U19880 (N_19880,N_14939,N_12681);
or U19881 (N_19881,N_13098,N_15266);
and U19882 (N_19882,N_12601,N_14406);
xor U19883 (N_19883,N_13354,N_15456);
xor U19884 (N_19884,N_14093,N_13394);
nand U19885 (N_19885,N_14921,N_13093);
nand U19886 (N_19886,N_15789,N_15473);
or U19887 (N_19887,N_12166,N_13923);
nor U19888 (N_19888,N_15808,N_13134);
nor U19889 (N_19889,N_12984,N_14857);
nor U19890 (N_19890,N_15995,N_13877);
nor U19891 (N_19891,N_12454,N_13306);
or U19892 (N_19892,N_15831,N_15700);
and U19893 (N_19893,N_12204,N_12856);
or U19894 (N_19894,N_13730,N_12857);
or U19895 (N_19895,N_12543,N_12057);
xor U19896 (N_19896,N_14479,N_13739);
nand U19897 (N_19897,N_12898,N_15637);
xor U19898 (N_19898,N_15008,N_13162);
nand U19899 (N_19899,N_13380,N_14795);
nand U19900 (N_19900,N_14047,N_14121);
or U19901 (N_19901,N_15849,N_13853);
and U19902 (N_19902,N_13389,N_15021);
or U19903 (N_19903,N_13589,N_13792);
or U19904 (N_19904,N_14348,N_14342);
nor U19905 (N_19905,N_14389,N_15220);
or U19906 (N_19906,N_15730,N_14367);
nor U19907 (N_19907,N_12122,N_12496);
or U19908 (N_19908,N_14911,N_15989);
and U19909 (N_19909,N_13769,N_12495);
or U19910 (N_19910,N_12021,N_14695);
nor U19911 (N_19911,N_14008,N_13144);
or U19912 (N_19912,N_15037,N_13607);
xor U19913 (N_19913,N_13426,N_12749);
and U19914 (N_19914,N_12737,N_13161);
nor U19915 (N_19915,N_15667,N_15547);
or U19916 (N_19916,N_12317,N_14746);
or U19917 (N_19917,N_12742,N_12372);
and U19918 (N_19918,N_13740,N_15210);
and U19919 (N_19919,N_14129,N_15218);
and U19920 (N_19920,N_13152,N_14415);
and U19921 (N_19921,N_13497,N_13506);
xnor U19922 (N_19922,N_14522,N_15674);
nand U19923 (N_19923,N_12585,N_12223);
nand U19924 (N_19924,N_12578,N_13450);
and U19925 (N_19925,N_15952,N_13890);
or U19926 (N_19926,N_15138,N_15776);
nor U19927 (N_19927,N_13823,N_14069);
nor U19928 (N_19928,N_12810,N_13987);
nand U19929 (N_19929,N_15153,N_13459);
or U19930 (N_19930,N_15685,N_13950);
or U19931 (N_19931,N_15659,N_13750);
or U19932 (N_19932,N_14608,N_14904);
or U19933 (N_19933,N_15397,N_12072);
nand U19934 (N_19934,N_14135,N_15356);
xor U19935 (N_19935,N_15087,N_13396);
nor U19936 (N_19936,N_12917,N_14428);
nand U19937 (N_19937,N_15317,N_14591);
and U19938 (N_19938,N_12623,N_12065);
nand U19939 (N_19939,N_15117,N_14138);
or U19940 (N_19940,N_15723,N_14362);
nand U19941 (N_19941,N_14816,N_14373);
or U19942 (N_19942,N_14398,N_13019);
or U19943 (N_19943,N_13695,N_15165);
nand U19944 (N_19944,N_15867,N_15622);
nor U19945 (N_19945,N_13624,N_13535);
nand U19946 (N_19946,N_14603,N_13864);
xor U19947 (N_19947,N_12338,N_13411);
and U19948 (N_19948,N_12142,N_12458);
nor U19949 (N_19949,N_12913,N_14014);
or U19950 (N_19950,N_13507,N_13251);
or U19951 (N_19951,N_12080,N_12832);
nor U19952 (N_19952,N_14509,N_12788);
nor U19953 (N_19953,N_13213,N_12766);
nor U19954 (N_19954,N_13027,N_15364);
and U19955 (N_19955,N_12946,N_13076);
nor U19956 (N_19956,N_13165,N_15936);
and U19957 (N_19957,N_12114,N_15616);
and U19958 (N_19958,N_14548,N_14809);
and U19959 (N_19959,N_15896,N_12873);
xor U19960 (N_19960,N_15841,N_14016);
and U19961 (N_19961,N_14457,N_14773);
nor U19962 (N_19962,N_14901,N_12993);
nand U19963 (N_19963,N_14300,N_13486);
nand U19964 (N_19964,N_12179,N_15903);
nor U19965 (N_19965,N_13386,N_13423);
nand U19966 (N_19966,N_14546,N_14643);
nor U19967 (N_19967,N_14960,N_13520);
xnor U19968 (N_19968,N_14238,N_15425);
nand U19969 (N_19969,N_12390,N_12623);
and U19970 (N_19970,N_14081,N_15554);
or U19971 (N_19971,N_15003,N_13060);
nor U19972 (N_19972,N_12383,N_12279);
and U19973 (N_19973,N_12958,N_12777);
or U19974 (N_19974,N_15335,N_13904);
or U19975 (N_19975,N_13286,N_15127);
or U19976 (N_19976,N_14425,N_15070);
xor U19977 (N_19977,N_13790,N_14733);
or U19978 (N_19978,N_13114,N_14756);
or U19979 (N_19979,N_15775,N_12571);
nor U19980 (N_19980,N_13743,N_14215);
nor U19981 (N_19981,N_15509,N_15047);
nand U19982 (N_19982,N_15920,N_15908);
and U19983 (N_19983,N_15285,N_15279);
nand U19984 (N_19984,N_14804,N_14181);
nor U19985 (N_19985,N_13936,N_12515);
nand U19986 (N_19986,N_12558,N_13623);
nor U19987 (N_19987,N_14525,N_14550);
or U19988 (N_19988,N_13405,N_14484);
nor U19989 (N_19989,N_12411,N_12528);
and U19990 (N_19990,N_15582,N_15260);
nor U19991 (N_19991,N_15214,N_15300);
or U19992 (N_19992,N_14616,N_13721);
and U19993 (N_19993,N_14202,N_13012);
nand U19994 (N_19994,N_14637,N_14678);
and U19995 (N_19995,N_14151,N_13516);
or U19996 (N_19996,N_12883,N_15536);
and U19997 (N_19997,N_13895,N_13220);
and U19998 (N_19998,N_15171,N_12725);
or U19999 (N_19999,N_14254,N_14996);
and UO_0 (O_0,N_19392,N_16029);
nor UO_1 (O_1,N_17238,N_17414);
or UO_2 (O_2,N_19547,N_18413);
or UO_3 (O_3,N_16292,N_18759);
nand UO_4 (O_4,N_19162,N_16228);
or UO_5 (O_5,N_16499,N_17733);
or UO_6 (O_6,N_18960,N_17861);
and UO_7 (O_7,N_16712,N_16011);
and UO_8 (O_8,N_19287,N_19596);
xor UO_9 (O_9,N_17185,N_19490);
nor UO_10 (O_10,N_18239,N_19860);
and UO_11 (O_11,N_17977,N_16922);
nand UO_12 (O_12,N_18581,N_19109);
nor UO_13 (O_13,N_18766,N_18039);
nand UO_14 (O_14,N_19632,N_17135);
nor UO_15 (O_15,N_17691,N_17374);
nor UO_16 (O_16,N_16757,N_17894);
or UO_17 (O_17,N_19743,N_19731);
xor UO_18 (O_18,N_19300,N_17525);
nor UO_19 (O_19,N_17795,N_19655);
nor UO_20 (O_20,N_19229,N_16854);
and UO_21 (O_21,N_19619,N_19948);
and UO_22 (O_22,N_19480,N_16999);
and UO_23 (O_23,N_16503,N_17754);
or UO_24 (O_24,N_17944,N_17488);
nand UO_25 (O_25,N_16995,N_17448);
nand UO_26 (O_26,N_18320,N_19177);
nand UO_27 (O_27,N_19918,N_17781);
or UO_28 (O_28,N_17785,N_18476);
xor UO_29 (O_29,N_17317,N_19096);
and UO_30 (O_30,N_16479,N_16792);
nor UO_31 (O_31,N_18227,N_17292);
and UO_32 (O_32,N_18285,N_17101);
and UO_33 (O_33,N_17653,N_16629);
xnor UO_34 (O_34,N_19355,N_17320);
and UO_35 (O_35,N_17847,N_17665);
and UO_36 (O_36,N_16789,N_18262);
nor UO_37 (O_37,N_19118,N_16458);
nor UO_38 (O_38,N_18448,N_17729);
or UO_39 (O_39,N_18196,N_17336);
or UO_40 (O_40,N_18078,N_19947);
and UO_41 (O_41,N_16406,N_18809);
nand UO_42 (O_42,N_19302,N_19774);
nand UO_43 (O_43,N_18100,N_19822);
and UO_44 (O_44,N_16282,N_17145);
nand UO_45 (O_45,N_19757,N_19156);
nor UO_46 (O_46,N_17848,N_19361);
nor UO_47 (O_47,N_16148,N_17255);
nor UO_48 (O_48,N_19911,N_16035);
or UO_49 (O_49,N_17108,N_17730);
and UO_50 (O_50,N_18040,N_17158);
nor UO_51 (O_51,N_17065,N_18543);
and UO_52 (O_52,N_17554,N_19325);
nor UO_53 (O_53,N_16997,N_18670);
or UO_54 (O_54,N_19310,N_16442);
or UO_55 (O_55,N_16304,N_16663);
xnor UO_56 (O_56,N_17631,N_18188);
xnor UO_57 (O_57,N_18477,N_16071);
xnor UO_58 (O_58,N_19227,N_17204);
or UO_59 (O_59,N_17557,N_18138);
nor UO_60 (O_60,N_18662,N_18342);
nor UO_61 (O_61,N_16937,N_17984);
xnor UO_62 (O_62,N_19435,N_16756);
and UO_63 (O_63,N_19925,N_16865);
nor UO_64 (O_64,N_19992,N_18771);
nand UO_65 (O_65,N_17810,N_17028);
and UO_66 (O_66,N_17304,N_18212);
xor UO_67 (O_67,N_18159,N_16489);
and UO_68 (O_68,N_16335,N_18938);
or UO_69 (O_69,N_16085,N_19613);
nand UO_70 (O_70,N_19854,N_16917);
nand UO_71 (O_71,N_18190,N_17353);
and UO_72 (O_72,N_19236,N_18324);
and UO_73 (O_73,N_17079,N_16332);
and UO_74 (O_74,N_19359,N_19523);
nor UO_75 (O_75,N_18683,N_19403);
xor UO_76 (O_76,N_17408,N_18385);
and UO_77 (O_77,N_18592,N_18723);
nand UO_78 (O_78,N_18207,N_19061);
xor UO_79 (O_79,N_16943,N_19638);
nor UO_80 (O_80,N_18487,N_17684);
xor UO_81 (O_81,N_19982,N_16001);
and UO_82 (O_82,N_17714,N_18594);
and UO_83 (O_83,N_16258,N_17744);
and UO_84 (O_84,N_18902,N_19777);
xnor UO_85 (O_85,N_18254,N_16519);
nand UO_86 (O_86,N_18620,N_16630);
and UO_87 (O_87,N_16413,N_16869);
nor UO_88 (O_88,N_18922,N_17860);
or UO_89 (O_89,N_16967,N_19512);
and UO_90 (O_90,N_19189,N_18483);
and UO_91 (O_91,N_16463,N_18005);
nor UO_92 (O_92,N_19183,N_17503);
and UO_93 (O_93,N_19123,N_18945);
nand UO_94 (O_94,N_19168,N_19117);
nor UO_95 (O_95,N_16154,N_16650);
or UO_96 (O_96,N_17950,N_19015);
nand UO_97 (O_97,N_19536,N_16565);
or UO_98 (O_98,N_18497,N_18804);
nor UO_99 (O_99,N_19405,N_17712);
or UO_100 (O_100,N_16984,N_18094);
xnor UO_101 (O_101,N_18618,N_18454);
xor UO_102 (O_102,N_16748,N_16184);
or UO_103 (O_103,N_19961,N_16488);
xor UO_104 (O_104,N_19328,N_18251);
and UO_105 (O_105,N_17772,N_16369);
or UO_106 (O_106,N_17721,N_18905);
nor UO_107 (O_107,N_17090,N_19919);
xor UO_108 (O_108,N_16086,N_16518);
or UO_109 (O_109,N_16752,N_16659);
and UO_110 (O_110,N_17958,N_17357);
and UO_111 (O_111,N_18724,N_16837);
or UO_112 (O_112,N_19668,N_17321);
xnor UO_113 (O_113,N_17583,N_19851);
nor UO_114 (O_114,N_16434,N_19569);
nand UO_115 (O_115,N_19553,N_16170);
nor UO_116 (O_116,N_19873,N_19381);
and UO_117 (O_117,N_18824,N_16446);
or UO_118 (O_118,N_19909,N_17989);
or UO_119 (O_119,N_16068,N_19308);
nand UO_120 (O_120,N_17254,N_19693);
nand UO_121 (O_121,N_19968,N_16061);
nand UO_122 (O_122,N_18979,N_18496);
nand UO_123 (O_123,N_18575,N_19217);
and UO_124 (O_124,N_17076,N_19494);
nand UO_125 (O_125,N_17617,N_19859);
and UO_126 (O_126,N_18810,N_17899);
nand UO_127 (O_127,N_16315,N_18803);
nand UO_128 (O_128,N_18919,N_18583);
or UO_129 (O_129,N_16520,N_18319);
nand UO_130 (O_130,N_16670,N_17107);
nor UO_131 (O_131,N_17981,N_18055);
nor UO_132 (O_132,N_16008,N_18181);
nand UO_133 (O_133,N_17946,N_19319);
xnor UO_134 (O_134,N_19510,N_19863);
and UO_135 (O_135,N_18479,N_18128);
or UO_136 (O_136,N_18537,N_18352);
or UO_137 (O_137,N_16323,N_18370);
or UO_138 (O_138,N_17490,N_19841);
nor UO_139 (O_139,N_17087,N_16283);
and UO_140 (O_140,N_17898,N_17632);
nand UO_141 (O_141,N_17912,N_18248);
nand UO_142 (O_142,N_16591,N_17278);
xnor UO_143 (O_143,N_17579,N_19049);
and UO_144 (O_144,N_16103,N_19175);
or UO_145 (O_145,N_17808,N_17480);
or UO_146 (O_146,N_16745,N_18240);
or UO_147 (O_147,N_16420,N_18193);
nor UO_148 (O_148,N_19294,N_18752);
nand UO_149 (O_149,N_17078,N_17610);
nor UO_150 (O_150,N_18591,N_17225);
and UO_151 (O_151,N_18253,N_16866);
and UO_152 (O_152,N_19993,N_18793);
nand UO_153 (O_153,N_16754,N_18283);
nor UO_154 (O_154,N_18561,N_19609);
or UO_155 (O_155,N_18050,N_18375);
nor UO_156 (O_156,N_18304,N_19820);
xnor UO_157 (O_157,N_19882,N_18402);
xnor UO_158 (O_158,N_19903,N_17156);
and UO_159 (O_159,N_17600,N_19402);
nand UO_160 (O_160,N_17792,N_16667);
and UO_161 (O_161,N_19267,N_16117);
nand UO_162 (O_162,N_18661,N_16422);
nand UO_163 (O_163,N_16447,N_18067);
xor UO_164 (O_164,N_19235,N_16437);
nor UO_165 (O_165,N_17911,N_19354);
nand UO_166 (O_166,N_18850,N_18520);
nor UO_167 (O_167,N_19566,N_17023);
and UO_168 (O_168,N_16370,N_17016);
xor UO_169 (O_169,N_16302,N_18224);
nand UO_170 (O_170,N_16906,N_17413);
and UO_171 (O_171,N_19709,N_19580);
and UO_172 (O_172,N_19631,N_16721);
nand UO_173 (O_173,N_19152,N_17493);
and UO_174 (O_174,N_18808,N_18422);
or UO_175 (O_175,N_16106,N_16825);
nand UO_176 (O_176,N_17869,N_19984);
and UO_177 (O_177,N_19541,N_18486);
nand UO_178 (O_178,N_16514,N_19912);
xnor UO_179 (O_179,N_19349,N_16094);
and UO_180 (O_180,N_17275,N_18644);
nor UO_181 (O_181,N_17831,N_18632);
or UO_182 (O_182,N_17945,N_19672);
and UO_183 (O_183,N_17205,N_19986);
and UO_184 (O_184,N_18812,N_17764);
and UO_185 (O_185,N_16524,N_17777);
nand UO_186 (O_186,N_16975,N_18186);
nand UO_187 (O_187,N_17990,N_19505);
nor UO_188 (O_188,N_18949,N_17259);
nand UO_189 (O_189,N_17951,N_17261);
xor UO_190 (O_190,N_17099,N_17816);
xor UO_191 (O_191,N_17900,N_16336);
nor UO_192 (O_192,N_18499,N_16940);
and UO_193 (O_193,N_18585,N_19900);
nand UO_194 (O_194,N_17774,N_19148);
and UO_195 (O_195,N_19884,N_17940);
nor UO_196 (O_196,N_19180,N_16073);
nor UO_197 (O_197,N_19238,N_18650);
and UO_198 (O_198,N_19249,N_16274);
nor UO_199 (O_199,N_19826,N_17309);
nand UO_200 (O_200,N_18119,N_19868);
and UO_201 (O_201,N_16321,N_18061);
xnor UO_202 (O_202,N_18947,N_17116);
nor UO_203 (O_203,N_17214,N_18237);
and UO_204 (O_204,N_16002,N_18171);
or UO_205 (O_205,N_16362,N_19511);
and UO_206 (O_206,N_16459,N_19926);
nand UO_207 (O_207,N_16130,N_16885);
nand UO_208 (O_208,N_17176,N_18018);
or UO_209 (O_209,N_16242,N_19833);
or UO_210 (O_210,N_18485,N_16423);
or UO_211 (O_211,N_16449,N_17932);
and UO_212 (O_212,N_17469,N_16541);
xnor UO_213 (O_213,N_19304,N_17526);
and UO_214 (O_214,N_17139,N_19726);
nand UO_215 (O_215,N_16562,N_16810);
nand UO_216 (O_216,N_16717,N_19342);
and UO_217 (O_217,N_18068,N_18435);
and UO_218 (O_218,N_16108,N_17882);
nor UO_219 (O_219,N_18893,N_19223);
nor UO_220 (O_220,N_16722,N_17709);
or UO_221 (O_221,N_19362,N_18028);
nand UO_222 (O_222,N_16875,N_19788);
or UO_223 (O_223,N_17578,N_16219);
nor UO_224 (O_224,N_16005,N_18731);
xnor UO_225 (O_225,N_17843,N_16234);
nand UO_226 (O_226,N_16121,N_18003);
or UO_227 (O_227,N_16768,N_19271);
nor UO_228 (O_228,N_18136,N_17456);
nor UO_229 (O_229,N_17701,N_16398);
nand UO_230 (O_230,N_18916,N_19973);
nor UO_231 (O_231,N_18876,N_17710);
and UO_232 (O_232,N_17359,N_19037);
nand UO_233 (O_233,N_16681,N_17715);
and UO_234 (O_234,N_19880,N_18436);
xor UO_235 (O_235,N_17089,N_19198);
xor UO_236 (O_236,N_16288,N_17114);
and UO_237 (O_237,N_17876,N_17479);
xor UO_238 (O_238,N_16870,N_17143);
and UO_239 (O_239,N_17546,N_17606);
or UO_240 (O_240,N_18587,N_18408);
and UO_241 (O_241,N_17608,N_19928);
nand UO_242 (O_242,N_16500,N_18617);
and UO_243 (O_243,N_18826,N_16763);
nor UO_244 (O_244,N_17818,N_16718);
nor UO_245 (O_245,N_18358,N_18480);
or UO_246 (O_246,N_16435,N_16773);
nor UO_247 (O_247,N_19472,N_17505);
or UO_248 (O_248,N_18711,N_17594);
nand UO_249 (O_249,N_17495,N_16063);
or UO_250 (O_250,N_18382,N_18406);
xor UO_251 (O_251,N_17763,N_16338);
or UO_252 (O_252,N_17804,N_18354);
or UO_253 (O_253,N_17192,N_19969);
and UO_254 (O_254,N_18700,N_19033);
or UO_255 (O_255,N_16122,N_18841);
nand UO_256 (O_256,N_16797,N_17838);
nor UO_257 (O_257,N_18574,N_16343);
or UO_258 (O_258,N_17858,N_18242);
and UO_259 (O_259,N_18524,N_19830);
nor UO_260 (O_260,N_19888,N_17095);
nor UO_261 (O_261,N_18547,N_17467);
or UO_262 (O_262,N_17293,N_19654);
nor UO_263 (O_263,N_16003,N_18709);
and UO_264 (O_264,N_16620,N_19088);
xor UO_265 (O_265,N_17438,N_17311);
nand UO_266 (O_266,N_16775,N_16666);
and UO_267 (O_267,N_18820,N_18705);
nand UO_268 (O_268,N_19920,N_19814);
and UO_269 (O_269,N_16521,N_16477);
nor UO_270 (O_270,N_17629,N_17906);
nor UO_271 (O_271,N_19185,N_17755);
xor UO_272 (O_272,N_17636,N_19414);
nor UO_273 (O_273,N_16824,N_16371);
nor UO_274 (O_274,N_18955,N_18492);
nand UO_275 (O_275,N_18441,N_19292);
or UO_276 (O_276,N_16075,N_17398);
nand UO_277 (O_277,N_18295,N_17252);
or UO_278 (O_278,N_19782,N_16511);
nand UO_279 (O_279,N_18223,N_17555);
nand UO_280 (O_280,N_18943,N_17697);
nand UO_281 (O_281,N_19315,N_19811);
or UO_282 (O_282,N_17171,N_19507);
or UO_283 (O_283,N_19462,N_19197);
xnor UO_284 (O_284,N_18481,N_16864);
nor UO_285 (O_285,N_18488,N_18570);
nand UO_286 (O_286,N_19058,N_19770);
or UO_287 (O_287,N_17313,N_16390);
nand UO_288 (O_288,N_16077,N_16595);
nand UO_289 (O_289,N_16091,N_18868);
or UO_290 (O_290,N_17794,N_16217);
or UO_291 (O_291,N_19172,N_17758);
and UO_292 (O_292,N_17406,N_16089);
and UO_293 (O_293,N_19627,N_16092);
or UO_294 (O_294,N_17072,N_18351);
and UO_295 (O_295,N_17197,N_19026);
nor UO_296 (O_296,N_19699,N_19714);
or UO_297 (O_297,N_17280,N_19681);
nor UO_298 (O_298,N_16015,N_16350);
nand UO_299 (O_299,N_18807,N_17532);
or UO_300 (O_300,N_19196,N_19815);
nor UO_301 (O_301,N_18162,N_17660);
nor UO_302 (O_302,N_16897,N_19913);
nor UO_303 (O_303,N_19520,N_19209);
and UO_304 (O_304,N_19230,N_18062);
or UO_305 (O_305,N_19112,N_19537);
and UO_306 (O_306,N_18639,N_18472);
xor UO_307 (O_307,N_18569,N_17350);
nand UO_308 (O_308,N_18869,N_17821);
and UO_309 (O_309,N_16613,N_17652);
and UO_310 (O_310,N_18118,N_17745);
and UO_311 (O_311,N_17923,N_18083);
or UO_312 (O_312,N_17635,N_16129);
or UO_313 (O_313,N_16761,N_17206);
nor UO_314 (O_314,N_17120,N_19802);
nor UO_315 (O_315,N_17459,N_16724);
and UO_316 (O_316,N_18802,N_18696);
nand UO_317 (O_317,N_16579,N_17559);
xnor UO_318 (O_318,N_19850,N_19543);
nor UO_319 (O_319,N_16504,N_17988);
nor UO_320 (O_320,N_16929,N_16786);
and UO_321 (O_321,N_19445,N_16767);
or UO_322 (O_322,N_16576,N_16855);
and UO_323 (O_323,N_19752,N_16549);
and UO_324 (O_324,N_16603,N_18187);
nand UO_325 (O_325,N_18727,N_18192);
nor UO_326 (O_326,N_18391,N_16583);
nand UO_327 (O_327,N_16515,N_18950);
and UO_328 (O_328,N_19044,N_17046);
nor UO_329 (O_329,N_18953,N_16244);
and UO_330 (O_330,N_19040,N_16349);
xnor UO_331 (O_331,N_18213,N_16218);
or UO_332 (O_332,N_18866,N_18498);
or UO_333 (O_333,N_18553,N_19396);
and UO_334 (O_334,N_17088,N_16739);
and UO_335 (O_335,N_18341,N_18090);
nor UO_336 (O_336,N_17622,N_19460);
nor UO_337 (O_337,N_18070,N_16705);
nand UO_338 (O_338,N_19704,N_19297);
and UO_339 (O_339,N_16607,N_19082);
nand UO_340 (O_340,N_16662,N_18234);
nand UO_341 (O_341,N_17801,N_18367);
nand UO_342 (O_342,N_16974,N_16537);
nand UO_343 (O_343,N_18403,N_19746);
nor UO_344 (O_344,N_18048,N_18649);
or UO_345 (O_345,N_18183,N_18029);
nor UO_346 (O_346,N_18322,N_18867);
nand UO_347 (O_347,N_19261,N_17683);
and UO_348 (O_348,N_19876,N_16564);
nor UO_349 (O_349,N_17068,N_16441);
or UO_350 (O_350,N_18501,N_17172);
nand UO_351 (O_351,N_18298,N_16533);
nand UO_352 (O_352,N_19182,N_18442);
nand UO_353 (O_353,N_18386,N_17337);
nand UO_354 (O_354,N_19639,N_18758);
xor UO_355 (O_355,N_16919,N_19397);
or UO_356 (O_356,N_19797,N_17713);
and UO_357 (O_357,N_19624,N_19215);
or UO_358 (O_358,N_17118,N_19094);
and UO_359 (O_359,N_18363,N_19901);
or UO_360 (O_360,N_19050,N_18806);
and UO_361 (O_361,N_18630,N_17437);
and UO_362 (O_362,N_19019,N_17022);
nor UO_363 (O_363,N_17690,N_16510);
nand UO_364 (O_364,N_18774,N_18629);
or UO_365 (O_365,N_18097,N_18468);
and UO_366 (O_366,N_17720,N_18823);
nor UO_367 (O_367,N_19531,N_16405);
xnor UO_368 (O_368,N_16374,N_18046);
nand UO_369 (O_369,N_16507,N_18527);
nor UO_370 (O_370,N_16078,N_17322);
xor UO_371 (O_371,N_17999,N_19419);
xor UO_372 (O_372,N_18228,N_17541);
xor UO_373 (O_373,N_18624,N_18348);
or UO_374 (O_374,N_16735,N_16112);
nor UO_375 (O_375,N_19975,N_16911);
nand UO_376 (O_376,N_19701,N_19821);
and UO_377 (O_377,N_16986,N_16365);
and UO_378 (O_378,N_18113,N_19207);
or UO_379 (O_379,N_16806,N_18800);
and UO_380 (O_380,N_17117,N_17982);
nand UO_381 (O_381,N_18131,N_17201);
and UO_382 (O_382,N_17236,N_18538);
nor UO_383 (O_383,N_16738,N_17338);
nor UO_384 (O_384,N_16083,N_19393);
or UO_385 (O_385,N_19338,N_17221);
xor UO_386 (O_386,N_16672,N_18238);
or UO_387 (O_387,N_16291,N_17431);
nand UO_388 (O_388,N_16570,N_18672);
nand UO_389 (O_389,N_19369,N_16776);
and UO_390 (O_390,N_18789,N_18350);
xor UO_391 (O_391,N_17105,N_16820);
or UO_392 (O_392,N_16054,N_18783);
nor UO_393 (O_393,N_18708,N_17805);
or UO_394 (O_394,N_17687,N_19253);
and UO_395 (O_395,N_18056,N_17991);
and UO_396 (O_396,N_16165,N_16225);
nand UO_397 (O_397,N_17036,N_18420);
or UO_398 (O_398,N_16544,N_17362);
xor UO_399 (O_399,N_17352,N_18658);
and UO_400 (O_400,N_16993,N_16925);
and UO_401 (O_401,N_18834,N_16725);
nor UO_402 (O_402,N_18034,N_19616);
and UO_403 (O_403,N_17674,N_16556);
nand UO_404 (O_404,N_16699,N_18918);
nand UO_405 (O_405,N_16399,N_18865);
or UO_406 (O_406,N_16578,N_19143);
xnor UO_407 (O_407,N_17442,N_16815);
or UO_408 (O_408,N_17434,N_19581);
or UO_409 (O_409,N_19771,N_19285);
and UO_410 (O_410,N_19358,N_17563);
and UO_411 (O_411,N_17196,N_19720);
or UO_412 (O_412,N_16568,N_16881);
or UO_413 (O_413,N_18270,N_19113);
nor UO_414 (O_414,N_19600,N_17884);
nor UO_415 (O_415,N_19705,N_19125);
nor UO_416 (O_416,N_18532,N_18356);
nor UO_417 (O_417,N_16044,N_17006);
and UO_418 (O_418,N_17512,N_19952);
nor UO_419 (O_419,N_16300,N_19590);
xnor UO_420 (O_420,N_19255,N_19719);
nor UO_421 (O_421,N_18719,N_17973);
xnor UO_422 (O_422,N_19495,N_17189);
and UO_423 (O_423,N_17859,N_18163);
nor UO_424 (O_424,N_18792,N_18857);
or UO_425 (O_425,N_16693,N_18556);
nor UO_426 (O_426,N_17696,N_17100);
xnor UO_427 (O_427,N_16923,N_17323);
and UO_428 (O_428,N_16539,N_17180);
or UO_429 (O_429,N_16661,N_17267);
nor UO_430 (O_430,N_18651,N_16638);
or UO_431 (O_431,N_17675,N_17427);
and UO_432 (O_432,N_19933,N_17411);
or UO_433 (O_433,N_18886,N_18885);
nor UO_434 (O_434,N_16115,N_18176);
nand UO_435 (O_435,N_19345,N_19649);
or UO_436 (O_436,N_17726,N_16769);
xnor UO_437 (O_437,N_17450,N_19137);
nor UO_438 (O_438,N_16654,N_18085);
nor UO_439 (O_439,N_18550,N_18060);
nand UO_440 (O_440,N_18859,N_19736);
and UO_441 (O_441,N_19716,N_18679);
nand UO_442 (O_442,N_18703,N_16691);
nor UO_443 (O_443,N_18677,N_18431);
or UO_444 (O_444,N_17743,N_18294);
nor UO_445 (O_445,N_18194,N_17222);
or UO_446 (O_446,N_19949,N_16918);
nand UO_447 (O_447,N_16469,N_17520);
and UO_448 (O_448,N_16577,N_18006);
and UO_449 (O_449,N_19930,N_17308);
xnor UO_450 (O_450,N_19650,N_18935);
nand UO_451 (O_451,N_17115,N_18530);
nand UO_452 (O_452,N_18787,N_18631);
nor UO_453 (O_453,N_18767,N_16272);
nor UO_454 (O_454,N_18044,N_19010);
and UO_455 (O_455,N_17356,N_19001);
nor UO_456 (O_456,N_19431,N_16857);
nor UO_457 (O_457,N_17786,N_17751);
and UO_458 (O_458,N_19957,N_18421);
xnor UO_459 (O_459,N_16114,N_16301);
nor UO_460 (O_460,N_19447,N_16146);
xnor UO_461 (O_461,N_19558,N_18475);
nor UO_462 (O_462,N_19781,N_19994);
or UO_463 (O_463,N_19905,N_17813);
nand UO_464 (O_464,N_17957,N_17966);
nand UO_465 (O_465,N_17399,N_18995);
or UO_466 (O_466,N_18558,N_16161);
or UO_467 (O_467,N_17596,N_16410);
nor UO_468 (O_468,N_19506,N_19312);
and UO_469 (O_469,N_16445,N_19382);
nand UO_470 (O_470,N_16840,N_19140);
nand UO_471 (O_471,N_19092,N_16303);
or UO_472 (O_472,N_17224,N_18621);
nor UO_473 (O_473,N_17530,N_18353);
or UO_474 (O_474,N_19108,N_16386);
and UO_475 (O_475,N_17478,N_19463);
and UO_476 (O_476,N_17699,N_16602);
or UO_477 (O_477,N_19576,N_16891);
and UO_478 (O_478,N_19907,N_16956);
xnor UO_479 (O_479,N_17487,N_16339);
nand UO_480 (O_480,N_17829,N_16606);
nor UO_481 (O_481,N_19767,N_17891);
nor UO_482 (O_482,N_16022,N_19931);
or UO_483 (O_483,N_18052,N_18712);
or UO_484 (O_484,N_18968,N_18858);
nand UO_485 (O_485,N_18278,N_16558);
nor UO_486 (O_486,N_16081,N_17266);
nor UO_487 (O_487,N_19922,N_16656);
and UO_488 (O_488,N_19356,N_17045);
nor UO_489 (O_489,N_18878,N_17949);
nand UO_490 (O_490,N_16941,N_16373);
nor UO_491 (O_491,N_16107,N_16596);
and UO_492 (O_492,N_19664,N_19351);
nand UO_493 (O_493,N_19211,N_17962);
nand UO_494 (O_494,N_19098,N_19067);
xnor UO_495 (O_495,N_16051,N_17878);
or UO_496 (O_496,N_16230,N_16356);
and UO_497 (O_497,N_16006,N_17986);
xnor UO_498 (O_498,N_19667,N_18389);
nand UO_499 (O_499,N_17778,N_19153);
nand UO_500 (O_500,N_19055,N_17239);
nor UO_501 (O_501,N_19430,N_17253);
nor UO_502 (O_502,N_18232,N_17144);
nand UO_503 (O_503,N_17200,N_16182);
nand UO_504 (O_504,N_18339,N_17473);
and UO_505 (O_505,N_18963,N_18439);
or UO_506 (O_506,N_17020,N_19458);
nor UO_507 (O_507,N_16366,N_16342);
xnor UO_508 (O_508,N_19545,N_19390);
and UO_509 (O_509,N_19158,N_19187);
nor UO_510 (O_510,N_19552,N_18552);
nor UO_511 (O_511,N_19628,N_18219);
nor UO_512 (O_512,N_16802,N_19891);
nor UO_513 (O_513,N_17689,N_18855);
nand UO_514 (O_514,N_18615,N_16702);
nand UO_515 (O_515,N_17383,N_16160);
xor UO_516 (O_516,N_19233,N_17749);
and UO_517 (O_517,N_19476,N_18280);
nor UO_518 (O_518,N_18948,N_16970);
or UO_519 (O_519,N_17166,N_19089);
nand UO_520 (O_520,N_19306,N_16788);
nand UO_521 (O_521,N_19035,N_19146);
or UO_522 (O_522,N_17640,N_17423);
nand UO_523 (O_523,N_19964,N_19320);
nand UO_524 (O_524,N_18531,N_19670);
or UO_525 (O_525,N_17595,N_19881);
or UO_526 (O_526,N_19823,N_19843);
nand UO_527 (O_527,N_18096,N_19885);
nand UO_528 (O_528,N_18268,N_17614);
nand UO_529 (O_529,N_16535,N_18013);
and UO_530 (O_530,N_19084,N_16169);
and UO_531 (O_531,N_18977,N_17811);
nor UO_532 (O_532,N_16803,N_17564);
xor UO_533 (O_533,N_18371,N_18980);
and UO_534 (O_534,N_18146,N_17570);
nand UO_535 (O_535,N_18444,N_16939);
nor UO_536 (O_536,N_17075,N_16559);
nor UO_537 (O_537,N_18216,N_16452);
xnor UO_538 (O_538,N_16785,N_19231);
nand UO_539 (O_539,N_17149,N_16293);
nor UO_540 (O_540,N_19344,N_16453);
and UO_541 (O_541,N_18045,N_18970);
and UO_542 (O_542,N_19456,N_17589);
xnor UO_543 (O_543,N_19091,N_19656);
nand UO_544 (O_544,N_18799,N_17179);
nand UO_545 (O_545,N_18199,N_16571);
nor UO_546 (O_546,N_18978,N_19174);
and UO_547 (O_547,N_16185,N_17992);
and UO_548 (O_548,N_18201,N_18545);
nor UO_549 (O_549,N_19924,N_16674);
nor UO_550 (O_550,N_17619,N_19839);
nor UO_551 (O_551,N_18656,N_18892);
or UO_552 (O_552,N_16992,N_17375);
or UO_553 (O_553,N_18753,N_19387);
and UO_554 (O_554,N_18437,N_19395);
and UO_555 (O_555,N_17871,N_17803);
nand UO_556 (O_556,N_19789,N_17397);
nor UO_557 (O_557,N_17879,N_19434);
nor UO_558 (O_558,N_16492,N_17857);
nand UO_559 (O_559,N_19519,N_18931);
and UO_560 (O_560,N_16977,N_19027);
and UO_561 (O_561,N_16618,N_19022);
and UO_562 (O_562,N_16019,N_19776);
or UO_563 (O_563,N_16004,N_18053);
nand UO_564 (O_564,N_18998,N_16700);
xor UO_565 (O_565,N_19685,N_18961);
or UO_566 (O_566,N_16552,N_19606);
and UO_567 (O_567,N_18484,N_18827);
nor UO_568 (O_568,N_16742,N_17227);
and UO_569 (O_569,N_19401,N_18814);
or UO_570 (O_570,N_18710,N_19150);
and UO_571 (O_571,N_16833,N_19245);
nor UO_572 (O_572,N_16222,N_18702);
or UO_573 (O_573,N_18775,N_18210);
or UO_574 (O_574,N_19090,N_18482);
and UO_575 (O_575,N_18445,N_17637);
or UO_576 (O_576,N_18059,N_19644);
xor UO_577 (O_577,N_16212,N_16836);
or UO_578 (O_578,N_18836,N_18519);
nor UO_579 (O_579,N_18726,N_16762);
nand UO_580 (O_580,N_17182,N_16155);
xnor UO_581 (O_581,N_19807,N_16104);
nand UO_582 (O_582,N_18080,N_19346);
or UO_583 (O_583,N_17937,N_18642);
and UO_584 (O_584,N_17603,N_16861);
nor UO_585 (O_585,N_18942,N_19728);
and UO_586 (O_586,N_17747,N_16162);
xor UO_587 (O_587,N_19425,N_19643);
or UO_588 (O_588,N_18830,N_16416);
nor UO_589 (O_589,N_18816,N_16538);
and UO_590 (O_590,N_18082,N_16683);
or UO_591 (O_591,N_17802,N_17418);
nor UO_592 (O_592,N_18965,N_18999);
nand UO_593 (O_593,N_18603,N_18637);
and UO_594 (O_594,N_17034,N_18263);
nand UO_595 (O_595,N_17866,N_18191);
nor UO_596 (O_596,N_19778,N_18981);
and UO_597 (O_597,N_19142,N_16847);
or UO_598 (O_598,N_18275,N_19908);
nor UO_599 (O_599,N_17662,N_16460);
nor UO_600 (O_600,N_17927,N_17127);
and UO_601 (O_601,N_17061,N_16266);
and UO_602 (O_602,N_16388,N_16750);
nor UO_603 (O_603,N_17716,N_17867);
nand UO_604 (O_604,N_18974,N_16604);
nand UO_605 (O_605,N_18564,N_19149);
nor UO_606 (O_606,N_16592,N_18145);
nand UO_607 (O_607,N_17630,N_19540);
and UO_608 (O_608,N_18526,N_17062);
nor UO_609 (O_609,N_18008,N_17654);
or UO_610 (O_610,N_16903,N_16096);
nand UO_611 (O_611,N_18172,N_18127);
nand UO_612 (O_612,N_16016,N_17363);
and UO_613 (O_613,N_19126,N_19465);
nor UO_614 (O_614,N_19222,N_17706);
or UO_615 (O_615,N_18103,N_17432);
xor UO_616 (O_616,N_16793,N_18409);
or UO_617 (O_617,N_17832,N_17897);
and UO_618 (O_618,N_16876,N_17700);
nor UO_619 (O_619,N_19047,N_19677);
and UO_620 (O_620,N_19134,N_17436);
nor UO_621 (O_621,N_17207,N_18414);
and UO_622 (O_622,N_19479,N_19684);
nor UO_623 (O_623,N_19983,N_18395);
and UO_624 (O_624,N_17573,N_17807);
nor UO_625 (O_625,N_19899,N_19595);
xnor UO_626 (O_626,N_17002,N_17765);
or UO_627 (O_627,N_18019,N_17645);
nor UO_628 (O_628,N_16069,N_17300);
or UO_629 (O_629,N_18593,N_16232);
nor UO_630 (O_630,N_17086,N_17823);
nor UO_631 (O_631,N_19516,N_17104);
nand UO_632 (O_632,N_19159,N_16196);
and UO_633 (O_633,N_17815,N_19784);
or UO_634 (O_634,N_16853,N_17331);
xnor UO_635 (O_635,N_18798,N_17620);
and UO_636 (O_636,N_16953,N_18274);
or UO_637 (O_637,N_19305,N_17486);
or UO_638 (O_638,N_17746,N_18451);
xnor UO_639 (O_639,N_17607,N_16340);
nand UO_640 (O_640,N_19513,N_16497);
nor UO_641 (O_641,N_17420,N_19131);
nor UO_642 (O_642,N_17552,N_18689);
nand UO_643 (O_643,N_18595,N_18739);
xor UO_644 (O_644,N_16214,N_19567);
nand UO_645 (O_645,N_16381,N_19625);
nand UO_646 (O_646,N_17245,N_19248);
and UO_647 (O_647,N_17510,N_18926);
and UO_648 (O_648,N_16448,N_16275);
nor UO_649 (O_649,N_19439,N_17820);
nand UO_650 (O_650,N_18106,N_16641);
nor UO_651 (O_651,N_18506,N_16010);
nand UO_652 (O_652,N_19852,N_17693);
nand UO_653 (O_653,N_17655,N_17188);
nor UO_654 (O_654,N_19717,N_18197);
or UO_655 (O_655,N_17770,N_19412);
nand UO_656 (O_656,N_18158,N_16529);
nand UO_657 (O_657,N_17499,N_18474);
nand UO_658 (O_658,N_18001,N_16261);
nor UO_659 (O_659,N_16290,N_17500);
and UO_660 (O_660,N_19764,N_18390);
and UO_661 (O_661,N_17297,N_16047);
nor UO_662 (O_662,N_19028,N_19960);
nand UO_663 (O_663,N_16128,N_16850);
and UO_664 (O_664,N_17217,N_16731);
nor UO_665 (O_665,N_16076,N_16440);
nor UO_666 (O_666,N_17870,N_18665);
nand UO_667 (O_667,N_19858,N_19436);
and UO_668 (O_668,N_18845,N_18139);
and UO_669 (O_669,N_19645,N_18597);
nand UO_670 (O_670,N_19651,N_19034);
nor UO_671 (O_671,N_16631,N_18906);
or UO_672 (O_672,N_16279,N_19598);
or UO_673 (O_673,N_19404,N_16046);
nand UO_674 (O_674,N_18897,N_17996);
and UO_675 (O_675,N_18725,N_18907);
nand UO_676 (O_676,N_19206,N_18657);
xnor UO_677 (O_677,N_16730,N_18560);
xnor UO_678 (O_678,N_19694,N_16254);
and UO_679 (O_679,N_17688,N_16243);
or UO_680 (O_680,N_16874,N_19164);
nand UO_681 (O_681,N_18794,N_19865);
nor UO_682 (O_682,N_19785,N_19442);
and UO_683 (O_683,N_19893,N_18025);
or UO_684 (O_684,N_18247,N_17790);
xor UO_685 (O_685,N_16701,N_19009);
nor UO_686 (O_686,N_17290,N_17123);
xnor UO_687 (O_687,N_16589,N_19703);
and UO_688 (O_688,N_17441,N_19564);
or UO_689 (O_689,N_19951,N_19186);
xor UO_690 (O_690,N_18737,N_17836);
xnor UO_691 (O_691,N_19497,N_18129);
nor UO_692 (O_692,N_19484,N_18720);
or UO_693 (O_693,N_18608,N_19429);
nand UO_694 (O_694,N_19665,N_16375);
or UO_695 (O_695,N_19840,N_19124);
or UO_696 (O_696,N_19834,N_17121);
or UO_697 (O_697,N_18847,N_18882);
or UO_698 (O_698,N_19538,N_19070);
or UO_699 (O_699,N_19138,N_18932);
or UO_700 (O_700,N_17351,N_18666);
xnor UO_701 (O_701,N_18860,N_16147);
nand UO_702 (O_702,N_18751,N_18625);
and UO_703 (O_703,N_17854,N_16888);
or UO_704 (O_704,N_18399,N_18598);
nand UO_705 (O_705,N_18323,N_17657);
and UO_706 (O_706,N_18790,N_16333);
nand UO_707 (O_707,N_16202,N_18054);
or UO_708 (O_708,N_17809,N_19932);
nand UO_709 (O_709,N_17769,N_17567);
xnor UO_710 (O_710,N_17421,N_19360);
and UO_711 (O_711,N_19524,N_18327);
and UO_712 (O_712,N_17283,N_18218);
nand UO_713 (O_713,N_16646,N_16741);
nor UO_714 (O_714,N_16688,N_17538);
nor UO_715 (O_715,N_19284,N_16780);
and UO_716 (O_716,N_19410,N_17494);
nor UO_717 (O_717,N_18578,N_16041);
nor UO_718 (O_718,N_17491,N_19542);
nand UO_719 (O_719,N_18300,N_16633);
or UO_720 (O_720,N_18494,N_16651);
nand UO_721 (O_721,N_18613,N_18331);
nor UO_722 (O_722,N_16120,N_18452);
nand UO_723 (O_723,N_18453,N_18010);
or UO_724 (O_724,N_17647,N_19181);
or UO_725 (O_725,N_17430,N_19237);
nor UO_726 (O_726,N_17163,N_18469);
and UO_727 (O_727,N_17366,N_19641);
nor UO_728 (O_728,N_18132,N_16844);
and UO_729 (O_729,N_18401,N_18817);
nand UO_730 (O_730,N_19388,N_17522);
nor UO_731 (O_731,N_17106,N_19157);
xor UO_732 (O_732,N_16527,N_18762);
nor UO_733 (O_733,N_18681,N_18393);
and UO_734 (O_734,N_18688,N_17668);
and UO_735 (O_735,N_19097,N_16969);
nor UO_736 (O_736,N_17994,N_19093);
xnor UO_737 (O_737,N_16851,N_16125);
and UO_738 (O_738,N_18110,N_16892);
xnor UO_739 (O_739,N_17575,N_19482);
and UO_740 (O_740,N_18889,N_19054);
nor UO_741 (O_741,N_17671,N_16550);
nand UO_742 (O_742,N_16271,N_16697);
or UO_743 (O_743,N_19483,N_16787);
or UO_744 (O_744,N_19039,N_19810);
xor UO_745 (O_745,N_18966,N_16496);
and UO_746 (O_746,N_16884,N_19621);
nor UO_747 (O_747,N_19769,N_19466);
and UO_748 (O_748,N_19499,N_18470);
or UO_749 (O_749,N_16421,N_16126);
nor UO_750 (O_750,N_16942,N_19587);
nand UO_751 (O_751,N_17943,N_17031);
or UO_752 (O_752,N_17681,N_18122);
or UO_753 (O_753,N_19972,N_19470);
and UO_754 (O_754,N_18588,N_16635);
nor UO_755 (O_755,N_18715,N_17511);
nand UO_756 (O_756,N_18160,N_16252);
and UO_757 (O_757,N_17928,N_19468);
nor UO_758 (O_758,N_17621,N_19014);
nor UO_759 (O_759,N_16201,N_17226);
nand UO_760 (O_760,N_18757,N_17910);
and UO_761 (O_761,N_19981,N_18911);
xor UO_762 (O_762,N_16322,N_19008);
xnor UO_763 (O_763,N_16394,N_16326);
or UO_764 (O_764,N_17365,N_19675);
nor UO_765 (O_765,N_17814,N_18337);
and UO_766 (O_766,N_16259,N_16588);
nor UO_767 (O_767,N_17718,N_19161);
or UO_768 (O_768,N_16947,N_17667);
and UO_769 (O_769,N_19075,N_19389);
nor UO_770 (O_770,N_17367,N_19713);
xnor UO_771 (O_771,N_19264,N_16059);
xor UO_772 (O_772,N_19514,N_17470);
nor UO_773 (O_773,N_17740,N_19079);
nor UO_774 (O_774,N_17468,N_18539);
nor UO_775 (O_775,N_19582,N_17628);
nor UO_776 (O_776,N_19321,N_17965);
nand UO_777 (O_777,N_19228,N_19129);
or UO_778 (O_778,N_17312,N_19060);
or UO_779 (O_779,N_16883,N_16601);
nand UO_780 (O_780,N_19825,N_17119);
nand UO_781 (O_781,N_16877,N_19000);
or UO_782 (O_782,N_17704,N_18064);
and UO_783 (O_783,N_18260,N_18584);
and UO_784 (O_784,N_17529,N_16064);
and UO_785 (O_785,N_18038,N_19653);
nor UO_786 (O_786,N_18909,N_19671);
nand UO_787 (O_787,N_18338,N_18923);
and UO_788 (O_788,N_16348,N_16110);
or UO_789 (O_789,N_19399,N_16099);
xnor UO_790 (O_790,N_17404,N_16560);
nand UO_791 (O_791,N_17644,N_19330);
nand UO_792 (O_792,N_19130,N_18256);
or UO_793 (O_793,N_16971,N_19110);
nand UO_794 (O_794,N_17880,N_18189);
xor UO_795 (O_795,N_19842,N_18554);
or UO_796 (O_796,N_17440,N_16540);
and UO_797 (O_797,N_17523,N_17533);
nand UO_798 (O_798,N_18733,N_19415);
or UO_799 (O_799,N_19828,N_16425);
and UO_800 (O_800,N_19357,N_17893);
or UO_801 (O_801,N_17348,N_18743);
or UO_802 (O_802,N_16909,N_18842);
nand UO_803 (O_803,N_16868,N_19317);
and UO_804 (O_804,N_17160,N_16819);
or UO_805 (O_805,N_16175,N_17753);
xor UO_806 (O_806,N_19554,N_17272);
or UO_807 (O_807,N_17000,N_16968);
and UO_808 (O_808,N_16152,N_16194);
and UO_809 (O_809,N_17274,N_18465);
nand UO_810 (O_810,N_16345,N_18231);
nor UO_811 (O_811,N_19491,N_17676);
nand UO_812 (O_812,N_19742,N_18208);
and UO_813 (O_813,N_18017,N_19690);
and UO_814 (O_814,N_19059,N_17465);
nand UO_815 (O_815,N_18840,N_16843);
and UO_816 (O_816,N_17800,N_18929);
nor UO_817 (O_817,N_17760,N_16097);
nand UO_818 (O_818,N_16021,N_18020);
xor UO_819 (O_819,N_16916,N_19855);
and UO_820 (O_820,N_19326,N_16610);
nor UO_821 (O_821,N_19874,N_17669);
nor UO_822 (O_822,N_16501,N_19103);
or UO_823 (O_823,N_19464,N_18284);
nand UO_824 (O_824,N_19734,N_16584);
and UO_825 (O_825,N_17798,N_16313);
nor UO_826 (O_826,N_16657,N_18315);
or UO_827 (O_827,N_16632,N_19607);
or UO_828 (O_828,N_17917,N_16944);
nand UO_829 (O_829,N_19646,N_19698);
nor UO_830 (O_830,N_16238,N_16575);
nor UO_831 (O_831,N_16391,N_16759);
xnor UO_832 (O_832,N_16782,N_17451);
and UO_833 (O_833,N_19428,N_17010);
nor UO_834 (O_834,N_18984,N_17433);
nand UO_835 (O_835,N_17841,N_19579);
xor UO_836 (O_836,N_17624,N_16744);
xor UO_837 (O_837,N_18879,N_17109);
nand UO_838 (O_838,N_16189,N_18092);
nand UO_839 (O_839,N_18596,N_16058);
nor UO_840 (O_840,N_18249,N_17386);
xor UO_841 (O_841,N_18141,N_18073);
or UO_842 (O_842,N_17388,N_19759);
nand UO_843 (O_843,N_16842,N_16400);
and UO_844 (O_844,N_16172,N_19391);
and UO_845 (O_845,N_16643,N_17230);
or UO_846 (O_846,N_16972,N_18333);
xor UO_847 (O_847,N_19692,N_18646);
xor UO_848 (O_848,N_17634,N_19432);
nor UO_849 (O_849,N_18116,N_16359);
or UO_850 (O_850,N_17347,N_19178);
nor UO_851 (O_851,N_19944,N_19296);
xor UO_852 (O_852,N_18473,N_18117);
and UO_853 (O_853,N_16241,N_19799);
and UO_854 (O_854,N_17582,N_18379);
nand UO_855 (O_855,N_18996,N_16166);
nor UO_856 (O_856,N_19214,N_16007);
nand UO_857 (O_857,N_18921,N_18438);
or UO_858 (O_858,N_18058,N_19220);
xor UO_859 (O_859,N_18738,N_18104);
nor UO_860 (O_860,N_19659,N_16962);
and UO_861 (O_861,N_17345,N_16673);
or UO_862 (O_862,N_16753,N_17953);
and UO_863 (O_863,N_17342,N_18610);
and UO_864 (O_864,N_16615,N_19521);
nor UO_865 (O_865,N_18779,N_16706);
nand UO_866 (O_866,N_19678,N_16551);
xor UO_867 (O_867,N_16328,N_18007);
and UO_868 (O_868,N_18691,N_17410);
and UO_869 (O_869,N_18204,N_16933);
and UO_870 (O_870,N_18057,N_18831);
and UO_871 (O_871,N_19262,N_16325);
nand UO_872 (O_872,N_19657,N_16367);
nor UO_873 (O_873,N_19194,N_18023);
nand UO_874 (O_874,N_17611,N_16996);
nand UO_875 (O_875,N_18463,N_19577);
nand UO_876 (O_876,N_16317,N_19758);
nor UO_877 (O_877,N_16856,N_19452);
and UO_878 (O_878,N_16920,N_19829);
nand UO_879 (O_879,N_19739,N_16680);
nand UO_880 (O_880,N_19791,N_17707);
xor UO_881 (O_881,N_19555,N_16586);
xor UO_882 (O_882,N_18449,N_19706);
nor UO_883 (O_883,N_18383,N_17514);
or UO_884 (O_884,N_17247,N_17887);
nand UO_885 (O_885,N_16818,N_19052);
or UO_886 (O_886,N_16268,N_16102);
and UO_887 (O_887,N_19967,N_17327);
and UO_888 (O_888,N_17153,N_18303);
nand UO_889 (O_889,N_19879,N_19424);
xor UO_890 (O_890,N_18675,N_16622);
nor UO_891 (O_891,N_16978,N_16384);
nor UO_892 (O_892,N_19532,N_17995);
nor UO_893 (O_893,N_17661,N_18424);
nor UO_894 (O_894,N_17565,N_16119);
or UO_895 (O_895,N_18211,N_18936);
nor UO_896 (O_896,N_17128,N_18095);
xor UO_897 (O_897,N_16711,N_16696);
or UO_898 (O_898,N_19721,N_18265);
and UO_899 (O_899,N_19890,N_18357);
nand UO_900 (O_900,N_18297,N_19324);
or UO_901 (O_901,N_18508,N_17731);
or UO_902 (O_902,N_17175,N_19371);
or UO_903 (O_903,N_19336,N_18133);
nor UO_904 (O_904,N_18087,N_17346);
or UO_905 (O_905,N_19474,N_18467);
or UO_906 (O_906,N_16910,N_19557);
nand UO_907 (O_907,N_17601,N_19603);
nor UO_908 (O_908,N_16363,N_19041);
nand UO_909 (O_909,N_16814,N_16133);
nor UO_910 (O_910,N_16616,N_17402);
nor UO_911 (O_911,N_17517,N_19077);
nand UO_912 (O_912,N_17295,N_16462);
nand UO_913 (O_913,N_19838,N_19787);
nand UO_914 (O_914,N_18412,N_19534);
or UO_915 (O_915,N_16176,N_18565);
or UO_916 (O_916,N_17926,N_17960);
and UO_917 (O_917,N_19433,N_16417);
and UO_918 (O_918,N_16140,N_18368);
nand UO_919 (O_919,N_18423,N_16594);
and UO_920 (O_920,N_17150,N_19313);
or UO_921 (O_921,N_18555,N_16528);
nand UO_922 (O_922,N_18848,N_18108);
xor UO_923 (O_923,N_17341,N_17748);
and UO_924 (O_924,N_17651,N_18134);
nand UO_925 (O_925,N_18252,N_16164);
nor UO_926 (O_926,N_18035,N_17077);
and UO_927 (O_927,N_18744,N_16597);
nand UO_928 (O_928,N_17286,N_19083);
or UO_929 (O_929,N_19950,N_19921);
nor UO_930 (O_930,N_19636,N_19748);
nor UO_931 (O_931,N_19449,N_17501);
and UO_932 (O_932,N_17277,N_16694);
xnor UO_933 (O_933,N_18277,N_17474);
nand UO_934 (O_934,N_17577,N_18716);
nor UO_935 (O_935,N_18434,N_17605);
nor UO_936 (O_936,N_19700,N_18447);
and UO_937 (O_937,N_18167,N_17301);
nand UO_938 (O_938,N_18928,N_18032);
and UO_939 (O_939,N_18349,N_18881);
and UO_940 (O_940,N_18233,N_18245);
nor UO_941 (O_941,N_19475,N_19074);
and UO_942 (O_942,N_16207,N_18031);
and UO_943 (O_943,N_18975,N_16481);
xnor UO_944 (O_944,N_18175,N_18075);
nand UO_945 (O_945,N_18747,N_18503);
and UO_946 (O_946,N_18030,N_16260);
xor UO_947 (O_947,N_17844,N_19902);
nand UO_948 (O_948,N_17931,N_19372);
or UO_949 (O_949,N_19501,N_17208);
nand UO_950 (O_950,N_19747,N_17082);
or UO_951 (O_951,N_17581,N_18369);
or UO_952 (O_952,N_17613,N_19991);
nor UO_953 (O_953,N_16145,N_17504);
and UO_954 (O_954,N_19250,N_18440);
and UO_955 (O_955,N_16829,N_19003);
and UO_956 (O_956,N_17299,N_19265);
or UO_957 (O_957,N_18460,N_16530);
nor UO_958 (O_958,N_16138,N_17935);
or UO_959 (O_959,N_19421,N_19753);
xor UO_960 (O_960,N_17360,N_17385);
nor UO_961 (O_961,N_18768,N_19846);
or UO_962 (O_962,N_16896,N_16764);
nand UO_963 (O_963,N_17349,N_17098);
and UO_964 (O_964,N_18522,N_16048);
and UO_965 (O_965,N_16298,N_18433);
and UO_966 (O_966,N_16582,N_17766);
nand UO_967 (O_967,N_18535,N_19339);
and UO_968 (O_968,N_18491,N_18755);
or UO_969 (O_969,N_17741,N_18967);
nand UO_970 (O_970,N_16346,N_17219);
xnor UO_971 (O_971,N_17895,N_18805);
and UO_972 (O_972,N_17041,N_19145);
xnor UO_973 (O_973,N_18920,N_17310);
or UO_974 (O_974,N_18495,N_19179);
nor UO_975 (O_975,N_16728,N_18937);
and UO_976 (O_976,N_17381,N_18015);
or UO_977 (O_977,N_19917,N_18355);
or UO_978 (O_978,N_17515,N_17168);
nand UO_979 (O_979,N_17627,N_19755);
or UO_980 (O_980,N_19741,N_18730);
or UO_981 (O_981,N_16553,N_18417);
or UO_982 (O_982,N_19252,N_19191);
nand UO_983 (O_983,N_17796,N_18282);
and UO_984 (O_984,N_19959,N_19599);
nand UO_985 (O_985,N_17378,N_18301);
or UO_986 (O_986,N_17084,N_18296);
nand UO_987 (O_987,N_18884,N_16817);
nand UO_988 (O_988,N_17562,N_17678);
or UO_989 (O_989,N_17543,N_16430);
nor UO_990 (O_990,N_16376,N_19353);
xor UO_991 (O_991,N_16490,N_17916);
or UO_992 (O_992,N_17789,N_16101);
nand UO_993 (O_993,N_16118,N_19254);
and UO_994 (O_994,N_19144,N_17658);
or UO_995 (O_995,N_17314,N_18330);
nand UO_996 (O_996,N_19167,N_16801);
nand UO_997 (O_997,N_19836,N_17177);
or UO_998 (O_998,N_17377,N_18347);
and UO_999 (O_999,N_16221,N_17584);
and UO_1000 (O_1000,N_17839,N_19954);
and UO_1001 (O_1001,N_18500,N_17257);
nor UO_1002 (O_1002,N_18910,N_19337);
and UO_1003 (O_1003,N_19204,N_16100);
nor UO_1004 (O_1004,N_19517,N_19942);
or UO_1005 (O_1005,N_18154,N_17328);
nand UO_1006 (O_1006,N_17979,N_19244);
nor UO_1007 (O_1007,N_17903,N_19169);
and UO_1008 (O_1008,N_17819,N_19623);
nor UO_1009 (O_1009,N_18042,N_16360);
nor UO_1010 (O_1010,N_19559,N_19280);
and UO_1011 (O_1011,N_19487,N_17929);
nor UO_1012 (O_1012,N_17137,N_19128);
nand UO_1013 (O_1013,N_18388,N_16186);
nand UO_1014 (O_1014,N_18734,N_19676);
nor UO_1015 (O_1015,N_19384,N_18912);
nand UO_1016 (O_1016,N_18081,N_16580);
nor UO_1017 (O_1017,N_17025,N_19422);
xor UO_1018 (O_1018,N_18987,N_17334);
nor UO_1019 (O_1019,N_19635,N_16211);
nand UO_1020 (O_1020,N_17650,N_17980);
nand UO_1021 (O_1021,N_19896,N_19804);
xnor UO_1022 (O_1022,N_18664,N_16546);
nand UO_1023 (O_1023,N_16628,N_16849);
nand UO_1024 (O_1024,N_17722,N_19444);
or UO_1025 (O_1025,N_19119,N_17056);
nand UO_1026 (O_1026,N_19166,N_16466);
or UO_1027 (O_1027,N_18021,N_18471);
nor UO_1028 (O_1028,N_19946,N_18915);
or UO_1029 (O_1029,N_16457,N_19383);
nand UO_1030 (O_1030,N_18120,N_18769);
or UO_1031 (O_1031,N_17318,N_19943);
xnor UO_1032 (O_1032,N_17502,N_17220);
nor UO_1033 (O_1033,N_17435,N_17968);
nor UO_1034 (O_1034,N_19958,N_18706);
nor UO_1035 (O_1035,N_18924,N_16822);
nor UO_1036 (O_1036,N_19020,N_17779);
or UO_1037 (O_1037,N_16432,N_16932);
nor UO_1038 (O_1038,N_17048,N_16547);
nor UO_1039 (O_1039,N_18432,N_19046);
xor UO_1040 (O_1040,N_19831,N_17550);
nor UO_1041 (O_1041,N_16707,N_16408);
and UO_1042 (O_1042,N_18335,N_17886);
nor UO_1043 (O_1043,N_19005,N_17269);
nand UO_1044 (O_1044,N_18648,N_17703);
nand UO_1045 (O_1045,N_18997,N_16327);
or UO_1046 (O_1046,N_19104,N_18900);
xnor UO_1047 (O_1047,N_17231,N_18002);
or UO_1048 (O_1048,N_18178,N_16136);
nand UO_1049 (O_1049,N_16900,N_19724);
nor UO_1050 (O_1050,N_18143,N_19772);
nand UO_1051 (O_1051,N_17039,N_18528);
and UO_1052 (O_1052,N_17242,N_18115);
or UO_1053 (O_1053,N_18099,N_18161);
nor UO_1054 (O_1054,N_18701,N_19279);
or UO_1055 (O_1055,N_18209,N_18718);
nand UO_1056 (O_1056,N_18394,N_16403);
nor UO_1057 (O_1057,N_16278,N_17851);
or UO_1058 (O_1058,N_19666,N_16020);
and UO_1059 (O_1059,N_18036,N_19953);
and UO_1060 (O_1060,N_17933,N_19416);
xor UO_1061 (O_1061,N_17027,N_17865);
or UO_1062 (O_1062,N_16886,N_16838);
nand UO_1063 (O_1063,N_18667,N_18908);
nor UO_1064 (O_1064,N_19240,N_16637);
and UO_1065 (O_1065,N_19869,N_16832);
and UO_1066 (O_1066,N_16713,N_18626);
nor UO_1067 (O_1067,N_16959,N_17466);
nor UO_1068 (O_1068,N_17409,N_18004);
and UO_1069 (O_1069,N_19385,N_17361);
or UO_1070 (O_1070,N_19225,N_17604);
nand UO_1071 (O_1071,N_16808,N_18579);
or UO_1072 (O_1072,N_17485,N_19578);
nand UO_1073 (O_1073,N_19634,N_16506);
and UO_1074 (O_1074,N_17694,N_16779);
xor UO_1075 (O_1075,N_17680,N_19268);
or UO_1076 (O_1076,N_16858,N_16311);
or UO_1077 (O_1077,N_17235,N_17677);
or UO_1078 (O_1078,N_19800,N_16192);
nor UO_1079 (O_1079,N_17574,N_18457);
and UO_1080 (O_1080,N_18397,N_16344);
nand UO_1081 (O_1081,N_18316,N_19105);
or UO_1082 (O_1082,N_19687,N_19386);
nand UO_1083 (O_1083,N_16987,N_18589);
nor UO_1084 (O_1084,N_19443,N_19256);
or UO_1085 (O_1085,N_16070,N_19715);
and UO_1086 (O_1086,N_16383,N_19955);
and UO_1087 (O_1087,N_18694,N_16805);
and UO_1088 (O_1088,N_19350,N_19469);
nor UO_1089 (O_1089,N_18959,N_16428);
nor UO_1090 (O_1090,N_19408,N_16566);
nand UO_1091 (O_1091,N_16611,N_19761);
and UO_1092 (O_1092,N_17161,N_16795);
and UO_1093 (O_1093,N_16960,N_18071);
and UO_1094 (O_1094,N_16784,N_18663);
nand UO_1095 (O_1095,N_19017,N_19331);
or UO_1096 (O_1096,N_19498,N_18009);
or UO_1097 (O_1097,N_18721,N_18041);
and UO_1098 (O_1098,N_18568,N_18818);
and UO_1099 (O_1099,N_18518,N_16772);
nand UO_1100 (O_1100,N_17260,N_16056);
nor UO_1101 (O_1101,N_16660,N_17159);
nor UO_1102 (O_1102,N_16862,N_17643);
nor UO_1103 (O_1103,N_16894,N_16543);
and UO_1104 (O_1104,N_19293,N_16812);
nor UO_1105 (O_1105,N_17905,N_18741);
nor UO_1106 (O_1106,N_18988,N_16928);
xor UO_1107 (O_1107,N_17155,N_18443);
nand UO_1108 (O_1108,N_17124,N_19116);
and UO_1109 (O_1109,N_18722,N_18985);
nor UO_1110 (O_1110,N_18184,N_17288);
and UO_1111 (O_1111,N_16625,N_18609);
nor UO_1112 (O_1112,N_19114,N_18387);
and UO_1113 (O_1113,N_17140,N_19935);
nand UO_1114 (O_1114,N_17194,N_17997);
xor UO_1115 (O_1115,N_16640,N_17742);
nand UO_1116 (O_1116,N_19561,N_19155);
or UO_1117 (O_1117,N_19199,N_19486);
nor UO_1118 (O_1118,N_18572,N_16055);
xor UO_1119 (O_1119,N_19132,N_17638);
nor UO_1120 (O_1120,N_17302,N_19867);
nand UO_1121 (O_1121,N_16915,N_17508);
or UO_1122 (O_1122,N_18325,N_19133);
and UO_1123 (O_1123,N_17516,N_18740);
and UO_1124 (O_1124,N_18415,N_19793);
nor UO_1125 (O_1125,N_18628,N_19263);
and UO_1126 (O_1126,N_16023,N_18124);
nor UO_1127 (O_1127,N_17279,N_18891);
or UO_1128 (O_1128,N_17395,N_17443);
and UO_1129 (O_1129,N_19894,N_17390);
nor UO_1130 (O_1130,N_18047,N_19999);
and UO_1131 (O_1131,N_18946,N_18016);
nor UO_1132 (O_1132,N_19875,N_16912);
nor UO_1133 (O_1133,N_17771,N_16395);
and UO_1134 (O_1134,N_17913,N_19963);
and UO_1135 (O_1135,N_18493,N_19373);
nand UO_1136 (O_1136,N_17416,N_18674);
or UO_1137 (O_1137,N_18225,N_16299);
or UO_1138 (O_1138,N_16057,N_16382);
and UO_1139 (O_1139,N_18149,N_16804);
nand UO_1140 (O_1140,N_16755,N_18971);
nand UO_1141 (O_1141,N_16475,N_18652);
and UO_1142 (O_1142,N_17602,N_16124);
nand UO_1143 (O_1143,N_17590,N_18536);
or UO_1144 (O_1144,N_17248,N_17181);
nand UO_1145 (O_1145,N_17711,N_18102);
and UO_1146 (O_1146,N_16931,N_18089);
xor UO_1147 (O_1147,N_17074,N_17358);
nor UO_1148 (O_1148,N_16050,N_17379);
nor UO_1149 (O_1149,N_16281,N_16914);
or UO_1150 (O_1150,N_18264,N_16397);
and UO_1151 (O_1151,N_16305,N_17174);
nor UO_1152 (O_1152,N_19160,N_18551);
or UO_1153 (O_1153,N_17021,N_19154);
and UO_1154 (O_1154,N_16935,N_19794);
nor UO_1155 (O_1155,N_16678,N_17332);
or UO_1156 (O_1156,N_17394,N_17011);
and UO_1157 (O_1157,N_18511,N_19805);
nor UO_1158 (O_1158,N_19556,N_18925);
xnor UO_1159 (O_1159,N_17837,N_17210);
and UO_1160 (O_1160,N_17666,N_18411);
xor UO_1161 (O_1161,N_16480,N_17842);
and UO_1162 (O_1162,N_16605,N_19572);
and UO_1163 (O_1163,N_19334,N_19333);
or UO_1164 (O_1164,N_18728,N_18875);
or UO_1165 (O_1165,N_16623,N_19533);
and UO_1166 (O_1166,N_16392,N_19451);
nor UO_1167 (O_1167,N_17195,N_19866);
nand UO_1168 (O_1168,N_18000,N_16043);
nand UO_1169 (O_1169,N_17193,N_17476);
nor UO_1170 (O_1170,N_16355,N_19376);
nand UO_1171 (O_1171,N_18821,N_17032);
and UO_1172 (O_1172,N_18266,N_18384);
and UO_1173 (O_1173,N_17298,N_16353);
nor UO_1174 (O_1174,N_19374,N_19492);
nor UO_1175 (O_1175,N_18236,N_19272);
or UO_1176 (O_1176,N_17892,N_17213);
nor UO_1177 (O_1177,N_19407,N_17521);
nor UO_1178 (O_1178,N_16830,N_17093);
nor UO_1179 (O_1179,N_19845,N_16312);
nand UO_1180 (O_1180,N_17042,N_17639);
and UO_1181 (O_1181,N_18546,N_17717);
nor UO_1182 (O_1182,N_18870,N_17679);
nor UO_1183 (O_1183,N_19591,N_18287);
and UO_1184 (O_1184,N_19493,N_19697);
nor UO_1185 (O_1185,N_19147,N_19689);
nand UO_1186 (O_1186,N_16240,N_16796);
and UO_1187 (O_1187,N_18220,N_17646);
nor UO_1188 (O_1188,N_18835,N_17489);
or UO_1189 (O_1189,N_16957,N_17705);
nand UO_1190 (O_1190,N_17136,N_19779);
nor UO_1191 (O_1191,N_19288,N_17908);
nand UO_1192 (O_1192,N_18014,N_18684);
or UO_1193 (O_1193,N_17806,N_18405);
nand UO_1194 (O_1194,N_18269,N_19363);
or UO_1195 (O_1195,N_17692,N_16505);
nand UO_1196 (O_1196,N_17507,N_18760);
and UO_1197 (O_1197,N_16235,N_16966);
nand UO_1198 (O_1198,N_16095,N_17735);
xor UO_1199 (O_1199,N_17737,N_19877);
or UO_1200 (O_1200,N_18844,N_18562);
and UO_1201 (O_1201,N_16961,N_18861);
nor UO_1202 (O_1202,N_16026,N_17909);
xnor UO_1203 (O_1203,N_19295,N_19246);
or UO_1204 (O_1204,N_19347,N_19266);
or UO_1205 (O_1205,N_17382,N_16289);
nand UO_1206 (O_1206,N_18311,N_17773);
nand UO_1207 (O_1207,N_19184,N_16704);
nor UO_1208 (O_1208,N_16734,N_19997);
and UO_1209 (O_1209,N_19798,N_16828);
and UO_1210 (O_1210,N_17561,N_17553);
nand UO_1211 (O_1211,N_18043,N_16190);
nor UO_1212 (O_1212,N_16749,N_16498);
or UO_1213 (O_1213,N_18930,N_16555);
nor UO_1214 (O_1214,N_18428,N_17281);
nand UO_1215 (O_1215,N_19508,N_19718);
nand UO_1216 (O_1216,N_19971,N_19996);
or UO_1217 (O_1217,N_16017,N_16156);
nor UO_1218 (O_1218,N_19340,N_16229);
or UO_1219 (O_1219,N_19216,N_19043);
nor UO_1220 (O_1220,N_18934,N_16246);
or UO_1221 (O_1221,N_19394,N_19673);
and UO_1222 (O_1222,N_17768,N_18012);
and UO_1223 (O_1223,N_16484,N_19348);
nor UO_1224 (O_1224,N_17216,N_19763);
nor UO_1225 (O_1225,N_18230,N_19176);
nand UO_1226 (O_1226,N_19024,N_16036);
nand UO_1227 (O_1227,N_16454,N_19122);
nor UO_1228 (O_1228,N_17663,N_16223);
or UO_1229 (O_1229,N_17975,N_18829);
and UO_1230 (O_1230,N_16052,N_17464);
nand UO_1231 (O_1231,N_19370,N_19500);
and UO_1232 (O_1232,N_16765,N_16200);
nand UO_1233 (O_1233,N_16396,N_19895);
xor UO_1234 (O_1234,N_19239,N_16545);
and UO_1235 (O_1235,N_16436,N_19832);
and UO_1236 (O_1236,N_19210,N_18398);
nand UO_1237 (O_1237,N_16439,N_17122);
nand UO_1238 (O_1238,N_18525,N_19013);
nand UO_1239 (O_1239,N_18308,N_18166);
and UO_1240 (O_1240,N_19377,N_16158);
and UO_1241 (O_1241,N_19939,N_16871);
and UO_1242 (O_1242,N_18880,N_17094);
nand UO_1243 (O_1243,N_18871,N_16309);
or UO_1244 (O_1244,N_16351,N_19605);
and UO_1245 (O_1245,N_18713,N_19998);
or UO_1246 (O_1246,N_16982,N_19380);
and UO_1247 (O_1247,N_16467,N_16139);
nor UO_1248 (O_1248,N_19515,N_19987);
nand UO_1249 (O_1249,N_17058,N_19906);
and UO_1250 (O_1250,N_17648,N_17384);
xor UO_1251 (O_1251,N_19551,N_19688);
nand UO_1252 (O_1252,N_19612,N_16698);
nand UO_1253 (O_1253,N_18109,N_16841);
nand UO_1254 (O_1254,N_17615,N_17890);
nand UO_1255 (O_1255,N_17066,N_17183);
or UO_1256 (O_1256,N_18815,N_18306);
and UO_1257 (O_1257,N_16816,N_19190);
nand UO_1258 (O_1258,N_18027,N_19448);
xor UO_1259 (O_1259,N_18376,N_16921);
nand UO_1260 (O_1260,N_16581,N_16319);
nand UO_1261 (O_1261,N_16686,N_17330);
nor UO_1262 (O_1262,N_19029,N_18828);
xnor UO_1263 (O_1263,N_19563,N_18795);
and UO_1264 (O_1264,N_17558,N_18853);
or UO_1265 (O_1265,N_17154,N_19081);
and UO_1266 (O_1266,N_19398,N_16619);
nand UO_1267 (O_1267,N_16649,N_19744);
nand UO_1268 (O_1268,N_16687,N_17463);
or UO_1269 (O_1269,N_19200,N_16116);
nor UO_1270 (O_1270,N_19341,N_16593);
nor UO_1271 (O_1271,N_19427,N_19011);
and UO_1272 (O_1272,N_18259,N_17961);
and UO_1273 (O_1273,N_16178,N_17452);
and UO_1274 (O_1274,N_16131,N_16671);
nand UO_1275 (O_1275,N_19530,N_16991);
xor UO_1276 (O_1276,N_17826,N_16168);
nor UO_1277 (O_1277,N_19611,N_17203);
or UO_1278 (O_1278,N_16364,N_19277);
nand UO_1279 (O_1279,N_17426,N_17914);
xor UO_1280 (O_1280,N_18614,N_19661);
nor UO_1281 (O_1281,N_18066,N_17354);
xor UO_1282 (O_1282,N_17750,N_16976);
and UO_1283 (O_1283,N_16415,N_17173);
and UO_1284 (O_1284,N_18153,N_17264);
and UO_1285 (O_1285,N_16197,N_19750);
nand UO_1286 (O_1286,N_16563,N_17369);
nor UO_1287 (O_1287,N_16173,N_16143);
nand UO_1288 (O_1288,N_19343,N_17191);
or UO_1289 (O_1289,N_17828,N_17064);
nand UO_1290 (O_1290,N_16379,N_16554);
or UO_1291 (O_1291,N_18992,N_16180);
nand UO_1292 (O_1292,N_18590,N_17371);
xnor UO_1293 (O_1293,N_18144,N_17572);
or UO_1294 (O_1294,N_17727,N_19976);
and UO_1295 (O_1295,N_17134,N_17053);
or UO_1296 (O_1296,N_19702,N_18226);
nand UO_1297 (O_1297,N_18343,N_18291);
or UO_1298 (O_1298,N_16372,N_17018);
nand UO_1299 (O_1299,N_17444,N_18899);
xnor UO_1300 (O_1300,N_19234,N_17372);
and UO_1301 (O_1301,N_17190,N_16314);
xor UO_1302 (O_1302,N_16609,N_17471);
and UO_1303 (O_1303,N_16587,N_19737);
nor UO_1304 (O_1304,N_18272,N_17862);
and UO_1305 (O_1305,N_18450,N_17043);
and UO_1306 (O_1306,N_19171,N_18904);
nand UO_1307 (O_1307,N_17326,N_19224);
or UO_1308 (O_1308,N_19765,N_17319);
xnor UO_1309 (O_1309,N_17306,N_19205);
nand UO_1310 (O_1310,N_17618,N_18235);
nand UO_1311 (O_1311,N_16072,N_16774);
or UO_1312 (O_1312,N_18557,N_17364);
or UO_1313 (O_1313,N_18607,N_16231);
and UO_1314 (O_1314,N_19792,N_18130);
xor UO_1315 (O_1315,N_18458,N_16034);
nor UO_1316 (O_1316,N_18761,N_18490);
nor UO_1317 (O_1317,N_17761,N_19522);
nor UO_1318 (O_1318,N_18459,N_16424);
or UO_1319 (O_1319,N_16901,N_18430);
or UO_1320 (O_1320,N_16220,N_16598);
nand UO_1321 (O_1321,N_18346,N_16468);
xor UO_1322 (O_1322,N_16989,N_19078);
nand UO_1323 (O_1323,N_16600,N_18796);
nor UO_1324 (O_1324,N_17237,N_16419);
or UO_1325 (O_1325,N_18206,N_16655);
nand UO_1326 (O_1326,N_16608,N_19817);
and UO_1327 (O_1327,N_18773,N_17670);
nand UO_1328 (O_1328,N_17883,N_18427);
nor UO_1329 (O_1329,N_19686,N_19218);
nand UO_1330 (O_1330,N_18514,N_19574);
or UO_1331 (O_1331,N_19219,N_19018);
nor UO_1332 (O_1332,N_16746,N_19418);
nand UO_1333 (O_1333,N_16798,N_19682);
nor UO_1334 (O_1334,N_17864,N_19413);
and UO_1335 (O_1335,N_17539,N_19525);
xnor UO_1336 (O_1336,N_18314,N_18765);
nor UO_1337 (O_1337,N_17455,N_17566);
nor UO_1338 (O_1338,N_16478,N_19618);
nor UO_1339 (O_1339,N_16226,N_18516);
nor UO_1340 (O_1340,N_17151,N_16491);
or UO_1341 (O_1341,N_17047,N_16531);
and UO_1342 (O_1342,N_16998,N_18309);
or UO_1343 (O_1343,N_18152,N_17925);
or UO_1344 (O_1344,N_19722,N_16732);
nand UO_1345 (O_1345,N_19242,N_16512);
and UO_1346 (O_1346,N_16895,N_19441);
or UO_1347 (O_1347,N_18944,N_17003);
nand UO_1348 (O_1348,N_16648,N_18157);
or UO_1349 (O_1349,N_18693,N_18135);
nand UO_1350 (O_1350,N_17896,N_18682);
xor UO_1351 (O_1351,N_19915,N_18976);
nor UO_1352 (O_1352,N_19813,N_18680);
and UO_1353 (O_1353,N_16464,N_18137);
or UO_1354 (O_1354,N_17568,N_19849);
xor UO_1355 (O_1355,N_17017,N_18407);
nor UO_1356 (O_1356,N_18735,N_16483);
or UO_1357 (O_1357,N_18647,N_19485);
and UO_1358 (O_1358,N_17492,N_17481);
or UO_1359 (O_1359,N_19652,N_16429);
nand UO_1360 (O_1360,N_16548,N_16150);
nand UO_1361 (O_1361,N_16474,N_19647);
and UO_1362 (O_1362,N_18359,N_16296);
or UO_1363 (O_1363,N_16799,N_17447);
or UO_1364 (O_1364,N_16310,N_18927);
nor UO_1365 (O_1365,N_19790,N_18673);
nand UO_1366 (O_1366,N_16179,N_17146);
or UO_1367 (O_1367,N_16267,N_16280);
nor UO_1368 (O_1368,N_16024,N_19213);
and UO_1369 (O_1369,N_17152,N_18627);
and UO_1370 (O_1370,N_18540,N_16859);
nor UO_1371 (O_1371,N_18659,N_16471);
or UO_1372 (O_1372,N_18616,N_16209);
and UO_1373 (O_1373,N_19503,N_18690);
and UO_1374 (O_1374,N_16297,N_17112);
nand UO_1375 (O_1375,N_19740,N_16174);
xnor UO_1376 (O_1376,N_16087,N_19773);
xor UO_1377 (O_1377,N_18634,N_16358);
xor UO_1378 (O_1378,N_18641,N_19786);
nor UO_1379 (O_1379,N_17548,N_17919);
nor UO_1380 (O_1380,N_18299,N_18736);
nand UO_1381 (O_1381,N_16950,N_19471);
and UO_1382 (O_1382,N_17518,N_18521);
and UO_1383 (O_1383,N_17877,N_16455);
nor UO_1384 (O_1384,N_19837,N_16066);
and UO_1385 (O_1385,N_16664,N_17387);
and UO_1386 (O_1386,N_18872,N_16709);
xnor UO_1387 (O_1387,N_18217,N_16522);
xnor UO_1388 (O_1388,N_16647,N_17251);
nor UO_1389 (O_1389,N_16905,N_16411);
or UO_1390 (O_1390,N_17162,N_19461);
and UO_1391 (O_1391,N_16747,N_16890);
xnor UO_1392 (O_1392,N_17889,N_16472);
or UO_1393 (O_1393,N_16249,N_19738);
and UO_1394 (O_1394,N_18655,N_17262);
nor UO_1395 (O_1395,N_18913,N_17775);
and UO_1396 (O_1396,N_19322,N_16320);
xor UO_1397 (O_1397,N_16216,N_16210);
nor UO_1398 (O_1398,N_17868,N_16783);
nor UO_1399 (O_1399,N_19857,N_16294);
nor UO_1400 (O_1400,N_16387,N_17963);
or UO_1401 (O_1401,N_16013,N_19202);
nor UO_1402 (O_1402,N_16636,N_17524);
nor UO_1403 (O_1403,N_18185,N_18037);
xor UO_1404 (O_1404,N_18566,N_19289);
and UO_1405 (O_1405,N_16159,N_18686);
nor UO_1406 (O_1406,N_16624,N_17598);
xnor UO_1407 (O_1407,N_17113,N_17544);
nor UO_1408 (O_1408,N_19069,N_16341);
nand UO_1409 (O_1409,N_16714,N_17142);
nand UO_1410 (O_1410,N_16590,N_17825);
nand UO_1411 (O_1411,N_17040,N_17403);
or UO_1412 (O_1412,N_16206,N_18856);
and UO_1413 (O_1413,N_19025,N_18507);
nand UO_1414 (O_1414,N_16751,N_19745);
nand UO_1415 (O_1415,N_16690,N_17852);
nor UO_1416 (O_1416,N_18026,N_18241);
nor UO_1417 (O_1417,N_16389,N_16287);
or UO_1418 (O_1418,N_16270,N_18635);
or UO_1419 (O_1419,N_16038,N_16324);
nand UO_1420 (O_1420,N_17186,N_16031);
nor UO_1421 (O_1421,N_16573,N_19291);
nor UO_1422 (O_1422,N_17947,N_17333);
and UO_1423 (O_1423,N_18895,N_17612);
and UO_1424 (O_1424,N_19819,N_18599);
and UO_1425 (O_1425,N_19914,N_16740);
and UO_1426 (O_1426,N_18380,N_16256);
nand UO_1427 (O_1427,N_18605,N_16639);
and UO_1428 (O_1428,N_19844,N_17863);
xor UO_1429 (O_1429,N_19106,N_16927);
and UO_1430 (O_1430,N_17461,N_18410);
or UO_1431 (O_1431,N_16981,N_19016);
nand UO_1432 (O_1432,N_16811,N_16028);
or UO_1433 (O_1433,N_16167,N_18559);
nor UO_1434 (O_1434,N_18748,N_16018);
and UO_1435 (O_1435,N_19073,N_16385);
and UO_1436 (O_1436,N_17969,N_16277);
and UO_1437 (O_1437,N_17080,N_17797);
nor UO_1438 (O_1438,N_16177,N_17739);
xor UO_1439 (O_1439,N_18839,N_16951);
and UO_1440 (O_1440,N_17659,N_17623);
nor UO_1441 (O_1441,N_16493,N_16227);
nand UO_1442 (O_1442,N_18426,N_17412);
or UO_1443 (O_1443,N_19473,N_17987);
and UO_1444 (O_1444,N_16269,N_19111);
and UO_1445 (O_1445,N_17276,N_16357);
or UO_1446 (O_1446,N_17738,N_18404);
or UO_1447 (O_1447,N_19063,N_16863);
and UO_1448 (O_1448,N_17964,N_19455);
nor UO_1449 (O_1449,N_18849,N_16924);
nor UO_1450 (O_1450,N_17484,N_18229);
or UO_1451 (O_1451,N_16247,N_17924);
or UO_1452 (O_1452,N_16949,N_18378);
or UO_1453 (O_1453,N_19127,N_17549);
xnor UO_1454 (O_1454,N_17641,N_16948);
xnor UO_1455 (O_1455,N_16098,N_18126);
nor UO_1456 (O_1456,N_16879,N_18782);
nand UO_1457 (O_1457,N_17215,N_19733);
or UO_1458 (O_1458,N_17976,N_16617);
nand UO_1459 (O_1459,N_18777,N_19303);
and UO_1460 (O_1460,N_18887,N_18464);
xnor UO_1461 (O_1461,N_16193,N_17948);
nand UO_1462 (O_1462,N_19978,N_19417);
nand UO_1463 (O_1463,N_19929,N_19299);
nor UO_1464 (O_1464,N_18750,N_19571);
xnor UO_1465 (O_1465,N_17787,N_19270);
or UO_1466 (O_1466,N_19004,N_19965);
xnor UO_1467 (O_1467,N_18898,N_17424);
nand UO_1468 (O_1468,N_17212,N_19311);
nor UO_1469 (O_1469,N_18653,N_19298);
and UO_1470 (O_1470,N_17527,N_19509);
nand UO_1471 (O_1471,N_18745,N_19640);
nor UO_1472 (O_1472,N_18024,N_18362);
and UO_1473 (O_1473,N_16109,N_17998);
nand UO_1474 (O_1474,N_16224,N_18510);
and UO_1475 (O_1475,N_19897,N_18544);
nand UO_1476 (O_1476,N_18505,N_16032);
nor UO_1477 (O_1477,N_16934,N_19535);
or UO_1478 (O_1478,N_17875,N_18833);
nand UO_1479 (O_1479,N_17256,N_17209);
or UO_1480 (O_1480,N_18305,N_18819);
nor UO_1481 (O_1481,N_18364,N_16354);
nor UO_1482 (O_1482,N_19691,N_19332);
or UO_1483 (O_1483,N_18611,N_16821);
xor UO_1484 (O_1484,N_17901,N_19856);
nor UO_1485 (O_1485,N_19862,N_16393);
and UO_1486 (O_1486,N_16163,N_18669);
or UO_1487 (O_1487,N_19910,N_16264);
nand UO_1488 (O_1488,N_17970,N_18534);
or UO_1489 (O_1489,N_19990,N_17014);
or UO_1490 (O_1490,N_16807,N_17593);
nand UO_1491 (O_1491,N_16012,N_18571);
nand UO_1492 (O_1492,N_17686,N_18200);
or UO_1493 (O_1493,N_16494,N_16627);
or UO_1494 (O_1494,N_19012,N_17850);
nand UO_1495 (O_1495,N_18215,N_17055);
nor UO_1496 (O_1496,N_19608,N_18074);
nor UO_1497 (O_1497,N_17482,N_16248);
and UO_1498 (O_1498,N_18093,N_18340);
or UO_1499 (O_1499,N_16567,N_17915);
and UO_1500 (O_1500,N_16286,N_16495);
nand UO_1501 (O_1501,N_17289,N_16902);
and UO_1502 (O_1502,N_16502,N_18170);
nor UO_1503 (O_1503,N_18466,N_19045);
xor UO_1504 (O_1504,N_19459,N_17551);
and UO_1505 (O_1505,N_16414,N_18365);
or UO_1506 (O_1506,N_19307,N_17767);
nand UO_1507 (O_1507,N_16542,N_17396);
nor UO_1508 (O_1508,N_18051,N_16945);
and UO_1509 (O_1509,N_16337,N_16653);
xnor UO_1510 (O_1510,N_18292,N_17695);
nor UO_1511 (O_1511,N_16958,N_18307);
nor UO_1512 (O_1512,N_17496,N_17130);
and UO_1513 (O_1513,N_19562,N_17799);
and UO_1514 (O_1514,N_16074,N_18643);
xnor UO_1515 (O_1515,N_19062,N_18917);
and UO_1516 (O_1516,N_19808,N_18619);
nor UO_1517 (O_1517,N_16485,N_16839);
nand UO_1518 (O_1518,N_19165,N_18896);
or UO_1519 (O_1519,N_18334,N_18515);
nor UO_1520 (O_1520,N_16526,N_19796);
and UO_1521 (O_1521,N_16111,N_17392);
and UO_1522 (O_1522,N_17855,N_18381);
and UO_1523 (O_1523,N_16572,N_18361);
xnor UO_1524 (O_1524,N_18336,N_18788);
nand UO_1525 (O_1525,N_17232,N_17597);
or UO_1526 (O_1526,N_16963,N_16195);
xnor UO_1527 (O_1527,N_17817,N_17757);
and UO_1528 (O_1528,N_17067,N_19751);
nor UO_1529 (O_1529,N_19980,N_17664);
or UO_1530 (O_1530,N_17534,N_19729);
and UO_1531 (O_1531,N_18121,N_18195);
and UO_1532 (O_1532,N_16668,N_17439);
or UO_1533 (O_1533,N_17536,N_18203);
nand UO_1534 (O_1534,N_16409,N_16994);
nand UO_1535 (O_1535,N_19379,N_19756);
nor UO_1536 (O_1536,N_16237,N_17229);
and UO_1537 (O_1537,N_19173,N_18502);
or UO_1538 (O_1538,N_17569,N_19496);
nand UO_1539 (O_1539,N_17540,N_18822);
nand UO_1540 (O_1540,N_19488,N_19727);
xor UO_1541 (O_1541,N_19053,N_18111);
nor UO_1542 (O_1542,N_18685,N_17822);
or UO_1543 (O_1543,N_18142,N_19835);
and UO_1544 (O_1544,N_18084,N_18392);
nor UO_1545 (O_1545,N_19107,N_17776);
nor UO_1546 (O_1546,N_17708,N_19818);
xnor UO_1547 (O_1547,N_19163,N_19301);
nor UO_1548 (O_1548,N_17405,N_16307);
and UO_1549 (O_1549,N_16513,N_16045);
xnor UO_1550 (O_1550,N_18168,N_18377);
nand UO_1551 (O_1551,N_16800,N_17063);
nand UO_1552 (O_1552,N_16134,N_19927);
or UO_1553 (O_1553,N_18290,N_18456);
and UO_1554 (O_1554,N_17682,N_19259);
xor UO_1555 (O_1555,N_19406,N_19314);
and UO_1556 (O_1556,N_16318,N_16401);
nor UO_1557 (O_1557,N_16988,N_18749);
and UO_1558 (O_1558,N_18504,N_19780);
and UO_1559 (O_1559,N_17044,N_17059);
nand UO_1560 (O_1560,N_19352,N_16964);
nand UO_1561 (O_1561,N_18022,N_19453);
nor UO_1562 (O_1562,N_18105,N_16450);
xnor UO_1563 (O_1563,N_17268,N_18890);
xor UO_1564 (O_1564,N_19593,N_19683);
and UO_1565 (O_1565,N_17092,N_16000);
nand UO_1566 (O_1566,N_16427,N_17234);
or UO_1567 (O_1567,N_17344,N_17592);
nand UO_1568 (O_1568,N_18255,N_19725);
nand UO_1569 (O_1569,N_18933,N_19696);
and UO_1570 (O_1570,N_17069,N_18077);
nor UO_1571 (O_1571,N_16239,N_16979);
xnor UO_1572 (O_1572,N_16137,N_18785);
nor UO_1573 (O_1573,N_19518,N_17993);
nor UO_1574 (O_1574,N_18214,N_17170);
nand UO_1575 (O_1575,N_19732,N_19622);
or UO_1576 (O_1576,N_16191,N_17284);
nand UO_1577 (O_1577,N_18372,N_16284);
or UO_1578 (O_1578,N_19539,N_16037);
nor UO_1579 (O_1579,N_19573,N_19007);
or UO_1580 (O_1580,N_18072,N_16273);
or UO_1581 (O_1581,N_18489,N_18101);
and UO_1582 (O_1582,N_17287,N_18697);
and UO_1583 (O_1583,N_18837,N_17972);
nor UO_1584 (O_1584,N_19193,N_19100);
or UO_1585 (O_1585,N_19768,N_17872);
nand UO_1586 (O_1586,N_16377,N_19065);
and UO_1587 (O_1587,N_18994,N_16835);
nor UO_1588 (O_1588,N_16250,N_18852);
or UO_1589 (O_1589,N_19615,N_19812);
and UO_1590 (O_1590,N_19170,N_16473);
or UO_1591 (O_1591,N_16983,N_16352);
nor UO_1592 (O_1592,N_18983,N_17907);
or UO_1593 (O_1593,N_18478,N_18843);
nor UO_1594 (O_1594,N_18638,N_18732);
nand UO_1595 (O_1595,N_16685,N_17885);
and UO_1596 (O_1596,N_19680,N_17462);
nor UO_1597 (O_1597,N_16658,N_17085);
and UO_1598 (O_1598,N_17983,N_17609);
nor UO_1599 (O_1599,N_19870,N_17812);
nor UO_1600 (O_1600,N_17148,N_17784);
or UO_1601 (O_1601,N_19002,N_16265);
nor UO_1602 (O_1602,N_18973,N_18811);
nand UO_1603 (O_1603,N_17240,N_19707);
and UO_1604 (O_1604,N_17591,N_17307);
and UO_1605 (O_1605,N_16955,N_17132);
nor UO_1606 (O_1606,N_17335,N_17324);
nor UO_1607 (O_1607,N_16039,N_18326);
nor UO_1608 (O_1608,N_17199,N_16585);
or UO_1609 (O_1609,N_18366,N_17545);
nor UO_1610 (O_1610,N_17370,N_17249);
xnor UO_1611 (O_1611,N_17415,N_19620);
xor UO_1612 (O_1612,N_18825,N_17537);
xnor UO_1613 (O_1613,N_18098,N_16614);
xor UO_1614 (O_1614,N_17054,N_16938);
or UO_1615 (O_1615,N_17296,N_16361);
nand UO_1616 (O_1616,N_16067,N_16285);
and UO_1617 (O_1617,N_18317,N_19695);
nand UO_1618 (O_1618,N_16692,N_16198);
and UO_1619 (O_1619,N_18088,N_16262);
nand UO_1620 (O_1620,N_16777,N_17576);
xor UO_1621 (O_1621,N_17051,N_17157);
nand UO_1622 (O_1622,N_17902,N_19066);
nor UO_1623 (O_1623,N_19589,N_17449);
nand UO_1624 (O_1624,N_16426,N_17904);
nand UO_1625 (O_1625,N_18257,N_19749);
nand UO_1626 (O_1626,N_17167,N_16695);
or UO_1627 (O_1627,N_18563,N_17547);
nor UO_1628 (O_1628,N_17934,N_19323);
nand UO_1629 (O_1629,N_19801,N_19101);
nor UO_1630 (O_1630,N_16062,N_19241);
or UO_1631 (O_1631,N_16487,N_17723);
nand UO_1632 (O_1632,N_19614,N_16188);
nand UO_1633 (O_1633,N_18698,N_16794);
xor UO_1634 (O_1634,N_16033,N_17029);
or UO_1635 (O_1635,N_19712,N_19549);
nand UO_1636 (O_1636,N_17759,N_17725);
nor UO_1637 (O_1637,N_18633,N_17782);
nor UO_1638 (O_1638,N_17164,N_19273);
nand UO_1639 (O_1639,N_18329,N_17355);
nor UO_1640 (O_1640,N_16049,N_16880);
nand UO_1641 (O_1641,N_16727,N_17202);
nor UO_1642 (O_1642,N_17368,N_17294);
or UO_1643 (O_1643,N_17187,N_16465);
nor UO_1644 (O_1644,N_19136,N_19283);
nand UO_1645 (O_1645,N_17673,N_18957);
nand UO_1646 (O_1646,N_18151,N_19995);
and UO_1647 (O_1647,N_19260,N_16093);
and UO_1648 (O_1648,N_16157,N_17030);
nor UO_1649 (O_1649,N_18786,N_16065);
or UO_1650 (O_1650,N_19023,N_19438);
and UO_1651 (O_1651,N_18541,N_18958);
nor UO_1652 (O_1652,N_16486,N_17586);
nand UO_1653 (O_1653,N_19316,N_16852);
nor UO_1654 (O_1654,N_19251,N_16470);
nor UO_1655 (O_1655,N_19243,N_16860);
or UO_1656 (O_1656,N_19597,N_18549);
or UO_1657 (O_1657,N_18509,N_17793);
xnor UO_1658 (O_1658,N_17835,N_18267);
xor UO_1659 (O_1659,N_19985,N_17519);
and UO_1660 (O_1660,N_17380,N_17052);
and UO_1661 (O_1661,N_18864,N_19276);
nor UO_1662 (O_1662,N_16523,N_16082);
nor UO_1663 (O_1663,N_16079,N_17376);
or UO_1664 (O_1664,N_19660,N_18586);
nor UO_1665 (O_1665,N_17007,N_16329);
nand UO_1666 (O_1666,N_18221,N_18877);
and UO_1667 (O_1667,N_19038,N_17458);
nor UO_1668 (O_1668,N_19723,N_16675);
xor UO_1669 (O_1669,N_18114,N_16316);
or UO_1670 (O_1670,N_17874,N_18273);
and UO_1671 (O_1671,N_17340,N_18962);
nor UO_1672 (O_1672,N_17325,N_18360);
nand UO_1673 (O_1673,N_19366,N_19212);
and UO_1674 (O_1674,N_18446,N_16645);
and UO_1675 (O_1675,N_16042,N_19923);
xnor UO_1676 (O_1676,N_19630,N_17849);
and UO_1677 (O_1677,N_19208,N_18778);
or UO_1678 (O_1678,N_17542,N_18281);
and UO_1679 (O_1679,N_17830,N_17454);
nand UO_1680 (O_1680,N_19080,N_17633);
and UO_1681 (O_1681,N_17918,N_18302);
nand UO_1682 (O_1682,N_18606,N_19188);
nor UO_1683 (O_1683,N_19945,N_19546);
or UO_1684 (O_1684,N_18993,N_16715);
nand UO_1685 (O_1685,N_17271,N_17024);
nand UO_1686 (O_1686,N_19203,N_19365);
and UO_1687 (O_1687,N_17967,N_17460);
nor UO_1688 (O_1688,N_18986,N_19662);
nand UO_1689 (O_1689,N_18729,N_17856);
xor UO_1690 (O_1690,N_18148,N_19115);
or UO_1691 (O_1691,N_19735,N_17791);
nand UO_1692 (O_1692,N_19674,N_16679);
or UO_1693 (O_1693,N_18513,N_16899);
and UO_1694 (O_1694,N_17556,N_18939);
nand UO_1695 (O_1695,N_19030,N_18512);
and UO_1696 (O_1696,N_16149,N_17407);
or UO_1697 (O_1697,N_16215,N_18567);
nor UO_1698 (O_1698,N_17428,N_16084);
xor UO_1699 (O_1699,N_18622,N_18951);
nand UO_1700 (O_1700,N_17425,N_17273);
nand UO_1701 (O_1701,N_19629,N_16245);
or UO_1702 (O_1702,N_18704,N_17873);
and UO_1703 (O_1703,N_19378,N_16080);
xnor UO_1704 (O_1704,N_18164,N_18462);
nor UO_1705 (O_1705,N_18956,N_16183);
xnor UO_1706 (O_1706,N_18396,N_17672);
and UO_1707 (O_1707,N_16557,N_16809);
nand UO_1708 (O_1708,N_18049,N_16985);
nand UO_1709 (O_1709,N_17922,N_16676);
and UO_1710 (O_1710,N_19864,N_16682);
nor UO_1711 (O_1711,N_18797,N_17938);
nand UO_1712 (O_1712,N_17126,N_17026);
and UO_1713 (O_1713,N_19626,N_16476);
nand UO_1714 (O_1714,N_16144,N_18772);
or UO_1715 (O_1715,N_16236,N_16710);
or UO_1716 (O_1716,N_18011,N_16898);
nor UO_1717 (O_1717,N_18707,N_19570);
xor UO_1718 (O_1718,N_17457,N_16781);
and UO_1719 (O_1719,N_16141,N_16090);
nor UO_1720 (O_1720,N_16703,N_19095);
nand UO_1721 (O_1721,N_16946,N_17263);
or UO_1722 (O_1722,N_16444,N_18604);
and UO_1723 (O_1723,N_19368,N_19633);
nand UO_1724 (O_1724,N_17445,N_19446);
and UO_1725 (O_1725,N_19454,N_19824);
nand UO_1726 (O_1726,N_18246,N_18332);
nor UO_1727 (O_1727,N_18063,N_17070);
nand UO_1728 (O_1728,N_17732,N_16893);
nand UO_1729 (O_1729,N_17888,N_19481);
or UO_1730 (O_1730,N_17477,N_18313);
nor UO_1731 (O_1731,N_16536,N_19528);
and UO_1732 (O_1732,N_17941,N_16407);
or UO_1733 (O_1733,N_18874,N_16181);
xnor UO_1734 (O_1734,N_18756,N_18243);
or UO_1735 (O_1735,N_17228,N_17840);
nor UO_1736 (O_1736,N_18776,N_18940);
nand UO_1737 (O_1737,N_19318,N_17736);
and UO_1738 (O_1738,N_17178,N_17788);
nor UO_1739 (O_1739,N_17974,N_17446);
or UO_1740 (O_1740,N_19892,N_19648);
or UO_1741 (O_1741,N_18418,N_19275);
or UO_1742 (O_1742,N_16766,N_18079);
and UO_1743 (O_1743,N_16708,N_17102);
nand UO_1744 (O_1744,N_18156,N_18529);
nor UO_1745 (O_1745,N_19904,N_18636);
nand UO_1746 (O_1746,N_17265,N_17057);
nor UO_1747 (O_1747,N_17936,N_17642);
nor UO_1748 (O_1748,N_17783,N_16030);
nor UO_1749 (O_1749,N_16644,N_16199);
and UO_1750 (O_1750,N_19036,N_17560);
nand UO_1751 (O_1751,N_19853,N_16733);
or UO_1752 (O_1752,N_16990,N_17141);
and UO_1753 (O_1753,N_17305,N_19710);
xnor UO_1754 (O_1754,N_19610,N_16846);
xor UO_1755 (O_1755,N_16380,N_19806);
and UO_1756 (O_1756,N_18888,N_17649);
nor UO_1757 (O_1757,N_17131,N_18699);
nand UO_1758 (O_1758,N_19526,N_19042);
nor UO_1759 (O_1759,N_17585,N_16848);
nor UO_1760 (O_1760,N_19085,N_16451);
nor UO_1761 (O_1761,N_17724,N_16791);
and UO_1762 (O_1762,N_18182,N_18901);
xnor UO_1763 (O_1763,N_19192,N_17050);
nor UO_1764 (O_1764,N_16626,N_16378);
nand UO_1765 (O_1765,N_17587,N_19309);
or UO_1766 (O_1766,N_16827,N_19221);
nor UO_1767 (O_1767,N_18846,N_17389);
and UO_1768 (O_1768,N_18429,N_16105);
nand UO_1769 (O_1769,N_16509,N_19601);
nand UO_1770 (O_1770,N_17702,N_19064);
or UO_1771 (O_1771,N_19938,N_19281);
and UO_1772 (O_1772,N_17921,N_17111);
nor UO_1773 (O_1773,N_18033,N_19102);
xnor UO_1774 (O_1774,N_16930,N_19032);
nor UO_1775 (O_1775,N_18813,N_19099);
nand UO_1776 (O_1776,N_17198,N_18671);
nor UO_1777 (O_1777,N_19021,N_16402);
nand UO_1778 (O_1778,N_17853,N_19604);
nor UO_1779 (O_1779,N_19278,N_17019);
nor UO_1780 (O_1780,N_19135,N_16334);
nand UO_1781 (O_1781,N_16276,N_16823);
nand UO_1782 (O_1782,N_18791,N_19450);
and UO_1783 (O_1783,N_19871,N_19327);
xor UO_1784 (O_1784,N_16845,N_18416);
or UO_1785 (O_1785,N_16135,N_19584);
xor UO_1786 (O_1786,N_17401,N_16913);
or UO_1787 (O_1787,N_16736,N_16737);
and UO_1788 (O_1788,N_18548,N_19934);
or UO_1789 (O_1789,N_16213,N_19400);
and UO_1790 (O_1790,N_17419,N_17258);
nor UO_1791 (O_1791,N_19056,N_19679);
nor UO_1792 (O_1792,N_19550,N_19548);
xnor UO_1793 (O_1793,N_18770,N_18851);
nor UO_1794 (O_1794,N_18517,N_16778);
nand UO_1795 (O_1795,N_19195,N_19916);
nor UO_1796 (O_1796,N_18576,N_17081);
xor UO_1797 (O_1797,N_17013,N_16404);
or UO_1798 (O_1798,N_19803,N_17599);
or UO_1799 (O_1799,N_16040,N_17506);
and UO_1800 (O_1800,N_17728,N_16826);
nand UO_1801 (O_1801,N_18654,N_17497);
nor UO_1802 (O_1802,N_16926,N_17285);
and UO_1803 (O_1803,N_19367,N_18086);
or UO_1804 (O_1804,N_17316,N_18784);
nand UO_1805 (O_1805,N_19051,N_16123);
nand UO_1806 (O_1806,N_16171,N_17417);
and UO_1807 (O_1807,N_17133,N_16980);
and UO_1808 (O_1808,N_17037,N_16665);
nand UO_1809 (O_1809,N_19057,N_16669);
and UO_1810 (O_1810,N_17241,N_17531);
and UO_1811 (O_1811,N_16438,N_16127);
nor UO_1812 (O_1812,N_18173,N_16060);
or UO_1813 (O_1813,N_16263,N_19887);
or UO_1814 (O_1814,N_16965,N_19711);
nor UO_1815 (O_1815,N_17881,N_19816);
xnor UO_1816 (O_1816,N_18600,N_18112);
or UO_1817 (O_1817,N_17780,N_18180);
and UO_1818 (O_1818,N_16689,N_19588);
and UO_1819 (O_1819,N_16014,N_16257);
and UO_1820 (O_1820,N_16771,N_17001);
and UO_1821 (O_1821,N_18523,N_19575);
nand UO_1822 (O_1822,N_19544,N_18258);
and UO_1823 (O_1823,N_16368,N_18374);
and UO_1824 (O_1824,N_16534,N_17978);
nor UO_1825 (O_1825,N_18107,N_18276);
nor UO_1826 (O_1826,N_19375,N_17956);
xnor UO_1827 (O_1827,N_17250,N_19290);
nand UO_1828 (O_1828,N_19411,N_19602);
and UO_1829 (O_1829,N_17138,N_18198);
nor UO_1830 (O_1830,N_16834,N_17756);
nor UO_1831 (O_1831,N_19663,N_17165);
nand UO_1832 (O_1832,N_17509,N_17291);
or UO_1833 (O_1833,N_16612,N_17580);
xor UO_1834 (O_1834,N_16867,N_17103);
nor UO_1835 (O_1835,N_17125,N_19586);
nand UO_1836 (O_1836,N_18801,N_18982);
and UO_1837 (O_1837,N_16306,N_17071);
and UO_1838 (O_1838,N_16973,N_18780);
xnor UO_1839 (O_1839,N_16482,N_18150);
nor UO_1840 (O_1840,N_17528,N_17719);
or UO_1841 (O_1841,N_19423,N_18310);
xor UO_1842 (O_1842,N_18455,N_19988);
and UO_1843 (O_1843,N_16720,N_17218);
nand UO_1844 (O_1844,N_18065,N_19861);
and UO_1845 (O_1845,N_18261,N_19120);
or UO_1846 (O_1846,N_17110,N_18147);
nor UO_1847 (O_1847,N_19258,N_19730);
xor UO_1848 (O_1848,N_18289,N_17955);
nand UO_1849 (O_1849,N_16634,N_17656);
or UO_1850 (O_1850,N_19977,N_17985);
or UO_1851 (O_1851,N_17233,N_18400);
or UO_1852 (O_1852,N_18293,N_18754);
nand UO_1853 (O_1853,N_18746,N_19086);
and UO_1854 (O_1854,N_19979,N_18419);
or UO_1855 (O_1855,N_19504,N_16443);
xor UO_1856 (O_1856,N_19760,N_18952);
nand UO_1857 (O_1857,N_18271,N_17429);
or UO_1858 (O_1858,N_18222,N_16142);
and UO_1859 (O_1859,N_16889,N_18991);
nand UO_1860 (O_1860,N_17939,N_18692);
nand UO_1861 (O_1861,N_17015,N_17223);
or UO_1862 (O_1862,N_18174,N_17244);
or UO_1863 (O_1863,N_17246,N_18580);
nand UO_1864 (O_1864,N_17060,N_19883);
nand UO_1865 (O_1865,N_16516,N_17930);
and UO_1866 (O_1866,N_19076,N_17008);
nand UO_1867 (O_1867,N_18781,N_19565);
nor UO_1868 (O_1868,N_18832,N_16652);
nand UO_1869 (O_1869,N_16525,N_16203);
or UO_1870 (O_1870,N_18318,N_16952);
nand UO_1871 (O_1871,N_19795,N_17734);
and UO_1872 (O_1872,N_18678,N_17097);
or UO_1873 (O_1873,N_19437,N_19658);
xnor UO_1874 (O_1874,N_19637,N_16456);
nand UO_1875 (O_1875,N_19502,N_17483);
nor UO_1876 (O_1876,N_17373,N_19775);
nand UO_1877 (O_1877,N_16461,N_17315);
or UO_1878 (O_1878,N_18169,N_18687);
nand UO_1879 (O_1879,N_16726,N_18373);
xnor UO_1880 (O_1880,N_17834,N_16347);
and UO_1881 (O_1881,N_17588,N_17035);
or UO_1882 (O_1882,N_17147,N_16719);
or UO_1883 (O_1883,N_18425,N_17129);
nor UO_1884 (O_1884,N_19594,N_16908);
or UO_1885 (O_1885,N_19878,N_19962);
nor UO_1886 (O_1886,N_18250,N_19754);
and UO_1887 (O_1887,N_18941,N_18069);
or UO_1888 (O_1888,N_17959,N_16770);
and UO_1889 (O_1889,N_18714,N_19809);
or UO_1890 (O_1890,N_16723,N_16882);
nand UO_1891 (O_1891,N_19457,N_16716);
and UO_1892 (O_1892,N_18288,N_17698);
nand UO_1893 (O_1893,N_16295,N_17616);
or UO_1894 (O_1894,N_17422,N_16642);
or UO_1895 (O_1895,N_19151,N_19708);
or UO_1896 (O_1896,N_17091,N_17400);
nor UO_1897 (O_1897,N_16532,N_19937);
nand UO_1898 (O_1898,N_17833,N_19583);
and UO_1899 (O_1899,N_19121,N_18972);
and UO_1900 (O_1900,N_19847,N_16813);
or UO_1901 (O_1901,N_19898,N_17169);
nor UO_1902 (O_1902,N_18763,N_16758);
nor UO_1903 (O_1903,N_19783,N_17282);
nand UO_1904 (O_1904,N_16009,N_18838);
and UO_1905 (O_1905,N_16153,N_18582);
nand UO_1906 (O_1906,N_16684,N_19886);
nand UO_1907 (O_1907,N_17453,N_17005);
nand UO_1908 (O_1908,N_19642,N_19071);
nor UO_1909 (O_1909,N_18244,N_17513);
and UO_1910 (O_1910,N_17391,N_19592);
or UO_1911 (O_1911,N_18542,N_19560);
nor UO_1912 (O_1912,N_17685,N_16508);
or UO_1913 (O_1913,N_18125,N_18742);
nand UO_1914 (O_1914,N_18954,N_16760);
nand UO_1915 (O_1915,N_16574,N_18573);
nor UO_1916 (O_1916,N_19409,N_17571);
and UO_1917 (O_1917,N_18123,N_18312);
xnor UO_1918 (O_1918,N_19072,N_16053);
and UO_1919 (O_1919,N_18964,N_19568);
and UO_1920 (O_1920,N_17184,N_17762);
or UO_1921 (O_1921,N_17343,N_16251);
xnor UO_1922 (O_1922,N_18717,N_19966);
and UO_1923 (O_1923,N_18533,N_19329);
nor UO_1924 (O_1924,N_19827,N_18903);
nand UO_1925 (O_1925,N_16561,N_16431);
xnor UO_1926 (O_1926,N_19141,N_19048);
and UO_1927 (O_1927,N_16331,N_17004);
or UO_1928 (O_1928,N_17243,N_17393);
nor UO_1929 (O_1929,N_19031,N_16132);
or UO_1930 (O_1930,N_18764,N_16907);
nand UO_1931 (O_1931,N_17329,N_18602);
xnor UO_1932 (O_1932,N_17012,N_18165);
and UO_1933 (O_1933,N_17270,N_17096);
or UO_1934 (O_1934,N_19848,N_17920);
nand UO_1935 (O_1935,N_16621,N_16204);
nor UO_1936 (O_1936,N_18155,N_19426);
and UO_1937 (O_1937,N_18179,N_16205);
nor UO_1938 (O_1938,N_19617,N_19201);
nand UO_1939 (O_1939,N_17752,N_18668);
nand UO_1940 (O_1940,N_18862,N_17472);
or UO_1941 (O_1941,N_18286,N_18914);
nand UO_1942 (O_1942,N_19335,N_17038);
nor UO_1943 (O_1943,N_16088,N_17535);
or UO_1944 (O_1944,N_17073,N_19286);
or UO_1945 (O_1945,N_19936,N_16904);
xor UO_1946 (O_1946,N_18854,N_19139);
nand UO_1947 (O_1947,N_18601,N_16330);
or UO_1948 (O_1948,N_18140,N_16729);
or UO_1949 (O_1949,N_17625,N_18091);
or UO_1950 (O_1950,N_16831,N_19364);
nor UO_1951 (O_1951,N_17971,N_19282);
or UO_1952 (O_1952,N_16954,N_16878);
xnor UO_1953 (O_1953,N_17211,N_18076);
nor UO_1954 (O_1954,N_17009,N_19478);
nand UO_1955 (O_1955,N_19989,N_16887);
nor UO_1956 (O_1956,N_18345,N_19477);
nor UO_1957 (O_1957,N_19529,N_17475);
and UO_1958 (O_1958,N_19940,N_18344);
nand UO_1959 (O_1959,N_16255,N_19956);
nor UO_1960 (O_1960,N_19585,N_17339);
nor UO_1961 (O_1961,N_18695,N_19232);
and UO_1962 (O_1962,N_19762,N_19970);
nor UO_1963 (O_1963,N_16208,N_18969);
or UO_1964 (O_1964,N_19274,N_17954);
and UO_1965 (O_1965,N_17824,N_16873);
or UO_1966 (O_1966,N_19941,N_17626);
xnor UO_1967 (O_1967,N_19257,N_18883);
or UO_1968 (O_1968,N_19087,N_18612);
xnor UO_1969 (O_1969,N_18461,N_16743);
nand UO_1970 (O_1970,N_18645,N_16936);
or UO_1971 (O_1971,N_18177,N_16872);
nand UO_1972 (O_1972,N_18321,N_19269);
xor UO_1973 (O_1973,N_16308,N_18863);
and UO_1974 (O_1974,N_16569,N_16418);
nand UO_1975 (O_1975,N_18205,N_16517);
and UO_1976 (O_1976,N_19467,N_17083);
nand UO_1977 (O_1977,N_17827,N_18989);
nand UO_1978 (O_1978,N_16253,N_17049);
xnor UO_1979 (O_1979,N_17033,N_18623);
nand UO_1980 (O_1980,N_19974,N_16599);
nand UO_1981 (O_1981,N_18577,N_19889);
nor UO_1982 (O_1982,N_16677,N_16433);
nand UO_1983 (O_1983,N_17845,N_16025);
or UO_1984 (O_1984,N_19006,N_19527);
nand UO_1985 (O_1985,N_18873,N_18640);
xnor UO_1986 (O_1986,N_17498,N_18676);
or UO_1987 (O_1987,N_17942,N_18990);
nand UO_1988 (O_1988,N_18328,N_16790);
nand UO_1989 (O_1989,N_19872,N_16113);
or UO_1990 (O_1990,N_17846,N_16151);
and UO_1991 (O_1991,N_18279,N_19247);
or UO_1992 (O_1992,N_16187,N_18894);
nor UO_1993 (O_1993,N_17952,N_16412);
nand UO_1994 (O_1994,N_19420,N_19766);
nor UO_1995 (O_1995,N_19068,N_16027);
nand UO_1996 (O_1996,N_18660,N_19440);
nor UO_1997 (O_1997,N_17303,N_16233);
or UO_1998 (O_1998,N_18202,N_19226);
or UO_1999 (O_1999,N_19669,N_19489);
and UO_2000 (O_2000,N_16540,N_18810);
or UO_2001 (O_2001,N_19654,N_19759);
and UO_2002 (O_2002,N_16721,N_17170);
or UO_2003 (O_2003,N_18596,N_18537);
nor UO_2004 (O_2004,N_19345,N_16289);
xor UO_2005 (O_2005,N_18587,N_18298);
and UO_2006 (O_2006,N_17867,N_18766);
nor UO_2007 (O_2007,N_16538,N_19390);
and UO_2008 (O_2008,N_19919,N_16015);
xnor UO_2009 (O_2009,N_18740,N_18959);
or UO_2010 (O_2010,N_18076,N_16559);
xor UO_2011 (O_2011,N_19418,N_19722);
nand UO_2012 (O_2012,N_18500,N_19108);
nand UO_2013 (O_2013,N_16469,N_18942);
or UO_2014 (O_2014,N_16899,N_16128);
nand UO_2015 (O_2015,N_17951,N_18279);
and UO_2016 (O_2016,N_18356,N_19073);
xor UO_2017 (O_2017,N_17002,N_18353);
nand UO_2018 (O_2018,N_16321,N_18660);
xor UO_2019 (O_2019,N_18863,N_18760);
and UO_2020 (O_2020,N_18874,N_18422);
xnor UO_2021 (O_2021,N_19836,N_17316);
nand UO_2022 (O_2022,N_17726,N_17451);
nor UO_2023 (O_2023,N_18284,N_19933);
nor UO_2024 (O_2024,N_18147,N_19647);
xor UO_2025 (O_2025,N_18998,N_19401);
nand UO_2026 (O_2026,N_19521,N_19324);
xor UO_2027 (O_2027,N_16381,N_16261);
nor UO_2028 (O_2028,N_19767,N_19837);
nand UO_2029 (O_2029,N_18509,N_17184);
xor UO_2030 (O_2030,N_19063,N_16660);
xnor UO_2031 (O_2031,N_17248,N_18447);
nor UO_2032 (O_2032,N_18378,N_19151);
nor UO_2033 (O_2033,N_16883,N_17030);
nand UO_2034 (O_2034,N_18018,N_18765);
or UO_2035 (O_2035,N_17107,N_19170);
nand UO_2036 (O_2036,N_17740,N_18851);
and UO_2037 (O_2037,N_19522,N_16733);
or UO_2038 (O_2038,N_17076,N_19103);
nor UO_2039 (O_2039,N_19970,N_17090);
nor UO_2040 (O_2040,N_19917,N_16618);
or UO_2041 (O_2041,N_16029,N_18722);
and UO_2042 (O_2042,N_18805,N_18011);
or UO_2043 (O_2043,N_18628,N_17199);
and UO_2044 (O_2044,N_18965,N_17306);
nor UO_2045 (O_2045,N_17294,N_16291);
xnor UO_2046 (O_2046,N_19047,N_19672);
or UO_2047 (O_2047,N_18713,N_19621);
and UO_2048 (O_2048,N_16270,N_16814);
nor UO_2049 (O_2049,N_16270,N_18982);
and UO_2050 (O_2050,N_18484,N_18580);
xnor UO_2051 (O_2051,N_18717,N_18394);
nor UO_2052 (O_2052,N_19102,N_16973);
nand UO_2053 (O_2053,N_17759,N_16209);
xor UO_2054 (O_2054,N_17557,N_16733);
nor UO_2055 (O_2055,N_18537,N_16392);
nor UO_2056 (O_2056,N_17815,N_18628);
xor UO_2057 (O_2057,N_17140,N_17446);
nor UO_2058 (O_2058,N_19707,N_19095);
nand UO_2059 (O_2059,N_18674,N_16422);
or UO_2060 (O_2060,N_16950,N_19178);
nor UO_2061 (O_2061,N_18211,N_16656);
or UO_2062 (O_2062,N_18191,N_17260);
nor UO_2063 (O_2063,N_17034,N_17983);
nand UO_2064 (O_2064,N_17129,N_18944);
or UO_2065 (O_2065,N_18677,N_18957);
nor UO_2066 (O_2066,N_18192,N_19056);
nor UO_2067 (O_2067,N_19802,N_17883);
or UO_2068 (O_2068,N_16866,N_19124);
xor UO_2069 (O_2069,N_17554,N_16903);
and UO_2070 (O_2070,N_16960,N_18487);
nor UO_2071 (O_2071,N_17664,N_16718);
or UO_2072 (O_2072,N_19088,N_16019);
or UO_2073 (O_2073,N_18282,N_18919);
or UO_2074 (O_2074,N_17303,N_19088);
nor UO_2075 (O_2075,N_19568,N_17198);
and UO_2076 (O_2076,N_18397,N_16316);
or UO_2077 (O_2077,N_19965,N_18334);
or UO_2078 (O_2078,N_19148,N_16236);
and UO_2079 (O_2079,N_18146,N_17464);
and UO_2080 (O_2080,N_19369,N_17852);
xor UO_2081 (O_2081,N_17653,N_17020);
nor UO_2082 (O_2082,N_19494,N_16072);
nand UO_2083 (O_2083,N_17014,N_18979);
nor UO_2084 (O_2084,N_18019,N_17850);
nand UO_2085 (O_2085,N_18631,N_18622);
and UO_2086 (O_2086,N_17563,N_18742);
xnor UO_2087 (O_2087,N_17025,N_16912);
or UO_2088 (O_2088,N_18915,N_17142);
nand UO_2089 (O_2089,N_18550,N_19472);
or UO_2090 (O_2090,N_17544,N_18843);
nor UO_2091 (O_2091,N_19410,N_17892);
nand UO_2092 (O_2092,N_16888,N_17048);
or UO_2093 (O_2093,N_16242,N_17763);
and UO_2094 (O_2094,N_19605,N_18917);
nor UO_2095 (O_2095,N_18278,N_18120);
and UO_2096 (O_2096,N_16875,N_18336);
or UO_2097 (O_2097,N_18821,N_16453);
or UO_2098 (O_2098,N_19713,N_18402);
and UO_2099 (O_2099,N_19676,N_16215);
and UO_2100 (O_2100,N_18015,N_17431);
or UO_2101 (O_2101,N_17144,N_19837);
and UO_2102 (O_2102,N_16288,N_19399);
nand UO_2103 (O_2103,N_18919,N_17108);
nor UO_2104 (O_2104,N_17253,N_17096);
nand UO_2105 (O_2105,N_16666,N_17255);
xor UO_2106 (O_2106,N_18958,N_18652);
and UO_2107 (O_2107,N_16580,N_19848);
xnor UO_2108 (O_2108,N_17389,N_16100);
xnor UO_2109 (O_2109,N_16551,N_17779);
nand UO_2110 (O_2110,N_19863,N_16689);
xnor UO_2111 (O_2111,N_18206,N_19760);
xnor UO_2112 (O_2112,N_19573,N_18244);
nor UO_2113 (O_2113,N_19358,N_19871);
xor UO_2114 (O_2114,N_19016,N_18978);
nor UO_2115 (O_2115,N_19133,N_19912);
xor UO_2116 (O_2116,N_17263,N_16767);
nor UO_2117 (O_2117,N_16026,N_18241);
nor UO_2118 (O_2118,N_16278,N_19597);
nor UO_2119 (O_2119,N_18349,N_19256);
or UO_2120 (O_2120,N_18358,N_18883);
xnor UO_2121 (O_2121,N_18752,N_16953);
and UO_2122 (O_2122,N_19722,N_17315);
and UO_2123 (O_2123,N_17250,N_17142);
and UO_2124 (O_2124,N_17505,N_19645);
or UO_2125 (O_2125,N_17957,N_19052);
nand UO_2126 (O_2126,N_19227,N_17862);
nand UO_2127 (O_2127,N_16104,N_17362);
xnor UO_2128 (O_2128,N_16521,N_16618);
xnor UO_2129 (O_2129,N_19372,N_17651);
or UO_2130 (O_2130,N_16984,N_18549);
nor UO_2131 (O_2131,N_18723,N_18646);
or UO_2132 (O_2132,N_17888,N_19514);
nor UO_2133 (O_2133,N_19534,N_18693);
nand UO_2134 (O_2134,N_16196,N_19422);
nand UO_2135 (O_2135,N_17023,N_17362);
and UO_2136 (O_2136,N_16722,N_18507);
or UO_2137 (O_2137,N_19962,N_18809);
nand UO_2138 (O_2138,N_19555,N_17348);
nor UO_2139 (O_2139,N_19300,N_19011);
nor UO_2140 (O_2140,N_18487,N_18699);
or UO_2141 (O_2141,N_17348,N_19208);
or UO_2142 (O_2142,N_18245,N_17684);
or UO_2143 (O_2143,N_17867,N_17917);
and UO_2144 (O_2144,N_18583,N_16249);
or UO_2145 (O_2145,N_17762,N_17532);
nor UO_2146 (O_2146,N_16580,N_16861);
nor UO_2147 (O_2147,N_17110,N_16676);
nand UO_2148 (O_2148,N_16019,N_16275);
nand UO_2149 (O_2149,N_18876,N_19556);
or UO_2150 (O_2150,N_19434,N_16294);
xor UO_2151 (O_2151,N_17085,N_18300);
and UO_2152 (O_2152,N_16164,N_16633);
nand UO_2153 (O_2153,N_16657,N_18414);
and UO_2154 (O_2154,N_18148,N_16766);
nor UO_2155 (O_2155,N_16143,N_16497);
xnor UO_2156 (O_2156,N_18265,N_18570);
or UO_2157 (O_2157,N_17717,N_19265);
xnor UO_2158 (O_2158,N_18401,N_19478);
or UO_2159 (O_2159,N_16181,N_16742);
nand UO_2160 (O_2160,N_19004,N_17968);
xnor UO_2161 (O_2161,N_16049,N_17345);
nand UO_2162 (O_2162,N_18875,N_18897);
nand UO_2163 (O_2163,N_16311,N_17589);
or UO_2164 (O_2164,N_18705,N_16000);
nand UO_2165 (O_2165,N_18611,N_16000);
nor UO_2166 (O_2166,N_19039,N_18184);
and UO_2167 (O_2167,N_19742,N_17529);
or UO_2168 (O_2168,N_17501,N_16007);
nor UO_2169 (O_2169,N_18063,N_19705);
xor UO_2170 (O_2170,N_19622,N_16886);
nand UO_2171 (O_2171,N_16562,N_19282);
nand UO_2172 (O_2172,N_16561,N_16416);
and UO_2173 (O_2173,N_16789,N_17603);
and UO_2174 (O_2174,N_19578,N_17934);
xnor UO_2175 (O_2175,N_16311,N_18481);
nor UO_2176 (O_2176,N_18666,N_16484);
and UO_2177 (O_2177,N_19225,N_19326);
and UO_2178 (O_2178,N_16005,N_16220);
xnor UO_2179 (O_2179,N_19691,N_19383);
nor UO_2180 (O_2180,N_18818,N_19182);
and UO_2181 (O_2181,N_18889,N_19216);
or UO_2182 (O_2182,N_18075,N_19076);
and UO_2183 (O_2183,N_16542,N_16652);
nor UO_2184 (O_2184,N_18331,N_17859);
nor UO_2185 (O_2185,N_17280,N_17464);
nor UO_2186 (O_2186,N_17441,N_16062);
nor UO_2187 (O_2187,N_17612,N_18507);
and UO_2188 (O_2188,N_17183,N_19079);
nor UO_2189 (O_2189,N_17878,N_18343);
nor UO_2190 (O_2190,N_17451,N_19258);
nor UO_2191 (O_2191,N_16542,N_18929);
xor UO_2192 (O_2192,N_18493,N_18777);
nand UO_2193 (O_2193,N_19297,N_18266);
nor UO_2194 (O_2194,N_18302,N_19638);
nor UO_2195 (O_2195,N_17014,N_18370);
or UO_2196 (O_2196,N_18564,N_17475);
xnor UO_2197 (O_2197,N_19824,N_18745);
and UO_2198 (O_2198,N_19711,N_18511);
or UO_2199 (O_2199,N_18252,N_16187);
and UO_2200 (O_2200,N_16375,N_17490);
or UO_2201 (O_2201,N_16120,N_17327);
nand UO_2202 (O_2202,N_18803,N_19808);
or UO_2203 (O_2203,N_17344,N_19314);
xor UO_2204 (O_2204,N_16058,N_18408);
nor UO_2205 (O_2205,N_18218,N_17423);
nand UO_2206 (O_2206,N_16819,N_18354);
nand UO_2207 (O_2207,N_16816,N_19016);
nand UO_2208 (O_2208,N_19838,N_17333);
nor UO_2209 (O_2209,N_16595,N_19754);
nand UO_2210 (O_2210,N_18456,N_19505);
nand UO_2211 (O_2211,N_16556,N_19550);
nand UO_2212 (O_2212,N_17680,N_18989);
and UO_2213 (O_2213,N_18566,N_17238);
nor UO_2214 (O_2214,N_17652,N_16648);
xnor UO_2215 (O_2215,N_19195,N_17426);
nand UO_2216 (O_2216,N_16096,N_18923);
and UO_2217 (O_2217,N_16639,N_18301);
nor UO_2218 (O_2218,N_16536,N_18244);
or UO_2219 (O_2219,N_16129,N_17473);
or UO_2220 (O_2220,N_19571,N_19080);
nor UO_2221 (O_2221,N_17362,N_18438);
nand UO_2222 (O_2222,N_17156,N_16832);
xnor UO_2223 (O_2223,N_19663,N_17987);
nand UO_2224 (O_2224,N_17552,N_17561);
nand UO_2225 (O_2225,N_16182,N_16707);
xor UO_2226 (O_2226,N_17315,N_17338);
nand UO_2227 (O_2227,N_16662,N_17156);
and UO_2228 (O_2228,N_19426,N_19607);
nor UO_2229 (O_2229,N_17097,N_18407);
and UO_2230 (O_2230,N_17371,N_17729);
nand UO_2231 (O_2231,N_18440,N_18673);
nand UO_2232 (O_2232,N_19897,N_18444);
nand UO_2233 (O_2233,N_18924,N_17857);
and UO_2234 (O_2234,N_16595,N_17489);
nor UO_2235 (O_2235,N_17589,N_16346);
nand UO_2236 (O_2236,N_16178,N_17481);
or UO_2237 (O_2237,N_17297,N_19482);
nand UO_2238 (O_2238,N_18953,N_18183);
nor UO_2239 (O_2239,N_18215,N_16797);
nor UO_2240 (O_2240,N_16238,N_18125);
and UO_2241 (O_2241,N_16621,N_16810);
xor UO_2242 (O_2242,N_17915,N_18391);
and UO_2243 (O_2243,N_18165,N_19180);
xor UO_2244 (O_2244,N_18601,N_18401);
and UO_2245 (O_2245,N_17259,N_18120);
nand UO_2246 (O_2246,N_19014,N_17594);
nor UO_2247 (O_2247,N_16539,N_18375);
or UO_2248 (O_2248,N_18300,N_16973);
nor UO_2249 (O_2249,N_19192,N_19468);
nor UO_2250 (O_2250,N_16748,N_17201);
nor UO_2251 (O_2251,N_16240,N_18234);
and UO_2252 (O_2252,N_19644,N_16615);
nor UO_2253 (O_2253,N_19390,N_19079);
nand UO_2254 (O_2254,N_18681,N_17579);
nand UO_2255 (O_2255,N_17139,N_19143);
nor UO_2256 (O_2256,N_16240,N_16747);
xor UO_2257 (O_2257,N_18655,N_17991);
xor UO_2258 (O_2258,N_16871,N_16840);
and UO_2259 (O_2259,N_16044,N_18686);
and UO_2260 (O_2260,N_16655,N_16457);
nor UO_2261 (O_2261,N_16659,N_16521);
nand UO_2262 (O_2262,N_19466,N_19732);
xnor UO_2263 (O_2263,N_17882,N_16331);
nand UO_2264 (O_2264,N_18137,N_18789);
nor UO_2265 (O_2265,N_19306,N_17084);
and UO_2266 (O_2266,N_17319,N_19701);
nand UO_2267 (O_2267,N_19215,N_16504);
or UO_2268 (O_2268,N_16446,N_18473);
nand UO_2269 (O_2269,N_18030,N_16595);
xor UO_2270 (O_2270,N_19395,N_17635);
nand UO_2271 (O_2271,N_18309,N_16282);
nor UO_2272 (O_2272,N_18992,N_19213);
or UO_2273 (O_2273,N_19528,N_18009);
nand UO_2274 (O_2274,N_19323,N_17901);
xor UO_2275 (O_2275,N_19047,N_19730);
or UO_2276 (O_2276,N_18030,N_16265);
nand UO_2277 (O_2277,N_19615,N_19263);
xnor UO_2278 (O_2278,N_16430,N_19422);
or UO_2279 (O_2279,N_19773,N_19600);
and UO_2280 (O_2280,N_17730,N_18457);
nand UO_2281 (O_2281,N_19458,N_16231);
or UO_2282 (O_2282,N_17486,N_19603);
nand UO_2283 (O_2283,N_18142,N_18636);
and UO_2284 (O_2284,N_19417,N_16904);
or UO_2285 (O_2285,N_19597,N_18982);
nor UO_2286 (O_2286,N_16602,N_18470);
nand UO_2287 (O_2287,N_17344,N_18247);
nor UO_2288 (O_2288,N_19769,N_16117);
nand UO_2289 (O_2289,N_17174,N_17408);
nand UO_2290 (O_2290,N_18051,N_17512);
and UO_2291 (O_2291,N_17794,N_18845);
nor UO_2292 (O_2292,N_17225,N_19271);
and UO_2293 (O_2293,N_17469,N_19895);
or UO_2294 (O_2294,N_18889,N_18137);
nor UO_2295 (O_2295,N_16330,N_16491);
nand UO_2296 (O_2296,N_16638,N_18669);
xor UO_2297 (O_2297,N_17565,N_17407);
nand UO_2298 (O_2298,N_17846,N_19012);
nor UO_2299 (O_2299,N_19580,N_16009);
nor UO_2300 (O_2300,N_18495,N_18003);
nor UO_2301 (O_2301,N_19502,N_18731);
nor UO_2302 (O_2302,N_18942,N_18601);
xnor UO_2303 (O_2303,N_17502,N_16496);
nand UO_2304 (O_2304,N_19155,N_17903);
nand UO_2305 (O_2305,N_18830,N_19272);
or UO_2306 (O_2306,N_17901,N_18865);
nor UO_2307 (O_2307,N_16824,N_17411);
and UO_2308 (O_2308,N_19139,N_16065);
and UO_2309 (O_2309,N_16382,N_17036);
nand UO_2310 (O_2310,N_17328,N_18463);
nand UO_2311 (O_2311,N_18743,N_19731);
nor UO_2312 (O_2312,N_17085,N_17782);
nor UO_2313 (O_2313,N_16787,N_18059);
nand UO_2314 (O_2314,N_17204,N_17551);
xor UO_2315 (O_2315,N_18177,N_16904);
or UO_2316 (O_2316,N_18677,N_18918);
nor UO_2317 (O_2317,N_18279,N_16503);
nor UO_2318 (O_2318,N_16767,N_18168);
nand UO_2319 (O_2319,N_19801,N_19367);
nor UO_2320 (O_2320,N_19472,N_17419);
or UO_2321 (O_2321,N_19911,N_16536);
xnor UO_2322 (O_2322,N_17936,N_16612);
and UO_2323 (O_2323,N_16606,N_17716);
nor UO_2324 (O_2324,N_19065,N_16301);
nand UO_2325 (O_2325,N_17555,N_18194);
nor UO_2326 (O_2326,N_19396,N_19825);
nor UO_2327 (O_2327,N_18812,N_17502);
and UO_2328 (O_2328,N_19651,N_19501);
or UO_2329 (O_2329,N_17899,N_19863);
nor UO_2330 (O_2330,N_18352,N_18139);
nand UO_2331 (O_2331,N_17732,N_18248);
nor UO_2332 (O_2332,N_16526,N_19376);
and UO_2333 (O_2333,N_17286,N_19505);
or UO_2334 (O_2334,N_16815,N_17560);
nand UO_2335 (O_2335,N_16574,N_19220);
nand UO_2336 (O_2336,N_16938,N_17681);
nand UO_2337 (O_2337,N_16285,N_16012);
nand UO_2338 (O_2338,N_16597,N_18869);
or UO_2339 (O_2339,N_18111,N_16674);
or UO_2340 (O_2340,N_18645,N_19886);
and UO_2341 (O_2341,N_18683,N_18646);
xor UO_2342 (O_2342,N_16280,N_17647);
or UO_2343 (O_2343,N_19952,N_18915);
xnor UO_2344 (O_2344,N_18961,N_16448);
or UO_2345 (O_2345,N_18103,N_17452);
xnor UO_2346 (O_2346,N_16495,N_19042);
nor UO_2347 (O_2347,N_19227,N_17151);
nand UO_2348 (O_2348,N_17177,N_19913);
nand UO_2349 (O_2349,N_17705,N_18996);
nand UO_2350 (O_2350,N_16256,N_19597);
nor UO_2351 (O_2351,N_19071,N_18579);
or UO_2352 (O_2352,N_19795,N_16801);
nor UO_2353 (O_2353,N_17551,N_18290);
and UO_2354 (O_2354,N_18141,N_17833);
nor UO_2355 (O_2355,N_19334,N_16926);
or UO_2356 (O_2356,N_17544,N_16706);
and UO_2357 (O_2357,N_19325,N_17182);
or UO_2358 (O_2358,N_18101,N_19076);
nor UO_2359 (O_2359,N_18224,N_18617);
xor UO_2360 (O_2360,N_19170,N_16744);
nor UO_2361 (O_2361,N_19058,N_17162);
nand UO_2362 (O_2362,N_16366,N_16641);
nand UO_2363 (O_2363,N_19429,N_19866);
or UO_2364 (O_2364,N_16218,N_17895);
or UO_2365 (O_2365,N_17361,N_17787);
xnor UO_2366 (O_2366,N_17122,N_18773);
or UO_2367 (O_2367,N_17364,N_19905);
nor UO_2368 (O_2368,N_18130,N_17854);
nand UO_2369 (O_2369,N_18929,N_17382);
nor UO_2370 (O_2370,N_18871,N_16269);
or UO_2371 (O_2371,N_16665,N_17976);
and UO_2372 (O_2372,N_17154,N_16469);
nor UO_2373 (O_2373,N_17574,N_16887);
xnor UO_2374 (O_2374,N_19542,N_16584);
nand UO_2375 (O_2375,N_19935,N_19398);
or UO_2376 (O_2376,N_16174,N_19974);
or UO_2377 (O_2377,N_19677,N_18745);
nor UO_2378 (O_2378,N_19604,N_18343);
or UO_2379 (O_2379,N_16418,N_19781);
nor UO_2380 (O_2380,N_18406,N_17813);
or UO_2381 (O_2381,N_18633,N_18203);
nor UO_2382 (O_2382,N_18504,N_17741);
and UO_2383 (O_2383,N_16603,N_18515);
and UO_2384 (O_2384,N_19290,N_17625);
or UO_2385 (O_2385,N_18106,N_18957);
nand UO_2386 (O_2386,N_17573,N_18074);
nor UO_2387 (O_2387,N_18515,N_17862);
and UO_2388 (O_2388,N_17557,N_16526);
nor UO_2389 (O_2389,N_17212,N_18067);
nor UO_2390 (O_2390,N_17790,N_16677);
and UO_2391 (O_2391,N_19699,N_18620);
nor UO_2392 (O_2392,N_19060,N_17089);
or UO_2393 (O_2393,N_19036,N_17189);
and UO_2394 (O_2394,N_17385,N_19441);
or UO_2395 (O_2395,N_19575,N_16513);
nand UO_2396 (O_2396,N_19204,N_16740);
and UO_2397 (O_2397,N_18459,N_16618);
or UO_2398 (O_2398,N_18442,N_19049);
and UO_2399 (O_2399,N_17629,N_19259);
xnor UO_2400 (O_2400,N_19508,N_17703);
or UO_2401 (O_2401,N_19856,N_17476);
nor UO_2402 (O_2402,N_18349,N_19424);
and UO_2403 (O_2403,N_19330,N_19769);
and UO_2404 (O_2404,N_18103,N_19379);
and UO_2405 (O_2405,N_18674,N_16035);
nor UO_2406 (O_2406,N_18274,N_17800);
nor UO_2407 (O_2407,N_17491,N_19868);
xnor UO_2408 (O_2408,N_17531,N_18288);
and UO_2409 (O_2409,N_19366,N_18041);
or UO_2410 (O_2410,N_19483,N_16987);
nor UO_2411 (O_2411,N_19148,N_18605);
nor UO_2412 (O_2412,N_16149,N_16716);
nand UO_2413 (O_2413,N_16362,N_17995);
or UO_2414 (O_2414,N_17831,N_17253);
and UO_2415 (O_2415,N_18354,N_16692);
nand UO_2416 (O_2416,N_18478,N_16707);
and UO_2417 (O_2417,N_18767,N_19432);
xnor UO_2418 (O_2418,N_16182,N_17180);
and UO_2419 (O_2419,N_19459,N_16902);
and UO_2420 (O_2420,N_17082,N_16345);
or UO_2421 (O_2421,N_17707,N_19075);
xnor UO_2422 (O_2422,N_16402,N_19738);
xor UO_2423 (O_2423,N_17062,N_17232);
nor UO_2424 (O_2424,N_18501,N_18320);
and UO_2425 (O_2425,N_17888,N_16473);
nand UO_2426 (O_2426,N_19985,N_16505);
or UO_2427 (O_2427,N_19331,N_19454);
and UO_2428 (O_2428,N_17835,N_19206);
nor UO_2429 (O_2429,N_19932,N_16660);
nor UO_2430 (O_2430,N_19958,N_18741);
nand UO_2431 (O_2431,N_18108,N_17773);
xnor UO_2432 (O_2432,N_16115,N_19384);
and UO_2433 (O_2433,N_16517,N_17296);
or UO_2434 (O_2434,N_16336,N_19818);
or UO_2435 (O_2435,N_16284,N_16748);
or UO_2436 (O_2436,N_16443,N_16802);
or UO_2437 (O_2437,N_17991,N_18734);
and UO_2438 (O_2438,N_16904,N_16826);
and UO_2439 (O_2439,N_19923,N_16550);
or UO_2440 (O_2440,N_17519,N_19375);
xnor UO_2441 (O_2441,N_19821,N_16587);
xor UO_2442 (O_2442,N_19128,N_17908);
nor UO_2443 (O_2443,N_18213,N_19591);
nor UO_2444 (O_2444,N_16898,N_18274);
xnor UO_2445 (O_2445,N_17101,N_18775);
and UO_2446 (O_2446,N_16185,N_19284);
and UO_2447 (O_2447,N_19969,N_16222);
and UO_2448 (O_2448,N_19281,N_18402);
or UO_2449 (O_2449,N_19269,N_19111);
nand UO_2450 (O_2450,N_17700,N_17695);
or UO_2451 (O_2451,N_18011,N_17308);
or UO_2452 (O_2452,N_16879,N_19583);
nand UO_2453 (O_2453,N_18399,N_17825);
and UO_2454 (O_2454,N_17847,N_17058);
or UO_2455 (O_2455,N_17081,N_16454);
and UO_2456 (O_2456,N_17719,N_18453);
nor UO_2457 (O_2457,N_19252,N_19289);
nand UO_2458 (O_2458,N_19839,N_17638);
or UO_2459 (O_2459,N_17894,N_17759);
nand UO_2460 (O_2460,N_18346,N_18303);
nand UO_2461 (O_2461,N_18852,N_17364);
xnor UO_2462 (O_2462,N_16939,N_19422);
xnor UO_2463 (O_2463,N_18910,N_18285);
nor UO_2464 (O_2464,N_19148,N_17655);
nor UO_2465 (O_2465,N_18754,N_16241);
nand UO_2466 (O_2466,N_19396,N_19081);
nand UO_2467 (O_2467,N_19643,N_16673);
nand UO_2468 (O_2468,N_17115,N_19701);
nand UO_2469 (O_2469,N_16347,N_18819);
nor UO_2470 (O_2470,N_17309,N_18308);
nor UO_2471 (O_2471,N_17934,N_19563);
nand UO_2472 (O_2472,N_19235,N_17409);
or UO_2473 (O_2473,N_19704,N_17080);
and UO_2474 (O_2474,N_19175,N_17807);
or UO_2475 (O_2475,N_18543,N_19834);
and UO_2476 (O_2476,N_16254,N_19538);
or UO_2477 (O_2477,N_17924,N_19737);
or UO_2478 (O_2478,N_17241,N_18868);
or UO_2479 (O_2479,N_17955,N_16107);
and UO_2480 (O_2480,N_19170,N_19705);
nand UO_2481 (O_2481,N_19476,N_16809);
nor UO_2482 (O_2482,N_19530,N_17722);
or UO_2483 (O_2483,N_19344,N_17752);
or UO_2484 (O_2484,N_19666,N_16428);
or UO_2485 (O_2485,N_19322,N_19703);
nand UO_2486 (O_2486,N_19543,N_17790);
xnor UO_2487 (O_2487,N_19869,N_16799);
nand UO_2488 (O_2488,N_19038,N_17945);
or UO_2489 (O_2489,N_18854,N_18794);
and UO_2490 (O_2490,N_17897,N_19296);
or UO_2491 (O_2491,N_18167,N_17275);
and UO_2492 (O_2492,N_18460,N_17458);
nor UO_2493 (O_2493,N_16488,N_16738);
xor UO_2494 (O_2494,N_19930,N_17256);
and UO_2495 (O_2495,N_19783,N_16914);
xnor UO_2496 (O_2496,N_16691,N_16882);
or UO_2497 (O_2497,N_19343,N_18703);
nor UO_2498 (O_2498,N_17001,N_17904);
and UO_2499 (O_2499,N_16293,N_18259);
endmodule