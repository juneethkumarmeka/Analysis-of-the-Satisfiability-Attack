module basic_750_5000_1000_10_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_76,In_82);
nor U1 (N_1,In_578,In_245);
or U2 (N_2,In_207,In_404);
nand U3 (N_3,In_191,In_583);
nand U4 (N_4,In_406,In_584);
nor U5 (N_5,In_201,In_73);
nor U6 (N_6,In_87,In_74);
or U7 (N_7,In_546,In_239);
nor U8 (N_8,In_261,In_125);
nor U9 (N_9,In_374,In_375);
xnor U10 (N_10,In_695,In_124);
and U11 (N_11,In_480,In_250);
or U12 (N_12,In_506,In_420);
xnor U13 (N_13,In_351,In_711);
or U14 (N_14,In_320,In_220);
nor U15 (N_15,In_276,In_716);
nand U16 (N_16,In_29,In_52);
nand U17 (N_17,In_311,In_321);
or U18 (N_18,In_241,In_461);
and U19 (N_19,In_453,In_113);
nand U20 (N_20,In_408,In_660);
and U21 (N_21,In_413,In_447);
nor U22 (N_22,In_2,In_189);
and U23 (N_23,In_312,In_723);
or U24 (N_24,In_460,In_53);
and U25 (N_25,In_91,In_496);
and U26 (N_26,In_720,In_535);
and U27 (N_27,In_180,In_565);
or U28 (N_28,In_636,In_418);
or U29 (N_29,In_89,In_302);
nor U30 (N_30,In_146,In_649);
and U31 (N_31,In_121,In_463);
nand U32 (N_32,In_120,In_279);
and U33 (N_33,In_514,In_209);
nand U34 (N_34,In_254,In_140);
and U35 (N_35,In_267,In_203);
or U36 (N_36,In_541,In_448);
xor U37 (N_37,In_223,In_296);
nor U38 (N_38,In_611,In_15);
or U39 (N_39,In_627,In_145);
nand U40 (N_40,In_466,In_462);
and U41 (N_41,In_334,In_661);
or U42 (N_42,In_260,In_364);
and U43 (N_43,In_589,In_727);
or U44 (N_44,In_316,In_475);
or U45 (N_45,In_456,In_370);
nor U46 (N_46,In_603,In_28);
xnor U47 (N_47,In_542,In_679);
nor U48 (N_48,In_645,In_304);
and U49 (N_49,In_629,In_634);
nand U50 (N_50,In_118,In_687);
nor U51 (N_51,In_468,In_152);
nor U52 (N_52,In_739,In_188);
and U53 (N_53,In_104,In_652);
and U54 (N_54,In_299,In_508);
or U55 (N_55,In_459,In_534);
nand U56 (N_56,In_399,In_479);
nand U57 (N_57,In_333,In_740);
and U58 (N_58,In_536,In_30);
or U59 (N_59,In_33,In_186);
nor U60 (N_60,In_600,In_274);
nand U61 (N_61,In_748,In_693);
or U62 (N_62,In_582,In_544);
or U63 (N_63,In_150,In_114);
or U64 (N_64,In_577,In_19);
and U65 (N_65,In_81,In_439);
nand U66 (N_66,In_470,In_482);
nand U67 (N_67,In_651,In_379);
nor U68 (N_68,In_731,In_707);
or U69 (N_69,In_605,In_95);
or U70 (N_70,In_77,In_474);
or U71 (N_71,In_571,In_719);
nand U72 (N_72,In_623,In_292);
and U73 (N_73,In_366,In_510);
and U74 (N_74,In_289,In_182);
nor U75 (N_75,In_123,In_653);
or U76 (N_76,In_252,In_174);
nor U77 (N_77,In_458,In_561);
nor U78 (N_78,In_166,In_708);
or U79 (N_79,In_669,In_243);
nand U80 (N_80,In_197,In_255);
nand U81 (N_81,In_725,In_110);
nand U82 (N_82,In_92,In_18);
nor U83 (N_83,In_512,In_677);
xor U84 (N_84,In_103,In_56);
or U85 (N_85,In_643,In_338);
nor U86 (N_86,In_38,In_354);
nand U87 (N_87,In_200,In_49);
nand U88 (N_88,In_410,In_13);
xor U89 (N_89,In_230,In_607);
and U90 (N_90,In_69,In_412);
or U91 (N_91,In_240,In_171);
nor U92 (N_92,In_728,In_135);
nor U93 (N_93,In_131,In_79);
nor U94 (N_94,In_489,In_601);
nand U95 (N_95,In_397,In_105);
nor U96 (N_96,In_694,In_699);
nor U97 (N_97,In_390,In_175);
or U98 (N_98,In_3,In_327);
or U99 (N_99,In_88,In_684);
and U100 (N_100,In_268,In_342);
xnor U101 (N_101,In_386,In_628);
nand U102 (N_102,In_575,In_117);
nand U103 (N_103,In_360,In_293);
nand U104 (N_104,In_646,In_572);
nand U105 (N_105,In_216,In_663);
and U106 (N_106,In_564,In_516);
nor U107 (N_107,In_288,In_256);
xor U108 (N_108,In_648,In_503);
or U109 (N_109,In_291,In_185);
and U110 (N_110,In_560,In_372);
or U111 (N_111,In_116,In_137);
and U112 (N_112,In_437,In_11);
or U113 (N_113,In_706,In_586);
nand U114 (N_114,In_164,In_314);
nor U115 (N_115,In_501,In_637);
xnor U116 (N_116,In_407,In_734);
nor U117 (N_117,In_148,In_562);
and U118 (N_118,In_610,In_395);
nand U119 (N_119,In_259,In_184);
nand U120 (N_120,In_668,In_724);
or U121 (N_121,In_278,In_10);
or U122 (N_122,In_615,In_313);
nor U123 (N_123,In_635,In_157);
and U124 (N_124,In_242,In_672);
or U125 (N_125,In_445,In_570);
or U126 (N_126,In_402,In_322);
and U127 (N_127,In_494,In_234);
nand U128 (N_128,In_509,In_698);
and U129 (N_129,In_51,In_317);
nand U130 (N_130,In_48,In_68);
and U131 (N_131,In_323,In_27);
xor U132 (N_132,In_67,In_625);
xnor U133 (N_133,In_650,In_746);
xnor U134 (N_134,In_591,In_165);
xnor U135 (N_135,In_31,In_553);
and U136 (N_136,In_657,In_326);
and U137 (N_137,In_537,In_128);
nor U138 (N_138,In_225,In_490);
or U139 (N_139,In_294,In_219);
or U140 (N_140,In_282,In_613);
xnor U141 (N_141,In_232,In_331);
nand U142 (N_142,In_499,In_290);
or U143 (N_143,In_609,In_540);
nor U144 (N_144,In_45,In_674);
nor U145 (N_145,In_251,In_336);
nor U146 (N_146,In_99,In_396);
nand U147 (N_147,In_181,In_258);
xor U148 (N_148,In_658,In_446);
nor U149 (N_149,In_491,In_484);
and U150 (N_150,In_376,In_54);
and U151 (N_151,In_218,In_35);
xor U152 (N_152,In_692,In_384);
nand U153 (N_153,In_476,In_112);
or U154 (N_154,In_617,In_696);
and U155 (N_155,In_23,In_587);
and U156 (N_156,In_233,In_359);
and U157 (N_157,In_744,In_332);
xor U158 (N_158,In_271,In_743);
nand U159 (N_159,In_551,In_283);
and U160 (N_160,In_75,In_97);
or U161 (N_161,In_626,In_107);
and U162 (N_162,In_556,In_50);
nor U163 (N_163,In_210,In_214);
nor U164 (N_164,In_513,In_705);
nand U165 (N_165,In_738,In_688);
and U166 (N_166,In_249,In_83);
and U167 (N_167,In_43,In_524);
nand U168 (N_168,In_640,In_340);
xnor U169 (N_169,In_548,In_173);
nor U170 (N_170,In_409,In_170);
nor U171 (N_171,In_655,In_477);
or U172 (N_172,In_25,In_525);
and U173 (N_173,In_298,In_20);
or U174 (N_174,In_452,In_394);
and U175 (N_175,In_337,In_427);
nand U176 (N_176,In_63,In_388);
xor U177 (N_177,In_741,In_248);
nand U178 (N_178,In_574,In_523);
nor U179 (N_179,In_487,In_358);
and U180 (N_180,In_6,In_295);
or U181 (N_181,In_502,In_208);
or U182 (N_182,In_141,In_328);
nor U183 (N_183,In_193,In_57);
nand U184 (N_184,In_495,In_155);
and U185 (N_185,In_17,In_465);
or U186 (N_186,In_133,In_159);
nand U187 (N_187,In_391,In_66);
nor U188 (N_188,In_40,In_347);
nand U189 (N_189,In_659,In_675);
nand U190 (N_190,In_417,In_485);
or U191 (N_191,In_378,In_136);
nand U192 (N_192,In_9,In_401);
nand U193 (N_193,In_498,In_325);
nand U194 (N_194,In_127,In_156);
and U195 (N_195,In_425,In_139);
nor U196 (N_196,In_444,In_287);
xor U197 (N_197,In_265,In_212);
or U198 (N_198,In_481,In_455);
or U199 (N_199,In_472,In_576);
and U200 (N_200,In_163,In_377);
nor U201 (N_201,In_85,In_319);
nor U202 (N_202,In_62,In_567);
and U203 (N_203,In_202,In_639);
nand U204 (N_204,In_531,In_341);
or U205 (N_205,In_604,In_37);
xor U206 (N_206,In_533,In_348);
and U207 (N_207,In_528,In_65);
nand U208 (N_208,In_438,In_196);
xor U209 (N_209,In_573,In_700);
and U210 (N_210,In_579,In_64);
and U211 (N_211,In_729,In_735);
and U212 (N_212,In_606,In_400);
nor U213 (N_213,In_60,In_108);
nor U214 (N_214,In_682,In_428);
and U215 (N_215,In_365,In_593);
or U216 (N_216,In_78,In_500);
nand U217 (N_217,In_109,In_229);
nand U218 (N_218,In_547,In_690);
or U219 (N_219,In_227,In_36);
and U220 (N_220,In_151,In_493);
or U221 (N_221,In_622,In_147);
or U222 (N_222,In_471,In_46);
nand U223 (N_223,In_411,In_1);
xnor U224 (N_224,In_632,In_594);
nor U225 (N_225,In_12,In_596);
nand U226 (N_226,In_614,In_72);
or U227 (N_227,In_671,In_310);
nand U228 (N_228,In_329,In_722);
nand U229 (N_229,In_70,In_599);
and U230 (N_230,In_231,In_270);
and U231 (N_231,In_588,In_612);
and U232 (N_232,In_416,In_530);
or U233 (N_233,In_32,In_697);
nor U234 (N_234,In_733,In_205);
nor U235 (N_235,In_161,In_308);
and U236 (N_236,In_335,In_122);
or U237 (N_237,In_608,In_309);
or U238 (N_238,In_736,In_176);
nor U239 (N_239,In_177,In_264);
xnor U240 (N_240,In_507,In_221);
or U241 (N_241,In_247,In_14);
and U242 (N_242,In_442,In_190);
nor U243 (N_243,In_158,In_633);
nor U244 (N_244,In_297,In_478);
or U245 (N_245,In_59,In_642);
and U246 (N_246,In_415,In_443);
and U247 (N_247,In_419,In_620);
xnor U248 (N_248,In_681,In_747);
or U249 (N_249,In_630,In_689);
and U250 (N_250,In_539,In_520);
nand U251 (N_251,In_228,In_441);
or U252 (N_252,In_664,In_519);
nor U253 (N_253,In_450,In_262);
nand U254 (N_254,In_497,In_285);
nand U255 (N_255,In_616,In_430);
and U256 (N_256,In_621,In_4);
or U257 (N_257,In_488,In_300);
nor U258 (N_258,In_451,In_685);
nand U259 (N_259,In_44,In_80);
xnor U260 (N_260,In_701,In_5);
and U261 (N_261,In_143,In_8);
and U262 (N_262,In_580,In_550);
and U263 (N_263,In_144,In_730);
nor U264 (N_264,In_330,In_592);
nand U265 (N_265,In_709,In_115);
and U266 (N_266,In_71,In_432);
or U267 (N_267,In_492,In_126);
or U268 (N_268,In_387,In_380);
and U269 (N_269,In_710,In_263);
or U270 (N_270,In_449,In_538);
nor U271 (N_271,In_371,In_742);
and U272 (N_272,In_194,In_269);
or U273 (N_273,In_367,In_585);
nor U274 (N_274,In_119,In_713);
and U275 (N_275,In_486,In_686);
nand U276 (N_276,In_349,In_702);
xnor U277 (N_277,In_206,In_353);
nor U278 (N_278,In_426,In_369);
or U279 (N_279,In_324,In_745);
or U280 (N_280,In_315,In_597);
or U281 (N_281,In_673,In_26);
and U282 (N_282,In_22,In_339);
and U283 (N_283,In_421,In_93);
and U284 (N_284,In_41,In_715);
or U285 (N_285,In_244,In_134);
nand U286 (N_286,In_129,In_732);
nand U287 (N_287,In_281,In_718);
or U288 (N_288,In_721,In_467);
or U289 (N_289,In_667,In_624);
and U290 (N_290,In_0,In_368);
and U291 (N_291,In_142,In_350);
nor U292 (N_292,In_557,In_505);
nor U293 (N_293,In_153,In_187);
nor U294 (N_294,In_749,In_346);
nand U295 (N_295,In_101,In_138);
and U296 (N_296,In_383,In_47);
or U297 (N_297,In_96,In_195);
nand U298 (N_298,In_257,In_559);
nor U299 (N_299,In_435,In_618);
and U300 (N_300,In_464,In_381);
nand U301 (N_301,In_529,In_34);
and U302 (N_302,In_280,In_98);
nor U303 (N_303,In_393,In_273);
xnor U304 (N_304,In_179,In_222);
and U305 (N_305,In_566,In_130);
nand U306 (N_306,In_7,In_554);
xnor U307 (N_307,In_392,In_178);
nand U308 (N_308,In_457,In_215);
and U309 (N_309,In_301,In_86);
nand U310 (N_310,In_717,In_595);
or U311 (N_311,In_414,In_665);
or U312 (N_312,In_305,In_382);
and U313 (N_313,In_473,In_226);
nand U314 (N_314,In_198,In_363);
or U315 (N_315,In_211,In_581);
nor U316 (N_316,In_545,In_238);
or U317 (N_317,In_403,In_39);
and U318 (N_318,In_199,In_429);
or U319 (N_319,In_16,In_436);
nand U320 (N_320,In_106,In_527);
and U321 (N_321,In_84,In_355);
or U322 (N_322,In_100,In_431);
or U323 (N_323,In_555,In_680);
xnor U324 (N_324,In_726,In_666);
xor U325 (N_325,In_94,In_224);
or U326 (N_326,In_149,In_469);
nand U327 (N_327,In_306,In_602);
or U328 (N_328,In_483,In_24);
and U329 (N_329,In_237,In_504);
or U330 (N_330,In_638,In_284);
and U331 (N_331,In_286,In_517);
nor U332 (N_332,In_691,In_356);
or U333 (N_333,In_631,In_521);
and U334 (N_334,In_678,In_373);
or U335 (N_335,In_422,In_132);
xor U336 (N_336,In_204,In_357);
xnor U337 (N_337,In_213,In_307);
nand U338 (N_338,In_558,In_552);
and U339 (N_339,In_352,In_434);
xnor U340 (N_340,In_361,In_511);
nor U341 (N_341,In_303,In_102);
or U342 (N_342,In_42,In_569);
xnor U343 (N_343,In_235,In_568);
xnor U344 (N_344,In_160,In_162);
nor U345 (N_345,In_345,In_253);
nor U346 (N_346,In_440,In_590);
or U347 (N_347,In_670,In_169);
nand U348 (N_348,In_21,In_424);
or U349 (N_349,In_423,In_362);
or U350 (N_350,In_192,In_58);
nand U351 (N_351,In_389,In_714);
nand U352 (N_352,In_704,In_167);
xor U353 (N_353,In_236,In_676);
nor U354 (N_354,In_641,In_433);
nand U355 (N_355,In_61,In_277);
and U356 (N_356,In_662,In_737);
nor U357 (N_357,In_549,In_217);
nand U358 (N_358,In_385,In_522);
nor U359 (N_359,In_168,In_644);
nand U360 (N_360,In_454,In_172);
and U361 (N_361,In_55,In_154);
xor U362 (N_362,In_647,In_246);
nor U363 (N_363,In_272,In_654);
and U364 (N_364,In_275,In_598);
nor U365 (N_365,In_266,In_405);
and U366 (N_366,In_563,In_183);
or U367 (N_367,In_656,In_398);
or U368 (N_368,In_344,In_683);
or U369 (N_369,In_526,In_703);
xor U370 (N_370,In_712,In_518);
nand U371 (N_371,In_90,In_619);
nor U372 (N_372,In_543,In_318);
or U373 (N_373,In_532,In_515);
and U374 (N_374,In_343,In_111);
nand U375 (N_375,In_144,In_104);
or U376 (N_376,In_243,In_483);
nor U377 (N_377,In_91,In_112);
or U378 (N_378,In_433,In_163);
nand U379 (N_379,In_608,In_599);
xnor U380 (N_380,In_153,In_134);
and U381 (N_381,In_176,In_195);
and U382 (N_382,In_102,In_278);
xor U383 (N_383,In_679,In_42);
nor U384 (N_384,In_604,In_80);
nor U385 (N_385,In_256,In_632);
nor U386 (N_386,In_196,In_48);
and U387 (N_387,In_667,In_559);
xor U388 (N_388,In_182,In_569);
and U389 (N_389,In_507,In_544);
nor U390 (N_390,In_106,In_556);
xnor U391 (N_391,In_160,In_655);
nor U392 (N_392,In_292,In_712);
nand U393 (N_393,In_203,In_570);
nand U394 (N_394,In_185,In_363);
or U395 (N_395,In_606,In_201);
or U396 (N_396,In_609,In_305);
or U397 (N_397,In_700,In_273);
and U398 (N_398,In_3,In_79);
nor U399 (N_399,In_459,In_139);
nand U400 (N_400,In_375,In_476);
xnor U401 (N_401,In_442,In_149);
nor U402 (N_402,In_564,In_268);
and U403 (N_403,In_363,In_552);
or U404 (N_404,In_679,In_421);
and U405 (N_405,In_684,In_465);
nor U406 (N_406,In_192,In_374);
nor U407 (N_407,In_633,In_746);
or U408 (N_408,In_329,In_302);
and U409 (N_409,In_573,In_453);
or U410 (N_410,In_208,In_173);
nand U411 (N_411,In_697,In_331);
and U412 (N_412,In_439,In_549);
or U413 (N_413,In_724,In_161);
and U414 (N_414,In_561,In_703);
and U415 (N_415,In_111,In_286);
or U416 (N_416,In_122,In_493);
and U417 (N_417,In_311,In_165);
xnor U418 (N_418,In_726,In_385);
and U419 (N_419,In_521,In_556);
and U420 (N_420,In_457,In_23);
nand U421 (N_421,In_160,In_246);
nand U422 (N_422,In_51,In_432);
nor U423 (N_423,In_336,In_181);
xor U424 (N_424,In_191,In_484);
or U425 (N_425,In_160,In_347);
nand U426 (N_426,In_637,In_602);
and U427 (N_427,In_700,In_385);
nor U428 (N_428,In_584,In_503);
nand U429 (N_429,In_143,In_80);
and U430 (N_430,In_138,In_108);
and U431 (N_431,In_305,In_555);
and U432 (N_432,In_218,In_165);
or U433 (N_433,In_681,In_270);
nand U434 (N_434,In_403,In_312);
xnor U435 (N_435,In_193,In_14);
and U436 (N_436,In_351,In_543);
or U437 (N_437,In_505,In_135);
and U438 (N_438,In_20,In_10);
or U439 (N_439,In_691,In_521);
and U440 (N_440,In_246,In_610);
and U441 (N_441,In_584,In_94);
or U442 (N_442,In_42,In_646);
or U443 (N_443,In_538,In_542);
or U444 (N_444,In_215,In_640);
and U445 (N_445,In_61,In_8);
and U446 (N_446,In_589,In_520);
and U447 (N_447,In_560,In_409);
and U448 (N_448,In_679,In_273);
nor U449 (N_449,In_523,In_106);
or U450 (N_450,In_144,In_557);
nor U451 (N_451,In_299,In_217);
nand U452 (N_452,In_681,In_329);
nor U453 (N_453,In_733,In_450);
nor U454 (N_454,In_114,In_134);
and U455 (N_455,In_107,In_458);
and U456 (N_456,In_404,In_563);
xnor U457 (N_457,In_194,In_519);
nor U458 (N_458,In_65,In_49);
and U459 (N_459,In_466,In_414);
nor U460 (N_460,In_91,In_477);
nor U461 (N_461,In_511,In_737);
and U462 (N_462,In_679,In_293);
nand U463 (N_463,In_269,In_447);
or U464 (N_464,In_477,In_703);
and U465 (N_465,In_325,In_158);
nor U466 (N_466,In_503,In_688);
or U467 (N_467,In_423,In_290);
or U468 (N_468,In_337,In_695);
or U469 (N_469,In_682,In_580);
nor U470 (N_470,In_245,In_570);
or U471 (N_471,In_259,In_454);
or U472 (N_472,In_394,In_471);
nor U473 (N_473,In_149,In_146);
or U474 (N_474,In_83,In_578);
nor U475 (N_475,In_381,In_506);
or U476 (N_476,In_82,In_602);
or U477 (N_477,In_298,In_512);
nor U478 (N_478,In_322,In_73);
or U479 (N_479,In_540,In_192);
nor U480 (N_480,In_557,In_596);
nand U481 (N_481,In_120,In_609);
xor U482 (N_482,In_651,In_225);
nor U483 (N_483,In_180,In_267);
nand U484 (N_484,In_32,In_546);
xor U485 (N_485,In_573,In_365);
nor U486 (N_486,In_30,In_561);
and U487 (N_487,In_9,In_26);
or U488 (N_488,In_265,In_548);
nand U489 (N_489,In_304,In_550);
or U490 (N_490,In_551,In_584);
and U491 (N_491,In_726,In_657);
nand U492 (N_492,In_180,In_380);
nor U493 (N_493,In_103,In_305);
or U494 (N_494,In_116,In_666);
and U495 (N_495,In_228,In_39);
and U496 (N_496,In_456,In_306);
nand U497 (N_497,In_710,In_206);
nor U498 (N_498,In_628,In_464);
or U499 (N_499,In_89,In_457);
and U500 (N_500,N_69,N_225);
and U501 (N_501,N_143,N_48);
nor U502 (N_502,N_487,N_207);
nand U503 (N_503,N_95,N_286);
nor U504 (N_504,N_302,N_218);
nand U505 (N_505,N_114,N_250);
xor U506 (N_506,N_97,N_20);
and U507 (N_507,N_192,N_493);
nor U508 (N_508,N_240,N_312);
or U509 (N_509,N_41,N_392);
and U510 (N_510,N_117,N_247);
xnor U511 (N_511,N_172,N_0);
xor U512 (N_512,N_319,N_469);
or U513 (N_513,N_40,N_138);
nor U514 (N_514,N_127,N_309);
nand U515 (N_515,N_166,N_416);
nand U516 (N_516,N_132,N_287);
nand U517 (N_517,N_393,N_373);
nor U518 (N_518,N_191,N_60);
or U519 (N_519,N_261,N_456);
and U520 (N_520,N_496,N_499);
nor U521 (N_521,N_93,N_107);
nand U522 (N_522,N_300,N_386);
or U523 (N_523,N_85,N_420);
nor U524 (N_524,N_355,N_10);
nand U525 (N_525,N_123,N_324);
nand U526 (N_526,N_485,N_494);
or U527 (N_527,N_448,N_238);
xor U528 (N_528,N_36,N_42);
nand U529 (N_529,N_360,N_446);
and U530 (N_530,N_246,N_118);
nand U531 (N_531,N_167,N_465);
and U532 (N_532,N_72,N_285);
nand U533 (N_533,N_176,N_136);
nand U534 (N_534,N_344,N_361);
and U535 (N_535,N_149,N_144);
or U536 (N_536,N_199,N_325);
nor U537 (N_537,N_243,N_29);
nand U538 (N_538,N_390,N_134);
nor U539 (N_539,N_466,N_337);
and U540 (N_540,N_327,N_347);
nand U541 (N_541,N_340,N_180);
nor U542 (N_542,N_489,N_55);
nand U543 (N_543,N_339,N_202);
nor U544 (N_544,N_151,N_258);
or U545 (N_545,N_230,N_46);
or U546 (N_546,N_495,N_220);
nand U547 (N_547,N_100,N_193);
nand U548 (N_548,N_184,N_183);
or U549 (N_549,N_375,N_450);
xnor U550 (N_550,N_307,N_231);
and U551 (N_551,N_451,N_275);
or U552 (N_552,N_256,N_387);
or U553 (N_553,N_237,N_61);
and U554 (N_554,N_162,N_471);
xor U555 (N_555,N_484,N_105);
and U556 (N_556,N_241,N_262);
nor U557 (N_557,N_81,N_457);
or U558 (N_558,N_379,N_370);
and U559 (N_559,N_481,N_27);
nand U560 (N_560,N_273,N_146);
or U561 (N_561,N_215,N_318);
nand U562 (N_562,N_388,N_259);
or U563 (N_563,N_188,N_413);
nor U564 (N_564,N_417,N_137);
nor U565 (N_565,N_98,N_263);
nand U566 (N_566,N_303,N_217);
nor U567 (N_567,N_89,N_242);
and U568 (N_568,N_77,N_179);
or U569 (N_569,N_122,N_251);
or U570 (N_570,N_43,N_236);
nand U571 (N_571,N_395,N_298);
nor U572 (N_572,N_75,N_274);
nand U573 (N_573,N_406,N_492);
nand U574 (N_574,N_78,N_56);
xor U575 (N_575,N_228,N_394);
and U576 (N_576,N_362,N_314);
or U577 (N_577,N_135,N_445);
or U578 (N_578,N_473,N_227);
xnor U579 (N_579,N_4,N_32);
or U580 (N_580,N_491,N_374);
nand U581 (N_581,N_226,N_99);
and U582 (N_582,N_21,N_208);
nand U583 (N_583,N_24,N_205);
xnor U584 (N_584,N_455,N_338);
nor U585 (N_585,N_443,N_358);
and U586 (N_586,N_234,N_345);
or U587 (N_587,N_64,N_354);
nand U588 (N_588,N_266,N_174);
nand U589 (N_589,N_15,N_350);
and U590 (N_590,N_197,N_323);
nand U591 (N_591,N_343,N_12);
and U592 (N_592,N_82,N_68);
nor U593 (N_593,N_164,N_433);
or U594 (N_594,N_201,N_463);
nor U595 (N_595,N_411,N_31);
xnor U596 (N_596,N_322,N_71);
or U597 (N_597,N_175,N_342);
xor U598 (N_598,N_67,N_128);
nor U599 (N_599,N_66,N_76);
nand U600 (N_600,N_313,N_356);
xor U601 (N_601,N_18,N_336);
xor U602 (N_602,N_235,N_378);
xnor U603 (N_603,N_497,N_131);
and U604 (N_604,N_468,N_434);
and U605 (N_605,N_369,N_139);
nor U606 (N_606,N_264,N_317);
or U607 (N_607,N_52,N_423);
or U608 (N_608,N_96,N_216);
and U609 (N_609,N_292,N_58);
nand U610 (N_610,N_452,N_357);
and U611 (N_611,N_165,N_209);
and U612 (N_612,N_331,N_321);
nor U613 (N_613,N_315,N_70);
or U614 (N_614,N_346,N_16);
nand U615 (N_615,N_59,N_39);
nand U616 (N_616,N_441,N_204);
and U617 (N_617,N_190,N_480);
nand U618 (N_618,N_133,N_163);
nor U619 (N_619,N_116,N_87);
nand U620 (N_620,N_383,N_25);
nor U621 (N_621,N_368,N_291);
or U622 (N_622,N_474,N_8);
nand U623 (N_623,N_173,N_245);
or U624 (N_624,N_414,N_341);
nor U625 (N_625,N_92,N_442);
nor U626 (N_626,N_129,N_156);
nor U627 (N_627,N_294,N_429);
or U628 (N_628,N_410,N_115);
and U629 (N_629,N_419,N_301);
nor U630 (N_630,N_83,N_399);
or U631 (N_631,N_408,N_308);
nand U632 (N_632,N_73,N_425);
nor U633 (N_633,N_203,N_380);
xnor U634 (N_634,N_145,N_295);
xnor U635 (N_635,N_415,N_289);
nand U636 (N_636,N_351,N_65);
nand U637 (N_637,N_224,N_35);
or U638 (N_638,N_112,N_11);
nor U639 (N_639,N_462,N_372);
xnor U640 (N_640,N_185,N_57);
or U641 (N_641,N_439,N_293);
and U642 (N_642,N_44,N_470);
or U643 (N_643,N_283,N_219);
and U644 (N_644,N_424,N_158);
xor U645 (N_645,N_421,N_498);
xnor U646 (N_646,N_282,N_459);
or U647 (N_647,N_486,N_189);
nor U648 (N_648,N_169,N_161);
nor U649 (N_649,N_402,N_430);
nand U650 (N_650,N_53,N_460);
nand U651 (N_651,N_353,N_104);
and U652 (N_652,N_221,N_329);
nand U653 (N_653,N_80,N_453);
and U654 (N_654,N_147,N_148);
xor U655 (N_655,N_14,N_458);
nor U656 (N_656,N_454,N_2);
and U657 (N_657,N_478,N_349);
and U658 (N_658,N_479,N_63);
nor U659 (N_659,N_120,N_38);
and U660 (N_660,N_384,N_400);
nor U661 (N_661,N_299,N_196);
or U662 (N_662,N_348,N_332);
nand U663 (N_663,N_113,N_124);
nand U664 (N_664,N_271,N_428);
or U665 (N_665,N_49,N_396);
or U666 (N_666,N_9,N_385);
and U667 (N_667,N_13,N_320);
and U668 (N_668,N_270,N_449);
nor U669 (N_669,N_277,N_160);
or U670 (N_670,N_391,N_33);
nor U671 (N_671,N_440,N_381);
nand U672 (N_672,N_22,N_377);
and U673 (N_673,N_126,N_418);
and U674 (N_674,N_267,N_19);
nand U675 (N_675,N_382,N_244);
or U676 (N_676,N_106,N_367);
xor U677 (N_677,N_426,N_482);
nor U678 (N_678,N_28,N_488);
and U679 (N_679,N_431,N_407);
or U680 (N_680,N_141,N_476);
and U681 (N_681,N_279,N_3);
nor U682 (N_682,N_194,N_50);
nand U683 (N_683,N_306,N_290);
xor U684 (N_684,N_397,N_252);
and U685 (N_685,N_51,N_310);
or U686 (N_686,N_376,N_437);
and U687 (N_687,N_109,N_86);
or U688 (N_688,N_359,N_154);
nor U689 (N_689,N_371,N_366);
nand U690 (N_690,N_444,N_363);
and U691 (N_691,N_278,N_422);
nor U692 (N_692,N_88,N_30);
and U693 (N_693,N_90,N_281);
nor U694 (N_694,N_438,N_404);
xnor U695 (N_695,N_206,N_125);
nor U696 (N_696,N_435,N_171);
and U697 (N_697,N_436,N_405);
xor U698 (N_698,N_157,N_467);
and U699 (N_699,N_178,N_398);
nor U700 (N_700,N_79,N_26);
nand U701 (N_701,N_47,N_182);
nand U702 (N_702,N_74,N_364);
nor U703 (N_703,N_260,N_5);
nor U704 (N_704,N_365,N_181);
and U705 (N_705,N_311,N_326);
xor U706 (N_706,N_153,N_297);
nand U707 (N_707,N_239,N_475);
nand U708 (N_708,N_142,N_200);
or U709 (N_709,N_229,N_140);
nor U710 (N_710,N_130,N_54);
nand U711 (N_711,N_211,N_401);
and U712 (N_712,N_37,N_62);
and U713 (N_713,N_472,N_17);
nor U714 (N_714,N_102,N_272);
and U715 (N_715,N_152,N_233);
and U716 (N_716,N_403,N_269);
nor U717 (N_717,N_352,N_432);
and U718 (N_718,N_409,N_177);
and U719 (N_719,N_150,N_84);
nand U720 (N_720,N_335,N_255);
or U721 (N_721,N_296,N_257);
xor U722 (N_722,N_305,N_121);
and U723 (N_723,N_108,N_254);
nand U724 (N_724,N_111,N_333);
and U725 (N_725,N_170,N_119);
or U726 (N_726,N_198,N_34);
nand U727 (N_727,N_101,N_23);
and U728 (N_728,N_212,N_248);
nor U729 (N_729,N_284,N_483);
nor U730 (N_730,N_276,N_223);
and U731 (N_731,N_155,N_249);
nand U732 (N_732,N_330,N_213);
nor U733 (N_733,N_6,N_490);
and U734 (N_734,N_412,N_447);
or U735 (N_735,N_461,N_210);
nand U736 (N_736,N_1,N_477);
or U737 (N_737,N_328,N_288);
nor U738 (N_738,N_186,N_232);
nand U739 (N_739,N_304,N_103);
xnor U740 (N_740,N_168,N_94);
nor U741 (N_741,N_389,N_187);
or U742 (N_742,N_253,N_464);
nor U743 (N_743,N_280,N_45);
xor U744 (N_744,N_222,N_91);
nor U745 (N_745,N_195,N_265);
xor U746 (N_746,N_334,N_7);
or U747 (N_747,N_159,N_268);
nand U748 (N_748,N_214,N_316);
nand U749 (N_749,N_427,N_110);
and U750 (N_750,N_178,N_23);
nand U751 (N_751,N_74,N_391);
nor U752 (N_752,N_279,N_474);
xor U753 (N_753,N_13,N_265);
or U754 (N_754,N_162,N_88);
nor U755 (N_755,N_272,N_160);
nor U756 (N_756,N_205,N_486);
nand U757 (N_757,N_466,N_441);
xnor U758 (N_758,N_447,N_242);
nand U759 (N_759,N_284,N_300);
and U760 (N_760,N_366,N_223);
nand U761 (N_761,N_230,N_305);
xor U762 (N_762,N_88,N_248);
nor U763 (N_763,N_57,N_133);
nand U764 (N_764,N_29,N_492);
nor U765 (N_765,N_185,N_470);
or U766 (N_766,N_30,N_54);
nor U767 (N_767,N_422,N_207);
or U768 (N_768,N_201,N_173);
nor U769 (N_769,N_131,N_68);
nand U770 (N_770,N_383,N_15);
nor U771 (N_771,N_110,N_499);
nand U772 (N_772,N_163,N_36);
nor U773 (N_773,N_390,N_102);
nand U774 (N_774,N_177,N_69);
or U775 (N_775,N_255,N_111);
or U776 (N_776,N_351,N_105);
or U777 (N_777,N_418,N_146);
nand U778 (N_778,N_25,N_26);
nor U779 (N_779,N_153,N_12);
nand U780 (N_780,N_319,N_326);
xnor U781 (N_781,N_218,N_400);
nand U782 (N_782,N_323,N_174);
nor U783 (N_783,N_193,N_22);
nand U784 (N_784,N_480,N_259);
xnor U785 (N_785,N_349,N_352);
nand U786 (N_786,N_288,N_369);
xnor U787 (N_787,N_35,N_254);
or U788 (N_788,N_54,N_183);
xnor U789 (N_789,N_457,N_453);
or U790 (N_790,N_113,N_417);
or U791 (N_791,N_248,N_351);
or U792 (N_792,N_118,N_435);
nor U793 (N_793,N_301,N_237);
nor U794 (N_794,N_225,N_103);
nor U795 (N_795,N_369,N_119);
nor U796 (N_796,N_4,N_482);
or U797 (N_797,N_301,N_236);
nand U798 (N_798,N_114,N_439);
nand U799 (N_799,N_318,N_52);
or U800 (N_800,N_107,N_32);
or U801 (N_801,N_421,N_131);
nand U802 (N_802,N_205,N_52);
nand U803 (N_803,N_195,N_162);
nor U804 (N_804,N_261,N_339);
or U805 (N_805,N_159,N_261);
nor U806 (N_806,N_135,N_248);
nand U807 (N_807,N_133,N_16);
or U808 (N_808,N_114,N_279);
nor U809 (N_809,N_165,N_252);
nand U810 (N_810,N_78,N_25);
or U811 (N_811,N_5,N_45);
and U812 (N_812,N_278,N_26);
nand U813 (N_813,N_377,N_103);
nand U814 (N_814,N_410,N_339);
nand U815 (N_815,N_17,N_401);
and U816 (N_816,N_417,N_204);
and U817 (N_817,N_28,N_45);
or U818 (N_818,N_251,N_68);
nor U819 (N_819,N_470,N_265);
or U820 (N_820,N_426,N_257);
nor U821 (N_821,N_248,N_442);
and U822 (N_822,N_5,N_448);
and U823 (N_823,N_303,N_344);
nand U824 (N_824,N_219,N_498);
or U825 (N_825,N_450,N_171);
nor U826 (N_826,N_107,N_303);
nand U827 (N_827,N_415,N_12);
nor U828 (N_828,N_327,N_382);
nor U829 (N_829,N_316,N_477);
nor U830 (N_830,N_24,N_168);
or U831 (N_831,N_168,N_480);
xnor U832 (N_832,N_76,N_198);
or U833 (N_833,N_210,N_376);
nand U834 (N_834,N_211,N_44);
or U835 (N_835,N_76,N_163);
nor U836 (N_836,N_391,N_468);
nand U837 (N_837,N_396,N_294);
xor U838 (N_838,N_216,N_146);
nor U839 (N_839,N_161,N_316);
xnor U840 (N_840,N_360,N_10);
xnor U841 (N_841,N_163,N_148);
nand U842 (N_842,N_462,N_84);
or U843 (N_843,N_357,N_325);
nor U844 (N_844,N_364,N_158);
nor U845 (N_845,N_50,N_460);
xnor U846 (N_846,N_313,N_80);
and U847 (N_847,N_355,N_211);
nor U848 (N_848,N_285,N_221);
and U849 (N_849,N_451,N_47);
nor U850 (N_850,N_118,N_139);
and U851 (N_851,N_82,N_413);
nor U852 (N_852,N_71,N_397);
or U853 (N_853,N_67,N_20);
and U854 (N_854,N_203,N_455);
or U855 (N_855,N_53,N_181);
and U856 (N_856,N_276,N_181);
and U857 (N_857,N_483,N_31);
xnor U858 (N_858,N_404,N_474);
xor U859 (N_859,N_49,N_245);
nor U860 (N_860,N_450,N_322);
nor U861 (N_861,N_441,N_446);
or U862 (N_862,N_206,N_226);
and U863 (N_863,N_378,N_232);
and U864 (N_864,N_267,N_327);
nor U865 (N_865,N_448,N_364);
nor U866 (N_866,N_256,N_422);
nor U867 (N_867,N_85,N_166);
nand U868 (N_868,N_304,N_181);
nor U869 (N_869,N_245,N_386);
and U870 (N_870,N_146,N_150);
nand U871 (N_871,N_182,N_283);
xnor U872 (N_872,N_115,N_193);
nor U873 (N_873,N_123,N_302);
nor U874 (N_874,N_305,N_70);
and U875 (N_875,N_476,N_173);
and U876 (N_876,N_398,N_143);
nand U877 (N_877,N_133,N_137);
nand U878 (N_878,N_450,N_14);
xnor U879 (N_879,N_130,N_478);
or U880 (N_880,N_221,N_10);
xnor U881 (N_881,N_323,N_400);
nor U882 (N_882,N_84,N_166);
nand U883 (N_883,N_14,N_152);
nor U884 (N_884,N_363,N_474);
or U885 (N_885,N_426,N_140);
nand U886 (N_886,N_154,N_72);
or U887 (N_887,N_124,N_411);
nor U888 (N_888,N_46,N_115);
or U889 (N_889,N_242,N_64);
xnor U890 (N_890,N_422,N_478);
and U891 (N_891,N_378,N_149);
xor U892 (N_892,N_480,N_10);
or U893 (N_893,N_0,N_230);
nor U894 (N_894,N_476,N_77);
nand U895 (N_895,N_230,N_283);
or U896 (N_896,N_45,N_367);
or U897 (N_897,N_338,N_495);
nor U898 (N_898,N_365,N_388);
and U899 (N_899,N_341,N_419);
nand U900 (N_900,N_171,N_108);
nand U901 (N_901,N_396,N_9);
nand U902 (N_902,N_177,N_238);
nand U903 (N_903,N_238,N_382);
nand U904 (N_904,N_109,N_120);
nor U905 (N_905,N_430,N_408);
or U906 (N_906,N_75,N_52);
nor U907 (N_907,N_169,N_34);
nand U908 (N_908,N_430,N_413);
xor U909 (N_909,N_119,N_489);
nor U910 (N_910,N_471,N_316);
nand U911 (N_911,N_458,N_135);
or U912 (N_912,N_474,N_453);
nor U913 (N_913,N_217,N_59);
and U914 (N_914,N_378,N_483);
nand U915 (N_915,N_203,N_312);
nor U916 (N_916,N_96,N_450);
or U917 (N_917,N_421,N_138);
nand U918 (N_918,N_42,N_154);
or U919 (N_919,N_167,N_57);
and U920 (N_920,N_362,N_338);
and U921 (N_921,N_179,N_487);
or U922 (N_922,N_416,N_335);
or U923 (N_923,N_467,N_268);
or U924 (N_924,N_129,N_303);
and U925 (N_925,N_43,N_207);
or U926 (N_926,N_476,N_351);
xor U927 (N_927,N_190,N_110);
and U928 (N_928,N_182,N_246);
and U929 (N_929,N_296,N_326);
and U930 (N_930,N_288,N_188);
nand U931 (N_931,N_45,N_454);
nor U932 (N_932,N_417,N_279);
xnor U933 (N_933,N_288,N_248);
and U934 (N_934,N_10,N_402);
and U935 (N_935,N_36,N_269);
nor U936 (N_936,N_67,N_347);
or U937 (N_937,N_183,N_327);
and U938 (N_938,N_235,N_429);
or U939 (N_939,N_315,N_247);
xor U940 (N_940,N_13,N_47);
nand U941 (N_941,N_333,N_262);
or U942 (N_942,N_427,N_36);
nand U943 (N_943,N_314,N_366);
nand U944 (N_944,N_285,N_9);
and U945 (N_945,N_75,N_188);
xor U946 (N_946,N_109,N_244);
and U947 (N_947,N_401,N_361);
or U948 (N_948,N_378,N_396);
or U949 (N_949,N_29,N_63);
nor U950 (N_950,N_136,N_43);
or U951 (N_951,N_198,N_356);
nor U952 (N_952,N_257,N_345);
and U953 (N_953,N_138,N_268);
and U954 (N_954,N_77,N_453);
xor U955 (N_955,N_403,N_327);
and U956 (N_956,N_105,N_86);
nor U957 (N_957,N_440,N_466);
nand U958 (N_958,N_265,N_476);
and U959 (N_959,N_29,N_431);
nor U960 (N_960,N_451,N_100);
or U961 (N_961,N_242,N_310);
xnor U962 (N_962,N_487,N_131);
and U963 (N_963,N_378,N_16);
and U964 (N_964,N_494,N_314);
nor U965 (N_965,N_52,N_166);
xnor U966 (N_966,N_407,N_174);
and U967 (N_967,N_461,N_28);
or U968 (N_968,N_10,N_339);
and U969 (N_969,N_169,N_244);
and U970 (N_970,N_313,N_23);
or U971 (N_971,N_272,N_38);
and U972 (N_972,N_205,N_244);
nor U973 (N_973,N_155,N_40);
nor U974 (N_974,N_57,N_495);
nor U975 (N_975,N_272,N_391);
nor U976 (N_976,N_307,N_412);
nor U977 (N_977,N_117,N_206);
nand U978 (N_978,N_219,N_441);
or U979 (N_979,N_439,N_309);
or U980 (N_980,N_356,N_298);
nor U981 (N_981,N_10,N_414);
or U982 (N_982,N_222,N_236);
xnor U983 (N_983,N_401,N_61);
nor U984 (N_984,N_390,N_419);
and U985 (N_985,N_247,N_335);
or U986 (N_986,N_2,N_448);
nor U987 (N_987,N_173,N_171);
nand U988 (N_988,N_18,N_49);
nand U989 (N_989,N_456,N_123);
nor U990 (N_990,N_226,N_316);
or U991 (N_991,N_179,N_281);
nand U992 (N_992,N_389,N_346);
or U993 (N_993,N_13,N_72);
xor U994 (N_994,N_341,N_295);
nor U995 (N_995,N_339,N_95);
or U996 (N_996,N_251,N_370);
or U997 (N_997,N_465,N_421);
and U998 (N_998,N_221,N_57);
nand U999 (N_999,N_356,N_195);
or U1000 (N_1000,N_916,N_800);
nand U1001 (N_1001,N_857,N_785);
and U1002 (N_1002,N_940,N_909);
xor U1003 (N_1003,N_674,N_573);
and U1004 (N_1004,N_521,N_662);
nand U1005 (N_1005,N_641,N_983);
nor U1006 (N_1006,N_699,N_576);
nand U1007 (N_1007,N_654,N_982);
nor U1008 (N_1008,N_542,N_907);
nor U1009 (N_1009,N_946,N_726);
or U1010 (N_1010,N_891,N_759);
and U1011 (N_1011,N_739,N_701);
and U1012 (N_1012,N_688,N_997);
nor U1013 (N_1013,N_612,N_884);
nor U1014 (N_1014,N_790,N_936);
or U1015 (N_1015,N_778,N_547);
nor U1016 (N_1016,N_691,N_500);
nand U1017 (N_1017,N_823,N_735);
xor U1018 (N_1018,N_945,N_861);
and U1019 (N_1019,N_535,N_860);
and U1020 (N_1020,N_523,N_723);
nor U1021 (N_1021,N_586,N_622);
or U1022 (N_1022,N_718,N_947);
nor U1023 (N_1023,N_668,N_826);
and U1024 (N_1024,N_698,N_855);
nand U1025 (N_1025,N_705,N_927);
or U1026 (N_1026,N_744,N_959);
or U1027 (N_1027,N_679,N_779);
and U1028 (N_1028,N_702,N_693);
or U1029 (N_1029,N_614,N_561);
nor U1030 (N_1030,N_596,N_512);
nand U1031 (N_1031,N_648,N_848);
nor U1032 (N_1032,N_903,N_694);
nand U1033 (N_1033,N_917,N_977);
and U1034 (N_1034,N_799,N_644);
or U1035 (N_1035,N_922,N_620);
or U1036 (N_1036,N_920,N_738);
nor U1037 (N_1037,N_808,N_856);
or U1038 (N_1038,N_525,N_656);
or U1039 (N_1039,N_872,N_734);
and U1040 (N_1040,N_589,N_864);
or U1041 (N_1041,N_637,N_757);
and U1042 (N_1042,N_850,N_840);
or U1043 (N_1043,N_834,N_554);
or U1044 (N_1044,N_731,N_540);
and U1045 (N_1045,N_876,N_733);
or U1046 (N_1046,N_882,N_888);
nand U1047 (N_1047,N_514,N_803);
nand U1048 (N_1048,N_867,N_755);
nor U1049 (N_1049,N_601,N_788);
or U1050 (N_1050,N_883,N_818);
nand U1051 (N_1051,N_865,N_955);
xor U1052 (N_1052,N_615,N_776);
nand U1053 (N_1053,N_651,N_578);
or U1054 (N_1054,N_667,N_748);
nor U1055 (N_1055,N_974,N_846);
nor U1056 (N_1056,N_600,N_642);
or U1057 (N_1057,N_517,N_634);
nor U1058 (N_1058,N_937,N_791);
nand U1059 (N_1059,N_984,N_773);
and U1060 (N_1060,N_511,N_939);
and U1061 (N_1061,N_740,N_967);
nor U1062 (N_1062,N_809,N_722);
nand U1063 (N_1063,N_518,N_673);
and U1064 (N_1064,N_716,N_877);
nor U1065 (N_1065,N_802,N_798);
nor U1066 (N_1066,N_839,N_880);
nor U1067 (N_1067,N_870,N_611);
and U1068 (N_1068,N_599,N_685);
nand U1069 (N_1069,N_902,N_952);
nand U1070 (N_1070,N_836,N_948);
or U1071 (N_1071,N_817,N_780);
nand U1072 (N_1072,N_938,N_976);
and U1073 (N_1073,N_912,N_918);
and U1074 (N_1074,N_562,N_590);
nand U1075 (N_1075,N_968,N_957);
nor U1076 (N_1076,N_549,N_680);
nor U1077 (N_1077,N_796,N_566);
and U1078 (N_1078,N_534,N_717);
or U1079 (N_1079,N_528,N_510);
nand U1080 (N_1080,N_545,N_666);
and U1081 (N_1081,N_607,N_862);
nand U1082 (N_1082,N_859,N_661);
or U1083 (N_1083,N_822,N_714);
nor U1084 (N_1084,N_978,N_794);
and U1085 (N_1085,N_736,N_979);
nor U1086 (N_1086,N_531,N_892);
or U1087 (N_1087,N_606,N_921);
or U1088 (N_1088,N_502,N_527);
nand U1089 (N_1089,N_754,N_572);
nor U1090 (N_1090,N_533,N_595);
or U1091 (N_1091,N_819,N_943);
nor U1092 (N_1092,N_954,N_756);
nand U1093 (N_1093,N_505,N_697);
nand U1094 (N_1094,N_886,N_924);
nor U1095 (N_1095,N_746,N_663);
or U1096 (N_1096,N_925,N_571);
nand U1097 (N_1097,N_960,N_588);
nor U1098 (N_1098,N_949,N_526);
nor U1099 (N_1099,N_631,N_720);
nand U1100 (N_1100,N_889,N_724);
nand U1101 (N_1101,N_593,N_898);
nand U1102 (N_1102,N_618,N_989);
xnor U1103 (N_1103,N_993,N_609);
or U1104 (N_1104,N_919,N_706);
and U1105 (N_1105,N_820,N_712);
and U1106 (N_1106,N_793,N_929);
nor U1107 (N_1107,N_762,N_558);
nand U1108 (N_1108,N_653,N_557);
and U1109 (N_1109,N_670,N_831);
nand U1110 (N_1110,N_646,N_704);
xnor U1111 (N_1111,N_501,N_832);
xor U1112 (N_1112,N_941,N_782);
or U1113 (N_1113,N_690,N_553);
or U1114 (N_1114,N_626,N_905);
or U1115 (N_1115,N_841,N_583);
or U1116 (N_1116,N_594,N_963);
and U1117 (N_1117,N_672,N_753);
nor U1118 (N_1118,N_623,N_700);
xnor U1119 (N_1119,N_635,N_923);
or U1120 (N_1120,N_789,N_887);
nand U1121 (N_1121,N_908,N_950);
nand U1122 (N_1122,N_783,N_890);
nor U1123 (N_1123,N_732,N_853);
nor U1124 (N_1124,N_871,N_652);
and U1125 (N_1125,N_695,N_543);
and U1126 (N_1126,N_575,N_893);
nor U1127 (N_1127,N_786,N_524);
and U1128 (N_1128,N_942,N_765);
and U1129 (N_1129,N_928,N_763);
and U1130 (N_1130,N_866,N_582);
xor U1131 (N_1131,N_632,N_986);
or U1132 (N_1132,N_807,N_777);
nor U1133 (N_1133,N_741,N_639);
and U1134 (N_1134,N_873,N_675);
nand U1135 (N_1135,N_645,N_964);
nand U1136 (N_1136,N_781,N_682);
or U1137 (N_1137,N_830,N_895);
and U1138 (N_1138,N_849,N_750);
nand U1139 (N_1139,N_838,N_520);
and U1140 (N_1140,N_627,N_844);
and U1141 (N_1141,N_715,N_980);
nand U1142 (N_1142,N_727,N_617);
xnor U1143 (N_1143,N_971,N_858);
or U1144 (N_1144,N_657,N_970);
nand U1145 (N_1145,N_676,N_771);
or U1146 (N_1146,N_988,N_506);
and U1147 (N_1147,N_513,N_879);
xnor U1148 (N_1148,N_587,N_811);
nand U1149 (N_1149,N_851,N_604);
nor U1150 (N_1150,N_729,N_768);
nor U1151 (N_1151,N_999,N_863);
nand U1152 (N_1152,N_681,N_597);
nand U1153 (N_1153,N_911,N_835);
nor U1154 (N_1154,N_815,N_998);
nand U1155 (N_1155,N_544,N_825);
nor U1156 (N_1156,N_655,N_707);
nor U1157 (N_1157,N_689,N_625);
and U1158 (N_1158,N_962,N_581);
nor U1159 (N_1159,N_636,N_975);
nor U1160 (N_1160,N_730,N_539);
and U1161 (N_1161,N_965,N_958);
nand U1162 (N_1162,N_602,N_926);
nor U1163 (N_1163,N_814,N_621);
nor U1164 (N_1164,N_649,N_930);
or U1165 (N_1165,N_991,N_953);
or U1166 (N_1166,N_875,N_813);
xnor U1167 (N_1167,N_605,N_899);
and U1168 (N_1168,N_548,N_684);
or U1169 (N_1169,N_994,N_981);
or U1170 (N_1170,N_747,N_881);
and U1171 (N_1171,N_797,N_742);
nor U1172 (N_1172,N_529,N_845);
and U1173 (N_1173,N_532,N_795);
nand U1174 (N_1174,N_709,N_987);
nand U1175 (N_1175,N_810,N_737);
and U1176 (N_1176,N_760,N_961);
xnor U1177 (N_1177,N_546,N_843);
or U1178 (N_1178,N_752,N_538);
nand U1179 (N_1179,N_821,N_696);
xnor U1180 (N_1180,N_665,N_852);
nand U1181 (N_1181,N_564,N_770);
nor U1182 (N_1182,N_966,N_703);
or U1183 (N_1183,N_868,N_503);
or U1184 (N_1184,N_812,N_847);
nor U1185 (N_1185,N_630,N_944);
nor U1186 (N_1186,N_574,N_878);
and U1187 (N_1187,N_772,N_931);
nand U1188 (N_1188,N_585,N_805);
nor U1189 (N_1189,N_643,N_854);
nand U1190 (N_1190,N_563,N_671);
nor U1191 (N_1191,N_552,N_619);
and U1192 (N_1192,N_591,N_792);
nor U1193 (N_1193,N_577,N_565);
and U1194 (N_1194,N_713,N_551);
xnor U1195 (N_1195,N_677,N_592);
or U1196 (N_1196,N_784,N_935);
nor U1197 (N_1197,N_914,N_761);
or U1198 (N_1198,N_874,N_509);
or U1199 (N_1199,N_640,N_550);
or U1200 (N_1200,N_992,N_650);
nor U1201 (N_1201,N_624,N_568);
nor U1202 (N_1202,N_530,N_985);
nor U1203 (N_1203,N_824,N_913);
nand U1204 (N_1204,N_686,N_659);
and U1205 (N_1205,N_897,N_774);
and U1206 (N_1206,N_721,N_603);
xor U1207 (N_1207,N_719,N_633);
nor U1208 (N_1208,N_710,N_995);
nand U1209 (N_1209,N_990,N_537);
nor U1210 (N_1210,N_900,N_869);
or U1211 (N_1211,N_972,N_751);
or U1212 (N_1212,N_616,N_749);
nand U1213 (N_1213,N_613,N_629);
nor U1214 (N_1214,N_559,N_658);
nor U1215 (N_1215,N_934,N_664);
and U1216 (N_1216,N_969,N_669);
nor U1217 (N_1217,N_647,N_833);
and U1218 (N_1218,N_906,N_555);
nor U1219 (N_1219,N_660,N_515);
xnor U1220 (N_1220,N_687,N_828);
or U1221 (N_1221,N_842,N_896);
xor U1222 (N_1222,N_806,N_904);
nand U1223 (N_1223,N_910,N_775);
or U1224 (N_1224,N_767,N_804);
xor U1225 (N_1225,N_560,N_508);
or U1226 (N_1226,N_692,N_816);
nor U1227 (N_1227,N_956,N_516);
xnor U1228 (N_1228,N_541,N_610);
nand U1229 (N_1229,N_728,N_708);
or U1230 (N_1230,N_801,N_743);
or U1231 (N_1231,N_569,N_787);
nor U1232 (N_1232,N_519,N_598);
or U1233 (N_1233,N_827,N_567);
and U1234 (N_1234,N_638,N_894);
and U1235 (N_1235,N_769,N_504);
and U1236 (N_1236,N_996,N_678);
or U1237 (N_1237,N_901,N_885);
and U1238 (N_1238,N_683,N_580);
xnor U1239 (N_1239,N_711,N_932);
or U1240 (N_1240,N_608,N_584);
or U1241 (N_1241,N_766,N_556);
or U1242 (N_1242,N_522,N_933);
nand U1243 (N_1243,N_837,N_507);
nor U1244 (N_1244,N_579,N_758);
nor U1245 (N_1245,N_725,N_829);
nor U1246 (N_1246,N_951,N_536);
nor U1247 (N_1247,N_973,N_628);
and U1248 (N_1248,N_570,N_915);
or U1249 (N_1249,N_764,N_745);
nor U1250 (N_1250,N_811,N_640);
xor U1251 (N_1251,N_510,N_601);
and U1252 (N_1252,N_934,N_714);
nor U1253 (N_1253,N_759,N_793);
xnor U1254 (N_1254,N_630,N_666);
nand U1255 (N_1255,N_701,N_753);
xnor U1256 (N_1256,N_815,N_963);
nand U1257 (N_1257,N_621,N_876);
nand U1258 (N_1258,N_526,N_572);
and U1259 (N_1259,N_850,N_809);
or U1260 (N_1260,N_684,N_559);
or U1261 (N_1261,N_735,N_841);
or U1262 (N_1262,N_641,N_601);
nor U1263 (N_1263,N_980,N_999);
nor U1264 (N_1264,N_879,N_606);
and U1265 (N_1265,N_730,N_803);
or U1266 (N_1266,N_889,N_899);
or U1267 (N_1267,N_621,N_839);
and U1268 (N_1268,N_818,N_564);
or U1269 (N_1269,N_566,N_529);
xnor U1270 (N_1270,N_976,N_757);
xor U1271 (N_1271,N_873,N_992);
nand U1272 (N_1272,N_683,N_661);
xnor U1273 (N_1273,N_883,N_884);
nor U1274 (N_1274,N_933,N_795);
nor U1275 (N_1275,N_576,N_582);
nand U1276 (N_1276,N_533,N_878);
nor U1277 (N_1277,N_754,N_828);
and U1278 (N_1278,N_728,N_850);
nand U1279 (N_1279,N_978,N_634);
nand U1280 (N_1280,N_684,N_914);
nand U1281 (N_1281,N_797,N_701);
nor U1282 (N_1282,N_743,N_950);
nor U1283 (N_1283,N_898,N_520);
nand U1284 (N_1284,N_955,N_523);
or U1285 (N_1285,N_601,N_659);
and U1286 (N_1286,N_710,N_990);
nand U1287 (N_1287,N_930,N_971);
nor U1288 (N_1288,N_728,N_732);
nand U1289 (N_1289,N_817,N_522);
or U1290 (N_1290,N_891,N_853);
xnor U1291 (N_1291,N_506,N_787);
xnor U1292 (N_1292,N_745,N_627);
nor U1293 (N_1293,N_749,N_615);
nor U1294 (N_1294,N_719,N_733);
nand U1295 (N_1295,N_635,N_759);
nor U1296 (N_1296,N_685,N_935);
and U1297 (N_1297,N_808,N_677);
nor U1298 (N_1298,N_817,N_677);
and U1299 (N_1299,N_558,N_713);
nor U1300 (N_1300,N_527,N_941);
and U1301 (N_1301,N_593,N_678);
and U1302 (N_1302,N_607,N_889);
or U1303 (N_1303,N_749,N_531);
nand U1304 (N_1304,N_985,N_653);
nand U1305 (N_1305,N_585,N_533);
and U1306 (N_1306,N_965,N_617);
nor U1307 (N_1307,N_873,N_884);
or U1308 (N_1308,N_652,N_970);
or U1309 (N_1309,N_892,N_941);
nand U1310 (N_1310,N_678,N_950);
or U1311 (N_1311,N_643,N_578);
nand U1312 (N_1312,N_685,N_708);
nand U1313 (N_1313,N_742,N_628);
nor U1314 (N_1314,N_987,N_672);
and U1315 (N_1315,N_876,N_783);
nand U1316 (N_1316,N_848,N_962);
or U1317 (N_1317,N_805,N_526);
nor U1318 (N_1318,N_924,N_908);
and U1319 (N_1319,N_964,N_709);
nand U1320 (N_1320,N_651,N_595);
xnor U1321 (N_1321,N_654,N_668);
or U1322 (N_1322,N_974,N_582);
nor U1323 (N_1323,N_889,N_829);
xor U1324 (N_1324,N_890,N_849);
nor U1325 (N_1325,N_827,N_982);
nand U1326 (N_1326,N_502,N_568);
nor U1327 (N_1327,N_783,N_710);
or U1328 (N_1328,N_946,N_869);
and U1329 (N_1329,N_729,N_845);
nand U1330 (N_1330,N_921,N_722);
nor U1331 (N_1331,N_839,N_736);
nand U1332 (N_1332,N_729,N_632);
and U1333 (N_1333,N_505,N_500);
or U1334 (N_1334,N_563,N_612);
nand U1335 (N_1335,N_581,N_715);
and U1336 (N_1336,N_988,N_928);
nor U1337 (N_1337,N_585,N_686);
nand U1338 (N_1338,N_931,N_580);
nor U1339 (N_1339,N_624,N_605);
xnor U1340 (N_1340,N_587,N_573);
or U1341 (N_1341,N_777,N_926);
or U1342 (N_1342,N_803,N_787);
and U1343 (N_1343,N_628,N_770);
xor U1344 (N_1344,N_618,N_931);
and U1345 (N_1345,N_651,N_926);
or U1346 (N_1346,N_608,N_530);
or U1347 (N_1347,N_890,N_887);
nor U1348 (N_1348,N_647,N_581);
nand U1349 (N_1349,N_783,N_719);
and U1350 (N_1350,N_639,N_710);
and U1351 (N_1351,N_800,N_764);
or U1352 (N_1352,N_664,N_881);
or U1353 (N_1353,N_891,N_575);
and U1354 (N_1354,N_730,N_727);
xor U1355 (N_1355,N_630,N_683);
nor U1356 (N_1356,N_505,N_940);
or U1357 (N_1357,N_671,N_738);
nand U1358 (N_1358,N_698,N_585);
and U1359 (N_1359,N_744,N_619);
or U1360 (N_1360,N_783,N_566);
xnor U1361 (N_1361,N_859,N_512);
nand U1362 (N_1362,N_897,N_977);
and U1363 (N_1363,N_746,N_980);
nand U1364 (N_1364,N_589,N_711);
nand U1365 (N_1365,N_674,N_601);
nand U1366 (N_1366,N_543,N_767);
nor U1367 (N_1367,N_990,N_952);
and U1368 (N_1368,N_605,N_857);
and U1369 (N_1369,N_663,N_857);
xnor U1370 (N_1370,N_986,N_858);
nand U1371 (N_1371,N_506,N_734);
nor U1372 (N_1372,N_975,N_714);
or U1373 (N_1373,N_576,N_609);
or U1374 (N_1374,N_742,N_520);
nor U1375 (N_1375,N_562,N_972);
or U1376 (N_1376,N_521,N_892);
nor U1377 (N_1377,N_950,N_582);
or U1378 (N_1378,N_529,N_503);
nor U1379 (N_1379,N_559,N_646);
or U1380 (N_1380,N_523,N_516);
nor U1381 (N_1381,N_809,N_610);
and U1382 (N_1382,N_945,N_959);
xor U1383 (N_1383,N_939,N_735);
and U1384 (N_1384,N_634,N_769);
xor U1385 (N_1385,N_668,N_875);
or U1386 (N_1386,N_836,N_734);
nand U1387 (N_1387,N_880,N_645);
xnor U1388 (N_1388,N_564,N_976);
or U1389 (N_1389,N_547,N_571);
or U1390 (N_1390,N_810,N_661);
nor U1391 (N_1391,N_892,N_682);
nand U1392 (N_1392,N_646,N_791);
xnor U1393 (N_1393,N_998,N_563);
and U1394 (N_1394,N_572,N_816);
and U1395 (N_1395,N_998,N_916);
nor U1396 (N_1396,N_705,N_617);
and U1397 (N_1397,N_636,N_876);
nand U1398 (N_1398,N_939,N_804);
and U1399 (N_1399,N_901,N_735);
xnor U1400 (N_1400,N_998,N_732);
or U1401 (N_1401,N_783,N_699);
nand U1402 (N_1402,N_605,N_752);
and U1403 (N_1403,N_990,N_567);
xnor U1404 (N_1404,N_806,N_835);
or U1405 (N_1405,N_668,N_914);
and U1406 (N_1406,N_956,N_997);
nor U1407 (N_1407,N_876,N_943);
nand U1408 (N_1408,N_804,N_992);
and U1409 (N_1409,N_513,N_625);
or U1410 (N_1410,N_777,N_679);
nand U1411 (N_1411,N_589,N_921);
or U1412 (N_1412,N_751,N_912);
or U1413 (N_1413,N_932,N_736);
nor U1414 (N_1414,N_957,N_917);
nand U1415 (N_1415,N_795,N_672);
or U1416 (N_1416,N_819,N_865);
nand U1417 (N_1417,N_919,N_961);
nand U1418 (N_1418,N_792,N_848);
nor U1419 (N_1419,N_500,N_683);
and U1420 (N_1420,N_694,N_681);
or U1421 (N_1421,N_963,N_659);
nand U1422 (N_1422,N_882,N_883);
or U1423 (N_1423,N_955,N_660);
nand U1424 (N_1424,N_860,N_878);
or U1425 (N_1425,N_540,N_896);
nor U1426 (N_1426,N_600,N_603);
or U1427 (N_1427,N_980,N_670);
and U1428 (N_1428,N_918,N_688);
nor U1429 (N_1429,N_702,N_509);
or U1430 (N_1430,N_516,N_520);
and U1431 (N_1431,N_963,N_616);
nand U1432 (N_1432,N_766,N_749);
nor U1433 (N_1433,N_577,N_895);
xnor U1434 (N_1434,N_639,N_525);
xnor U1435 (N_1435,N_800,N_655);
nor U1436 (N_1436,N_593,N_569);
nand U1437 (N_1437,N_694,N_851);
nand U1438 (N_1438,N_596,N_731);
nor U1439 (N_1439,N_968,N_571);
and U1440 (N_1440,N_656,N_811);
and U1441 (N_1441,N_872,N_805);
xnor U1442 (N_1442,N_889,N_571);
or U1443 (N_1443,N_757,N_953);
nand U1444 (N_1444,N_970,N_729);
and U1445 (N_1445,N_898,N_735);
nand U1446 (N_1446,N_735,N_509);
and U1447 (N_1447,N_602,N_766);
nor U1448 (N_1448,N_792,N_811);
xor U1449 (N_1449,N_630,N_714);
and U1450 (N_1450,N_854,N_503);
and U1451 (N_1451,N_894,N_975);
nor U1452 (N_1452,N_691,N_903);
or U1453 (N_1453,N_512,N_760);
and U1454 (N_1454,N_885,N_541);
or U1455 (N_1455,N_614,N_916);
nor U1456 (N_1456,N_869,N_747);
and U1457 (N_1457,N_752,N_842);
xor U1458 (N_1458,N_599,N_684);
nand U1459 (N_1459,N_690,N_544);
nand U1460 (N_1460,N_720,N_990);
or U1461 (N_1461,N_613,N_797);
nor U1462 (N_1462,N_501,N_966);
or U1463 (N_1463,N_823,N_578);
and U1464 (N_1464,N_718,N_534);
nand U1465 (N_1465,N_855,N_586);
or U1466 (N_1466,N_818,N_603);
nor U1467 (N_1467,N_963,N_987);
xnor U1468 (N_1468,N_826,N_854);
or U1469 (N_1469,N_514,N_798);
nand U1470 (N_1470,N_825,N_800);
or U1471 (N_1471,N_641,N_623);
nand U1472 (N_1472,N_517,N_526);
nand U1473 (N_1473,N_583,N_704);
nand U1474 (N_1474,N_612,N_895);
nand U1475 (N_1475,N_772,N_643);
nor U1476 (N_1476,N_874,N_811);
and U1477 (N_1477,N_680,N_823);
or U1478 (N_1478,N_700,N_646);
or U1479 (N_1479,N_631,N_748);
or U1480 (N_1480,N_937,N_961);
or U1481 (N_1481,N_592,N_701);
and U1482 (N_1482,N_636,N_829);
nor U1483 (N_1483,N_573,N_709);
and U1484 (N_1484,N_570,N_878);
nand U1485 (N_1485,N_670,N_635);
nor U1486 (N_1486,N_891,N_852);
and U1487 (N_1487,N_715,N_783);
and U1488 (N_1488,N_944,N_537);
or U1489 (N_1489,N_698,N_628);
or U1490 (N_1490,N_903,N_640);
nor U1491 (N_1491,N_624,N_814);
xnor U1492 (N_1492,N_928,N_925);
and U1493 (N_1493,N_753,N_549);
or U1494 (N_1494,N_818,N_654);
xnor U1495 (N_1495,N_614,N_788);
nand U1496 (N_1496,N_639,N_597);
nand U1497 (N_1497,N_948,N_885);
xnor U1498 (N_1498,N_631,N_596);
nor U1499 (N_1499,N_742,N_965);
or U1500 (N_1500,N_1454,N_1158);
nor U1501 (N_1501,N_1422,N_1122);
nand U1502 (N_1502,N_1143,N_1476);
nand U1503 (N_1503,N_1222,N_1388);
and U1504 (N_1504,N_1091,N_1325);
nand U1505 (N_1505,N_1113,N_1443);
nor U1506 (N_1506,N_1394,N_1365);
nor U1507 (N_1507,N_1212,N_1322);
nor U1508 (N_1508,N_1280,N_1067);
and U1509 (N_1509,N_1306,N_1132);
nor U1510 (N_1510,N_1124,N_1286);
nor U1511 (N_1511,N_1344,N_1219);
xor U1512 (N_1512,N_1362,N_1066);
nor U1513 (N_1513,N_1237,N_1152);
or U1514 (N_1514,N_1358,N_1372);
nor U1515 (N_1515,N_1270,N_1228);
nand U1516 (N_1516,N_1075,N_1016);
xor U1517 (N_1517,N_1336,N_1009);
or U1518 (N_1518,N_1214,N_1201);
and U1519 (N_1519,N_1316,N_1044);
nand U1520 (N_1520,N_1240,N_1492);
and U1521 (N_1521,N_1456,N_1249);
nand U1522 (N_1522,N_1176,N_1490);
or U1523 (N_1523,N_1360,N_1188);
or U1524 (N_1524,N_1043,N_1072);
nor U1525 (N_1525,N_1100,N_1076);
and U1526 (N_1526,N_1131,N_1056);
xnor U1527 (N_1527,N_1022,N_1354);
and U1528 (N_1528,N_1485,N_1315);
nand U1529 (N_1529,N_1262,N_1256);
nand U1530 (N_1530,N_1384,N_1339);
or U1531 (N_1531,N_1037,N_1006);
nand U1532 (N_1532,N_1129,N_1120);
nor U1533 (N_1533,N_1215,N_1020);
nor U1534 (N_1534,N_1038,N_1294);
xnor U1535 (N_1535,N_1293,N_1431);
nor U1536 (N_1536,N_1082,N_1040);
and U1537 (N_1537,N_1455,N_1334);
nor U1538 (N_1538,N_1302,N_1493);
or U1539 (N_1539,N_1001,N_1332);
and U1540 (N_1540,N_1127,N_1265);
and U1541 (N_1541,N_1245,N_1216);
nand U1542 (N_1542,N_1218,N_1317);
and U1543 (N_1543,N_1287,N_1411);
and U1544 (N_1544,N_1496,N_1371);
and U1545 (N_1545,N_1271,N_1217);
or U1546 (N_1546,N_1200,N_1115);
nor U1547 (N_1547,N_1025,N_1346);
nand U1548 (N_1548,N_1057,N_1128);
or U1549 (N_1549,N_1199,N_1439);
xor U1550 (N_1550,N_1383,N_1474);
nand U1551 (N_1551,N_1226,N_1172);
nand U1552 (N_1552,N_1349,N_1327);
nor U1553 (N_1553,N_1376,N_1015);
or U1554 (N_1554,N_1425,N_1413);
or U1555 (N_1555,N_1130,N_1133);
or U1556 (N_1556,N_1300,N_1366);
nor U1557 (N_1557,N_1448,N_1489);
or U1558 (N_1558,N_1209,N_1162);
nand U1559 (N_1559,N_1207,N_1177);
and U1560 (N_1560,N_1343,N_1042);
and U1561 (N_1561,N_1225,N_1019);
xor U1562 (N_1562,N_1107,N_1080);
nor U1563 (N_1563,N_1429,N_1193);
nor U1564 (N_1564,N_1117,N_1033);
and U1565 (N_1565,N_1059,N_1399);
and U1566 (N_1566,N_1077,N_1460);
nor U1567 (N_1567,N_1364,N_1004);
nor U1568 (N_1568,N_1467,N_1375);
nand U1569 (N_1569,N_1463,N_1052);
nor U1570 (N_1570,N_1248,N_1141);
and U1571 (N_1571,N_1003,N_1449);
nor U1572 (N_1572,N_1373,N_1139);
and U1573 (N_1573,N_1161,N_1446);
nand U1574 (N_1574,N_1095,N_1355);
nand U1575 (N_1575,N_1285,N_1005);
and U1576 (N_1576,N_1442,N_1497);
nor U1577 (N_1577,N_1121,N_1054);
or U1578 (N_1578,N_1230,N_1254);
nand U1579 (N_1579,N_1331,N_1369);
or U1580 (N_1580,N_1094,N_1295);
nand U1581 (N_1581,N_1096,N_1466);
nor U1582 (N_1582,N_1278,N_1114);
nand U1583 (N_1583,N_1181,N_1260);
or U1584 (N_1584,N_1081,N_1039);
and U1585 (N_1585,N_1173,N_1031);
xor U1586 (N_1586,N_1488,N_1118);
or U1587 (N_1587,N_1481,N_1437);
nor U1588 (N_1588,N_1273,N_1169);
and U1589 (N_1589,N_1235,N_1447);
nand U1590 (N_1590,N_1397,N_1324);
and U1591 (N_1591,N_1427,N_1328);
or U1592 (N_1592,N_1105,N_1462);
nand U1593 (N_1593,N_1060,N_1180);
nor U1594 (N_1594,N_1164,N_1203);
nor U1595 (N_1595,N_1068,N_1368);
and U1596 (N_1596,N_1232,N_1348);
or U1597 (N_1597,N_1478,N_1421);
and U1598 (N_1598,N_1444,N_1171);
nand U1599 (N_1599,N_1284,N_1160);
or U1600 (N_1600,N_1277,N_1137);
and U1601 (N_1601,N_1291,N_1175);
and U1602 (N_1602,N_1189,N_1419);
or U1603 (N_1603,N_1312,N_1147);
nand U1604 (N_1604,N_1378,N_1389);
and U1605 (N_1605,N_1400,N_1409);
or U1606 (N_1606,N_1477,N_1392);
and U1607 (N_1607,N_1036,N_1318);
and U1608 (N_1608,N_1010,N_1473);
nand U1609 (N_1609,N_1403,N_1154);
or U1610 (N_1610,N_1320,N_1071);
or U1611 (N_1611,N_1035,N_1051);
or U1612 (N_1612,N_1157,N_1178);
and U1613 (N_1613,N_1426,N_1008);
nor U1614 (N_1614,N_1023,N_1024);
and U1615 (N_1615,N_1055,N_1459);
and U1616 (N_1616,N_1144,N_1184);
nand U1617 (N_1617,N_1404,N_1007);
nor U1618 (N_1618,N_1011,N_1102);
and U1619 (N_1619,N_1275,N_1182);
xor U1620 (N_1620,N_1029,N_1276);
or U1621 (N_1621,N_1445,N_1074);
and U1622 (N_1622,N_1367,N_1241);
xnor U1623 (N_1623,N_1387,N_1104);
nand U1624 (N_1624,N_1468,N_1380);
or U1625 (N_1625,N_1242,N_1111);
xor U1626 (N_1626,N_1148,N_1179);
or U1627 (N_1627,N_1494,N_1269);
or U1628 (N_1628,N_1483,N_1149);
nor U1629 (N_1629,N_1434,N_1138);
nor U1630 (N_1630,N_1085,N_1053);
nor U1631 (N_1631,N_1335,N_1436);
nor U1632 (N_1632,N_1109,N_1498);
nor U1633 (N_1633,N_1424,N_1027);
and U1634 (N_1634,N_1292,N_1359);
nor U1635 (N_1635,N_1002,N_1186);
and U1636 (N_1636,N_1309,N_1377);
and U1637 (N_1637,N_1391,N_1279);
nor U1638 (N_1638,N_1261,N_1079);
nor U1639 (N_1639,N_1450,N_1153);
nor U1640 (N_1640,N_1471,N_1415);
and U1641 (N_1641,N_1470,N_1099);
or U1642 (N_1642,N_1288,N_1311);
nand U1643 (N_1643,N_1382,N_1165);
nand U1644 (N_1644,N_1012,N_1183);
nor U1645 (N_1645,N_1101,N_1352);
xnor U1646 (N_1646,N_1440,N_1491);
nor U1647 (N_1647,N_1307,N_1319);
nor U1648 (N_1648,N_1026,N_1396);
xnor U1649 (N_1649,N_1398,N_1469);
nand U1650 (N_1650,N_1451,N_1345);
or U1651 (N_1651,N_1475,N_1374);
or U1652 (N_1652,N_1298,N_1103);
xor U1653 (N_1653,N_1014,N_1092);
or U1654 (N_1654,N_1457,N_1106);
and U1655 (N_1655,N_1234,N_1185);
or U1656 (N_1656,N_1406,N_1151);
xnor U1657 (N_1657,N_1112,N_1417);
or U1658 (N_1658,N_1070,N_1304);
nor U1659 (N_1659,N_1499,N_1244);
nor U1660 (N_1660,N_1464,N_1123);
or U1661 (N_1661,N_1195,N_1159);
nor U1662 (N_1662,N_1150,N_1281);
or U1663 (N_1663,N_1192,N_1337);
nor U1664 (N_1664,N_1323,N_1238);
or U1665 (N_1665,N_1089,N_1340);
and U1666 (N_1666,N_1402,N_1297);
or U1667 (N_1667,N_1236,N_1046);
or U1668 (N_1668,N_1090,N_1196);
nor U1669 (N_1669,N_1482,N_1453);
nand U1670 (N_1670,N_1206,N_1246);
nand U1671 (N_1671,N_1308,N_1155);
and U1672 (N_1672,N_1259,N_1299);
or U1673 (N_1673,N_1204,N_1050);
nor U1674 (N_1674,N_1423,N_1353);
nand U1675 (N_1675,N_1418,N_1205);
xor U1676 (N_1676,N_1083,N_1227);
and U1677 (N_1677,N_1379,N_1452);
nand U1678 (N_1678,N_1170,N_1168);
and U1679 (N_1679,N_1430,N_1303);
xnor U1680 (N_1680,N_1194,N_1156);
nor U1681 (N_1681,N_1486,N_1108);
nand U1682 (N_1682,N_1140,N_1093);
nor U1683 (N_1683,N_1441,N_1296);
xor U1684 (N_1684,N_1393,N_1058);
nor U1685 (N_1685,N_1047,N_1032);
and U1686 (N_1686,N_1229,N_1420);
or U1687 (N_1687,N_1480,N_1385);
or U1688 (N_1688,N_1330,N_1407);
and U1689 (N_1689,N_1069,N_1191);
nand U1690 (N_1690,N_1174,N_1041);
xor U1691 (N_1691,N_1305,N_1135);
and U1692 (N_1692,N_1472,N_1283);
xnor U1693 (N_1693,N_1465,N_1034);
or U1694 (N_1694,N_1251,N_1495);
and U1695 (N_1695,N_1428,N_1163);
or U1696 (N_1696,N_1145,N_1166);
nor U1697 (N_1697,N_1282,N_1125);
xor U1698 (N_1698,N_1146,N_1116);
xnor U1699 (N_1699,N_1408,N_1267);
nor U1700 (N_1700,N_1313,N_1410);
and U1701 (N_1701,N_1253,N_1314);
and U1702 (N_1702,N_1301,N_1414);
or U1703 (N_1703,N_1211,N_1272);
nand U1704 (N_1704,N_1487,N_1073);
or U1705 (N_1705,N_1333,N_1061);
and U1706 (N_1706,N_1432,N_1208);
xnor U1707 (N_1707,N_1326,N_1357);
or U1708 (N_1708,N_1381,N_1458);
xor U1709 (N_1709,N_1097,N_1119);
nand U1710 (N_1710,N_1134,N_1224);
and U1711 (N_1711,N_1401,N_1461);
and U1712 (N_1712,N_1030,N_1433);
or U1713 (N_1713,N_1045,N_1064);
or U1714 (N_1714,N_1087,N_1110);
and U1715 (N_1715,N_1000,N_1484);
and U1716 (N_1716,N_1198,N_1048);
nor U1717 (N_1717,N_1239,N_1126);
nand U1718 (N_1718,N_1086,N_1250);
nor U1719 (N_1719,N_1390,N_1136);
or U1720 (N_1720,N_1190,N_1405);
nand U1721 (N_1721,N_1049,N_1361);
nor U1722 (N_1722,N_1247,N_1351);
xnor U1723 (N_1723,N_1266,N_1338);
and U1724 (N_1724,N_1063,N_1395);
nor U1725 (N_1725,N_1062,N_1013);
xor U1726 (N_1726,N_1065,N_1213);
nor U1727 (N_1727,N_1274,N_1347);
xnor U1728 (N_1728,N_1341,N_1329);
nor U1729 (N_1729,N_1167,N_1258);
and U1730 (N_1730,N_1223,N_1263);
xor U1731 (N_1731,N_1210,N_1197);
nand U1732 (N_1732,N_1084,N_1438);
and U1733 (N_1733,N_1252,N_1021);
and U1734 (N_1734,N_1342,N_1356);
nor U1735 (N_1735,N_1202,N_1479);
and U1736 (N_1736,N_1268,N_1088);
nand U1737 (N_1737,N_1435,N_1370);
nor U1738 (N_1738,N_1233,N_1221);
nor U1739 (N_1739,N_1321,N_1018);
or U1740 (N_1740,N_1220,N_1350);
or U1741 (N_1741,N_1290,N_1098);
nor U1742 (N_1742,N_1386,N_1187);
nand U1743 (N_1743,N_1412,N_1416);
and U1744 (N_1744,N_1078,N_1028);
and U1745 (N_1745,N_1310,N_1257);
and U1746 (N_1746,N_1289,N_1142);
nand U1747 (N_1747,N_1017,N_1255);
nor U1748 (N_1748,N_1231,N_1363);
and U1749 (N_1749,N_1264,N_1243);
nand U1750 (N_1750,N_1274,N_1367);
nor U1751 (N_1751,N_1081,N_1499);
nand U1752 (N_1752,N_1076,N_1479);
nand U1753 (N_1753,N_1479,N_1312);
nor U1754 (N_1754,N_1159,N_1052);
nor U1755 (N_1755,N_1361,N_1038);
or U1756 (N_1756,N_1314,N_1039);
xnor U1757 (N_1757,N_1121,N_1494);
and U1758 (N_1758,N_1393,N_1482);
nand U1759 (N_1759,N_1358,N_1014);
nor U1760 (N_1760,N_1259,N_1099);
and U1761 (N_1761,N_1300,N_1292);
nand U1762 (N_1762,N_1307,N_1262);
or U1763 (N_1763,N_1065,N_1007);
nand U1764 (N_1764,N_1338,N_1136);
or U1765 (N_1765,N_1076,N_1212);
or U1766 (N_1766,N_1033,N_1180);
nor U1767 (N_1767,N_1056,N_1128);
and U1768 (N_1768,N_1274,N_1114);
and U1769 (N_1769,N_1057,N_1136);
or U1770 (N_1770,N_1294,N_1033);
and U1771 (N_1771,N_1023,N_1469);
nand U1772 (N_1772,N_1373,N_1186);
nor U1773 (N_1773,N_1477,N_1251);
and U1774 (N_1774,N_1341,N_1028);
and U1775 (N_1775,N_1046,N_1098);
and U1776 (N_1776,N_1218,N_1191);
nor U1777 (N_1777,N_1432,N_1259);
nor U1778 (N_1778,N_1052,N_1426);
nor U1779 (N_1779,N_1438,N_1135);
or U1780 (N_1780,N_1152,N_1068);
or U1781 (N_1781,N_1165,N_1123);
xnor U1782 (N_1782,N_1253,N_1432);
and U1783 (N_1783,N_1205,N_1067);
and U1784 (N_1784,N_1474,N_1423);
or U1785 (N_1785,N_1494,N_1259);
nand U1786 (N_1786,N_1014,N_1487);
nand U1787 (N_1787,N_1321,N_1216);
nor U1788 (N_1788,N_1062,N_1219);
nor U1789 (N_1789,N_1367,N_1225);
or U1790 (N_1790,N_1082,N_1124);
or U1791 (N_1791,N_1252,N_1016);
or U1792 (N_1792,N_1267,N_1076);
or U1793 (N_1793,N_1295,N_1000);
xnor U1794 (N_1794,N_1390,N_1315);
nor U1795 (N_1795,N_1386,N_1257);
and U1796 (N_1796,N_1327,N_1128);
and U1797 (N_1797,N_1380,N_1300);
and U1798 (N_1798,N_1281,N_1474);
or U1799 (N_1799,N_1040,N_1116);
nor U1800 (N_1800,N_1083,N_1211);
nand U1801 (N_1801,N_1004,N_1445);
and U1802 (N_1802,N_1060,N_1367);
and U1803 (N_1803,N_1028,N_1008);
nand U1804 (N_1804,N_1231,N_1479);
and U1805 (N_1805,N_1431,N_1183);
xnor U1806 (N_1806,N_1417,N_1003);
or U1807 (N_1807,N_1298,N_1262);
nand U1808 (N_1808,N_1064,N_1385);
or U1809 (N_1809,N_1122,N_1214);
or U1810 (N_1810,N_1133,N_1032);
and U1811 (N_1811,N_1479,N_1273);
or U1812 (N_1812,N_1029,N_1159);
nand U1813 (N_1813,N_1142,N_1484);
nor U1814 (N_1814,N_1186,N_1396);
and U1815 (N_1815,N_1295,N_1411);
and U1816 (N_1816,N_1333,N_1465);
nand U1817 (N_1817,N_1324,N_1278);
and U1818 (N_1818,N_1237,N_1322);
xor U1819 (N_1819,N_1181,N_1464);
nor U1820 (N_1820,N_1127,N_1358);
nand U1821 (N_1821,N_1146,N_1201);
or U1822 (N_1822,N_1105,N_1248);
nand U1823 (N_1823,N_1399,N_1162);
and U1824 (N_1824,N_1324,N_1070);
nor U1825 (N_1825,N_1343,N_1260);
xnor U1826 (N_1826,N_1259,N_1006);
nand U1827 (N_1827,N_1471,N_1305);
nand U1828 (N_1828,N_1048,N_1294);
xor U1829 (N_1829,N_1392,N_1394);
nor U1830 (N_1830,N_1479,N_1284);
xor U1831 (N_1831,N_1040,N_1031);
nand U1832 (N_1832,N_1138,N_1213);
and U1833 (N_1833,N_1073,N_1007);
nand U1834 (N_1834,N_1313,N_1090);
nor U1835 (N_1835,N_1091,N_1417);
nor U1836 (N_1836,N_1191,N_1490);
xor U1837 (N_1837,N_1105,N_1085);
nor U1838 (N_1838,N_1008,N_1201);
nor U1839 (N_1839,N_1472,N_1395);
nor U1840 (N_1840,N_1430,N_1188);
and U1841 (N_1841,N_1484,N_1333);
xnor U1842 (N_1842,N_1237,N_1415);
or U1843 (N_1843,N_1486,N_1218);
and U1844 (N_1844,N_1312,N_1182);
or U1845 (N_1845,N_1341,N_1007);
nand U1846 (N_1846,N_1359,N_1435);
xor U1847 (N_1847,N_1119,N_1300);
nand U1848 (N_1848,N_1127,N_1039);
nor U1849 (N_1849,N_1166,N_1148);
or U1850 (N_1850,N_1447,N_1204);
and U1851 (N_1851,N_1175,N_1429);
nand U1852 (N_1852,N_1294,N_1495);
xnor U1853 (N_1853,N_1013,N_1161);
nor U1854 (N_1854,N_1093,N_1443);
xor U1855 (N_1855,N_1255,N_1069);
nand U1856 (N_1856,N_1088,N_1260);
nand U1857 (N_1857,N_1248,N_1457);
and U1858 (N_1858,N_1190,N_1323);
xor U1859 (N_1859,N_1282,N_1413);
nor U1860 (N_1860,N_1317,N_1332);
or U1861 (N_1861,N_1228,N_1444);
nand U1862 (N_1862,N_1305,N_1470);
nand U1863 (N_1863,N_1007,N_1163);
nor U1864 (N_1864,N_1029,N_1183);
or U1865 (N_1865,N_1063,N_1423);
and U1866 (N_1866,N_1135,N_1182);
nor U1867 (N_1867,N_1084,N_1255);
nand U1868 (N_1868,N_1478,N_1353);
nand U1869 (N_1869,N_1020,N_1416);
nor U1870 (N_1870,N_1274,N_1464);
and U1871 (N_1871,N_1065,N_1279);
or U1872 (N_1872,N_1465,N_1065);
and U1873 (N_1873,N_1107,N_1282);
and U1874 (N_1874,N_1104,N_1098);
nor U1875 (N_1875,N_1025,N_1195);
nor U1876 (N_1876,N_1333,N_1392);
nor U1877 (N_1877,N_1328,N_1428);
and U1878 (N_1878,N_1357,N_1009);
nand U1879 (N_1879,N_1367,N_1394);
or U1880 (N_1880,N_1116,N_1338);
nor U1881 (N_1881,N_1218,N_1356);
or U1882 (N_1882,N_1239,N_1368);
nand U1883 (N_1883,N_1476,N_1262);
or U1884 (N_1884,N_1008,N_1248);
and U1885 (N_1885,N_1204,N_1039);
and U1886 (N_1886,N_1188,N_1046);
and U1887 (N_1887,N_1383,N_1495);
nand U1888 (N_1888,N_1496,N_1314);
nor U1889 (N_1889,N_1485,N_1217);
nor U1890 (N_1890,N_1047,N_1087);
nand U1891 (N_1891,N_1201,N_1316);
nand U1892 (N_1892,N_1015,N_1242);
or U1893 (N_1893,N_1351,N_1432);
and U1894 (N_1894,N_1047,N_1352);
and U1895 (N_1895,N_1486,N_1277);
or U1896 (N_1896,N_1224,N_1309);
or U1897 (N_1897,N_1130,N_1155);
nand U1898 (N_1898,N_1194,N_1277);
nand U1899 (N_1899,N_1435,N_1258);
and U1900 (N_1900,N_1051,N_1339);
and U1901 (N_1901,N_1323,N_1469);
and U1902 (N_1902,N_1387,N_1097);
nand U1903 (N_1903,N_1267,N_1172);
nor U1904 (N_1904,N_1101,N_1486);
or U1905 (N_1905,N_1192,N_1179);
nand U1906 (N_1906,N_1428,N_1189);
and U1907 (N_1907,N_1061,N_1015);
nand U1908 (N_1908,N_1164,N_1080);
or U1909 (N_1909,N_1164,N_1295);
nor U1910 (N_1910,N_1266,N_1230);
or U1911 (N_1911,N_1370,N_1089);
and U1912 (N_1912,N_1108,N_1386);
nand U1913 (N_1913,N_1383,N_1088);
nand U1914 (N_1914,N_1039,N_1098);
and U1915 (N_1915,N_1421,N_1282);
nand U1916 (N_1916,N_1206,N_1437);
nor U1917 (N_1917,N_1465,N_1172);
nor U1918 (N_1918,N_1003,N_1289);
or U1919 (N_1919,N_1017,N_1398);
nor U1920 (N_1920,N_1259,N_1384);
or U1921 (N_1921,N_1177,N_1395);
xnor U1922 (N_1922,N_1373,N_1272);
and U1923 (N_1923,N_1122,N_1339);
nand U1924 (N_1924,N_1473,N_1417);
nand U1925 (N_1925,N_1241,N_1113);
xor U1926 (N_1926,N_1077,N_1165);
nand U1927 (N_1927,N_1376,N_1016);
and U1928 (N_1928,N_1159,N_1462);
and U1929 (N_1929,N_1128,N_1044);
nor U1930 (N_1930,N_1484,N_1258);
or U1931 (N_1931,N_1064,N_1122);
nand U1932 (N_1932,N_1318,N_1457);
nor U1933 (N_1933,N_1036,N_1057);
and U1934 (N_1934,N_1177,N_1091);
or U1935 (N_1935,N_1214,N_1304);
and U1936 (N_1936,N_1306,N_1049);
and U1937 (N_1937,N_1336,N_1236);
nor U1938 (N_1938,N_1377,N_1068);
nor U1939 (N_1939,N_1479,N_1167);
and U1940 (N_1940,N_1072,N_1288);
nand U1941 (N_1941,N_1389,N_1316);
or U1942 (N_1942,N_1068,N_1337);
xor U1943 (N_1943,N_1116,N_1287);
and U1944 (N_1944,N_1268,N_1277);
nor U1945 (N_1945,N_1414,N_1437);
or U1946 (N_1946,N_1233,N_1159);
nor U1947 (N_1947,N_1387,N_1224);
or U1948 (N_1948,N_1031,N_1150);
and U1949 (N_1949,N_1084,N_1290);
nor U1950 (N_1950,N_1389,N_1274);
nand U1951 (N_1951,N_1294,N_1155);
nand U1952 (N_1952,N_1323,N_1104);
and U1953 (N_1953,N_1063,N_1404);
and U1954 (N_1954,N_1498,N_1410);
and U1955 (N_1955,N_1070,N_1431);
nand U1956 (N_1956,N_1143,N_1262);
nand U1957 (N_1957,N_1102,N_1250);
and U1958 (N_1958,N_1008,N_1142);
xnor U1959 (N_1959,N_1322,N_1090);
xor U1960 (N_1960,N_1385,N_1451);
and U1961 (N_1961,N_1215,N_1185);
nor U1962 (N_1962,N_1340,N_1264);
nand U1963 (N_1963,N_1131,N_1484);
nor U1964 (N_1964,N_1192,N_1471);
nand U1965 (N_1965,N_1227,N_1127);
nand U1966 (N_1966,N_1478,N_1136);
nor U1967 (N_1967,N_1215,N_1250);
nor U1968 (N_1968,N_1011,N_1149);
xnor U1969 (N_1969,N_1126,N_1300);
and U1970 (N_1970,N_1330,N_1307);
xor U1971 (N_1971,N_1455,N_1204);
nor U1972 (N_1972,N_1433,N_1197);
nor U1973 (N_1973,N_1249,N_1078);
and U1974 (N_1974,N_1381,N_1346);
xor U1975 (N_1975,N_1340,N_1497);
nand U1976 (N_1976,N_1035,N_1414);
xnor U1977 (N_1977,N_1060,N_1142);
nor U1978 (N_1978,N_1376,N_1032);
or U1979 (N_1979,N_1129,N_1460);
nor U1980 (N_1980,N_1455,N_1238);
or U1981 (N_1981,N_1078,N_1228);
xor U1982 (N_1982,N_1348,N_1495);
and U1983 (N_1983,N_1279,N_1471);
and U1984 (N_1984,N_1206,N_1432);
nor U1985 (N_1985,N_1187,N_1473);
nand U1986 (N_1986,N_1433,N_1469);
and U1987 (N_1987,N_1399,N_1281);
nor U1988 (N_1988,N_1085,N_1162);
nor U1989 (N_1989,N_1404,N_1498);
xnor U1990 (N_1990,N_1489,N_1367);
nor U1991 (N_1991,N_1477,N_1221);
nand U1992 (N_1992,N_1352,N_1139);
nor U1993 (N_1993,N_1243,N_1324);
or U1994 (N_1994,N_1491,N_1393);
nand U1995 (N_1995,N_1094,N_1322);
and U1996 (N_1996,N_1053,N_1260);
nand U1997 (N_1997,N_1403,N_1491);
xor U1998 (N_1998,N_1420,N_1369);
xor U1999 (N_1999,N_1112,N_1019);
and U2000 (N_2000,N_1971,N_1870);
nor U2001 (N_2001,N_1574,N_1851);
nor U2002 (N_2002,N_1620,N_1775);
nand U2003 (N_2003,N_1881,N_1756);
or U2004 (N_2004,N_1769,N_1644);
nand U2005 (N_2005,N_1680,N_1920);
xor U2006 (N_2006,N_1793,N_1580);
nor U2007 (N_2007,N_1992,N_1906);
nor U2008 (N_2008,N_1702,N_1777);
and U2009 (N_2009,N_1999,N_1751);
nand U2010 (N_2010,N_1658,N_1539);
and U2011 (N_2011,N_1507,N_1515);
and U2012 (N_2012,N_1944,N_1510);
nor U2013 (N_2013,N_1950,N_1958);
and U2014 (N_2014,N_1815,N_1930);
and U2015 (N_2015,N_1737,N_1599);
and U2016 (N_2016,N_1526,N_1879);
nor U2017 (N_2017,N_1970,N_1991);
xor U2018 (N_2018,N_1562,N_1577);
or U2019 (N_2019,N_1691,N_1509);
nand U2020 (N_2020,N_1759,N_1636);
nand U2021 (N_2021,N_1624,N_1901);
or U2022 (N_2022,N_1679,N_1742);
or U2023 (N_2023,N_1587,N_1969);
nor U2024 (N_2024,N_1734,N_1570);
nor U2025 (N_2025,N_1749,N_1607);
xnor U2026 (N_2026,N_1645,N_1728);
and U2027 (N_2027,N_1959,N_1546);
or U2028 (N_2028,N_1722,N_1779);
nor U2029 (N_2029,N_1905,N_1584);
nor U2030 (N_2030,N_1738,N_1614);
or U2031 (N_2031,N_1972,N_1834);
xor U2032 (N_2032,N_1836,N_1754);
nor U2033 (N_2033,N_1608,N_1976);
xor U2034 (N_2034,N_1572,N_1946);
or U2035 (N_2035,N_1990,N_1826);
nor U2036 (N_2036,N_1867,N_1513);
nand U2037 (N_2037,N_1505,N_1723);
and U2038 (N_2038,N_1925,N_1506);
nor U2039 (N_2039,N_1641,N_1592);
and U2040 (N_2040,N_1997,N_1922);
or U2041 (N_2041,N_1895,N_1907);
nor U2042 (N_2042,N_1886,N_1632);
xnor U2043 (N_2043,N_1852,N_1554);
nor U2044 (N_2044,N_1774,N_1838);
or U2045 (N_2045,N_1795,N_1831);
nor U2046 (N_2046,N_1618,N_1948);
nand U2047 (N_2047,N_1649,N_1800);
and U2048 (N_2048,N_1753,N_1880);
nor U2049 (N_2049,N_1571,N_1511);
xnor U2050 (N_2050,N_1604,N_1827);
or U2051 (N_2051,N_1974,N_1908);
nor U2052 (N_2052,N_1806,N_1504);
nand U2053 (N_2053,N_1935,N_1916);
or U2054 (N_2054,N_1830,N_1667);
nor U2055 (N_2055,N_1843,N_1809);
xor U2056 (N_2056,N_1537,N_1718);
or U2057 (N_2057,N_1522,N_1555);
nand U2058 (N_2058,N_1597,N_1824);
or U2059 (N_2059,N_1847,N_1663);
nand U2060 (N_2060,N_1651,N_1891);
and U2061 (N_2061,N_1730,N_1615);
nor U2062 (N_2062,N_1520,N_1594);
nand U2063 (N_2063,N_1811,N_1889);
xor U2064 (N_2064,N_1963,N_1564);
and U2065 (N_2065,N_1642,N_1671);
nand U2066 (N_2066,N_1817,N_1683);
or U2067 (N_2067,N_1763,N_1985);
nand U2068 (N_2068,N_1949,N_1979);
nor U2069 (N_2069,N_1813,N_1877);
or U2070 (N_2070,N_1794,N_1568);
and U2071 (N_2071,N_1732,N_1681);
xor U2072 (N_2072,N_1514,N_1525);
nor U2073 (N_2073,N_1839,N_1919);
nand U2074 (N_2074,N_1656,N_1954);
or U2075 (N_2075,N_1848,N_1996);
xnor U2076 (N_2076,N_1810,N_1967);
and U2077 (N_2077,N_1752,N_1558);
or U2078 (N_2078,N_1778,N_1589);
nand U2079 (N_2079,N_1676,N_1927);
and U2080 (N_2080,N_1892,N_1966);
nor U2081 (N_2081,N_1699,N_1943);
nor U2082 (N_2082,N_1726,N_1821);
nand U2083 (N_2083,N_1973,N_1524);
nor U2084 (N_2084,N_1605,N_1982);
nand U2085 (N_2085,N_1897,N_1819);
or U2086 (N_2086,N_1557,N_1915);
nor U2087 (N_2087,N_1686,N_1887);
nand U2088 (N_2088,N_1773,N_1903);
or U2089 (N_2089,N_1626,N_1637);
nor U2090 (N_2090,N_1647,N_1617);
nor U2091 (N_2091,N_1986,N_1850);
nand U2092 (N_2092,N_1713,N_1654);
or U2093 (N_2093,N_1914,N_1760);
and U2094 (N_2094,N_1657,N_1684);
xor U2095 (N_2095,N_1947,N_1720);
nor U2096 (N_2096,N_1573,N_1712);
xnor U2097 (N_2097,N_1833,N_1755);
nand U2098 (N_2098,N_1937,N_1782);
and U2099 (N_2099,N_1933,N_1655);
and U2100 (N_2100,N_1603,N_1725);
and U2101 (N_2101,N_1576,N_1805);
nand U2102 (N_2102,N_1508,N_1978);
or U2103 (N_2103,N_1998,N_1864);
nor U2104 (N_2104,N_1540,N_1674);
and U2105 (N_2105,N_1988,N_1899);
and U2106 (N_2106,N_1748,N_1670);
or U2107 (N_2107,N_1535,N_1547);
nand U2108 (N_2108,N_1701,N_1952);
and U2109 (N_2109,N_1758,N_1646);
xnor U2110 (N_2110,N_1548,N_1733);
nor U2111 (N_2111,N_1918,N_1567);
nor U2112 (N_2112,N_1660,N_1640);
nor U2113 (N_2113,N_1560,N_1648);
or U2114 (N_2114,N_1980,N_1531);
and U2115 (N_2115,N_1512,N_1706);
nand U2116 (N_2116,N_1695,N_1862);
or U2117 (N_2117,N_1823,N_1939);
and U2118 (N_2118,N_1638,N_1623);
xor U2119 (N_2119,N_1784,N_1521);
nor U2120 (N_2120,N_1766,N_1888);
nor U2121 (N_2121,N_1820,N_1705);
nor U2122 (N_2122,N_1904,N_1639);
nand U2123 (N_2123,N_1669,N_1581);
or U2124 (N_2124,N_1865,N_1764);
or U2125 (N_2125,N_1653,N_1662);
and U2126 (N_2126,N_1931,N_1714);
nor U2127 (N_2127,N_1791,N_1700);
xor U2128 (N_2128,N_1694,N_1551);
and U2129 (N_2129,N_1698,N_1715);
or U2130 (N_2130,N_1747,N_1534);
xor U2131 (N_2131,N_1583,N_1924);
xnor U2132 (N_2132,N_1566,N_1735);
nor U2133 (N_2133,N_1968,N_1828);
or U2134 (N_2134,N_1711,N_1709);
nor U2135 (N_2135,N_1668,N_1503);
nor U2136 (N_2136,N_1876,N_1703);
xnor U2137 (N_2137,N_1602,N_1743);
or U2138 (N_2138,N_1550,N_1767);
nand U2139 (N_2139,N_1801,N_1527);
nand U2140 (N_2140,N_1565,N_1627);
and U2141 (N_2141,N_1625,N_1523);
or U2142 (N_2142,N_1917,N_1692);
nor U2143 (N_2143,N_1629,N_1832);
nor U2144 (N_2144,N_1552,N_1929);
and U2145 (N_2145,N_1802,N_1942);
nor U2146 (N_2146,N_1708,N_1517);
nor U2147 (N_2147,N_1559,N_1501);
nor U2148 (N_2148,N_1951,N_1921);
and U2149 (N_2149,N_1772,N_1956);
nor U2150 (N_2150,N_1840,N_1872);
nand U2151 (N_2151,N_1588,N_1789);
nor U2152 (N_2152,N_1673,N_1871);
or U2153 (N_2153,N_1849,N_1893);
nor U2154 (N_2154,N_1873,N_1621);
xnor U2155 (N_2155,N_1808,N_1628);
nand U2156 (N_2156,N_1762,N_1635);
or U2157 (N_2157,N_1770,N_1875);
and U2158 (N_2158,N_1690,N_1545);
and U2159 (N_2159,N_1687,N_1541);
or U2160 (N_2160,N_1825,N_1788);
and U2161 (N_2161,N_1745,N_1781);
nor U2162 (N_2162,N_1556,N_1598);
and U2163 (N_2163,N_1807,N_1731);
and U2164 (N_2164,N_1600,N_1896);
nand U2165 (N_2165,N_1707,N_1797);
nor U2166 (N_2166,N_1884,N_1878);
and U2167 (N_2167,N_1874,N_1719);
nand U2168 (N_2168,N_1530,N_1936);
or U2169 (N_2169,N_1804,N_1859);
nor U2170 (N_2170,N_1582,N_1519);
or U2171 (N_2171,N_1606,N_1857);
or U2172 (N_2172,N_1923,N_1928);
nor U2173 (N_2173,N_1855,N_1902);
or U2174 (N_2174,N_1544,N_1696);
nor U2175 (N_2175,N_1664,N_1910);
and U2176 (N_2176,N_1650,N_1661);
nor U2177 (N_2177,N_1926,N_1866);
nand U2178 (N_2178,N_1746,N_1912);
or U2179 (N_2179,N_1724,N_1894);
xor U2180 (N_2180,N_1776,N_1961);
and U2181 (N_2181,N_1689,N_1622);
or U2182 (N_2182,N_1977,N_1563);
or U2183 (N_2183,N_1516,N_1957);
xnor U2184 (N_2184,N_1744,N_1586);
nor U2185 (N_2185,N_1578,N_1591);
or U2186 (N_2186,N_1672,N_1854);
and U2187 (N_2187,N_1717,N_1780);
or U2188 (N_2188,N_1652,N_1913);
nand U2189 (N_2189,N_1960,N_1765);
nand U2190 (N_2190,N_1538,N_1829);
and U2191 (N_2191,N_1736,N_1575);
and U2192 (N_2192,N_1613,N_1814);
nand U2193 (N_2193,N_1955,N_1909);
and U2194 (N_2194,N_1856,N_1643);
and U2195 (N_2195,N_1542,N_1863);
nand U2196 (N_2196,N_1853,N_1837);
nand U2197 (N_2197,N_1727,N_1585);
nor U2198 (N_2198,N_1685,N_1962);
or U2199 (N_2199,N_1822,N_1710);
and U2200 (N_2200,N_1693,N_1883);
nand U2201 (N_2201,N_1812,N_1569);
and U2202 (N_2202,N_1869,N_1900);
or U2203 (N_2203,N_1739,N_1502);
nand U2204 (N_2204,N_1835,N_1561);
or U2205 (N_2205,N_1945,N_1536);
nor U2206 (N_2206,N_1842,N_1678);
nor U2207 (N_2207,N_1729,N_1529);
or U2208 (N_2208,N_1579,N_1790);
nand U2209 (N_2209,N_1612,N_1771);
nor U2210 (N_2210,N_1665,N_1964);
or U2211 (N_2211,N_1938,N_1846);
or U2212 (N_2212,N_1987,N_1981);
and U2213 (N_2213,N_1596,N_1528);
nand U2214 (N_2214,N_1704,N_1630);
nor U2215 (N_2215,N_1792,N_1787);
and U2216 (N_2216,N_1697,N_1858);
or U2217 (N_2217,N_1590,N_1841);
or U2218 (N_2218,N_1716,N_1553);
nor U2219 (N_2219,N_1803,N_1989);
and U2220 (N_2220,N_1934,N_1543);
and U2221 (N_2221,N_1798,N_1533);
nor U2222 (N_2222,N_1595,N_1593);
nor U2223 (N_2223,N_1740,N_1796);
nor U2224 (N_2224,N_1890,N_1532);
nor U2225 (N_2225,N_1741,N_1610);
nor U2226 (N_2226,N_1616,N_1500);
nor U2227 (N_2227,N_1633,N_1941);
nor U2228 (N_2228,N_1634,N_1975);
nand U2229 (N_2229,N_1721,N_1611);
nand U2230 (N_2230,N_1631,N_1861);
nor U2231 (N_2231,N_1688,N_1995);
xor U2232 (N_2232,N_1601,N_1965);
or U2233 (N_2233,N_1799,N_1786);
nand U2234 (N_2234,N_1983,N_1953);
xor U2235 (N_2235,N_1818,N_1682);
or U2236 (N_2236,N_1845,N_1785);
xnor U2237 (N_2237,N_1844,N_1757);
xor U2238 (N_2238,N_1816,N_1768);
xor U2239 (N_2239,N_1994,N_1932);
xor U2240 (N_2240,N_1666,N_1984);
nand U2241 (N_2241,N_1761,N_1993);
and U2242 (N_2242,N_1518,N_1860);
and U2243 (N_2243,N_1940,N_1677);
nor U2244 (N_2244,N_1885,N_1619);
and U2245 (N_2245,N_1675,N_1783);
or U2246 (N_2246,N_1868,N_1549);
nor U2247 (N_2247,N_1609,N_1898);
or U2248 (N_2248,N_1659,N_1911);
or U2249 (N_2249,N_1882,N_1750);
nand U2250 (N_2250,N_1811,N_1524);
and U2251 (N_2251,N_1588,N_1868);
nor U2252 (N_2252,N_1891,N_1645);
and U2253 (N_2253,N_1536,N_1702);
and U2254 (N_2254,N_1837,N_1824);
nand U2255 (N_2255,N_1950,N_1685);
or U2256 (N_2256,N_1954,N_1862);
nand U2257 (N_2257,N_1647,N_1932);
xor U2258 (N_2258,N_1772,N_1977);
nor U2259 (N_2259,N_1781,N_1890);
or U2260 (N_2260,N_1680,N_1829);
and U2261 (N_2261,N_1781,N_1970);
xor U2262 (N_2262,N_1720,N_1707);
nand U2263 (N_2263,N_1980,N_1908);
nand U2264 (N_2264,N_1942,N_1896);
xnor U2265 (N_2265,N_1953,N_1951);
and U2266 (N_2266,N_1537,N_1912);
nand U2267 (N_2267,N_1780,N_1662);
nand U2268 (N_2268,N_1805,N_1791);
nand U2269 (N_2269,N_1970,N_1908);
or U2270 (N_2270,N_1501,N_1542);
nand U2271 (N_2271,N_1705,N_1999);
and U2272 (N_2272,N_1664,N_1996);
nor U2273 (N_2273,N_1704,N_1604);
nor U2274 (N_2274,N_1627,N_1606);
xnor U2275 (N_2275,N_1752,N_1874);
or U2276 (N_2276,N_1716,N_1678);
nor U2277 (N_2277,N_1931,N_1909);
or U2278 (N_2278,N_1604,N_1797);
xor U2279 (N_2279,N_1837,N_1804);
nor U2280 (N_2280,N_1614,N_1874);
xor U2281 (N_2281,N_1521,N_1925);
or U2282 (N_2282,N_1810,N_1501);
and U2283 (N_2283,N_1849,N_1560);
or U2284 (N_2284,N_1693,N_1791);
and U2285 (N_2285,N_1752,N_1955);
or U2286 (N_2286,N_1963,N_1637);
nor U2287 (N_2287,N_1640,N_1948);
nand U2288 (N_2288,N_1678,N_1535);
nand U2289 (N_2289,N_1981,N_1759);
or U2290 (N_2290,N_1710,N_1953);
nor U2291 (N_2291,N_1572,N_1912);
nand U2292 (N_2292,N_1852,N_1811);
xor U2293 (N_2293,N_1745,N_1619);
and U2294 (N_2294,N_1966,N_1972);
xnor U2295 (N_2295,N_1863,N_1886);
nor U2296 (N_2296,N_1891,N_1811);
xnor U2297 (N_2297,N_1897,N_1987);
xnor U2298 (N_2298,N_1956,N_1891);
and U2299 (N_2299,N_1947,N_1966);
nor U2300 (N_2300,N_1818,N_1788);
and U2301 (N_2301,N_1841,N_1730);
nor U2302 (N_2302,N_1500,N_1978);
and U2303 (N_2303,N_1644,N_1595);
or U2304 (N_2304,N_1784,N_1571);
nor U2305 (N_2305,N_1927,N_1695);
or U2306 (N_2306,N_1597,N_1802);
nor U2307 (N_2307,N_1622,N_1838);
or U2308 (N_2308,N_1982,N_1511);
and U2309 (N_2309,N_1971,N_1666);
nor U2310 (N_2310,N_1807,N_1580);
nor U2311 (N_2311,N_1989,N_1957);
nand U2312 (N_2312,N_1864,N_1799);
xor U2313 (N_2313,N_1778,N_1882);
and U2314 (N_2314,N_1985,N_1511);
or U2315 (N_2315,N_1987,N_1619);
nand U2316 (N_2316,N_1858,N_1671);
or U2317 (N_2317,N_1669,N_1552);
xnor U2318 (N_2318,N_1875,N_1545);
nor U2319 (N_2319,N_1902,N_1864);
nand U2320 (N_2320,N_1876,N_1503);
xor U2321 (N_2321,N_1534,N_1789);
and U2322 (N_2322,N_1925,N_1519);
and U2323 (N_2323,N_1829,N_1974);
nor U2324 (N_2324,N_1980,N_1732);
nor U2325 (N_2325,N_1555,N_1582);
xor U2326 (N_2326,N_1903,N_1960);
and U2327 (N_2327,N_1953,N_1799);
and U2328 (N_2328,N_1629,N_1601);
nand U2329 (N_2329,N_1651,N_1501);
xor U2330 (N_2330,N_1504,N_1546);
or U2331 (N_2331,N_1540,N_1561);
nand U2332 (N_2332,N_1918,N_1517);
xor U2333 (N_2333,N_1647,N_1793);
nor U2334 (N_2334,N_1639,N_1587);
or U2335 (N_2335,N_1652,N_1508);
xnor U2336 (N_2336,N_1554,N_1617);
nor U2337 (N_2337,N_1516,N_1690);
and U2338 (N_2338,N_1828,N_1679);
xor U2339 (N_2339,N_1865,N_1882);
nor U2340 (N_2340,N_1835,N_1558);
or U2341 (N_2341,N_1516,N_1564);
or U2342 (N_2342,N_1716,N_1834);
and U2343 (N_2343,N_1856,N_1722);
or U2344 (N_2344,N_1978,N_1699);
nand U2345 (N_2345,N_1673,N_1834);
xnor U2346 (N_2346,N_1517,N_1815);
or U2347 (N_2347,N_1718,N_1999);
or U2348 (N_2348,N_1836,N_1876);
nand U2349 (N_2349,N_1993,N_1754);
and U2350 (N_2350,N_1724,N_1833);
nor U2351 (N_2351,N_1982,N_1956);
nand U2352 (N_2352,N_1614,N_1560);
nand U2353 (N_2353,N_1829,N_1647);
and U2354 (N_2354,N_1780,N_1538);
and U2355 (N_2355,N_1666,N_1517);
nand U2356 (N_2356,N_1512,N_1622);
nand U2357 (N_2357,N_1948,N_1889);
xor U2358 (N_2358,N_1951,N_1645);
or U2359 (N_2359,N_1755,N_1824);
and U2360 (N_2360,N_1817,N_1800);
and U2361 (N_2361,N_1808,N_1982);
nand U2362 (N_2362,N_1783,N_1562);
or U2363 (N_2363,N_1973,N_1855);
and U2364 (N_2364,N_1576,N_1676);
nand U2365 (N_2365,N_1599,N_1699);
or U2366 (N_2366,N_1907,N_1555);
and U2367 (N_2367,N_1968,N_1997);
or U2368 (N_2368,N_1742,N_1514);
and U2369 (N_2369,N_1974,N_1953);
and U2370 (N_2370,N_1788,N_1594);
nand U2371 (N_2371,N_1680,N_1666);
or U2372 (N_2372,N_1907,N_1717);
or U2373 (N_2373,N_1522,N_1843);
and U2374 (N_2374,N_1545,N_1931);
and U2375 (N_2375,N_1559,N_1995);
nand U2376 (N_2376,N_1806,N_1943);
and U2377 (N_2377,N_1696,N_1933);
xnor U2378 (N_2378,N_1869,N_1864);
or U2379 (N_2379,N_1511,N_1560);
nand U2380 (N_2380,N_1955,N_1908);
or U2381 (N_2381,N_1551,N_1877);
nand U2382 (N_2382,N_1820,N_1657);
nor U2383 (N_2383,N_1705,N_1838);
and U2384 (N_2384,N_1980,N_1972);
or U2385 (N_2385,N_1716,N_1514);
nand U2386 (N_2386,N_1770,N_1748);
xor U2387 (N_2387,N_1805,N_1929);
nand U2388 (N_2388,N_1688,N_1516);
and U2389 (N_2389,N_1566,N_1965);
or U2390 (N_2390,N_1538,N_1765);
or U2391 (N_2391,N_1529,N_1547);
and U2392 (N_2392,N_1873,N_1957);
and U2393 (N_2393,N_1842,N_1611);
or U2394 (N_2394,N_1522,N_1947);
nor U2395 (N_2395,N_1531,N_1533);
nor U2396 (N_2396,N_1529,N_1692);
nand U2397 (N_2397,N_1657,N_1637);
or U2398 (N_2398,N_1506,N_1525);
or U2399 (N_2399,N_1866,N_1541);
or U2400 (N_2400,N_1654,N_1922);
and U2401 (N_2401,N_1592,N_1817);
or U2402 (N_2402,N_1894,N_1934);
and U2403 (N_2403,N_1641,N_1997);
nand U2404 (N_2404,N_1512,N_1648);
nand U2405 (N_2405,N_1557,N_1943);
xor U2406 (N_2406,N_1561,N_1991);
nand U2407 (N_2407,N_1516,N_1724);
xnor U2408 (N_2408,N_1571,N_1505);
and U2409 (N_2409,N_1901,N_1575);
or U2410 (N_2410,N_1757,N_1729);
nor U2411 (N_2411,N_1560,N_1610);
nand U2412 (N_2412,N_1548,N_1950);
and U2413 (N_2413,N_1846,N_1599);
nand U2414 (N_2414,N_1918,N_1546);
xnor U2415 (N_2415,N_1562,N_1810);
nand U2416 (N_2416,N_1572,N_1855);
nor U2417 (N_2417,N_1982,N_1692);
xor U2418 (N_2418,N_1585,N_1739);
xnor U2419 (N_2419,N_1680,N_1601);
nor U2420 (N_2420,N_1687,N_1964);
nor U2421 (N_2421,N_1659,N_1831);
or U2422 (N_2422,N_1556,N_1635);
or U2423 (N_2423,N_1530,N_1672);
nor U2424 (N_2424,N_1685,N_1668);
nand U2425 (N_2425,N_1660,N_1583);
nand U2426 (N_2426,N_1575,N_1953);
and U2427 (N_2427,N_1737,N_1987);
nor U2428 (N_2428,N_1916,N_1519);
xor U2429 (N_2429,N_1545,N_1560);
nor U2430 (N_2430,N_1938,N_1522);
and U2431 (N_2431,N_1654,N_1596);
nor U2432 (N_2432,N_1690,N_1827);
nand U2433 (N_2433,N_1704,N_1929);
or U2434 (N_2434,N_1721,N_1660);
nand U2435 (N_2435,N_1792,N_1624);
or U2436 (N_2436,N_1653,N_1945);
nand U2437 (N_2437,N_1749,N_1983);
nor U2438 (N_2438,N_1992,N_1781);
and U2439 (N_2439,N_1795,N_1692);
and U2440 (N_2440,N_1818,N_1519);
xnor U2441 (N_2441,N_1888,N_1984);
nor U2442 (N_2442,N_1834,N_1504);
nor U2443 (N_2443,N_1577,N_1664);
or U2444 (N_2444,N_1648,N_1596);
or U2445 (N_2445,N_1606,N_1690);
nor U2446 (N_2446,N_1522,N_1548);
nand U2447 (N_2447,N_1843,N_1909);
nor U2448 (N_2448,N_1977,N_1620);
or U2449 (N_2449,N_1605,N_1601);
and U2450 (N_2450,N_1880,N_1583);
xor U2451 (N_2451,N_1570,N_1880);
nand U2452 (N_2452,N_1655,N_1533);
and U2453 (N_2453,N_1804,N_1829);
xnor U2454 (N_2454,N_1769,N_1689);
nor U2455 (N_2455,N_1898,N_1592);
and U2456 (N_2456,N_1643,N_1576);
nor U2457 (N_2457,N_1553,N_1780);
nor U2458 (N_2458,N_1678,N_1764);
nor U2459 (N_2459,N_1842,N_1996);
or U2460 (N_2460,N_1621,N_1920);
and U2461 (N_2461,N_1580,N_1782);
nand U2462 (N_2462,N_1946,N_1782);
xnor U2463 (N_2463,N_1537,N_1872);
or U2464 (N_2464,N_1821,N_1590);
and U2465 (N_2465,N_1559,N_1503);
nand U2466 (N_2466,N_1586,N_1508);
nor U2467 (N_2467,N_1762,N_1555);
or U2468 (N_2468,N_1727,N_1576);
nand U2469 (N_2469,N_1651,N_1774);
or U2470 (N_2470,N_1714,N_1983);
nor U2471 (N_2471,N_1791,N_1613);
and U2472 (N_2472,N_1848,N_1648);
or U2473 (N_2473,N_1728,N_1858);
or U2474 (N_2474,N_1583,N_1605);
nor U2475 (N_2475,N_1712,N_1992);
and U2476 (N_2476,N_1790,N_1651);
nor U2477 (N_2477,N_1841,N_1650);
nor U2478 (N_2478,N_1942,N_1725);
or U2479 (N_2479,N_1827,N_1711);
or U2480 (N_2480,N_1560,N_1936);
xor U2481 (N_2481,N_1873,N_1505);
nand U2482 (N_2482,N_1914,N_1637);
nand U2483 (N_2483,N_1604,N_1705);
nor U2484 (N_2484,N_1740,N_1697);
and U2485 (N_2485,N_1580,N_1555);
nand U2486 (N_2486,N_1962,N_1798);
and U2487 (N_2487,N_1770,N_1541);
and U2488 (N_2488,N_1697,N_1956);
nor U2489 (N_2489,N_1765,N_1510);
xnor U2490 (N_2490,N_1565,N_1772);
nor U2491 (N_2491,N_1569,N_1802);
nor U2492 (N_2492,N_1624,N_1811);
or U2493 (N_2493,N_1608,N_1716);
and U2494 (N_2494,N_1836,N_1623);
nor U2495 (N_2495,N_1978,N_1846);
nand U2496 (N_2496,N_1799,N_1968);
and U2497 (N_2497,N_1597,N_1794);
and U2498 (N_2498,N_1536,N_1680);
and U2499 (N_2499,N_1840,N_1619);
or U2500 (N_2500,N_2478,N_2482);
nand U2501 (N_2501,N_2364,N_2230);
xor U2502 (N_2502,N_2167,N_2455);
xor U2503 (N_2503,N_2027,N_2054);
or U2504 (N_2504,N_2466,N_2127);
nand U2505 (N_2505,N_2302,N_2467);
and U2506 (N_2506,N_2222,N_2477);
and U2507 (N_2507,N_2052,N_2205);
nor U2508 (N_2508,N_2453,N_2069);
and U2509 (N_2509,N_2189,N_2298);
nand U2510 (N_2510,N_2125,N_2153);
or U2511 (N_2511,N_2074,N_2460);
nor U2512 (N_2512,N_2136,N_2324);
and U2513 (N_2513,N_2281,N_2045);
and U2514 (N_2514,N_2446,N_2315);
nor U2515 (N_2515,N_2030,N_2044);
nor U2516 (N_2516,N_2040,N_2490);
nand U2517 (N_2517,N_2140,N_2249);
nand U2518 (N_2518,N_2131,N_2461);
nor U2519 (N_2519,N_2252,N_2392);
nor U2520 (N_2520,N_2068,N_2458);
nand U2521 (N_2521,N_2350,N_2371);
xnor U2522 (N_2522,N_2411,N_2396);
nor U2523 (N_2523,N_2388,N_2076);
and U2524 (N_2524,N_2144,N_2137);
or U2525 (N_2525,N_2138,N_2261);
and U2526 (N_2526,N_2267,N_2025);
and U2527 (N_2527,N_2110,N_2250);
nor U2528 (N_2528,N_2151,N_2447);
nand U2529 (N_2529,N_2166,N_2026);
nand U2530 (N_2530,N_2154,N_2245);
nor U2531 (N_2531,N_2156,N_2257);
or U2532 (N_2532,N_2376,N_2119);
nand U2533 (N_2533,N_2418,N_2410);
nor U2534 (N_2534,N_2183,N_2062);
and U2535 (N_2535,N_2106,N_2193);
nor U2536 (N_2536,N_2090,N_2223);
xnor U2537 (N_2537,N_2115,N_2299);
nor U2538 (N_2538,N_2228,N_2117);
or U2539 (N_2539,N_2060,N_2277);
nor U2540 (N_2540,N_2024,N_2329);
xnor U2541 (N_2541,N_2464,N_2197);
xnor U2542 (N_2542,N_2171,N_2306);
nor U2543 (N_2543,N_2310,N_2462);
and U2544 (N_2544,N_2012,N_2336);
xnor U2545 (N_2545,N_2071,N_2425);
nor U2546 (N_2546,N_2155,N_2280);
or U2547 (N_2547,N_2322,N_2304);
and U2548 (N_2548,N_2242,N_2247);
nand U2549 (N_2549,N_2181,N_2255);
xnor U2550 (N_2550,N_2226,N_2358);
or U2551 (N_2551,N_2098,N_2009);
nand U2552 (N_2552,N_2483,N_2177);
and U2553 (N_2553,N_2192,N_2349);
nand U2554 (N_2554,N_2225,N_2493);
nor U2555 (N_2555,N_2473,N_2399);
nor U2556 (N_2556,N_2355,N_2390);
nor U2557 (N_2557,N_2382,N_2111);
and U2558 (N_2558,N_2476,N_2340);
xnor U2559 (N_2559,N_2269,N_2056);
and U2560 (N_2560,N_2449,N_2305);
or U2561 (N_2561,N_2199,N_2000);
or U2562 (N_2562,N_2170,N_2094);
and U2563 (N_2563,N_2073,N_2018);
or U2564 (N_2564,N_2178,N_2270);
nor U2565 (N_2565,N_2379,N_2161);
xor U2566 (N_2566,N_2229,N_2203);
xnor U2567 (N_2567,N_2375,N_2419);
or U2568 (N_2568,N_2129,N_2053);
and U2569 (N_2569,N_2179,N_2152);
or U2570 (N_2570,N_2283,N_2423);
or U2571 (N_2571,N_2377,N_2092);
or U2572 (N_2572,N_2198,N_2489);
nand U2573 (N_2573,N_2176,N_2149);
and U2574 (N_2574,N_2321,N_2331);
and U2575 (N_2575,N_2046,N_2217);
and U2576 (N_2576,N_2492,N_2211);
nand U2577 (N_2577,N_2437,N_2484);
or U2578 (N_2578,N_2133,N_2417);
or U2579 (N_2579,N_2470,N_2101);
and U2580 (N_2580,N_2370,N_2195);
nand U2581 (N_2581,N_2498,N_2172);
and U2582 (N_2582,N_2487,N_2288);
or U2583 (N_2583,N_2121,N_2327);
nand U2584 (N_2584,N_2312,N_2429);
nand U2585 (N_2585,N_2104,N_2415);
nor U2586 (N_2586,N_2290,N_2072);
and U2587 (N_2587,N_2356,N_2343);
nor U2588 (N_2588,N_2307,N_2134);
nor U2589 (N_2589,N_2235,N_2479);
nand U2590 (N_2590,N_2236,N_2282);
or U2591 (N_2591,N_2234,N_2362);
or U2592 (N_2592,N_2159,N_2440);
nand U2593 (N_2593,N_2293,N_2357);
or U2594 (N_2594,N_2031,N_2416);
or U2595 (N_2595,N_2278,N_2365);
or U2596 (N_2596,N_2318,N_2408);
nor U2597 (N_2597,N_2354,N_2471);
or U2598 (N_2598,N_2049,N_2442);
nand U2599 (N_2599,N_2480,N_2157);
nand U2600 (N_2600,N_2465,N_2294);
xor U2601 (N_2601,N_2180,N_2038);
nor U2602 (N_2602,N_2202,N_2126);
nor U2603 (N_2603,N_2058,N_2070);
nor U2604 (N_2604,N_2275,N_2116);
and U2605 (N_2605,N_2344,N_2082);
and U2606 (N_2606,N_2345,N_2241);
nor U2607 (N_2607,N_2488,N_2017);
or U2608 (N_2608,N_2201,N_2219);
and U2609 (N_2609,N_2006,N_2019);
nor U2610 (N_2610,N_2472,N_2118);
xor U2611 (N_2611,N_2491,N_2065);
xnor U2612 (N_2612,N_2139,N_2433);
and U2613 (N_2613,N_2457,N_2485);
xor U2614 (N_2614,N_2095,N_2268);
or U2615 (N_2615,N_2174,N_2407);
nand U2616 (N_2616,N_2227,N_2196);
nand U2617 (N_2617,N_2123,N_2093);
nand U2618 (N_2618,N_2296,N_2400);
nor U2619 (N_2619,N_2032,N_2373);
or U2620 (N_2620,N_2339,N_2286);
xor U2621 (N_2621,N_2285,N_2207);
or U2622 (N_2622,N_2158,N_2187);
and U2623 (N_2623,N_2454,N_2338);
and U2624 (N_2624,N_2035,N_2244);
nand U2625 (N_2625,N_2274,N_2401);
or U2626 (N_2626,N_2168,N_2313);
nor U2627 (N_2627,N_2436,N_2254);
or U2628 (N_2628,N_2004,N_2337);
nand U2629 (N_2629,N_2221,N_2445);
nor U2630 (N_2630,N_2055,N_2108);
or U2631 (N_2631,N_2438,N_2297);
nand U2632 (N_2632,N_2368,N_2367);
xor U2633 (N_2633,N_2165,N_2424);
and U2634 (N_2634,N_2220,N_2021);
and U2635 (N_2635,N_2287,N_2099);
xor U2636 (N_2636,N_2311,N_2409);
nand U2637 (N_2637,N_2120,N_2061);
nor U2638 (N_2638,N_2352,N_2173);
xor U2639 (N_2639,N_2050,N_2253);
nor U2640 (N_2640,N_2474,N_2435);
nor U2641 (N_2641,N_2214,N_2260);
nand U2642 (N_2642,N_2185,N_2206);
nand U2643 (N_2643,N_2325,N_2439);
nand U2644 (N_2644,N_2264,N_2014);
and U2645 (N_2645,N_2164,N_2499);
or U2646 (N_2646,N_2342,N_2463);
or U2647 (N_2647,N_2057,N_2289);
or U2648 (N_2648,N_2080,N_2361);
and U2649 (N_2649,N_2332,N_2091);
nor U2650 (N_2650,N_2406,N_2259);
and U2651 (N_2651,N_2495,N_2238);
or U2652 (N_2652,N_2064,N_2295);
nor U2653 (N_2653,N_2114,N_2146);
nand U2654 (N_2654,N_2142,N_2303);
nor U2655 (N_2655,N_2204,N_2216);
xnor U2656 (N_2656,N_2273,N_2328);
nor U2657 (N_2657,N_2243,N_2130);
and U2658 (N_2658,N_2405,N_2150);
nand U2659 (N_2659,N_2135,N_2039);
and U2660 (N_2660,N_2414,N_2097);
nand U2661 (N_2661,N_2320,N_2444);
and U2662 (N_2662,N_2430,N_2015);
and U2663 (N_2663,N_2420,N_2378);
and U2664 (N_2664,N_2319,N_2041);
and U2665 (N_2665,N_2341,N_2124);
or U2666 (N_2666,N_2231,N_2085);
nor U2667 (N_2667,N_2496,N_2494);
nor U2668 (N_2668,N_2148,N_2089);
nand U2669 (N_2669,N_2456,N_2107);
xor U2670 (N_2670,N_2386,N_2003);
or U2671 (N_2671,N_2326,N_2113);
and U2672 (N_2672,N_2194,N_2434);
or U2673 (N_2673,N_2347,N_2016);
and U2674 (N_2674,N_2200,N_2122);
and U2675 (N_2675,N_2224,N_2078);
xor U2676 (N_2676,N_2441,N_2316);
nor U2677 (N_2677,N_2308,N_2427);
nor U2678 (N_2678,N_2346,N_2047);
nand U2679 (N_2679,N_2334,N_2448);
xnor U2680 (N_2680,N_2486,N_2237);
nand U2681 (N_2681,N_2422,N_2452);
or U2682 (N_2682,N_2169,N_2087);
or U2683 (N_2683,N_2374,N_2186);
xor U2684 (N_2684,N_2301,N_2363);
nand U2685 (N_2685,N_2141,N_2239);
or U2686 (N_2686,N_2109,N_2208);
and U2687 (N_2687,N_2103,N_2210);
xnor U2688 (N_2688,N_2063,N_2459);
nand U2689 (N_2689,N_2147,N_2105);
and U2690 (N_2690,N_2209,N_2075);
or U2691 (N_2691,N_2212,N_2391);
or U2692 (N_2692,N_2385,N_2497);
nand U2693 (N_2693,N_2426,N_2443);
xnor U2694 (N_2694,N_2413,N_2013);
or U2695 (N_2695,N_2284,N_2246);
nand U2696 (N_2696,N_2309,N_2292);
or U2697 (N_2697,N_2271,N_2397);
nor U2698 (N_2698,N_2132,N_2394);
nor U2699 (N_2699,N_2393,N_2029);
nand U2700 (N_2700,N_2366,N_2317);
or U2701 (N_2701,N_2333,N_2145);
and U2702 (N_2702,N_2389,N_2233);
and U2703 (N_2703,N_2182,N_2010);
and U2704 (N_2704,N_2034,N_2383);
nor U2705 (N_2705,N_2353,N_2272);
nand U2706 (N_2706,N_2256,N_2395);
and U2707 (N_2707,N_2048,N_2380);
nand U2708 (N_2708,N_2213,N_2450);
or U2709 (N_2709,N_2083,N_2008);
xnor U2710 (N_2710,N_2266,N_2279);
and U2711 (N_2711,N_2096,N_2188);
and U2712 (N_2712,N_2323,N_2265);
xor U2713 (N_2713,N_2475,N_2191);
or U2714 (N_2714,N_2262,N_2020);
and U2715 (N_2715,N_2163,N_2036);
nor U2716 (N_2716,N_2258,N_2086);
xnor U2717 (N_2717,N_2043,N_2402);
nand U2718 (N_2718,N_2059,N_2412);
or U2719 (N_2719,N_2359,N_2007);
nor U2720 (N_2720,N_2081,N_2184);
nor U2721 (N_2721,N_2348,N_2403);
or U2722 (N_2722,N_2011,N_2381);
nor U2723 (N_2723,N_2084,N_2404);
xor U2724 (N_2724,N_2335,N_2102);
and U2725 (N_2725,N_2300,N_2028);
nor U2726 (N_2726,N_2240,N_2428);
nor U2727 (N_2727,N_2066,N_2251);
nor U2728 (N_2728,N_2022,N_2291);
xor U2729 (N_2729,N_2143,N_2218);
nand U2730 (N_2730,N_2037,N_2033);
and U2731 (N_2731,N_2067,N_2468);
and U2732 (N_2732,N_2387,N_2481);
and U2733 (N_2733,N_2175,N_2421);
or U2734 (N_2734,N_2384,N_2232);
or U2735 (N_2735,N_2451,N_2360);
or U2736 (N_2736,N_2372,N_2112);
and U2737 (N_2737,N_2162,N_2042);
nand U2738 (N_2738,N_2369,N_2432);
and U2739 (N_2739,N_2001,N_2088);
or U2740 (N_2740,N_2077,N_2051);
nor U2741 (N_2741,N_2190,N_2002);
nor U2742 (N_2742,N_2160,N_2128);
and U2743 (N_2743,N_2079,N_2215);
nor U2744 (N_2744,N_2100,N_2314);
nor U2745 (N_2745,N_2398,N_2431);
xnor U2746 (N_2746,N_2469,N_2005);
nor U2747 (N_2747,N_2351,N_2248);
and U2748 (N_2748,N_2330,N_2276);
or U2749 (N_2749,N_2263,N_2023);
nor U2750 (N_2750,N_2164,N_2461);
and U2751 (N_2751,N_2494,N_2374);
and U2752 (N_2752,N_2426,N_2358);
nor U2753 (N_2753,N_2152,N_2176);
xor U2754 (N_2754,N_2188,N_2055);
xor U2755 (N_2755,N_2314,N_2034);
and U2756 (N_2756,N_2238,N_2436);
nand U2757 (N_2757,N_2099,N_2105);
nand U2758 (N_2758,N_2324,N_2379);
or U2759 (N_2759,N_2484,N_2331);
and U2760 (N_2760,N_2484,N_2159);
nor U2761 (N_2761,N_2403,N_2111);
and U2762 (N_2762,N_2415,N_2274);
nor U2763 (N_2763,N_2079,N_2420);
or U2764 (N_2764,N_2365,N_2246);
and U2765 (N_2765,N_2119,N_2384);
nand U2766 (N_2766,N_2420,N_2198);
and U2767 (N_2767,N_2479,N_2477);
nor U2768 (N_2768,N_2098,N_2068);
and U2769 (N_2769,N_2425,N_2068);
and U2770 (N_2770,N_2127,N_2371);
and U2771 (N_2771,N_2330,N_2109);
and U2772 (N_2772,N_2305,N_2343);
and U2773 (N_2773,N_2183,N_2009);
nand U2774 (N_2774,N_2325,N_2329);
or U2775 (N_2775,N_2084,N_2105);
nand U2776 (N_2776,N_2279,N_2162);
or U2777 (N_2777,N_2227,N_2003);
or U2778 (N_2778,N_2080,N_2107);
nand U2779 (N_2779,N_2024,N_2286);
nand U2780 (N_2780,N_2221,N_2260);
or U2781 (N_2781,N_2046,N_2246);
or U2782 (N_2782,N_2389,N_2117);
and U2783 (N_2783,N_2443,N_2195);
and U2784 (N_2784,N_2398,N_2284);
nand U2785 (N_2785,N_2312,N_2230);
or U2786 (N_2786,N_2253,N_2258);
and U2787 (N_2787,N_2171,N_2105);
or U2788 (N_2788,N_2360,N_2477);
and U2789 (N_2789,N_2131,N_2244);
or U2790 (N_2790,N_2381,N_2073);
and U2791 (N_2791,N_2171,N_2240);
nor U2792 (N_2792,N_2499,N_2298);
and U2793 (N_2793,N_2183,N_2289);
and U2794 (N_2794,N_2155,N_2113);
nand U2795 (N_2795,N_2388,N_2048);
nor U2796 (N_2796,N_2025,N_2424);
and U2797 (N_2797,N_2081,N_2352);
xor U2798 (N_2798,N_2368,N_2400);
or U2799 (N_2799,N_2475,N_2154);
nor U2800 (N_2800,N_2274,N_2136);
or U2801 (N_2801,N_2202,N_2190);
nor U2802 (N_2802,N_2449,N_2326);
and U2803 (N_2803,N_2258,N_2405);
nor U2804 (N_2804,N_2081,N_2017);
and U2805 (N_2805,N_2282,N_2146);
and U2806 (N_2806,N_2122,N_2073);
or U2807 (N_2807,N_2137,N_2445);
nand U2808 (N_2808,N_2149,N_2306);
nor U2809 (N_2809,N_2462,N_2186);
and U2810 (N_2810,N_2080,N_2268);
or U2811 (N_2811,N_2067,N_2174);
or U2812 (N_2812,N_2420,N_2000);
nand U2813 (N_2813,N_2121,N_2398);
nor U2814 (N_2814,N_2080,N_2002);
and U2815 (N_2815,N_2430,N_2216);
nand U2816 (N_2816,N_2316,N_2160);
nor U2817 (N_2817,N_2124,N_2220);
xnor U2818 (N_2818,N_2026,N_2075);
or U2819 (N_2819,N_2077,N_2212);
and U2820 (N_2820,N_2021,N_2438);
or U2821 (N_2821,N_2340,N_2481);
nand U2822 (N_2822,N_2265,N_2422);
and U2823 (N_2823,N_2040,N_2265);
or U2824 (N_2824,N_2280,N_2188);
and U2825 (N_2825,N_2182,N_2280);
nand U2826 (N_2826,N_2337,N_2049);
xnor U2827 (N_2827,N_2178,N_2091);
and U2828 (N_2828,N_2220,N_2389);
nand U2829 (N_2829,N_2289,N_2211);
or U2830 (N_2830,N_2173,N_2218);
nor U2831 (N_2831,N_2430,N_2401);
and U2832 (N_2832,N_2205,N_2038);
nor U2833 (N_2833,N_2213,N_2391);
nor U2834 (N_2834,N_2333,N_2264);
nand U2835 (N_2835,N_2055,N_2007);
nor U2836 (N_2836,N_2326,N_2479);
or U2837 (N_2837,N_2074,N_2006);
or U2838 (N_2838,N_2053,N_2413);
nand U2839 (N_2839,N_2234,N_2004);
or U2840 (N_2840,N_2351,N_2387);
or U2841 (N_2841,N_2490,N_2298);
nand U2842 (N_2842,N_2181,N_2179);
nand U2843 (N_2843,N_2114,N_2106);
nand U2844 (N_2844,N_2130,N_2172);
and U2845 (N_2845,N_2065,N_2405);
xnor U2846 (N_2846,N_2338,N_2420);
nand U2847 (N_2847,N_2365,N_2217);
nand U2848 (N_2848,N_2496,N_2211);
and U2849 (N_2849,N_2223,N_2181);
nand U2850 (N_2850,N_2286,N_2136);
and U2851 (N_2851,N_2442,N_2198);
and U2852 (N_2852,N_2336,N_2210);
xor U2853 (N_2853,N_2258,N_2213);
nor U2854 (N_2854,N_2135,N_2491);
and U2855 (N_2855,N_2093,N_2291);
and U2856 (N_2856,N_2472,N_2376);
nand U2857 (N_2857,N_2118,N_2171);
or U2858 (N_2858,N_2134,N_2084);
nand U2859 (N_2859,N_2067,N_2199);
xnor U2860 (N_2860,N_2189,N_2230);
nor U2861 (N_2861,N_2188,N_2332);
nand U2862 (N_2862,N_2034,N_2451);
and U2863 (N_2863,N_2016,N_2029);
or U2864 (N_2864,N_2341,N_2051);
nand U2865 (N_2865,N_2402,N_2243);
nand U2866 (N_2866,N_2458,N_2064);
or U2867 (N_2867,N_2435,N_2467);
or U2868 (N_2868,N_2051,N_2225);
nand U2869 (N_2869,N_2235,N_2199);
and U2870 (N_2870,N_2073,N_2005);
and U2871 (N_2871,N_2160,N_2051);
nand U2872 (N_2872,N_2156,N_2172);
nor U2873 (N_2873,N_2300,N_2359);
xor U2874 (N_2874,N_2484,N_2275);
or U2875 (N_2875,N_2182,N_2150);
xor U2876 (N_2876,N_2186,N_2013);
nand U2877 (N_2877,N_2338,N_2337);
or U2878 (N_2878,N_2032,N_2262);
and U2879 (N_2879,N_2427,N_2433);
nand U2880 (N_2880,N_2351,N_2187);
and U2881 (N_2881,N_2343,N_2020);
and U2882 (N_2882,N_2170,N_2109);
nor U2883 (N_2883,N_2046,N_2331);
or U2884 (N_2884,N_2169,N_2430);
nand U2885 (N_2885,N_2124,N_2494);
nor U2886 (N_2886,N_2067,N_2354);
xnor U2887 (N_2887,N_2410,N_2360);
xnor U2888 (N_2888,N_2292,N_2394);
and U2889 (N_2889,N_2345,N_2064);
and U2890 (N_2890,N_2306,N_2329);
or U2891 (N_2891,N_2041,N_2084);
or U2892 (N_2892,N_2338,N_2125);
and U2893 (N_2893,N_2368,N_2138);
nand U2894 (N_2894,N_2065,N_2207);
xnor U2895 (N_2895,N_2463,N_2027);
nand U2896 (N_2896,N_2180,N_2494);
nor U2897 (N_2897,N_2056,N_2255);
nor U2898 (N_2898,N_2087,N_2270);
or U2899 (N_2899,N_2005,N_2198);
xor U2900 (N_2900,N_2490,N_2166);
nand U2901 (N_2901,N_2301,N_2498);
nor U2902 (N_2902,N_2236,N_2421);
xor U2903 (N_2903,N_2224,N_2316);
nand U2904 (N_2904,N_2202,N_2157);
nand U2905 (N_2905,N_2001,N_2143);
or U2906 (N_2906,N_2085,N_2125);
and U2907 (N_2907,N_2281,N_2475);
nor U2908 (N_2908,N_2041,N_2228);
nor U2909 (N_2909,N_2446,N_2009);
and U2910 (N_2910,N_2054,N_2251);
or U2911 (N_2911,N_2023,N_2413);
nor U2912 (N_2912,N_2060,N_2251);
or U2913 (N_2913,N_2051,N_2261);
and U2914 (N_2914,N_2194,N_2252);
nand U2915 (N_2915,N_2065,N_2086);
or U2916 (N_2916,N_2080,N_2001);
nand U2917 (N_2917,N_2059,N_2135);
and U2918 (N_2918,N_2439,N_2245);
or U2919 (N_2919,N_2425,N_2440);
nor U2920 (N_2920,N_2326,N_2126);
or U2921 (N_2921,N_2009,N_2398);
nor U2922 (N_2922,N_2368,N_2032);
nor U2923 (N_2923,N_2177,N_2493);
nor U2924 (N_2924,N_2459,N_2037);
or U2925 (N_2925,N_2467,N_2453);
nand U2926 (N_2926,N_2028,N_2483);
nand U2927 (N_2927,N_2045,N_2296);
nor U2928 (N_2928,N_2104,N_2336);
and U2929 (N_2929,N_2376,N_2482);
xnor U2930 (N_2930,N_2192,N_2027);
or U2931 (N_2931,N_2175,N_2487);
nand U2932 (N_2932,N_2062,N_2225);
or U2933 (N_2933,N_2139,N_2307);
and U2934 (N_2934,N_2052,N_2061);
nor U2935 (N_2935,N_2240,N_2257);
nor U2936 (N_2936,N_2341,N_2457);
nand U2937 (N_2937,N_2282,N_2244);
or U2938 (N_2938,N_2220,N_2419);
or U2939 (N_2939,N_2226,N_2077);
nand U2940 (N_2940,N_2229,N_2300);
or U2941 (N_2941,N_2056,N_2168);
nand U2942 (N_2942,N_2341,N_2194);
and U2943 (N_2943,N_2319,N_2005);
and U2944 (N_2944,N_2452,N_2402);
xnor U2945 (N_2945,N_2247,N_2222);
and U2946 (N_2946,N_2365,N_2368);
or U2947 (N_2947,N_2086,N_2234);
and U2948 (N_2948,N_2441,N_2467);
and U2949 (N_2949,N_2194,N_2224);
and U2950 (N_2950,N_2046,N_2324);
nand U2951 (N_2951,N_2371,N_2076);
and U2952 (N_2952,N_2330,N_2312);
and U2953 (N_2953,N_2250,N_2048);
nand U2954 (N_2954,N_2062,N_2213);
xnor U2955 (N_2955,N_2467,N_2277);
and U2956 (N_2956,N_2388,N_2454);
nand U2957 (N_2957,N_2129,N_2002);
and U2958 (N_2958,N_2260,N_2361);
and U2959 (N_2959,N_2128,N_2287);
and U2960 (N_2960,N_2361,N_2202);
nand U2961 (N_2961,N_2037,N_2348);
and U2962 (N_2962,N_2492,N_2259);
nand U2963 (N_2963,N_2209,N_2419);
nor U2964 (N_2964,N_2086,N_2023);
or U2965 (N_2965,N_2076,N_2352);
nand U2966 (N_2966,N_2231,N_2130);
nand U2967 (N_2967,N_2339,N_2341);
and U2968 (N_2968,N_2471,N_2226);
xnor U2969 (N_2969,N_2194,N_2219);
or U2970 (N_2970,N_2380,N_2190);
nor U2971 (N_2971,N_2056,N_2034);
xor U2972 (N_2972,N_2024,N_2363);
xnor U2973 (N_2973,N_2443,N_2060);
nand U2974 (N_2974,N_2450,N_2009);
nor U2975 (N_2975,N_2402,N_2014);
nand U2976 (N_2976,N_2371,N_2085);
nand U2977 (N_2977,N_2361,N_2009);
and U2978 (N_2978,N_2154,N_2449);
nor U2979 (N_2979,N_2139,N_2370);
xnor U2980 (N_2980,N_2252,N_2074);
nand U2981 (N_2981,N_2030,N_2490);
nand U2982 (N_2982,N_2405,N_2388);
and U2983 (N_2983,N_2477,N_2417);
and U2984 (N_2984,N_2466,N_2226);
nor U2985 (N_2985,N_2098,N_2206);
nor U2986 (N_2986,N_2169,N_2083);
nand U2987 (N_2987,N_2035,N_2002);
nand U2988 (N_2988,N_2222,N_2216);
xor U2989 (N_2989,N_2493,N_2026);
xnor U2990 (N_2990,N_2410,N_2234);
or U2991 (N_2991,N_2473,N_2267);
nand U2992 (N_2992,N_2036,N_2362);
nor U2993 (N_2993,N_2302,N_2187);
and U2994 (N_2994,N_2072,N_2300);
nor U2995 (N_2995,N_2368,N_2489);
nor U2996 (N_2996,N_2318,N_2422);
nor U2997 (N_2997,N_2102,N_2096);
or U2998 (N_2998,N_2149,N_2384);
and U2999 (N_2999,N_2293,N_2017);
or U3000 (N_3000,N_2993,N_2627);
nor U3001 (N_3001,N_2587,N_2671);
or U3002 (N_3002,N_2878,N_2711);
nand U3003 (N_3003,N_2669,N_2905);
or U3004 (N_3004,N_2638,N_2663);
or U3005 (N_3005,N_2557,N_2822);
or U3006 (N_3006,N_2592,N_2885);
nand U3007 (N_3007,N_2992,N_2629);
and U3008 (N_3008,N_2736,N_2668);
nor U3009 (N_3009,N_2730,N_2820);
and U3010 (N_3010,N_2771,N_2725);
and U3011 (N_3011,N_2862,N_2751);
and U3012 (N_3012,N_2677,N_2778);
nor U3013 (N_3013,N_2833,N_2781);
nor U3014 (N_3014,N_2787,N_2691);
nand U3015 (N_3015,N_2943,N_2721);
nor U3016 (N_3016,N_2966,N_2786);
nor U3017 (N_3017,N_2983,N_2731);
nor U3018 (N_3018,N_2869,N_2904);
nor U3019 (N_3019,N_2584,N_2750);
nand U3020 (N_3020,N_2648,N_2615);
and U3021 (N_3021,N_2875,N_2617);
and U3022 (N_3022,N_2957,N_2856);
nand U3023 (N_3023,N_2985,N_2623);
nand U3024 (N_3024,N_2806,N_2548);
and U3025 (N_3025,N_2998,N_2549);
nand U3026 (N_3026,N_2819,N_2792);
nor U3027 (N_3027,N_2956,N_2754);
nand U3028 (N_3028,N_2683,N_2760);
and U3029 (N_3029,N_2534,N_2612);
and U3030 (N_3030,N_2641,N_2670);
nand U3031 (N_3031,N_2618,N_2765);
xor U3032 (N_3032,N_2817,N_2915);
nand U3033 (N_3033,N_2673,N_2969);
xor U3034 (N_3034,N_2515,N_2928);
nor U3035 (N_3035,N_2883,N_2748);
nor U3036 (N_3036,N_2593,N_2766);
nand U3037 (N_3037,N_2934,N_2724);
and U3038 (N_3038,N_2620,N_2844);
nor U3039 (N_3039,N_2594,N_2961);
nand U3040 (N_3040,N_2718,N_2597);
nand U3041 (N_3041,N_2810,N_2968);
nor U3042 (N_3042,N_2890,N_2936);
or U3043 (N_3043,N_2954,N_2876);
and U3044 (N_3044,N_2995,N_2636);
or U3045 (N_3045,N_2520,N_2893);
or U3046 (N_3046,N_2749,N_2982);
nand U3047 (N_3047,N_2884,N_2632);
or U3048 (N_3048,N_2656,N_2588);
nor U3049 (N_3049,N_2811,N_2753);
xor U3050 (N_3050,N_2624,N_2797);
and U3051 (N_3051,N_2951,N_2897);
nor U3052 (N_3052,N_2855,N_2959);
nor U3053 (N_3053,N_2614,N_2681);
nor U3054 (N_3054,N_2772,N_2764);
nor U3055 (N_3055,N_2676,N_2963);
and U3056 (N_3056,N_2744,N_2733);
xnor U3057 (N_3057,N_2531,N_2794);
nor U3058 (N_3058,N_2907,N_2726);
and U3059 (N_3059,N_2901,N_2767);
and U3060 (N_3060,N_2542,N_2571);
and U3061 (N_3061,N_2740,N_2812);
xor U3062 (N_3062,N_2834,N_2729);
or U3063 (N_3063,N_2836,N_2927);
nand U3064 (N_3064,N_2821,N_2570);
or U3065 (N_3065,N_2581,N_2563);
nand U3066 (N_3066,N_2518,N_2840);
or U3067 (N_3067,N_2679,N_2761);
nor U3068 (N_3068,N_2888,N_2853);
and U3069 (N_3069,N_2860,N_2599);
nand U3070 (N_3070,N_2657,N_2947);
and U3071 (N_3071,N_2950,N_2949);
and U3072 (N_3072,N_2984,N_2756);
xor U3073 (N_3073,N_2607,N_2933);
nand U3074 (N_3074,N_2953,N_2872);
nor U3075 (N_3075,N_2573,N_2622);
nor U3076 (N_3076,N_2535,N_2835);
nor U3077 (N_3077,N_2757,N_2988);
or U3078 (N_3078,N_2654,N_2578);
nand U3079 (N_3079,N_2640,N_2604);
xnor U3080 (N_3080,N_2980,N_2521);
xnor U3081 (N_3081,N_2987,N_2831);
nand U3082 (N_3082,N_2560,N_2738);
nor U3083 (N_3083,N_2849,N_2500);
and U3084 (N_3084,N_2804,N_2805);
or U3085 (N_3085,N_2965,N_2802);
xnor U3086 (N_3086,N_2783,N_2637);
nand U3087 (N_3087,N_2868,N_2874);
nand U3088 (N_3088,N_2684,N_2867);
or U3089 (N_3089,N_2758,N_2643);
or U3090 (N_3090,N_2687,N_2559);
xnor U3091 (N_3091,N_2903,N_2938);
and U3092 (N_3092,N_2672,N_2715);
nor U3093 (N_3093,N_2958,N_2543);
nor U3094 (N_3094,N_2908,N_2782);
nand U3095 (N_3095,N_2539,N_2556);
and U3096 (N_3096,N_2707,N_2722);
nand U3097 (N_3097,N_2603,N_2871);
xnor U3098 (N_3098,N_2800,N_2839);
nor U3099 (N_3099,N_2913,N_2944);
xor U3100 (N_3100,N_2937,N_2553);
nor U3101 (N_3101,N_2680,N_2635);
xnor U3102 (N_3102,N_2659,N_2994);
nand U3103 (N_3103,N_2743,N_2658);
or U3104 (N_3104,N_2507,N_2986);
or U3105 (N_3105,N_2630,N_2894);
nor U3106 (N_3106,N_2864,N_2540);
or U3107 (N_3107,N_2583,N_2664);
or U3108 (N_3108,N_2526,N_2912);
or U3109 (N_3109,N_2523,N_2688);
and U3110 (N_3110,N_2837,N_2686);
or U3111 (N_3111,N_2935,N_2891);
nand U3112 (N_3112,N_2970,N_2705);
nor U3113 (N_3113,N_2973,N_2896);
and U3114 (N_3114,N_2512,N_2595);
nand U3115 (N_3115,N_2555,N_2914);
nand U3116 (N_3116,N_2841,N_2606);
nand U3117 (N_3117,N_2788,N_2698);
nor U3118 (N_3118,N_2880,N_2941);
nand U3119 (N_3119,N_2922,N_2533);
nand U3120 (N_3120,N_2703,N_2601);
nor U3121 (N_3121,N_2742,N_2784);
nand U3122 (N_3122,N_2530,N_2886);
nand U3123 (N_3123,N_2851,N_2706);
nand U3124 (N_3124,N_2785,N_2644);
xor U3125 (N_3125,N_2699,N_2911);
or U3126 (N_3126,N_2589,N_2979);
xor U3127 (N_3127,N_2946,N_2762);
or U3128 (N_3128,N_2974,N_2999);
and U3129 (N_3129,N_2900,N_2552);
nor U3130 (N_3130,N_2926,N_2532);
nor U3131 (N_3131,N_2895,N_2769);
or U3132 (N_3132,N_2972,N_2892);
nand U3133 (N_3133,N_2678,N_2824);
or U3134 (N_3134,N_2608,N_2651);
and U3135 (N_3135,N_2536,N_2793);
xnor U3136 (N_3136,N_2716,N_2924);
xor U3137 (N_3137,N_2858,N_2977);
and U3138 (N_3138,N_2675,N_2967);
nand U3139 (N_3139,N_2830,N_2546);
nor U3140 (N_3140,N_2777,N_2551);
nor U3141 (N_3141,N_2667,N_2501);
xnor U3142 (N_3142,N_2661,N_2976);
nand U3143 (N_3143,N_2565,N_2510);
or U3144 (N_3144,N_2791,N_2544);
and U3145 (N_3145,N_2550,N_2505);
nand U3146 (N_3146,N_2779,N_2879);
and U3147 (N_3147,N_2930,N_2650);
or U3148 (N_3148,N_2918,N_2889);
and U3149 (N_3149,N_2942,N_2741);
or U3150 (N_3150,N_2978,N_2865);
or U3151 (N_3151,N_2964,N_2613);
nor U3152 (N_3152,N_2734,N_2576);
and U3153 (N_3153,N_2780,N_2732);
or U3154 (N_3154,N_2932,N_2558);
or U3155 (N_3155,N_2859,N_2666);
or U3156 (N_3156,N_2713,N_2795);
nor U3157 (N_3157,N_2939,N_2720);
or U3158 (N_3158,N_2955,N_2665);
and U3159 (N_3159,N_2909,N_2971);
nor U3160 (N_3160,N_2598,N_2575);
or U3161 (N_3161,N_2633,N_2857);
nand U3162 (N_3162,N_2585,N_2642);
or U3163 (N_3163,N_2799,N_2517);
or U3164 (N_3164,N_2846,N_2682);
xnor U3165 (N_3165,N_2694,N_2631);
nor U3166 (N_3166,N_2990,N_2850);
xnor U3167 (N_3167,N_2823,N_2626);
and U3168 (N_3168,N_2747,N_2605);
nand U3169 (N_3169,N_2775,N_2996);
nand U3170 (N_3170,N_2728,N_2674);
nor U3171 (N_3171,N_2712,N_2768);
or U3172 (N_3172,N_2945,N_2528);
nand U3173 (N_3173,N_2649,N_2723);
nor U3174 (N_3174,N_2847,N_2801);
nand U3175 (N_3175,N_2991,N_2647);
or U3176 (N_3176,N_2541,N_2739);
and U3177 (N_3177,N_2899,N_2763);
or U3178 (N_3178,N_2848,N_2770);
xor U3179 (N_3179,N_2808,N_2975);
nand U3180 (N_3180,N_2610,N_2870);
nor U3181 (N_3181,N_2522,N_2561);
nor U3182 (N_3182,N_2816,N_2693);
xnor U3183 (N_3183,N_2828,N_2568);
nor U3184 (N_3184,N_2818,N_2745);
and U3185 (N_3185,N_2702,N_2696);
nand U3186 (N_3186,N_2514,N_2873);
xnor U3187 (N_3187,N_2809,N_2572);
or U3188 (N_3188,N_2685,N_2695);
and U3189 (N_3189,N_2815,N_2591);
or U3190 (N_3190,N_2602,N_2566);
and U3191 (N_3191,N_2746,N_2917);
nand U3192 (N_3192,N_2960,N_2519);
nand U3193 (N_3193,N_2628,N_2925);
or U3194 (N_3194,N_2652,N_2826);
or U3195 (N_3195,N_2537,N_2854);
or U3196 (N_3196,N_2827,N_2735);
nand U3197 (N_3197,N_2861,N_2655);
and U3198 (N_3198,N_2527,N_2852);
and U3199 (N_3199,N_2564,N_2940);
nand U3200 (N_3200,N_2887,N_2902);
or U3201 (N_3201,N_2653,N_2717);
nor U3202 (N_3202,N_2529,N_2727);
or U3203 (N_3203,N_2710,N_2962);
or U3204 (N_3204,N_2525,N_2863);
nand U3205 (N_3205,N_2919,N_2755);
or U3206 (N_3206,N_2577,N_2619);
or U3207 (N_3207,N_2759,N_2662);
nor U3208 (N_3208,N_2646,N_2590);
xnor U3209 (N_3209,N_2790,N_2814);
xnor U3210 (N_3210,N_2625,N_2952);
and U3211 (N_3211,N_2877,N_2600);
nor U3212 (N_3212,N_2838,N_2547);
or U3213 (N_3213,N_2586,N_2714);
or U3214 (N_3214,N_2773,N_2910);
nand U3215 (N_3215,N_2579,N_2832);
nor U3216 (N_3216,N_2916,N_2789);
or U3217 (N_3217,N_2803,N_2906);
xnor U3218 (N_3218,N_2708,N_2881);
nand U3219 (N_3219,N_2866,N_2511);
or U3220 (N_3220,N_2562,N_2639);
or U3221 (N_3221,N_2616,N_2660);
nand U3222 (N_3222,N_2538,N_2545);
or U3223 (N_3223,N_2989,N_2508);
nand U3224 (N_3224,N_2898,N_2574);
xor U3225 (N_3225,N_2524,N_2690);
and U3226 (N_3226,N_2621,N_2709);
nor U3227 (N_3227,N_2567,N_2813);
or U3228 (N_3228,N_2609,N_2645);
and U3229 (N_3229,N_2923,N_2843);
or U3230 (N_3230,N_2554,N_2774);
nand U3231 (N_3231,N_2506,N_2796);
nand U3232 (N_3232,N_2689,N_2504);
or U3233 (N_3233,N_2697,N_2502);
and U3234 (N_3234,N_2997,N_2845);
nor U3235 (N_3235,N_2737,N_2700);
and U3236 (N_3236,N_2825,N_2948);
and U3237 (N_3237,N_2634,N_2503);
nor U3238 (N_3238,N_2516,N_2829);
nand U3239 (N_3239,N_2704,N_2580);
and U3240 (N_3240,N_2929,N_2882);
and U3241 (N_3241,N_2692,N_2931);
nand U3242 (N_3242,N_2807,N_2719);
or U3243 (N_3243,N_2921,N_2582);
nor U3244 (N_3244,N_2596,N_2920);
nor U3245 (N_3245,N_2776,N_2981);
nor U3246 (N_3246,N_2752,N_2842);
and U3247 (N_3247,N_2513,N_2798);
nor U3248 (N_3248,N_2569,N_2611);
nor U3249 (N_3249,N_2509,N_2701);
nand U3250 (N_3250,N_2994,N_2851);
nand U3251 (N_3251,N_2941,N_2562);
or U3252 (N_3252,N_2834,N_2557);
or U3253 (N_3253,N_2709,N_2734);
nand U3254 (N_3254,N_2723,N_2781);
or U3255 (N_3255,N_2851,N_2911);
or U3256 (N_3256,N_2550,N_2588);
or U3257 (N_3257,N_2999,N_2936);
xor U3258 (N_3258,N_2888,N_2610);
and U3259 (N_3259,N_2819,N_2536);
and U3260 (N_3260,N_2634,N_2875);
or U3261 (N_3261,N_2930,N_2750);
and U3262 (N_3262,N_2690,N_2704);
and U3263 (N_3263,N_2887,N_2528);
and U3264 (N_3264,N_2868,N_2612);
or U3265 (N_3265,N_2622,N_2746);
or U3266 (N_3266,N_2761,N_2967);
nand U3267 (N_3267,N_2922,N_2969);
or U3268 (N_3268,N_2896,N_2544);
nor U3269 (N_3269,N_2706,N_2841);
nor U3270 (N_3270,N_2904,N_2914);
nand U3271 (N_3271,N_2800,N_2726);
xor U3272 (N_3272,N_2966,N_2977);
nand U3273 (N_3273,N_2534,N_2699);
or U3274 (N_3274,N_2543,N_2516);
nand U3275 (N_3275,N_2693,N_2690);
nor U3276 (N_3276,N_2918,N_2592);
or U3277 (N_3277,N_2687,N_2782);
and U3278 (N_3278,N_2923,N_2706);
nor U3279 (N_3279,N_2796,N_2987);
and U3280 (N_3280,N_2731,N_2613);
nor U3281 (N_3281,N_2885,N_2766);
nor U3282 (N_3282,N_2685,N_2564);
and U3283 (N_3283,N_2656,N_2741);
and U3284 (N_3284,N_2608,N_2785);
and U3285 (N_3285,N_2553,N_2756);
or U3286 (N_3286,N_2993,N_2924);
xor U3287 (N_3287,N_2634,N_2976);
and U3288 (N_3288,N_2693,N_2627);
and U3289 (N_3289,N_2560,N_2770);
and U3290 (N_3290,N_2822,N_2968);
xor U3291 (N_3291,N_2500,N_2614);
nor U3292 (N_3292,N_2539,N_2591);
or U3293 (N_3293,N_2502,N_2688);
and U3294 (N_3294,N_2767,N_2949);
or U3295 (N_3295,N_2527,N_2857);
xnor U3296 (N_3296,N_2719,N_2505);
and U3297 (N_3297,N_2776,N_2659);
nor U3298 (N_3298,N_2655,N_2668);
or U3299 (N_3299,N_2737,N_2816);
and U3300 (N_3300,N_2861,N_2958);
nor U3301 (N_3301,N_2555,N_2790);
nor U3302 (N_3302,N_2569,N_2612);
nand U3303 (N_3303,N_2569,N_2733);
nor U3304 (N_3304,N_2742,N_2807);
or U3305 (N_3305,N_2599,N_2953);
or U3306 (N_3306,N_2583,N_2916);
and U3307 (N_3307,N_2948,N_2671);
or U3308 (N_3308,N_2551,N_2906);
nand U3309 (N_3309,N_2653,N_2758);
nor U3310 (N_3310,N_2888,N_2657);
and U3311 (N_3311,N_2568,N_2991);
and U3312 (N_3312,N_2502,N_2940);
nor U3313 (N_3313,N_2516,N_2805);
nor U3314 (N_3314,N_2830,N_2615);
and U3315 (N_3315,N_2556,N_2773);
nand U3316 (N_3316,N_2691,N_2635);
nand U3317 (N_3317,N_2589,N_2972);
or U3318 (N_3318,N_2549,N_2919);
xnor U3319 (N_3319,N_2909,N_2812);
nand U3320 (N_3320,N_2892,N_2962);
nor U3321 (N_3321,N_2730,N_2695);
or U3322 (N_3322,N_2518,N_2602);
or U3323 (N_3323,N_2612,N_2524);
and U3324 (N_3324,N_2596,N_2858);
xor U3325 (N_3325,N_2592,N_2676);
nor U3326 (N_3326,N_2747,N_2552);
and U3327 (N_3327,N_2801,N_2613);
or U3328 (N_3328,N_2625,N_2951);
or U3329 (N_3329,N_2893,N_2786);
or U3330 (N_3330,N_2734,N_2877);
nand U3331 (N_3331,N_2807,N_2653);
or U3332 (N_3332,N_2554,N_2807);
and U3333 (N_3333,N_2514,N_2523);
or U3334 (N_3334,N_2879,N_2587);
nor U3335 (N_3335,N_2788,N_2529);
nand U3336 (N_3336,N_2572,N_2997);
nand U3337 (N_3337,N_2922,N_2949);
or U3338 (N_3338,N_2951,N_2626);
nor U3339 (N_3339,N_2942,N_2764);
nor U3340 (N_3340,N_2859,N_2991);
nor U3341 (N_3341,N_2807,N_2974);
and U3342 (N_3342,N_2636,N_2961);
nor U3343 (N_3343,N_2891,N_2957);
xor U3344 (N_3344,N_2593,N_2871);
nand U3345 (N_3345,N_2769,N_2560);
xor U3346 (N_3346,N_2684,N_2972);
and U3347 (N_3347,N_2755,N_2601);
and U3348 (N_3348,N_2538,N_2849);
nor U3349 (N_3349,N_2873,N_2565);
and U3350 (N_3350,N_2734,N_2524);
or U3351 (N_3351,N_2771,N_2678);
nand U3352 (N_3352,N_2943,N_2561);
nand U3353 (N_3353,N_2804,N_2683);
xor U3354 (N_3354,N_2987,N_2693);
or U3355 (N_3355,N_2756,N_2742);
or U3356 (N_3356,N_2573,N_2787);
nand U3357 (N_3357,N_2902,N_2804);
nor U3358 (N_3358,N_2548,N_2672);
nand U3359 (N_3359,N_2688,N_2777);
or U3360 (N_3360,N_2517,N_2924);
or U3361 (N_3361,N_2795,N_2528);
nor U3362 (N_3362,N_2872,N_2674);
xor U3363 (N_3363,N_2563,N_2556);
xnor U3364 (N_3364,N_2566,N_2654);
nand U3365 (N_3365,N_2626,N_2896);
or U3366 (N_3366,N_2525,N_2683);
nand U3367 (N_3367,N_2626,N_2946);
nor U3368 (N_3368,N_2881,N_2812);
and U3369 (N_3369,N_2737,N_2739);
nand U3370 (N_3370,N_2875,N_2821);
or U3371 (N_3371,N_2685,N_2623);
and U3372 (N_3372,N_2958,N_2502);
and U3373 (N_3373,N_2956,N_2643);
nand U3374 (N_3374,N_2763,N_2560);
and U3375 (N_3375,N_2806,N_2643);
nor U3376 (N_3376,N_2957,N_2675);
nand U3377 (N_3377,N_2696,N_2607);
nand U3378 (N_3378,N_2807,N_2863);
xor U3379 (N_3379,N_2964,N_2714);
nand U3380 (N_3380,N_2955,N_2730);
or U3381 (N_3381,N_2961,N_2643);
nand U3382 (N_3382,N_2853,N_2827);
and U3383 (N_3383,N_2919,N_2580);
or U3384 (N_3384,N_2993,N_2847);
nor U3385 (N_3385,N_2998,N_2858);
and U3386 (N_3386,N_2594,N_2993);
xnor U3387 (N_3387,N_2620,N_2820);
nor U3388 (N_3388,N_2516,N_2892);
nand U3389 (N_3389,N_2834,N_2674);
nand U3390 (N_3390,N_2864,N_2615);
nand U3391 (N_3391,N_2506,N_2645);
nor U3392 (N_3392,N_2605,N_2843);
nand U3393 (N_3393,N_2622,N_2987);
and U3394 (N_3394,N_2818,N_2674);
or U3395 (N_3395,N_2862,N_2926);
or U3396 (N_3396,N_2594,N_2617);
nor U3397 (N_3397,N_2679,N_2625);
or U3398 (N_3398,N_2923,N_2783);
nor U3399 (N_3399,N_2939,N_2793);
nor U3400 (N_3400,N_2973,N_2969);
nand U3401 (N_3401,N_2544,N_2852);
nand U3402 (N_3402,N_2516,N_2581);
and U3403 (N_3403,N_2595,N_2649);
and U3404 (N_3404,N_2632,N_2710);
nor U3405 (N_3405,N_2594,N_2684);
nor U3406 (N_3406,N_2515,N_2682);
and U3407 (N_3407,N_2665,N_2972);
nand U3408 (N_3408,N_2511,N_2910);
nand U3409 (N_3409,N_2625,N_2926);
nand U3410 (N_3410,N_2782,N_2565);
and U3411 (N_3411,N_2830,N_2929);
and U3412 (N_3412,N_2801,N_2568);
or U3413 (N_3413,N_2510,N_2969);
nor U3414 (N_3414,N_2566,N_2961);
nor U3415 (N_3415,N_2653,N_2510);
xor U3416 (N_3416,N_2555,N_2748);
nand U3417 (N_3417,N_2553,N_2880);
xor U3418 (N_3418,N_2889,N_2759);
nand U3419 (N_3419,N_2933,N_2858);
and U3420 (N_3420,N_2737,N_2710);
nor U3421 (N_3421,N_2824,N_2787);
nor U3422 (N_3422,N_2925,N_2546);
nand U3423 (N_3423,N_2678,N_2723);
and U3424 (N_3424,N_2935,N_2638);
nand U3425 (N_3425,N_2970,N_2905);
nand U3426 (N_3426,N_2701,N_2731);
nor U3427 (N_3427,N_2792,N_2658);
nand U3428 (N_3428,N_2574,N_2500);
nand U3429 (N_3429,N_2713,N_2988);
nor U3430 (N_3430,N_2964,N_2503);
nor U3431 (N_3431,N_2541,N_2850);
nor U3432 (N_3432,N_2748,N_2569);
and U3433 (N_3433,N_2841,N_2516);
or U3434 (N_3434,N_2805,N_2596);
and U3435 (N_3435,N_2824,N_2608);
or U3436 (N_3436,N_2768,N_2517);
nor U3437 (N_3437,N_2903,N_2622);
nor U3438 (N_3438,N_2707,N_2540);
or U3439 (N_3439,N_2550,N_2806);
and U3440 (N_3440,N_2806,N_2733);
nand U3441 (N_3441,N_2537,N_2955);
or U3442 (N_3442,N_2755,N_2981);
nor U3443 (N_3443,N_2909,N_2890);
and U3444 (N_3444,N_2904,N_2664);
and U3445 (N_3445,N_2610,N_2784);
and U3446 (N_3446,N_2836,N_2819);
and U3447 (N_3447,N_2705,N_2813);
nand U3448 (N_3448,N_2931,N_2828);
nor U3449 (N_3449,N_2538,N_2767);
nor U3450 (N_3450,N_2857,N_2740);
or U3451 (N_3451,N_2968,N_2931);
nand U3452 (N_3452,N_2588,N_2855);
and U3453 (N_3453,N_2718,N_2679);
nor U3454 (N_3454,N_2984,N_2619);
or U3455 (N_3455,N_2863,N_2741);
nor U3456 (N_3456,N_2832,N_2712);
and U3457 (N_3457,N_2908,N_2922);
nor U3458 (N_3458,N_2757,N_2627);
or U3459 (N_3459,N_2951,N_2738);
nor U3460 (N_3460,N_2667,N_2559);
or U3461 (N_3461,N_2819,N_2719);
nand U3462 (N_3462,N_2611,N_2550);
and U3463 (N_3463,N_2808,N_2659);
or U3464 (N_3464,N_2771,N_2510);
and U3465 (N_3465,N_2786,N_2793);
or U3466 (N_3466,N_2563,N_2605);
and U3467 (N_3467,N_2649,N_2771);
nor U3468 (N_3468,N_2762,N_2707);
or U3469 (N_3469,N_2560,N_2901);
nand U3470 (N_3470,N_2631,N_2563);
xor U3471 (N_3471,N_2866,N_2507);
or U3472 (N_3472,N_2745,N_2588);
nand U3473 (N_3473,N_2843,N_2716);
or U3474 (N_3474,N_2829,N_2950);
and U3475 (N_3475,N_2965,N_2982);
or U3476 (N_3476,N_2596,N_2738);
xor U3477 (N_3477,N_2656,N_2641);
or U3478 (N_3478,N_2591,N_2723);
nor U3479 (N_3479,N_2522,N_2596);
or U3480 (N_3480,N_2952,N_2659);
nor U3481 (N_3481,N_2676,N_2605);
and U3482 (N_3482,N_2505,N_2749);
nor U3483 (N_3483,N_2649,N_2945);
nor U3484 (N_3484,N_2667,N_2934);
xor U3485 (N_3485,N_2826,N_2655);
nor U3486 (N_3486,N_2522,N_2719);
xor U3487 (N_3487,N_2690,N_2760);
nand U3488 (N_3488,N_2731,N_2697);
and U3489 (N_3489,N_2599,N_2625);
nand U3490 (N_3490,N_2745,N_2975);
nor U3491 (N_3491,N_2631,N_2730);
and U3492 (N_3492,N_2829,N_2743);
nand U3493 (N_3493,N_2884,N_2997);
nor U3494 (N_3494,N_2770,N_2671);
nand U3495 (N_3495,N_2933,N_2689);
nor U3496 (N_3496,N_2883,N_2963);
nand U3497 (N_3497,N_2780,N_2702);
xor U3498 (N_3498,N_2642,N_2607);
or U3499 (N_3499,N_2710,N_2802);
or U3500 (N_3500,N_3055,N_3484);
nor U3501 (N_3501,N_3335,N_3401);
and U3502 (N_3502,N_3322,N_3446);
nand U3503 (N_3503,N_3179,N_3278);
and U3504 (N_3504,N_3052,N_3376);
and U3505 (N_3505,N_3234,N_3082);
nand U3506 (N_3506,N_3090,N_3425);
nand U3507 (N_3507,N_3256,N_3309);
or U3508 (N_3508,N_3147,N_3184);
and U3509 (N_3509,N_3222,N_3193);
xnor U3510 (N_3510,N_3451,N_3428);
and U3511 (N_3511,N_3421,N_3315);
nor U3512 (N_3512,N_3163,N_3036);
and U3513 (N_3513,N_3265,N_3028);
and U3514 (N_3514,N_3183,N_3151);
and U3515 (N_3515,N_3244,N_3392);
nor U3516 (N_3516,N_3268,N_3239);
nand U3517 (N_3517,N_3295,N_3248);
nand U3518 (N_3518,N_3060,N_3472);
or U3519 (N_3519,N_3370,N_3250);
or U3520 (N_3520,N_3161,N_3025);
or U3521 (N_3521,N_3020,N_3288);
or U3522 (N_3522,N_3152,N_3470);
or U3523 (N_3523,N_3026,N_3204);
nand U3524 (N_3524,N_3139,N_3226);
nand U3525 (N_3525,N_3479,N_3215);
nand U3526 (N_3526,N_3460,N_3396);
or U3527 (N_3527,N_3402,N_3348);
nand U3528 (N_3528,N_3415,N_3178);
nand U3529 (N_3529,N_3084,N_3488);
or U3530 (N_3530,N_3086,N_3216);
and U3531 (N_3531,N_3398,N_3491);
nand U3532 (N_3532,N_3306,N_3005);
nor U3533 (N_3533,N_3326,N_3010);
nor U3534 (N_3534,N_3349,N_3158);
or U3535 (N_3535,N_3373,N_3499);
or U3536 (N_3536,N_3308,N_3462);
nand U3537 (N_3537,N_3403,N_3124);
and U3538 (N_3538,N_3380,N_3382);
or U3539 (N_3539,N_3375,N_3476);
or U3540 (N_3540,N_3455,N_3471);
nand U3541 (N_3541,N_3467,N_3283);
nor U3542 (N_3542,N_3397,N_3177);
and U3543 (N_3543,N_3317,N_3214);
nor U3544 (N_3544,N_3343,N_3141);
xnor U3545 (N_3545,N_3079,N_3384);
nand U3546 (N_3546,N_3127,N_3280);
nand U3547 (N_3547,N_3182,N_3218);
xor U3548 (N_3548,N_3024,N_3217);
and U3549 (N_3549,N_3063,N_3180);
and U3550 (N_3550,N_3135,N_3138);
nor U3551 (N_3551,N_3071,N_3300);
nor U3552 (N_3552,N_3153,N_3498);
and U3553 (N_3553,N_3112,N_3203);
nor U3554 (N_3554,N_3013,N_3262);
nand U3555 (N_3555,N_3292,N_3378);
nand U3556 (N_3556,N_3047,N_3437);
nor U3557 (N_3557,N_3123,N_3482);
nand U3558 (N_3558,N_3046,N_3496);
and U3559 (N_3559,N_3076,N_3048);
nor U3560 (N_3560,N_3209,N_3230);
xor U3561 (N_3561,N_3088,N_3424);
or U3562 (N_3562,N_3417,N_3128);
or U3563 (N_3563,N_3101,N_3121);
and U3564 (N_3564,N_3253,N_3388);
and U3565 (N_3565,N_3255,N_3031);
and U3566 (N_3566,N_3312,N_3159);
or U3567 (N_3567,N_3438,N_3241);
nor U3568 (N_3568,N_3399,N_3469);
xor U3569 (N_3569,N_3175,N_3225);
and U3570 (N_3570,N_3385,N_3212);
nor U3571 (N_3571,N_3365,N_3087);
nand U3572 (N_3572,N_3347,N_3129);
nor U3573 (N_3573,N_3166,N_3078);
and U3574 (N_3574,N_3196,N_3439);
nand U3575 (N_3575,N_3233,N_3085);
or U3576 (N_3576,N_3468,N_3126);
nor U3577 (N_3577,N_3259,N_3390);
nand U3578 (N_3578,N_3236,N_3346);
and U3579 (N_3579,N_3474,N_3369);
or U3580 (N_3580,N_3423,N_3386);
nor U3581 (N_3581,N_3172,N_3430);
nor U3582 (N_3582,N_3277,N_3334);
nand U3583 (N_3583,N_3420,N_3045);
nand U3584 (N_3584,N_3165,N_3220);
nor U3585 (N_3585,N_3211,N_3477);
nor U3586 (N_3586,N_3068,N_3251);
nand U3587 (N_3587,N_3272,N_3188);
nand U3588 (N_3588,N_3458,N_3395);
or U3589 (N_3589,N_3050,N_3014);
or U3590 (N_3590,N_3174,N_3033);
nor U3591 (N_3591,N_3270,N_3461);
or U3592 (N_3592,N_3206,N_3168);
nand U3593 (N_3593,N_3342,N_3333);
and U3594 (N_3594,N_3302,N_3091);
or U3595 (N_3595,N_3328,N_3007);
nand U3596 (N_3596,N_3387,N_3298);
xor U3597 (N_3597,N_3100,N_3310);
nor U3598 (N_3598,N_3150,N_3249);
xor U3599 (N_3599,N_3064,N_3015);
nand U3600 (N_3600,N_3453,N_3412);
and U3601 (N_3601,N_3246,N_3271);
or U3602 (N_3602,N_3235,N_3017);
nand U3603 (N_3603,N_3113,N_3232);
xnor U3604 (N_3604,N_3266,N_3379);
and U3605 (N_3605,N_3098,N_3116);
nor U3606 (N_3606,N_3441,N_3173);
nand U3607 (N_3607,N_3229,N_3459);
xor U3608 (N_3608,N_3105,N_3301);
nor U3609 (N_3609,N_3314,N_3407);
nand U3610 (N_3610,N_3355,N_3044);
or U3611 (N_3611,N_3311,N_3497);
nor U3612 (N_3612,N_3160,N_3115);
nand U3613 (N_3613,N_3092,N_3006);
or U3614 (N_3614,N_3210,N_3318);
or U3615 (N_3615,N_3016,N_3039);
nor U3616 (N_3616,N_3372,N_3494);
nand U3617 (N_3617,N_3103,N_3035);
xnor U3618 (N_3618,N_3185,N_3449);
and U3619 (N_3619,N_3452,N_3436);
nand U3620 (N_3620,N_3104,N_3029);
or U3621 (N_3621,N_3463,N_3406);
nor U3622 (N_3622,N_3190,N_3287);
nor U3623 (N_3623,N_3022,N_3276);
nor U3624 (N_3624,N_3457,N_3057);
or U3625 (N_3625,N_3197,N_3120);
or U3626 (N_3626,N_3483,N_3238);
nor U3627 (N_3627,N_3356,N_3409);
nand U3628 (N_3628,N_3434,N_3245);
and U3629 (N_3629,N_3359,N_3337);
xor U3630 (N_3630,N_3109,N_3321);
nor U3631 (N_3631,N_3008,N_3073);
nor U3632 (N_3632,N_3202,N_3191);
and U3633 (N_3633,N_3454,N_3426);
nor U3634 (N_3634,N_3187,N_3487);
and U3635 (N_3635,N_3358,N_3074);
or U3636 (N_3636,N_3243,N_3205);
or U3637 (N_3637,N_3081,N_3072);
nand U3638 (N_3638,N_3329,N_3340);
nor U3639 (N_3639,N_3267,N_3341);
nand U3640 (N_3640,N_3289,N_3383);
nor U3641 (N_3641,N_3133,N_3061);
or U3642 (N_3642,N_3040,N_3350);
or U3643 (N_3643,N_3065,N_3227);
and U3644 (N_3644,N_3058,N_3170);
nand U3645 (N_3645,N_3069,N_3381);
or U3646 (N_3646,N_3332,N_3192);
or U3647 (N_3647,N_3374,N_3368);
nand U3648 (N_3648,N_3012,N_3286);
nand U3649 (N_3649,N_3466,N_3201);
or U3650 (N_3650,N_3140,N_3433);
or U3651 (N_3651,N_3075,N_3456);
and U3652 (N_3652,N_3108,N_3228);
nor U3653 (N_3653,N_3319,N_3281);
xnor U3654 (N_3654,N_3207,N_3169);
nor U3655 (N_3655,N_3194,N_3110);
nor U3656 (N_3656,N_3331,N_3320);
or U3657 (N_3657,N_3030,N_3275);
xnor U3658 (N_3658,N_3299,N_3053);
and U3659 (N_3659,N_3070,N_3450);
nor U3660 (N_3660,N_3237,N_3231);
and U3661 (N_3661,N_3221,N_3413);
or U3662 (N_3662,N_3464,N_3264);
and U3663 (N_3663,N_3181,N_3293);
nand U3664 (N_3664,N_3445,N_3431);
nand U3665 (N_3665,N_3478,N_3223);
nor U3666 (N_3666,N_3132,N_3327);
nand U3667 (N_3667,N_3367,N_3200);
nand U3668 (N_3668,N_3167,N_3480);
or U3669 (N_3669,N_3258,N_3297);
and U3670 (N_3670,N_3134,N_3142);
or U3671 (N_3671,N_3486,N_3418);
xnor U3672 (N_3672,N_3473,N_3389);
and U3673 (N_3673,N_3408,N_3186);
or U3674 (N_3674,N_3018,N_3303);
or U3675 (N_3675,N_3224,N_3001);
xnor U3676 (N_3676,N_3465,N_3023);
xnor U3677 (N_3677,N_3213,N_3261);
and U3678 (N_3678,N_3344,N_3049);
xnor U3679 (N_3679,N_3404,N_3419);
nor U3680 (N_3680,N_3489,N_3146);
or U3681 (N_3681,N_3144,N_3037);
and U3682 (N_3682,N_3432,N_3111);
or U3683 (N_3683,N_3162,N_3354);
nand U3684 (N_3684,N_3125,N_3034);
or U3685 (N_3685,N_3492,N_3291);
nor U3686 (N_3686,N_3361,N_3156);
nor U3687 (N_3687,N_3011,N_3493);
and U3688 (N_3688,N_3038,N_3357);
nand U3689 (N_3689,N_3304,N_3323);
or U3690 (N_3690,N_3282,N_3066);
xor U3691 (N_3691,N_3485,N_3360);
or U3692 (N_3692,N_3208,N_3095);
or U3693 (N_3693,N_3416,N_3440);
and U3694 (N_3694,N_3481,N_3447);
or U3695 (N_3695,N_3490,N_3000);
nor U3696 (N_3696,N_3394,N_3003);
and U3697 (N_3697,N_3366,N_3325);
and U3698 (N_3698,N_3393,N_3427);
nor U3699 (N_3699,N_3444,N_3313);
nor U3700 (N_3700,N_3019,N_3257);
nor U3701 (N_3701,N_3102,N_3093);
and U3702 (N_3702,N_3189,N_3099);
nand U3703 (N_3703,N_3269,N_3149);
nor U3704 (N_3704,N_3435,N_3119);
nor U3705 (N_3705,N_3296,N_3279);
nand U3706 (N_3706,N_3154,N_3363);
and U3707 (N_3707,N_3145,N_3391);
and U3708 (N_3708,N_3351,N_3056);
nand U3709 (N_3709,N_3219,N_3274);
nand U3710 (N_3710,N_3032,N_3155);
or U3711 (N_3711,N_3054,N_3106);
nor U3712 (N_3712,N_3254,N_3021);
nand U3713 (N_3713,N_3294,N_3131);
xor U3714 (N_3714,N_3002,N_3353);
and U3715 (N_3715,N_3442,N_3157);
and U3716 (N_3716,N_3284,N_3067);
and U3717 (N_3717,N_3260,N_3004);
xor U3718 (N_3718,N_3118,N_3448);
or U3719 (N_3719,N_3405,N_3352);
nand U3720 (N_3720,N_3475,N_3240);
and U3721 (N_3721,N_3171,N_3117);
nand U3722 (N_3722,N_3330,N_3164);
or U3723 (N_3723,N_3362,N_3495);
nor U3724 (N_3724,N_3137,N_3414);
nand U3725 (N_3725,N_3089,N_3336);
and U3726 (N_3726,N_3042,N_3429);
nand U3727 (N_3727,N_3077,N_3339);
and U3728 (N_3728,N_3094,N_3136);
nand U3729 (N_3729,N_3410,N_3411);
nand U3730 (N_3730,N_3338,N_3148);
nand U3731 (N_3731,N_3080,N_3345);
nor U3732 (N_3732,N_3107,N_3009);
xor U3733 (N_3733,N_3371,N_3059);
nand U3734 (N_3734,N_3324,N_3043);
nor U3735 (N_3735,N_3114,N_3252);
nor U3736 (N_3736,N_3027,N_3051);
or U3737 (N_3737,N_3247,N_3307);
nand U3738 (N_3738,N_3364,N_3062);
xnor U3739 (N_3739,N_3195,N_3176);
nand U3740 (N_3740,N_3316,N_3290);
or U3741 (N_3741,N_3422,N_3130);
and U3742 (N_3742,N_3242,N_3097);
nor U3743 (N_3743,N_3096,N_3199);
or U3744 (N_3744,N_3377,N_3143);
nand U3745 (N_3745,N_3285,N_3305);
nand U3746 (N_3746,N_3083,N_3041);
nor U3747 (N_3747,N_3122,N_3198);
and U3748 (N_3748,N_3443,N_3263);
xor U3749 (N_3749,N_3400,N_3273);
nor U3750 (N_3750,N_3161,N_3386);
and U3751 (N_3751,N_3255,N_3240);
nand U3752 (N_3752,N_3267,N_3128);
or U3753 (N_3753,N_3438,N_3319);
nor U3754 (N_3754,N_3469,N_3314);
or U3755 (N_3755,N_3426,N_3052);
and U3756 (N_3756,N_3389,N_3203);
nand U3757 (N_3757,N_3220,N_3317);
nand U3758 (N_3758,N_3037,N_3122);
nand U3759 (N_3759,N_3130,N_3154);
nor U3760 (N_3760,N_3387,N_3441);
nand U3761 (N_3761,N_3375,N_3278);
nor U3762 (N_3762,N_3000,N_3029);
nand U3763 (N_3763,N_3495,N_3263);
or U3764 (N_3764,N_3080,N_3021);
nor U3765 (N_3765,N_3309,N_3051);
or U3766 (N_3766,N_3202,N_3210);
xor U3767 (N_3767,N_3211,N_3290);
and U3768 (N_3768,N_3190,N_3440);
nor U3769 (N_3769,N_3359,N_3076);
nor U3770 (N_3770,N_3114,N_3282);
and U3771 (N_3771,N_3109,N_3289);
and U3772 (N_3772,N_3100,N_3221);
or U3773 (N_3773,N_3299,N_3361);
nand U3774 (N_3774,N_3178,N_3421);
nand U3775 (N_3775,N_3193,N_3458);
nor U3776 (N_3776,N_3125,N_3362);
or U3777 (N_3777,N_3463,N_3383);
or U3778 (N_3778,N_3307,N_3103);
xor U3779 (N_3779,N_3031,N_3277);
and U3780 (N_3780,N_3162,N_3442);
or U3781 (N_3781,N_3275,N_3336);
or U3782 (N_3782,N_3476,N_3336);
or U3783 (N_3783,N_3069,N_3061);
and U3784 (N_3784,N_3397,N_3278);
or U3785 (N_3785,N_3361,N_3472);
nor U3786 (N_3786,N_3425,N_3442);
and U3787 (N_3787,N_3476,N_3037);
or U3788 (N_3788,N_3389,N_3145);
and U3789 (N_3789,N_3417,N_3069);
nor U3790 (N_3790,N_3418,N_3452);
nand U3791 (N_3791,N_3181,N_3090);
or U3792 (N_3792,N_3295,N_3326);
nand U3793 (N_3793,N_3332,N_3266);
nand U3794 (N_3794,N_3092,N_3085);
or U3795 (N_3795,N_3284,N_3458);
nand U3796 (N_3796,N_3017,N_3477);
xnor U3797 (N_3797,N_3400,N_3393);
nor U3798 (N_3798,N_3262,N_3078);
xnor U3799 (N_3799,N_3138,N_3180);
nand U3800 (N_3800,N_3483,N_3347);
or U3801 (N_3801,N_3300,N_3399);
nand U3802 (N_3802,N_3466,N_3379);
xnor U3803 (N_3803,N_3385,N_3257);
or U3804 (N_3804,N_3105,N_3275);
or U3805 (N_3805,N_3104,N_3030);
and U3806 (N_3806,N_3091,N_3198);
and U3807 (N_3807,N_3060,N_3386);
nor U3808 (N_3808,N_3136,N_3271);
and U3809 (N_3809,N_3290,N_3087);
nand U3810 (N_3810,N_3053,N_3255);
nand U3811 (N_3811,N_3172,N_3105);
nor U3812 (N_3812,N_3235,N_3281);
nand U3813 (N_3813,N_3154,N_3174);
nand U3814 (N_3814,N_3348,N_3171);
nor U3815 (N_3815,N_3394,N_3367);
and U3816 (N_3816,N_3312,N_3199);
and U3817 (N_3817,N_3000,N_3346);
nor U3818 (N_3818,N_3446,N_3139);
nor U3819 (N_3819,N_3323,N_3091);
nor U3820 (N_3820,N_3354,N_3484);
nand U3821 (N_3821,N_3044,N_3354);
nand U3822 (N_3822,N_3212,N_3014);
nand U3823 (N_3823,N_3271,N_3281);
and U3824 (N_3824,N_3236,N_3187);
nand U3825 (N_3825,N_3153,N_3450);
xor U3826 (N_3826,N_3031,N_3434);
nor U3827 (N_3827,N_3459,N_3133);
nand U3828 (N_3828,N_3250,N_3073);
or U3829 (N_3829,N_3460,N_3317);
xnor U3830 (N_3830,N_3265,N_3455);
and U3831 (N_3831,N_3276,N_3351);
or U3832 (N_3832,N_3197,N_3308);
nand U3833 (N_3833,N_3462,N_3052);
xor U3834 (N_3834,N_3089,N_3400);
nor U3835 (N_3835,N_3450,N_3145);
nor U3836 (N_3836,N_3107,N_3121);
or U3837 (N_3837,N_3181,N_3337);
xor U3838 (N_3838,N_3491,N_3337);
and U3839 (N_3839,N_3103,N_3345);
nor U3840 (N_3840,N_3140,N_3160);
or U3841 (N_3841,N_3408,N_3063);
nand U3842 (N_3842,N_3467,N_3439);
nand U3843 (N_3843,N_3322,N_3451);
and U3844 (N_3844,N_3029,N_3201);
or U3845 (N_3845,N_3170,N_3370);
nand U3846 (N_3846,N_3256,N_3333);
nor U3847 (N_3847,N_3367,N_3178);
and U3848 (N_3848,N_3372,N_3161);
nor U3849 (N_3849,N_3371,N_3290);
or U3850 (N_3850,N_3110,N_3393);
nand U3851 (N_3851,N_3261,N_3116);
nor U3852 (N_3852,N_3397,N_3394);
nand U3853 (N_3853,N_3157,N_3109);
or U3854 (N_3854,N_3168,N_3372);
and U3855 (N_3855,N_3091,N_3049);
or U3856 (N_3856,N_3466,N_3343);
or U3857 (N_3857,N_3478,N_3102);
or U3858 (N_3858,N_3460,N_3003);
nor U3859 (N_3859,N_3415,N_3243);
xor U3860 (N_3860,N_3014,N_3395);
and U3861 (N_3861,N_3396,N_3008);
nor U3862 (N_3862,N_3062,N_3253);
and U3863 (N_3863,N_3383,N_3411);
or U3864 (N_3864,N_3418,N_3344);
and U3865 (N_3865,N_3478,N_3093);
or U3866 (N_3866,N_3027,N_3118);
nor U3867 (N_3867,N_3134,N_3123);
and U3868 (N_3868,N_3312,N_3057);
nor U3869 (N_3869,N_3485,N_3008);
and U3870 (N_3870,N_3041,N_3386);
and U3871 (N_3871,N_3156,N_3270);
and U3872 (N_3872,N_3320,N_3001);
or U3873 (N_3873,N_3296,N_3436);
or U3874 (N_3874,N_3445,N_3390);
nor U3875 (N_3875,N_3355,N_3118);
or U3876 (N_3876,N_3056,N_3002);
or U3877 (N_3877,N_3413,N_3169);
nor U3878 (N_3878,N_3348,N_3068);
or U3879 (N_3879,N_3497,N_3459);
or U3880 (N_3880,N_3332,N_3375);
nor U3881 (N_3881,N_3170,N_3399);
and U3882 (N_3882,N_3389,N_3246);
nor U3883 (N_3883,N_3414,N_3189);
or U3884 (N_3884,N_3086,N_3463);
or U3885 (N_3885,N_3471,N_3472);
nand U3886 (N_3886,N_3312,N_3125);
or U3887 (N_3887,N_3033,N_3406);
nand U3888 (N_3888,N_3247,N_3009);
and U3889 (N_3889,N_3016,N_3101);
and U3890 (N_3890,N_3375,N_3044);
nor U3891 (N_3891,N_3108,N_3315);
nor U3892 (N_3892,N_3417,N_3489);
and U3893 (N_3893,N_3462,N_3337);
and U3894 (N_3894,N_3387,N_3360);
or U3895 (N_3895,N_3236,N_3414);
and U3896 (N_3896,N_3201,N_3434);
or U3897 (N_3897,N_3172,N_3243);
nor U3898 (N_3898,N_3403,N_3216);
or U3899 (N_3899,N_3388,N_3196);
nor U3900 (N_3900,N_3379,N_3350);
and U3901 (N_3901,N_3469,N_3042);
nor U3902 (N_3902,N_3292,N_3494);
or U3903 (N_3903,N_3227,N_3027);
and U3904 (N_3904,N_3254,N_3144);
or U3905 (N_3905,N_3113,N_3139);
nand U3906 (N_3906,N_3370,N_3087);
nand U3907 (N_3907,N_3267,N_3069);
and U3908 (N_3908,N_3378,N_3064);
nand U3909 (N_3909,N_3211,N_3402);
and U3910 (N_3910,N_3206,N_3143);
and U3911 (N_3911,N_3166,N_3452);
or U3912 (N_3912,N_3349,N_3332);
nand U3913 (N_3913,N_3096,N_3271);
nand U3914 (N_3914,N_3155,N_3192);
or U3915 (N_3915,N_3453,N_3445);
and U3916 (N_3916,N_3026,N_3264);
or U3917 (N_3917,N_3127,N_3016);
and U3918 (N_3918,N_3458,N_3390);
or U3919 (N_3919,N_3321,N_3418);
or U3920 (N_3920,N_3027,N_3429);
or U3921 (N_3921,N_3060,N_3105);
or U3922 (N_3922,N_3411,N_3009);
nor U3923 (N_3923,N_3194,N_3191);
and U3924 (N_3924,N_3420,N_3430);
nor U3925 (N_3925,N_3043,N_3317);
nor U3926 (N_3926,N_3107,N_3113);
nor U3927 (N_3927,N_3088,N_3120);
or U3928 (N_3928,N_3090,N_3249);
or U3929 (N_3929,N_3364,N_3043);
xnor U3930 (N_3930,N_3009,N_3299);
nor U3931 (N_3931,N_3249,N_3124);
nor U3932 (N_3932,N_3499,N_3498);
xnor U3933 (N_3933,N_3204,N_3318);
and U3934 (N_3934,N_3368,N_3110);
and U3935 (N_3935,N_3026,N_3223);
and U3936 (N_3936,N_3025,N_3313);
and U3937 (N_3937,N_3079,N_3199);
or U3938 (N_3938,N_3109,N_3407);
nor U3939 (N_3939,N_3006,N_3381);
nand U3940 (N_3940,N_3186,N_3303);
nor U3941 (N_3941,N_3327,N_3117);
nor U3942 (N_3942,N_3149,N_3142);
or U3943 (N_3943,N_3451,N_3209);
or U3944 (N_3944,N_3105,N_3057);
nor U3945 (N_3945,N_3347,N_3376);
nor U3946 (N_3946,N_3278,N_3440);
xnor U3947 (N_3947,N_3344,N_3365);
and U3948 (N_3948,N_3007,N_3306);
xor U3949 (N_3949,N_3411,N_3187);
nand U3950 (N_3950,N_3023,N_3408);
or U3951 (N_3951,N_3353,N_3080);
xor U3952 (N_3952,N_3247,N_3005);
nand U3953 (N_3953,N_3040,N_3062);
nand U3954 (N_3954,N_3222,N_3435);
xor U3955 (N_3955,N_3094,N_3145);
or U3956 (N_3956,N_3029,N_3116);
or U3957 (N_3957,N_3454,N_3058);
nor U3958 (N_3958,N_3212,N_3384);
or U3959 (N_3959,N_3224,N_3459);
nand U3960 (N_3960,N_3432,N_3240);
nor U3961 (N_3961,N_3216,N_3225);
nor U3962 (N_3962,N_3494,N_3045);
nor U3963 (N_3963,N_3335,N_3182);
or U3964 (N_3964,N_3245,N_3182);
or U3965 (N_3965,N_3053,N_3265);
xnor U3966 (N_3966,N_3353,N_3395);
nand U3967 (N_3967,N_3493,N_3478);
nor U3968 (N_3968,N_3264,N_3262);
or U3969 (N_3969,N_3494,N_3314);
and U3970 (N_3970,N_3147,N_3425);
xor U3971 (N_3971,N_3321,N_3400);
xnor U3972 (N_3972,N_3460,N_3043);
or U3973 (N_3973,N_3448,N_3338);
and U3974 (N_3974,N_3406,N_3096);
and U3975 (N_3975,N_3441,N_3009);
or U3976 (N_3976,N_3194,N_3125);
or U3977 (N_3977,N_3439,N_3262);
or U3978 (N_3978,N_3113,N_3456);
and U3979 (N_3979,N_3478,N_3182);
nand U3980 (N_3980,N_3403,N_3207);
and U3981 (N_3981,N_3238,N_3418);
and U3982 (N_3982,N_3499,N_3273);
or U3983 (N_3983,N_3362,N_3229);
and U3984 (N_3984,N_3138,N_3208);
nand U3985 (N_3985,N_3205,N_3395);
and U3986 (N_3986,N_3314,N_3184);
nor U3987 (N_3987,N_3438,N_3253);
nor U3988 (N_3988,N_3437,N_3459);
or U3989 (N_3989,N_3337,N_3466);
and U3990 (N_3990,N_3439,N_3254);
nor U3991 (N_3991,N_3143,N_3237);
or U3992 (N_3992,N_3203,N_3108);
nand U3993 (N_3993,N_3394,N_3065);
nor U3994 (N_3994,N_3271,N_3340);
or U3995 (N_3995,N_3257,N_3145);
and U3996 (N_3996,N_3094,N_3352);
and U3997 (N_3997,N_3291,N_3340);
and U3998 (N_3998,N_3281,N_3218);
or U3999 (N_3999,N_3313,N_3022);
and U4000 (N_4000,N_3940,N_3815);
or U4001 (N_4001,N_3694,N_3991);
nor U4002 (N_4002,N_3697,N_3797);
nor U4003 (N_4003,N_3730,N_3700);
nor U4004 (N_4004,N_3541,N_3679);
and U4005 (N_4005,N_3512,N_3959);
and U4006 (N_4006,N_3593,N_3916);
nor U4007 (N_4007,N_3767,N_3814);
nor U4008 (N_4008,N_3937,N_3821);
or U4009 (N_4009,N_3586,N_3880);
or U4010 (N_4010,N_3854,N_3590);
or U4011 (N_4011,N_3985,N_3754);
xor U4012 (N_4012,N_3841,N_3670);
or U4013 (N_4013,N_3933,N_3912);
or U4014 (N_4014,N_3921,N_3832);
or U4015 (N_4015,N_3805,N_3846);
nand U4016 (N_4016,N_3999,N_3974);
xnor U4017 (N_4017,N_3981,N_3594);
nand U4018 (N_4018,N_3717,N_3827);
and U4019 (N_4019,N_3672,N_3877);
and U4020 (N_4020,N_3806,N_3629);
nor U4021 (N_4021,N_3655,N_3547);
xor U4022 (N_4022,N_3711,N_3558);
nor U4023 (N_4023,N_3851,N_3607);
nor U4024 (N_4024,N_3600,N_3637);
and U4025 (N_4025,N_3755,N_3719);
xnor U4026 (N_4026,N_3731,N_3869);
or U4027 (N_4027,N_3964,N_3707);
xnor U4028 (N_4028,N_3968,N_3901);
or U4029 (N_4029,N_3918,N_3534);
nand U4030 (N_4030,N_3750,N_3660);
or U4031 (N_4031,N_3631,N_3524);
or U4032 (N_4032,N_3626,N_3992);
nand U4033 (N_4033,N_3894,N_3885);
and U4034 (N_4034,N_3966,N_3520);
or U4035 (N_4035,N_3501,N_3780);
nor U4036 (N_4036,N_3963,N_3625);
and U4037 (N_4037,N_3828,N_3681);
and U4038 (N_4038,N_3680,N_3721);
or U4039 (N_4039,N_3764,N_3930);
xnor U4040 (N_4040,N_3633,N_3953);
and U4041 (N_4041,N_3561,N_3812);
and U4042 (N_4042,N_3920,N_3613);
nand U4043 (N_4043,N_3733,N_3663);
or U4044 (N_4044,N_3566,N_3636);
nand U4045 (N_4045,N_3888,N_3983);
and U4046 (N_4046,N_3913,N_3500);
or U4047 (N_4047,N_3544,N_3905);
nor U4048 (N_4048,N_3861,N_3917);
nand U4049 (N_4049,N_3824,N_3745);
xnor U4050 (N_4050,N_3927,N_3509);
nor U4051 (N_4051,N_3615,N_3849);
nand U4052 (N_4052,N_3896,N_3659);
nand U4053 (N_4053,N_3870,N_3687);
or U4054 (N_4054,N_3906,N_3708);
nor U4055 (N_4055,N_3645,N_3732);
nand U4056 (N_4056,N_3638,N_3688);
xor U4057 (N_4057,N_3619,N_3528);
or U4058 (N_4058,N_3954,N_3587);
or U4059 (N_4059,N_3602,N_3871);
xor U4060 (N_4060,N_3951,N_3511);
xnor U4061 (N_4061,N_3521,N_3903);
nor U4062 (N_4062,N_3902,N_3542);
or U4063 (N_4063,N_3642,N_3858);
or U4064 (N_4064,N_3654,N_3793);
and U4065 (N_4065,N_3519,N_3575);
xor U4066 (N_4066,N_3839,N_3662);
nor U4067 (N_4067,N_3787,N_3908);
nor U4068 (N_4068,N_3706,N_3976);
and U4069 (N_4069,N_3749,N_3897);
and U4070 (N_4070,N_3924,N_3726);
nor U4071 (N_4071,N_3859,N_3855);
and U4072 (N_4072,N_3523,N_3965);
nor U4073 (N_4073,N_3508,N_3865);
xnor U4074 (N_4074,N_3932,N_3984);
xor U4075 (N_4075,N_3746,N_3843);
nor U4076 (N_4076,N_3955,N_3549);
nor U4077 (N_4077,N_3893,N_3747);
nor U4078 (N_4078,N_3971,N_3866);
or U4079 (N_4079,N_3585,N_3819);
and U4080 (N_4080,N_3786,N_3588);
or U4081 (N_4081,N_3550,N_3958);
and U4082 (N_4082,N_3571,N_3853);
nand U4083 (N_4083,N_3702,N_3518);
nand U4084 (N_4084,N_3979,N_3522);
xnor U4085 (N_4085,N_3591,N_3830);
nor U4086 (N_4086,N_3551,N_3712);
nor U4087 (N_4087,N_3833,N_3624);
nor U4088 (N_4088,N_3683,N_3502);
nor U4089 (N_4089,N_3682,N_3847);
or U4090 (N_4090,N_3825,N_3639);
nor U4091 (N_4091,N_3695,N_3601);
or U4092 (N_4092,N_3796,N_3527);
nand U4093 (N_4093,N_3540,N_3775);
and U4094 (N_4094,N_3704,N_3986);
or U4095 (N_4095,N_3889,N_3898);
or U4096 (N_4096,N_3513,N_3857);
and U4097 (N_4097,N_3989,N_3945);
nor U4098 (N_4098,N_3569,N_3627);
xnor U4099 (N_4099,N_3818,N_3644);
nand U4100 (N_4100,N_3650,N_3729);
or U4101 (N_4101,N_3568,N_3612);
or U4102 (N_4102,N_3635,N_3890);
nor U4103 (N_4103,N_3505,N_3879);
nor U4104 (N_4104,N_3864,N_3781);
nor U4105 (N_4105,N_3884,N_3532);
xor U4106 (N_4106,N_3826,N_3554);
or U4107 (N_4107,N_3752,N_3582);
or U4108 (N_4108,N_3577,N_3943);
and U4109 (N_4109,N_3882,N_3763);
xnor U4110 (N_4110,N_3715,N_3572);
or U4111 (N_4111,N_3993,N_3678);
nor U4112 (N_4112,N_3623,N_3603);
nor U4113 (N_4113,N_3589,N_3507);
nand U4114 (N_4114,N_3962,N_3852);
nand U4115 (N_4115,N_3641,N_3620);
nor U4116 (N_4116,N_3868,N_3768);
nand U4117 (N_4117,N_3649,N_3565);
nand U4118 (N_4118,N_3674,N_3515);
nor U4119 (N_4119,N_3790,N_3929);
or U4120 (N_4120,N_3560,N_3584);
and U4121 (N_4121,N_3709,N_3611);
nor U4122 (N_4122,N_3840,N_3684);
and U4123 (N_4123,N_3808,N_3952);
or U4124 (N_4124,N_3811,N_3967);
xnor U4125 (N_4125,N_3722,N_3530);
xor U4126 (N_4126,N_3608,N_3552);
and U4127 (N_4127,N_3701,N_3794);
nor U4128 (N_4128,N_3673,N_3848);
nor U4129 (N_4129,N_3516,N_3876);
or U4130 (N_4130,N_3664,N_3947);
or U4131 (N_4131,N_3891,N_3758);
or U4132 (N_4132,N_3980,N_3807);
and U4133 (N_4133,N_3961,N_3872);
xor U4134 (N_4134,N_3677,N_3904);
and U4135 (N_4135,N_3616,N_3705);
nor U4136 (N_4136,N_3630,N_3881);
and U4137 (N_4137,N_3783,N_3735);
nor U4138 (N_4138,N_3987,N_3835);
or U4139 (N_4139,N_3765,N_3658);
nand U4140 (N_4140,N_3696,N_3922);
or U4141 (N_4141,N_3784,N_3648);
nor U4142 (N_4142,N_3564,N_3716);
or U4143 (N_4143,N_3666,N_3531);
or U4144 (N_4144,N_3606,N_3751);
and U4145 (N_4145,N_3628,N_3517);
and U4146 (N_4146,N_3718,N_3973);
nand U4147 (N_4147,N_3759,N_3977);
or U4148 (N_4148,N_3647,N_3693);
nand U4149 (N_4149,N_3900,N_3776);
nand U4150 (N_4150,N_3997,N_3838);
and U4151 (N_4151,N_3911,N_3652);
or U4152 (N_4152,N_3567,N_3720);
or U4153 (N_4153,N_3939,N_3526);
and U4154 (N_4154,N_3609,N_3914);
nor U4155 (N_4155,N_3949,N_3873);
nand U4156 (N_4156,N_3771,N_3779);
or U4157 (N_4157,N_3982,N_3632);
nand U4158 (N_4158,N_3621,N_3686);
nor U4159 (N_4159,N_3756,N_3543);
nand U4160 (N_4160,N_3909,N_3867);
nor U4161 (N_4161,N_3948,N_3533);
nand U4162 (N_4162,N_3570,N_3944);
xor U4163 (N_4163,N_3960,N_3777);
xnor U4164 (N_4164,N_3691,N_3850);
or U4165 (N_4165,N_3845,N_3895);
or U4166 (N_4166,N_3975,N_3837);
xor U4167 (N_4167,N_3725,N_3823);
nand U4168 (N_4168,N_3809,N_3676);
and U4169 (N_4169,N_3618,N_3675);
nand U4170 (N_4170,N_3789,N_3559);
and U4171 (N_4171,N_3772,N_3799);
nor U4172 (N_4172,N_3535,N_3723);
or U4173 (N_4173,N_3583,N_3669);
nor U4174 (N_4174,N_3892,N_3978);
nand U4175 (N_4175,N_3785,N_3651);
nor U4176 (N_4176,N_3820,N_3646);
and U4177 (N_4177,N_3605,N_3657);
or U4178 (N_4178,N_3813,N_3698);
nor U4179 (N_4179,N_3555,N_3822);
or U4180 (N_4180,N_3574,N_3801);
or U4181 (N_4181,N_3548,N_3795);
nand U4182 (N_4182,N_3553,N_3856);
and U4183 (N_4183,N_3546,N_3599);
nor U4184 (N_4184,N_3862,N_3580);
nor U4185 (N_4185,N_3692,N_3970);
and U4186 (N_4186,N_3860,N_3685);
nor U4187 (N_4187,N_3998,N_3878);
xnor U4188 (N_4188,N_3802,N_3668);
and U4189 (N_4189,N_3748,N_3539);
nand U4190 (N_4190,N_3934,N_3710);
or U4191 (N_4191,N_3741,N_3757);
nor U4192 (N_4192,N_3875,N_3923);
or U4193 (N_4193,N_3899,N_3703);
xor U4194 (N_4194,N_3689,N_3562);
nor U4195 (N_4195,N_3836,N_3969);
nand U4196 (N_4196,N_3665,N_3537);
nand U4197 (N_4197,N_3592,N_3671);
nand U4198 (N_4198,N_3503,N_3595);
or U4199 (N_4199,N_3931,N_3831);
xnor U4200 (N_4200,N_3738,N_3614);
nand U4201 (N_4201,N_3727,N_3817);
nor U4202 (N_4202,N_3538,N_3690);
xor U4203 (N_4203,N_3778,N_3829);
nand U4204 (N_4204,N_3557,N_3742);
nor U4205 (N_4205,N_3788,N_3950);
nand U4206 (N_4206,N_3842,N_3597);
xnor U4207 (N_4207,N_3640,N_3728);
nor U4208 (N_4208,N_3762,N_3643);
or U4209 (N_4209,N_3529,N_3990);
and U4210 (N_4210,N_3834,N_3816);
xor U4211 (N_4211,N_3510,N_3525);
nor U4212 (N_4212,N_3760,N_3791);
nor U4213 (N_4213,N_3942,N_3804);
nand U4214 (N_4214,N_3744,N_3941);
nor U4215 (N_4215,N_3972,N_3928);
xor U4216 (N_4216,N_3740,N_3886);
nand U4217 (N_4217,N_3946,N_3770);
nand U4218 (N_4218,N_3910,N_3573);
or U4219 (N_4219,N_3504,N_3734);
and U4220 (N_4220,N_3994,N_3536);
nor U4221 (N_4221,N_3844,N_3736);
and U4222 (N_4222,N_3661,N_3610);
xnor U4223 (N_4223,N_3936,N_3935);
xor U4224 (N_4224,N_3761,N_3792);
or U4225 (N_4225,N_3556,N_3667);
nand U4226 (N_4226,N_3737,N_3996);
nor U4227 (N_4227,N_3995,N_3753);
and U4228 (N_4228,N_3925,N_3545);
nor U4229 (N_4229,N_3604,N_3634);
or U4230 (N_4230,N_3810,N_3766);
and U4231 (N_4231,N_3926,N_3798);
nand U4232 (N_4232,N_3938,N_3743);
nor U4233 (N_4233,N_3724,N_3656);
or U4234 (N_4234,N_3578,N_3988);
xnor U4235 (N_4235,N_3907,N_3739);
or U4236 (N_4236,N_3714,N_3622);
nor U4237 (N_4237,N_3769,N_3887);
and U4238 (N_4238,N_3915,N_3803);
nor U4239 (N_4239,N_3800,N_3874);
nor U4240 (N_4240,N_3514,N_3506);
xnor U4241 (N_4241,N_3956,N_3774);
xnor U4242 (N_4242,N_3653,N_3919);
nand U4243 (N_4243,N_3581,N_3596);
nor U4244 (N_4244,N_3699,N_3598);
nand U4245 (N_4245,N_3617,N_3863);
xor U4246 (N_4246,N_3713,N_3957);
or U4247 (N_4247,N_3576,N_3773);
nand U4248 (N_4248,N_3782,N_3883);
or U4249 (N_4249,N_3563,N_3579);
or U4250 (N_4250,N_3763,N_3825);
nand U4251 (N_4251,N_3978,N_3760);
nand U4252 (N_4252,N_3912,N_3892);
nand U4253 (N_4253,N_3877,N_3714);
or U4254 (N_4254,N_3603,N_3946);
xnor U4255 (N_4255,N_3848,N_3719);
nand U4256 (N_4256,N_3799,N_3590);
or U4257 (N_4257,N_3539,N_3552);
and U4258 (N_4258,N_3704,N_3859);
nor U4259 (N_4259,N_3805,N_3610);
or U4260 (N_4260,N_3664,N_3605);
xnor U4261 (N_4261,N_3764,N_3697);
nor U4262 (N_4262,N_3531,N_3808);
and U4263 (N_4263,N_3822,N_3740);
nand U4264 (N_4264,N_3958,N_3815);
nand U4265 (N_4265,N_3991,N_3553);
nor U4266 (N_4266,N_3754,N_3998);
nor U4267 (N_4267,N_3746,N_3649);
and U4268 (N_4268,N_3906,N_3573);
and U4269 (N_4269,N_3892,N_3624);
and U4270 (N_4270,N_3644,N_3522);
or U4271 (N_4271,N_3793,N_3768);
nand U4272 (N_4272,N_3956,N_3912);
and U4273 (N_4273,N_3965,N_3725);
xnor U4274 (N_4274,N_3852,N_3796);
nor U4275 (N_4275,N_3612,N_3753);
and U4276 (N_4276,N_3985,N_3869);
and U4277 (N_4277,N_3901,N_3956);
nor U4278 (N_4278,N_3945,N_3885);
xor U4279 (N_4279,N_3748,N_3830);
and U4280 (N_4280,N_3662,N_3799);
nand U4281 (N_4281,N_3890,N_3885);
and U4282 (N_4282,N_3633,N_3939);
or U4283 (N_4283,N_3931,N_3631);
nand U4284 (N_4284,N_3788,N_3817);
nor U4285 (N_4285,N_3555,N_3838);
xor U4286 (N_4286,N_3686,N_3548);
nor U4287 (N_4287,N_3998,N_3986);
or U4288 (N_4288,N_3899,N_3621);
nor U4289 (N_4289,N_3724,N_3761);
nor U4290 (N_4290,N_3613,N_3896);
nor U4291 (N_4291,N_3660,N_3743);
or U4292 (N_4292,N_3900,N_3697);
or U4293 (N_4293,N_3659,N_3932);
and U4294 (N_4294,N_3853,N_3692);
and U4295 (N_4295,N_3710,N_3947);
or U4296 (N_4296,N_3789,N_3654);
nor U4297 (N_4297,N_3955,N_3651);
nor U4298 (N_4298,N_3595,N_3544);
nand U4299 (N_4299,N_3642,N_3644);
nand U4300 (N_4300,N_3655,N_3773);
nand U4301 (N_4301,N_3765,N_3692);
or U4302 (N_4302,N_3563,N_3524);
and U4303 (N_4303,N_3865,N_3698);
nor U4304 (N_4304,N_3913,N_3634);
or U4305 (N_4305,N_3618,N_3512);
or U4306 (N_4306,N_3904,N_3557);
and U4307 (N_4307,N_3801,N_3697);
and U4308 (N_4308,N_3791,N_3649);
nor U4309 (N_4309,N_3612,N_3779);
and U4310 (N_4310,N_3637,N_3561);
and U4311 (N_4311,N_3862,N_3874);
or U4312 (N_4312,N_3587,N_3965);
nor U4313 (N_4313,N_3790,N_3610);
and U4314 (N_4314,N_3882,N_3931);
xnor U4315 (N_4315,N_3574,N_3876);
and U4316 (N_4316,N_3988,N_3874);
xor U4317 (N_4317,N_3608,N_3996);
xnor U4318 (N_4318,N_3939,N_3693);
nor U4319 (N_4319,N_3719,N_3789);
or U4320 (N_4320,N_3795,N_3973);
or U4321 (N_4321,N_3530,N_3963);
or U4322 (N_4322,N_3707,N_3767);
and U4323 (N_4323,N_3802,N_3530);
xor U4324 (N_4324,N_3591,N_3516);
nor U4325 (N_4325,N_3876,N_3828);
and U4326 (N_4326,N_3938,N_3844);
or U4327 (N_4327,N_3669,N_3803);
nor U4328 (N_4328,N_3688,N_3894);
nor U4329 (N_4329,N_3501,N_3622);
and U4330 (N_4330,N_3767,N_3784);
nor U4331 (N_4331,N_3566,N_3856);
nand U4332 (N_4332,N_3670,N_3847);
nor U4333 (N_4333,N_3579,N_3709);
nor U4334 (N_4334,N_3656,N_3812);
nand U4335 (N_4335,N_3681,N_3852);
or U4336 (N_4336,N_3701,N_3596);
nor U4337 (N_4337,N_3626,N_3690);
or U4338 (N_4338,N_3957,N_3716);
nand U4339 (N_4339,N_3541,N_3672);
nor U4340 (N_4340,N_3890,N_3586);
nor U4341 (N_4341,N_3610,N_3982);
nand U4342 (N_4342,N_3787,N_3547);
xor U4343 (N_4343,N_3698,N_3941);
nand U4344 (N_4344,N_3910,N_3825);
or U4345 (N_4345,N_3597,N_3583);
nand U4346 (N_4346,N_3695,N_3981);
nor U4347 (N_4347,N_3641,N_3963);
xnor U4348 (N_4348,N_3750,N_3788);
nand U4349 (N_4349,N_3541,N_3698);
and U4350 (N_4350,N_3589,N_3827);
nand U4351 (N_4351,N_3901,N_3828);
nor U4352 (N_4352,N_3810,N_3536);
and U4353 (N_4353,N_3562,N_3585);
or U4354 (N_4354,N_3574,N_3645);
nor U4355 (N_4355,N_3750,N_3962);
nand U4356 (N_4356,N_3656,N_3887);
nand U4357 (N_4357,N_3567,N_3773);
nand U4358 (N_4358,N_3994,N_3871);
nor U4359 (N_4359,N_3655,N_3749);
and U4360 (N_4360,N_3988,N_3810);
nand U4361 (N_4361,N_3831,N_3527);
or U4362 (N_4362,N_3539,N_3607);
nor U4363 (N_4363,N_3696,N_3685);
xnor U4364 (N_4364,N_3997,N_3925);
nor U4365 (N_4365,N_3551,N_3510);
and U4366 (N_4366,N_3895,N_3830);
xor U4367 (N_4367,N_3580,N_3835);
and U4368 (N_4368,N_3567,N_3800);
or U4369 (N_4369,N_3770,N_3996);
nor U4370 (N_4370,N_3595,N_3635);
or U4371 (N_4371,N_3727,N_3898);
nor U4372 (N_4372,N_3917,N_3738);
or U4373 (N_4373,N_3812,N_3661);
xnor U4374 (N_4374,N_3852,N_3870);
and U4375 (N_4375,N_3536,N_3665);
nor U4376 (N_4376,N_3883,N_3803);
and U4377 (N_4377,N_3576,N_3612);
xnor U4378 (N_4378,N_3517,N_3534);
nand U4379 (N_4379,N_3512,N_3549);
xor U4380 (N_4380,N_3842,N_3862);
nor U4381 (N_4381,N_3994,N_3537);
and U4382 (N_4382,N_3526,N_3694);
and U4383 (N_4383,N_3542,N_3550);
nor U4384 (N_4384,N_3577,N_3662);
or U4385 (N_4385,N_3538,N_3754);
nor U4386 (N_4386,N_3926,N_3563);
or U4387 (N_4387,N_3685,N_3586);
or U4388 (N_4388,N_3796,N_3873);
or U4389 (N_4389,N_3693,N_3548);
xnor U4390 (N_4390,N_3564,N_3748);
and U4391 (N_4391,N_3717,N_3623);
nand U4392 (N_4392,N_3894,N_3559);
nor U4393 (N_4393,N_3593,N_3686);
nor U4394 (N_4394,N_3923,N_3633);
or U4395 (N_4395,N_3787,N_3565);
or U4396 (N_4396,N_3908,N_3951);
nor U4397 (N_4397,N_3769,N_3513);
or U4398 (N_4398,N_3634,N_3927);
and U4399 (N_4399,N_3980,N_3901);
or U4400 (N_4400,N_3731,N_3515);
nand U4401 (N_4401,N_3558,N_3826);
nor U4402 (N_4402,N_3598,N_3685);
or U4403 (N_4403,N_3762,N_3616);
or U4404 (N_4404,N_3875,N_3917);
and U4405 (N_4405,N_3873,N_3848);
and U4406 (N_4406,N_3659,N_3988);
nand U4407 (N_4407,N_3564,N_3758);
and U4408 (N_4408,N_3803,N_3565);
or U4409 (N_4409,N_3634,N_3759);
and U4410 (N_4410,N_3586,N_3778);
or U4411 (N_4411,N_3965,N_3570);
or U4412 (N_4412,N_3957,N_3998);
xnor U4413 (N_4413,N_3900,N_3711);
and U4414 (N_4414,N_3596,N_3634);
nand U4415 (N_4415,N_3853,N_3846);
nor U4416 (N_4416,N_3922,N_3584);
nor U4417 (N_4417,N_3790,N_3504);
nand U4418 (N_4418,N_3878,N_3782);
and U4419 (N_4419,N_3771,N_3980);
nand U4420 (N_4420,N_3751,N_3921);
nand U4421 (N_4421,N_3514,N_3867);
nand U4422 (N_4422,N_3772,N_3723);
xor U4423 (N_4423,N_3520,N_3885);
nor U4424 (N_4424,N_3912,N_3900);
or U4425 (N_4425,N_3625,N_3662);
and U4426 (N_4426,N_3949,N_3548);
nand U4427 (N_4427,N_3978,N_3821);
or U4428 (N_4428,N_3985,N_3605);
nand U4429 (N_4429,N_3928,N_3910);
nand U4430 (N_4430,N_3620,N_3982);
or U4431 (N_4431,N_3708,N_3623);
nand U4432 (N_4432,N_3532,N_3752);
or U4433 (N_4433,N_3975,N_3643);
nor U4434 (N_4434,N_3901,N_3589);
and U4435 (N_4435,N_3601,N_3986);
nand U4436 (N_4436,N_3891,N_3530);
nor U4437 (N_4437,N_3804,N_3988);
nor U4438 (N_4438,N_3807,N_3542);
or U4439 (N_4439,N_3698,N_3770);
or U4440 (N_4440,N_3613,N_3878);
nor U4441 (N_4441,N_3780,N_3629);
and U4442 (N_4442,N_3677,N_3711);
nor U4443 (N_4443,N_3817,N_3900);
nand U4444 (N_4444,N_3783,N_3838);
xnor U4445 (N_4445,N_3914,N_3896);
or U4446 (N_4446,N_3985,N_3817);
nand U4447 (N_4447,N_3826,N_3697);
or U4448 (N_4448,N_3879,N_3979);
nor U4449 (N_4449,N_3999,N_3852);
or U4450 (N_4450,N_3725,N_3687);
nor U4451 (N_4451,N_3857,N_3535);
or U4452 (N_4452,N_3513,N_3967);
or U4453 (N_4453,N_3617,N_3938);
nor U4454 (N_4454,N_3588,N_3854);
nand U4455 (N_4455,N_3576,N_3667);
nor U4456 (N_4456,N_3940,N_3955);
nand U4457 (N_4457,N_3872,N_3848);
or U4458 (N_4458,N_3538,N_3895);
nor U4459 (N_4459,N_3527,N_3585);
and U4460 (N_4460,N_3636,N_3580);
and U4461 (N_4461,N_3570,N_3726);
and U4462 (N_4462,N_3743,N_3632);
nand U4463 (N_4463,N_3621,N_3901);
nand U4464 (N_4464,N_3628,N_3980);
and U4465 (N_4465,N_3631,N_3663);
nand U4466 (N_4466,N_3748,N_3572);
nand U4467 (N_4467,N_3917,N_3951);
and U4468 (N_4468,N_3855,N_3633);
or U4469 (N_4469,N_3595,N_3722);
and U4470 (N_4470,N_3506,N_3725);
xor U4471 (N_4471,N_3681,N_3996);
or U4472 (N_4472,N_3815,N_3687);
or U4473 (N_4473,N_3841,N_3965);
nand U4474 (N_4474,N_3719,N_3903);
and U4475 (N_4475,N_3557,N_3833);
nor U4476 (N_4476,N_3685,N_3875);
nor U4477 (N_4477,N_3786,N_3848);
and U4478 (N_4478,N_3988,N_3669);
and U4479 (N_4479,N_3944,N_3703);
and U4480 (N_4480,N_3512,N_3761);
or U4481 (N_4481,N_3568,N_3547);
nand U4482 (N_4482,N_3503,N_3942);
and U4483 (N_4483,N_3916,N_3863);
nand U4484 (N_4484,N_3774,N_3699);
or U4485 (N_4485,N_3820,N_3725);
nor U4486 (N_4486,N_3591,N_3957);
and U4487 (N_4487,N_3582,N_3626);
xnor U4488 (N_4488,N_3937,N_3805);
xor U4489 (N_4489,N_3547,N_3700);
nand U4490 (N_4490,N_3580,N_3690);
nor U4491 (N_4491,N_3606,N_3625);
nand U4492 (N_4492,N_3916,N_3691);
and U4493 (N_4493,N_3668,N_3686);
nor U4494 (N_4494,N_3754,N_3977);
xor U4495 (N_4495,N_3647,N_3558);
or U4496 (N_4496,N_3798,N_3766);
or U4497 (N_4497,N_3573,N_3991);
nor U4498 (N_4498,N_3884,N_3825);
xor U4499 (N_4499,N_3696,N_3525);
and U4500 (N_4500,N_4453,N_4189);
or U4501 (N_4501,N_4455,N_4293);
nor U4502 (N_4502,N_4406,N_4324);
nand U4503 (N_4503,N_4031,N_4125);
nor U4504 (N_4504,N_4145,N_4113);
and U4505 (N_4505,N_4090,N_4120);
and U4506 (N_4506,N_4404,N_4191);
nor U4507 (N_4507,N_4354,N_4396);
nor U4508 (N_4508,N_4359,N_4115);
nand U4509 (N_4509,N_4273,N_4248);
nor U4510 (N_4510,N_4195,N_4035);
nor U4511 (N_4511,N_4496,N_4445);
or U4512 (N_4512,N_4152,N_4190);
nand U4513 (N_4513,N_4274,N_4384);
and U4514 (N_4514,N_4425,N_4175);
and U4515 (N_4515,N_4071,N_4499);
nor U4516 (N_4516,N_4114,N_4441);
or U4517 (N_4517,N_4122,N_4421);
or U4518 (N_4518,N_4270,N_4172);
nor U4519 (N_4519,N_4267,N_4200);
nand U4520 (N_4520,N_4217,N_4291);
xnor U4521 (N_4521,N_4146,N_4194);
nand U4522 (N_4522,N_4302,N_4032);
nor U4523 (N_4523,N_4297,N_4084);
nor U4524 (N_4524,N_4424,N_4048);
xor U4525 (N_4525,N_4207,N_4340);
or U4526 (N_4526,N_4362,N_4062);
nor U4527 (N_4527,N_4403,N_4161);
and U4528 (N_4528,N_4014,N_4276);
or U4529 (N_4529,N_4167,N_4299);
nand U4530 (N_4530,N_4454,N_4350);
nand U4531 (N_4531,N_4147,N_4021);
nand U4532 (N_4532,N_4349,N_4236);
nand U4533 (N_4533,N_4108,N_4458);
and U4534 (N_4534,N_4437,N_4215);
nor U4535 (N_4535,N_4080,N_4164);
and U4536 (N_4536,N_4344,N_4402);
and U4537 (N_4537,N_4295,N_4294);
and U4538 (N_4538,N_4156,N_4180);
and U4539 (N_4539,N_4352,N_4104);
xnor U4540 (N_4540,N_4173,N_4305);
or U4541 (N_4541,N_4321,N_4000);
or U4542 (N_4542,N_4472,N_4093);
nand U4543 (N_4543,N_4361,N_4105);
or U4544 (N_4544,N_4205,N_4485);
nand U4545 (N_4545,N_4464,N_4330);
xor U4546 (N_4546,N_4256,N_4002);
or U4547 (N_4547,N_4475,N_4360);
or U4548 (N_4548,N_4422,N_4068);
nand U4549 (N_4549,N_4363,N_4366);
nand U4550 (N_4550,N_4351,N_4466);
xnor U4551 (N_4551,N_4039,N_4202);
and U4552 (N_4552,N_4368,N_4316);
or U4553 (N_4553,N_4058,N_4467);
and U4554 (N_4554,N_4369,N_4420);
or U4555 (N_4555,N_4436,N_4301);
nand U4556 (N_4556,N_4252,N_4017);
and U4557 (N_4557,N_4240,N_4414);
nand U4558 (N_4558,N_4036,N_4280);
and U4559 (N_4559,N_4231,N_4386);
nor U4560 (N_4560,N_4254,N_4086);
nor U4561 (N_4561,N_4281,N_4313);
and U4562 (N_4562,N_4381,N_4199);
or U4563 (N_4563,N_4459,N_4444);
and U4564 (N_4564,N_4133,N_4491);
nor U4565 (N_4565,N_4409,N_4395);
nor U4566 (N_4566,N_4495,N_4337);
nand U4567 (N_4567,N_4006,N_4059);
nor U4568 (N_4568,N_4010,N_4116);
nand U4569 (N_4569,N_4192,N_4348);
or U4570 (N_4570,N_4271,N_4374);
or U4571 (N_4571,N_4498,N_4038);
nand U4572 (N_4572,N_4226,N_4083);
nand U4573 (N_4573,N_4182,N_4245);
and U4574 (N_4574,N_4233,N_4438);
nand U4575 (N_4575,N_4096,N_4155);
nor U4576 (N_4576,N_4132,N_4338);
nor U4577 (N_4577,N_4335,N_4311);
nand U4578 (N_4578,N_4061,N_4244);
nor U4579 (N_4579,N_4442,N_4397);
or U4580 (N_4580,N_4243,N_4110);
nand U4581 (N_4581,N_4051,N_4140);
xnor U4582 (N_4582,N_4377,N_4144);
xnor U4583 (N_4583,N_4450,N_4430);
nand U4584 (N_4584,N_4264,N_4290);
and U4585 (N_4585,N_4181,N_4221);
nor U4586 (N_4586,N_4385,N_4027);
xor U4587 (N_4587,N_4007,N_4228);
or U4588 (N_4588,N_4187,N_4213);
nor U4589 (N_4589,N_4149,N_4004);
or U4590 (N_4590,N_4364,N_4411);
or U4591 (N_4591,N_4435,N_4312);
nand U4592 (N_4592,N_4262,N_4085);
and U4593 (N_4593,N_4001,N_4204);
or U4594 (N_4594,N_4306,N_4206);
nand U4595 (N_4595,N_4428,N_4022);
or U4596 (N_4596,N_4296,N_4148);
nand U4597 (N_4597,N_4426,N_4072);
or U4598 (N_4598,N_4009,N_4353);
and U4599 (N_4599,N_4470,N_4179);
and U4600 (N_4600,N_4123,N_4465);
and U4601 (N_4601,N_4469,N_4484);
nor U4602 (N_4602,N_4432,N_4098);
nor U4603 (N_4603,N_4102,N_4183);
xor U4604 (N_4604,N_4358,N_4355);
nor U4605 (N_4605,N_4033,N_4250);
nand U4606 (N_4606,N_4124,N_4117);
or U4607 (N_4607,N_4052,N_4253);
nor U4608 (N_4608,N_4143,N_4188);
or U4609 (N_4609,N_4166,N_4079);
and U4610 (N_4610,N_4488,N_4480);
nand U4611 (N_4611,N_4493,N_4387);
nand U4612 (N_4612,N_4408,N_4037);
or U4613 (N_4613,N_4412,N_4284);
nand U4614 (N_4614,N_4269,N_4433);
nor U4615 (N_4615,N_4107,N_4429);
nor U4616 (N_4616,N_4456,N_4208);
nor U4617 (N_4617,N_4268,N_4212);
and U4618 (N_4618,N_4081,N_4139);
xnor U4619 (N_4619,N_4497,N_4242);
nand U4620 (N_4620,N_4440,N_4030);
or U4621 (N_4621,N_4092,N_4272);
nand U4622 (N_4622,N_4398,N_4066);
or U4623 (N_4623,N_4091,N_4157);
nor U4624 (N_4624,N_4057,N_4121);
nand U4625 (N_4625,N_4492,N_4103);
xnor U4626 (N_4626,N_4319,N_4288);
or U4627 (N_4627,N_4334,N_4448);
or U4628 (N_4628,N_4201,N_4238);
nand U4629 (N_4629,N_4278,N_4232);
nand U4630 (N_4630,N_4449,N_4023);
xnor U4631 (N_4631,N_4154,N_4044);
and U4632 (N_4632,N_4317,N_4400);
and U4633 (N_4633,N_4060,N_4382);
nor U4634 (N_4634,N_4378,N_4130);
nand U4635 (N_4635,N_4041,N_4249);
or U4636 (N_4636,N_4367,N_4094);
nand U4637 (N_4637,N_4418,N_4451);
and U4638 (N_4638,N_4136,N_4342);
or U4639 (N_4639,N_4169,N_4478);
nor U4640 (N_4640,N_4111,N_4356);
nor U4641 (N_4641,N_4141,N_4246);
xnor U4642 (N_4642,N_4018,N_4118);
nor U4643 (N_4643,N_4261,N_4375);
and U4644 (N_4644,N_4235,N_4119);
or U4645 (N_4645,N_4314,N_4447);
nand U4646 (N_4646,N_4309,N_4285);
xor U4647 (N_4647,N_4223,N_4128);
nor U4648 (N_4648,N_4127,N_4013);
and U4649 (N_4649,N_4069,N_4042);
and U4650 (N_4650,N_4494,N_4176);
nand U4651 (N_4651,N_4347,N_4332);
xor U4652 (N_4652,N_4186,N_4076);
and U4653 (N_4653,N_4135,N_4196);
nand U4654 (N_4654,N_4265,N_4477);
nand U4655 (N_4655,N_4266,N_4315);
and U4656 (N_4656,N_4333,N_4417);
and U4657 (N_4657,N_4327,N_4222);
xnor U4658 (N_4658,N_4399,N_4339);
nor U4659 (N_4659,N_4325,N_4292);
nand U4660 (N_4660,N_4431,N_4286);
or U4661 (N_4661,N_4029,N_4298);
and U4662 (N_4662,N_4461,N_4210);
or U4663 (N_4663,N_4357,N_4024);
nor U4664 (N_4664,N_4322,N_4331);
or U4665 (N_4665,N_4008,N_4198);
nor U4666 (N_4666,N_4405,N_4005);
and U4667 (N_4667,N_4415,N_4345);
or U4668 (N_4668,N_4416,N_4391);
and U4669 (N_4669,N_4075,N_4241);
or U4670 (N_4670,N_4320,N_4336);
and U4671 (N_4671,N_4073,N_4476);
nand U4672 (N_4672,N_4218,N_4452);
nand U4673 (N_4673,N_4462,N_4054);
nor U4674 (N_4674,N_4434,N_4065);
or U4675 (N_4675,N_4043,N_4482);
or U4676 (N_4676,N_4487,N_4251);
xnor U4677 (N_4677,N_4471,N_4479);
nand U4678 (N_4678,N_4063,N_4049);
nor U4679 (N_4679,N_4011,N_4394);
or U4680 (N_4680,N_4277,N_4318);
nand U4681 (N_4681,N_4390,N_4401);
or U4682 (N_4682,N_4056,N_4040);
nand U4683 (N_4683,N_4070,N_4383);
or U4684 (N_4684,N_4279,N_4165);
and U4685 (N_4685,N_4287,N_4372);
nor U4686 (N_4686,N_4388,N_4224);
and U4687 (N_4687,N_4178,N_4260);
or U4688 (N_4688,N_4185,N_4025);
and U4689 (N_4689,N_4087,N_4239);
nor U4690 (N_4690,N_4171,N_4389);
nand U4691 (N_4691,N_4197,N_4304);
and U4692 (N_4692,N_4308,N_4393);
and U4693 (N_4693,N_4275,N_4112);
or U4694 (N_4694,N_4160,N_4392);
and U4695 (N_4695,N_4015,N_4481);
and U4696 (N_4696,N_4234,N_4050);
xnor U4697 (N_4697,N_4126,N_4211);
nand U4698 (N_4698,N_4443,N_4474);
xnor U4699 (N_4699,N_4163,N_4341);
nand U4700 (N_4700,N_4106,N_4323);
and U4701 (N_4701,N_4219,N_4046);
and U4702 (N_4702,N_4078,N_4203);
nor U4703 (N_4703,N_4151,N_4427);
xnor U4704 (N_4704,N_4159,N_4129);
nor U4705 (N_4705,N_4214,N_4174);
nand U4706 (N_4706,N_4486,N_4184);
or U4707 (N_4707,N_4074,N_4019);
and U4708 (N_4708,N_4413,N_4150);
and U4709 (N_4709,N_4067,N_4257);
nand U4710 (N_4710,N_4439,N_4158);
or U4711 (N_4711,N_4101,N_4346);
and U4712 (N_4712,N_4097,N_4225);
or U4713 (N_4713,N_4343,N_4100);
xor U4714 (N_4714,N_4255,N_4258);
nor U4715 (N_4715,N_4373,N_4468);
or U4716 (N_4716,N_4473,N_4170);
and U4717 (N_4717,N_4247,N_4300);
or U4718 (N_4718,N_4282,N_4229);
and U4719 (N_4719,N_4329,N_4283);
or U4720 (N_4720,N_4003,N_4380);
or U4721 (N_4721,N_4016,N_4370);
or U4722 (N_4722,N_4162,N_4303);
xnor U4723 (N_4723,N_4289,N_4483);
or U4724 (N_4724,N_4055,N_4237);
nand U4725 (N_4725,N_4371,N_4379);
nand U4726 (N_4726,N_4307,N_4089);
or U4727 (N_4727,N_4082,N_4168);
or U4728 (N_4728,N_4020,N_4423);
and U4729 (N_4729,N_4142,N_4077);
nand U4730 (N_4730,N_4376,N_4153);
nand U4731 (N_4731,N_4365,N_4220);
or U4732 (N_4732,N_4263,N_4227);
nand U4733 (N_4733,N_4064,N_4034);
or U4734 (N_4734,N_4326,N_4489);
or U4735 (N_4735,N_4137,N_4460);
and U4736 (N_4736,N_4463,N_4310);
or U4737 (N_4737,N_4328,N_4045);
or U4738 (N_4738,N_4088,N_4230);
nor U4739 (N_4739,N_4138,N_4109);
nand U4740 (N_4740,N_4457,N_4134);
and U4741 (N_4741,N_4259,N_4490);
and U4742 (N_4742,N_4446,N_4209);
or U4743 (N_4743,N_4047,N_4131);
nor U4744 (N_4744,N_4012,N_4095);
xor U4745 (N_4745,N_4099,N_4216);
and U4746 (N_4746,N_4028,N_4026);
nor U4747 (N_4747,N_4410,N_4177);
nand U4748 (N_4748,N_4407,N_4193);
or U4749 (N_4749,N_4419,N_4053);
xnor U4750 (N_4750,N_4251,N_4017);
nand U4751 (N_4751,N_4136,N_4126);
and U4752 (N_4752,N_4030,N_4225);
and U4753 (N_4753,N_4403,N_4076);
nand U4754 (N_4754,N_4199,N_4143);
nand U4755 (N_4755,N_4314,N_4290);
or U4756 (N_4756,N_4203,N_4368);
and U4757 (N_4757,N_4327,N_4475);
or U4758 (N_4758,N_4394,N_4433);
xor U4759 (N_4759,N_4100,N_4309);
nand U4760 (N_4760,N_4223,N_4478);
nor U4761 (N_4761,N_4207,N_4282);
nand U4762 (N_4762,N_4414,N_4113);
nand U4763 (N_4763,N_4450,N_4365);
nor U4764 (N_4764,N_4390,N_4477);
nand U4765 (N_4765,N_4315,N_4404);
or U4766 (N_4766,N_4378,N_4335);
nand U4767 (N_4767,N_4103,N_4014);
or U4768 (N_4768,N_4149,N_4155);
nor U4769 (N_4769,N_4326,N_4446);
and U4770 (N_4770,N_4146,N_4226);
nor U4771 (N_4771,N_4485,N_4102);
or U4772 (N_4772,N_4212,N_4062);
or U4773 (N_4773,N_4344,N_4080);
nand U4774 (N_4774,N_4060,N_4339);
nor U4775 (N_4775,N_4105,N_4115);
nor U4776 (N_4776,N_4072,N_4034);
xor U4777 (N_4777,N_4149,N_4475);
or U4778 (N_4778,N_4019,N_4315);
nor U4779 (N_4779,N_4109,N_4180);
or U4780 (N_4780,N_4344,N_4408);
or U4781 (N_4781,N_4363,N_4247);
or U4782 (N_4782,N_4135,N_4177);
nand U4783 (N_4783,N_4291,N_4453);
or U4784 (N_4784,N_4348,N_4060);
nor U4785 (N_4785,N_4240,N_4381);
and U4786 (N_4786,N_4234,N_4486);
or U4787 (N_4787,N_4140,N_4457);
or U4788 (N_4788,N_4147,N_4229);
nor U4789 (N_4789,N_4415,N_4196);
nor U4790 (N_4790,N_4276,N_4043);
nand U4791 (N_4791,N_4215,N_4326);
nand U4792 (N_4792,N_4006,N_4062);
xnor U4793 (N_4793,N_4217,N_4096);
nor U4794 (N_4794,N_4267,N_4353);
and U4795 (N_4795,N_4116,N_4061);
nor U4796 (N_4796,N_4067,N_4182);
or U4797 (N_4797,N_4301,N_4363);
nor U4798 (N_4798,N_4256,N_4429);
nand U4799 (N_4799,N_4294,N_4431);
nor U4800 (N_4800,N_4190,N_4268);
nand U4801 (N_4801,N_4133,N_4407);
nand U4802 (N_4802,N_4383,N_4423);
or U4803 (N_4803,N_4438,N_4404);
and U4804 (N_4804,N_4100,N_4050);
or U4805 (N_4805,N_4167,N_4268);
nor U4806 (N_4806,N_4073,N_4102);
nand U4807 (N_4807,N_4449,N_4303);
nor U4808 (N_4808,N_4051,N_4085);
or U4809 (N_4809,N_4273,N_4166);
or U4810 (N_4810,N_4251,N_4420);
xor U4811 (N_4811,N_4321,N_4448);
nand U4812 (N_4812,N_4365,N_4052);
or U4813 (N_4813,N_4197,N_4157);
xnor U4814 (N_4814,N_4035,N_4471);
and U4815 (N_4815,N_4390,N_4197);
or U4816 (N_4816,N_4008,N_4060);
nand U4817 (N_4817,N_4013,N_4442);
nand U4818 (N_4818,N_4244,N_4088);
or U4819 (N_4819,N_4224,N_4320);
nand U4820 (N_4820,N_4027,N_4486);
nand U4821 (N_4821,N_4326,N_4419);
nand U4822 (N_4822,N_4030,N_4183);
or U4823 (N_4823,N_4118,N_4292);
or U4824 (N_4824,N_4114,N_4242);
xor U4825 (N_4825,N_4379,N_4496);
and U4826 (N_4826,N_4142,N_4130);
and U4827 (N_4827,N_4267,N_4176);
nor U4828 (N_4828,N_4471,N_4316);
or U4829 (N_4829,N_4155,N_4432);
or U4830 (N_4830,N_4393,N_4215);
or U4831 (N_4831,N_4228,N_4387);
nand U4832 (N_4832,N_4461,N_4140);
and U4833 (N_4833,N_4434,N_4476);
and U4834 (N_4834,N_4142,N_4400);
xnor U4835 (N_4835,N_4417,N_4252);
nand U4836 (N_4836,N_4189,N_4454);
or U4837 (N_4837,N_4345,N_4164);
and U4838 (N_4838,N_4366,N_4237);
and U4839 (N_4839,N_4159,N_4327);
and U4840 (N_4840,N_4352,N_4264);
nor U4841 (N_4841,N_4152,N_4002);
nand U4842 (N_4842,N_4074,N_4287);
and U4843 (N_4843,N_4214,N_4432);
or U4844 (N_4844,N_4042,N_4284);
nor U4845 (N_4845,N_4437,N_4289);
or U4846 (N_4846,N_4221,N_4495);
or U4847 (N_4847,N_4060,N_4132);
nor U4848 (N_4848,N_4115,N_4355);
or U4849 (N_4849,N_4118,N_4016);
nor U4850 (N_4850,N_4112,N_4264);
nor U4851 (N_4851,N_4493,N_4087);
nand U4852 (N_4852,N_4097,N_4149);
and U4853 (N_4853,N_4160,N_4147);
or U4854 (N_4854,N_4121,N_4289);
and U4855 (N_4855,N_4124,N_4055);
nand U4856 (N_4856,N_4243,N_4435);
nand U4857 (N_4857,N_4489,N_4298);
or U4858 (N_4858,N_4281,N_4176);
xor U4859 (N_4859,N_4304,N_4440);
or U4860 (N_4860,N_4220,N_4444);
nor U4861 (N_4861,N_4376,N_4367);
or U4862 (N_4862,N_4000,N_4345);
nor U4863 (N_4863,N_4289,N_4120);
xor U4864 (N_4864,N_4382,N_4234);
nor U4865 (N_4865,N_4023,N_4097);
xnor U4866 (N_4866,N_4306,N_4377);
or U4867 (N_4867,N_4130,N_4031);
nor U4868 (N_4868,N_4334,N_4470);
or U4869 (N_4869,N_4118,N_4080);
xor U4870 (N_4870,N_4243,N_4384);
nand U4871 (N_4871,N_4241,N_4400);
nor U4872 (N_4872,N_4313,N_4046);
nor U4873 (N_4873,N_4336,N_4492);
or U4874 (N_4874,N_4069,N_4167);
nor U4875 (N_4875,N_4464,N_4352);
nand U4876 (N_4876,N_4204,N_4254);
nor U4877 (N_4877,N_4157,N_4438);
nand U4878 (N_4878,N_4450,N_4273);
and U4879 (N_4879,N_4377,N_4198);
xor U4880 (N_4880,N_4490,N_4002);
xnor U4881 (N_4881,N_4243,N_4128);
nor U4882 (N_4882,N_4067,N_4005);
nor U4883 (N_4883,N_4342,N_4484);
nand U4884 (N_4884,N_4261,N_4071);
and U4885 (N_4885,N_4158,N_4071);
nor U4886 (N_4886,N_4075,N_4126);
nand U4887 (N_4887,N_4101,N_4015);
nand U4888 (N_4888,N_4314,N_4037);
and U4889 (N_4889,N_4320,N_4425);
or U4890 (N_4890,N_4043,N_4300);
nand U4891 (N_4891,N_4042,N_4324);
or U4892 (N_4892,N_4140,N_4258);
and U4893 (N_4893,N_4003,N_4335);
nand U4894 (N_4894,N_4122,N_4275);
and U4895 (N_4895,N_4041,N_4102);
xnor U4896 (N_4896,N_4496,N_4395);
or U4897 (N_4897,N_4193,N_4033);
nor U4898 (N_4898,N_4225,N_4178);
xor U4899 (N_4899,N_4356,N_4183);
nand U4900 (N_4900,N_4254,N_4082);
nand U4901 (N_4901,N_4455,N_4274);
or U4902 (N_4902,N_4219,N_4359);
nand U4903 (N_4903,N_4170,N_4221);
xor U4904 (N_4904,N_4415,N_4168);
or U4905 (N_4905,N_4021,N_4249);
nor U4906 (N_4906,N_4394,N_4266);
nand U4907 (N_4907,N_4372,N_4461);
nand U4908 (N_4908,N_4454,N_4476);
and U4909 (N_4909,N_4294,N_4414);
or U4910 (N_4910,N_4096,N_4039);
nor U4911 (N_4911,N_4353,N_4438);
nor U4912 (N_4912,N_4173,N_4111);
xnor U4913 (N_4913,N_4309,N_4001);
nor U4914 (N_4914,N_4220,N_4142);
nor U4915 (N_4915,N_4344,N_4353);
nand U4916 (N_4916,N_4234,N_4287);
or U4917 (N_4917,N_4141,N_4168);
or U4918 (N_4918,N_4250,N_4358);
and U4919 (N_4919,N_4314,N_4179);
nand U4920 (N_4920,N_4340,N_4396);
nand U4921 (N_4921,N_4348,N_4314);
and U4922 (N_4922,N_4499,N_4013);
or U4923 (N_4923,N_4414,N_4084);
nor U4924 (N_4924,N_4115,N_4112);
nand U4925 (N_4925,N_4456,N_4369);
and U4926 (N_4926,N_4227,N_4116);
nor U4927 (N_4927,N_4001,N_4141);
and U4928 (N_4928,N_4225,N_4057);
nand U4929 (N_4929,N_4290,N_4270);
and U4930 (N_4930,N_4306,N_4115);
nand U4931 (N_4931,N_4003,N_4497);
and U4932 (N_4932,N_4279,N_4340);
or U4933 (N_4933,N_4429,N_4315);
and U4934 (N_4934,N_4455,N_4087);
and U4935 (N_4935,N_4244,N_4361);
xor U4936 (N_4936,N_4287,N_4240);
xnor U4937 (N_4937,N_4321,N_4385);
or U4938 (N_4938,N_4332,N_4260);
nand U4939 (N_4939,N_4334,N_4093);
nor U4940 (N_4940,N_4186,N_4485);
nor U4941 (N_4941,N_4213,N_4291);
nand U4942 (N_4942,N_4234,N_4110);
or U4943 (N_4943,N_4437,N_4001);
nor U4944 (N_4944,N_4027,N_4049);
and U4945 (N_4945,N_4423,N_4062);
and U4946 (N_4946,N_4075,N_4490);
nand U4947 (N_4947,N_4306,N_4447);
nand U4948 (N_4948,N_4038,N_4141);
or U4949 (N_4949,N_4305,N_4315);
or U4950 (N_4950,N_4191,N_4122);
nor U4951 (N_4951,N_4223,N_4459);
or U4952 (N_4952,N_4001,N_4025);
or U4953 (N_4953,N_4095,N_4017);
or U4954 (N_4954,N_4433,N_4348);
or U4955 (N_4955,N_4040,N_4253);
xnor U4956 (N_4956,N_4400,N_4233);
nor U4957 (N_4957,N_4269,N_4196);
and U4958 (N_4958,N_4421,N_4351);
nor U4959 (N_4959,N_4497,N_4276);
nor U4960 (N_4960,N_4183,N_4347);
or U4961 (N_4961,N_4297,N_4003);
or U4962 (N_4962,N_4254,N_4250);
xnor U4963 (N_4963,N_4471,N_4476);
or U4964 (N_4964,N_4360,N_4263);
or U4965 (N_4965,N_4405,N_4354);
nand U4966 (N_4966,N_4402,N_4165);
or U4967 (N_4967,N_4312,N_4377);
xor U4968 (N_4968,N_4298,N_4200);
and U4969 (N_4969,N_4102,N_4454);
or U4970 (N_4970,N_4149,N_4062);
nand U4971 (N_4971,N_4258,N_4198);
and U4972 (N_4972,N_4363,N_4308);
xor U4973 (N_4973,N_4074,N_4080);
xor U4974 (N_4974,N_4396,N_4473);
or U4975 (N_4975,N_4294,N_4119);
and U4976 (N_4976,N_4177,N_4133);
or U4977 (N_4977,N_4053,N_4486);
or U4978 (N_4978,N_4389,N_4367);
nor U4979 (N_4979,N_4198,N_4461);
or U4980 (N_4980,N_4272,N_4476);
and U4981 (N_4981,N_4143,N_4043);
and U4982 (N_4982,N_4258,N_4191);
nor U4983 (N_4983,N_4253,N_4443);
nand U4984 (N_4984,N_4362,N_4466);
nor U4985 (N_4985,N_4394,N_4478);
and U4986 (N_4986,N_4240,N_4382);
or U4987 (N_4987,N_4253,N_4269);
nor U4988 (N_4988,N_4397,N_4055);
nor U4989 (N_4989,N_4451,N_4008);
nor U4990 (N_4990,N_4224,N_4070);
nand U4991 (N_4991,N_4085,N_4420);
nor U4992 (N_4992,N_4267,N_4455);
nand U4993 (N_4993,N_4149,N_4268);
or U4994 (N_4994,N_4402,N_4202);
nand U4995 (N_4995,N_4131,N_4388);
nand U4996 (N_4996,N_4485,N_4328);
or U4997 (N_4997,N_4320,N_4388);
or U4998 (N_4998,N_4050,N_4035);
nand U4999 (N_4999,N_4154,N_4324);
nor UO_0 (O_0,N_4776,N_4519);
nand UO_1 (O_1,N_4678,N_4758);
or UO_2 (O_2,N_4906,N_4989);
xor UO_3 (O_3,N_4879,N_4871);
nor UO_4 (O_4,N_4817,N_4825);
nor UO_5 (O_5,N_4530,N_4539);
nand UO_6 (O_6,N_4861,N_4522);
and UO_7 (O_7,N_4851,N_4595);
or UO_8 (O_8,N_4729,N_4752);
nor UO_9 (O_9,N_4762,N_4669);
or UO_10 (O_10,N_4596,N_4676);
nor UO_11 (O_11,N_4800,N_4746);
nand UO_12 (O_12,N_4505,N_4860);
or UO_13 (O_13,N_4532,N_4659);
or UO_14 (O_14,N_4545,N_4883);
and UO_15 (O_15,N_4690,N_4699);
or UO_16 (O_16,N_4930,N_4534);
nand UO_17 (O_17,N_4938,N_4587);
and UO_18 (O_18,N_4740,N_4797);
and UO_19 (O_19,N_4869,N_4943);
nor UO_20 (O_20,N_4865,N_4891);
nand UO_21 (O_21,N_4858,N_4567);
or UO_22 (O_22,N_4759,N_4514);
nand UO_23 (O_23,N_4820,N_4512);
nor UO_24 (O_24,N_4633,N_4630);
or UO_25 (O_25,N_4753,N_4908);
xor UO_26 (O_26,N_4953,N_4834);
nand UO_27 (O_27,N_4626,N_4772);
nand UO_28 (O_28,N_4742,N_4824);
or UO_29 (O_29,N_4896,N_4809);
nor UO_30 (O_30,N_4830,N_4510);
or UO_31 (O_31,N_4836,N_4538);
nor UO_32 (O_32,N_4582,N_4981);
nand UO_33 (O_33,N_4638,N_4639);
or UO_34 (O_34,N_4875,N_4673);
or UO_35 (O_35,N_4917,N_4700);
or UO_36 (O_36,N_4620,N_4501);
or UO_37 (O_37,N_4507,N_4806);
and UO_38 (O_38,N_4611,N_4573);
nor UO_39 (O_39,N_4666,N_4764);
and UO_40 (O_40,N_4947,N_4798);
nor UO_41 (O_41,N_4625,N_4963);
nor UO_42 (O_42,N_4617,N_4980);
and UO_43 (O_43,N_4572,N_4781);
or UO_44 (O_44,N_4999,N_4614);
nor UO_45 (O_45,N_4502,N_4855);
and UO_46 (O_46,N_4914,N_4763);
xnor UO_47 (O_47,N_4897,N_4744);
or UO_48 (O_48,N_4523,N_4535);
or UO_49 (O_49,N_4844,N_4782);
nor UO_50 (O_50,N_4585,N_4702);
and UO_51 (O_51,N_4656,N_4928);
xor UO_52 (O_52,N_4819,N_4863);
nand UO_53 (O_53,N_4648,N_4542);
or UO_54 (O_54,N_4951,N_4878);
or UO_55 (O_55,N_4650,N_4706);
and UO_56 (O_56,N_4504,N_4885);
nor UO_57 (O_57,N_4707,N_4672);
xnor UO_58 (O_58,N_4708,N_4827);
nor UO_59 (O_59,N_4992,N_4795);
xor UO_60 (O_60,N_4870,N_4894);
nand UO_61 (O_61,N_4619,N_4660);
and UO_62 (O_62,N_4559,N_4662);
or UO_63 (O_63,N_4727,N_4900);
or UO_64 (O_64,N_4605,N_4886);
nor UO_65 (O_65,N_4540,N_4622);
nor UO_66 (O_66,N_4590,N_4760);
nor UO_67 (O_67,N_4598,N_4747);
nor UO_68 (O_68,N_4786,N_4592);
and UO_69 (O_69,N_4826,N_4730);
and UO_70 (O_70,N_4718,N_4985);
or UO_71 (O_71,N_4548,N_4899);
xnor UO_72 (O_72,N_4687,N_4960);
or UO_73 (O_73,N_4848,N_4681);
or UO_74 (O_74,N_4881,N_4667);
or UO_75 (O_75,N_4518,N_4516);
and UO_76 (O_76,N_4839,N_4868);
nor UO_77 (O_77,N_4832,N_4815);
nand UO_78 (O_78,N_4964,N_4962);
and UO_79 (O_79,N_4558,N_4631);
or UO_80 (O_80,N_4779,N_4884);
nor UO_81 (O_81,N_4850,N_4997);
or UO_82 (O_82,N_4805,N_4922);
nand UO_83 (O_83,N_4921,N_4998);
or UO_84 (O_84,N_4768,N_4649);
nor UO_85 (O_85,N_4647,N_4841);
nand UO_86 (O_86,N_4682,N_4694);
and UO_87 (O_87,N_4551,N_4643);
and UO_88 (O_88,N_4887,N_4932);
and UO_89 (O_89,N_4529,N_4688);
nor UO_90 (O_90,N_4578,N_4679);
nand UO_91 (O_91,N_4916,N_4720);
and UO_92 (O_92,N_4701,N_4791);
and UO_93 (O_93,N_4948,N_4618);
nor UO_94 (O_94,N_4968,N_4586);
or UO_95 (O_95,N_4623,N_4569);
and UO_96 (O_96,N_4577,N_4628);
nor UO_97 (O_97,N_4712,N_4565);
nor UO_98 (O_98,N_4793,N_4944);
or UO_99 (O_99,N_4789,N_4893);
nor UO_100 (O_100,N_4831,N_4517);
xnor UO_101 (O_101,N_4500,N_4949);
or UO_102 (O_102,N_4554,N_4895);
or UO_103 (O_103,N_4515,N_4695);
nand UO_104 (O_104,N_4696,N_4550);
or UO_105 (O_105,N_4710,N_4993);
or UO_106 (O_106,N_4571,N_4579);
nor UO_107 (O_107,N_4835,N_4840);
nor UO_108 (O_108,N_4693,N_4645);
nor UO_109 (O_109,N_4597,N_4686);
nand UO_110 (O_110,N_4683,N_4866);
nor UO_111 (O_111,N_4864,N_4801);
nor UO_112 (O_112,N_4988,N_4777);
nand UO_113 (O_113,N_4608,N_4799);
nor UO_114 (O_114,N_4580,N_4979);
or UO_115 (O_115,N_4602,N_4506);
xnor UO_116 (O_116,N_4684,N_4549);
or UO_117 (O_117,N_4913,N_4967);
nor UO_118 (O_118,N_4823,N_4936);
or UO_119 (O_119,N_4588,N_4765);
nand UO_120 (O_120,N_4721,N_4561);
and UO_121 (O_121,N_4990,N_4942);
and UO_122 (O_122,N_4796,N_4788);
and UO_123 (O_123,N_4837,N_4509);
nor UO_124 (O_124,N_4632,N_4775);
nand UO_125 (O_125,N_4594,N_4874);
nor UO_126 (O_126,N_4748,N_4911);
nor UO_127 (O_127,N_4735,N_4905);
nor UO_128 (O_128,N_4902,N_4526);
or UO_129 (O_129,N_4803,N_4739);
and UO_130 (O_130,N_4954,N_4600);
nor UO_131 (O_131,N_4593,N_4521);
nor UO_132 (O_132,N_4959,N_4876);
nand UO_133 (O_133,N_4636,N_4661);
and UO_134 (O_134,N_4889,N_4603);
or UO_135 (O_135,N_4845,N_4704);
or UO_136 (O_136,N_4670,N_4890);
xor UO_137 (O_137,N_4641,N_4555);
or UO_138 (O_138,N_4698,N_4969);
nand UO_139 (O_139,N_4674,N_4527);
or UO_140 (O_140,N_4543,N_4970);
and UO_141 (O_141,N_4652,N_4725);
xnor UO_142 (O_142,N_4520,N_4931);
nand UO_143 (O_143,N_4918,N_4552);
xor UO_144 (O_144,N_4562,N_4536);
and UO_145 (O_145,N_4734,N_4640);
or UO_146 (O_146,N_4731,N_4945);
and UO_147 (O_147,N_4615,N_4713);
nor UO_148 (O_148,N_4978,N_4783);
xor UO_149 (O_149,N_4743,N_4958);
nand UO_150 (O_150,N_4961,N_4898);
and UO_151 (O_151,N_4787,N_4852);
nor UO_152 (O_152,N_4723,N_4508);
nor UO_153 (O_153,N_4737,N_4750);
and UO_154 (O_154,N_4637,N_4880);
nand UO_155 (O_155,N_4877,N_4941);
and UO_156 (O_156,N_4816,N_4675);
or UO_157 (O_157,N_4654,N_4849);
and UO_158 (O_158,N_4655,N_4745);
or UO_159 (O_159,N_4599,N_4726);
nand UO_160 (O_160,N_4564,N_4829);
xnor UO_161 (O_161,N_4584,N_4991);
and UO_162 (O_162,N_4818,N_4946);
or UO_163 (O_163,N_4856,N_4925);
nand UO_164 (O_164,N_4955,N_4872);
and UO_165 (O_165,N_4644,N_4929);
and UO_166 (O_166,N_4717,N_4581);
and UO_167 (O_167,N_4814,N_4755);
or UO_168 (O_168,N_4901,N_4663);
or UO_169 (O_169,N_4665,N_4972);
nand UO_170 (O_170,N_4923,N_4627);
nand UO_171 (O_171,N_4533,N_4570);
and UO_172 (O_172,N_4774,N_4910);
nor UO_173 (O_173,N_4790,N_4807);
nor UO_174 (O_174,N_4859,N_4828);
and UO_175 (O_175,N_4525,N_4811);
nor UO_176 (O_176,N_4996,N_4904);
nor UO_177 (O_177,N_4761,N_4987);
nor UO_178 (O_178,N_4915,N_4591);
and UO_179 (O_179,N_4767,N_4892);
nand UO_180 (O_180,N_4566,N_4738);
nor UO_181 (O_181,N_4715,N_4935);
or UO_182 (O_182,N_4984,N_4741);
nor UO_183 (O_183,N_4813,N_4537);
and UO_184 (O_184,N_4503,N_4616);
and UO_185 (O_185,N_4986,N_4808);
nand UO_186 (O_186,N_4927,N_4719);
and UO_187 (O_187,N_4965,N_4524);
nor UO_188 (O_188,N_4784,N_4589);
nand UO_189 (O_189,N_4604,N_4771);
nor UO_190 (O_190,N_4976,N_4711);
xnor UO_191 (O_191,N_4677,N_4853);
or UO_192 (O_192,N_4933,N_4629);
nor UO_193 (O_193,N_4940,N_4822);
or UO_194 (O_194,N_4671,N_4642);
or UO_195 (O_195,N_4692,N_4653);
nand UO_196 (O_196,N_4934,N_4691);
and UO_197 (O_197,N_4714,N_4724);
xnor UO_198 (O_198,N_4689,N_4709);
nor UO_199 (O_199,N_4556,N_4977);
and UO_200 (O_200,N_4624,N_4780);
or UO_201 (O_201,N_4802,N_4854);
nor UO_202 (O_202,N_4994,N_4664);
nand UO_203 (O_203,N_4651,N_4847);
nand UO_204 (O_204,N_4557,N_4939);
or UO_205 (O_205,N_4975,N_4956);
nor UO_206 (O_206,N_4574,N_4792);
nand UO_207 (O_207,N_4751,N_4754);
nor UO_208 (O_208,N_4912,N_4513);
nor UO_209 (O_209,N_4685,N_4544);
xor UO_210 (O_210,N_4563,N_4560);
nor UO_211 (O_211,N_4924,N_4888);
xnor UO_212 (O_212,N_4606,N_4546);
or UO_213 (O_213,N_4804,N_4680);
nor UO_214 (O_214,N_4612,N_4733);
nor UO_215 (O_215,N_4757,N_4531);
nor UO_216 (O_216,N_4974,N_4635);
or UO_217 (O_217,N_4995,N_4770);
nor UO_218 (O_218,N_4576,N_4722);
or UO_219 (O_219,N_4541,N_4610);
or UO_220 (O_220,N_4634,N_4862);
nor UO_221 (O_221,N_4736,N_4842);
and UO_222 (O_222,N_4846,N_4821);
and UO_223 (O_223,N_4838,N_4971);
nand UO_224 (O_224,N_4833,N_4926);
xor UO_225 (O_225,N_4607,N_4950);
nand UO_226 (O_226,N_4657,N_4903);
and UO_227 (O_227,N_4873,N_4547);
xnor UO_228 (O_228,N_4810,N_4812);
nand UO_229 (O_229,N_4716,N_4857);
nand UO_230 (O_230,N_4646,N_4983);
and UO_231 (O_231,N_4583,N_4528);
xor UO_232 (O_232,N_4785,N_4957);
and UO_233 (O_233,N_4601,N_4778);
or UO_234 (O_234,N_4756,N_4511);
nor UO_235 (O_235,N_4794,N_4920);
xnor UO_236 (O_236,N_4705,N_4697);
nor UO_237 (O_237,N_4867,N_4749);
and UO_238 (O_238,N_4773,N_4728);
or UO_239 (O_239,N_4703,N_4553);
nand UO_240 (O_240,N_4613,N_4973);
nor UO_241 (O_241,N_4658,N_4621);
or UO_242 (O_242,N_4732,N_4966);
or UO_243 (O_243,N_4882,N_4668);
and UO_244 (O_244,N_4909,N_4843);
and UO_245 (O_245,N_4766,N_4769);
nand UO_246 (O_246,N_4907,N_4919);
or UO_247 (O_247,N_4575,N_4982);
and UO_248 (O_248,N_4952,N_4609);
nand UO_249 (O_249,N_4937,N_4568);
or UO_250 (O_250,N_4863,N_4798);
nand UO_251 (O_251,N_4833,N_4592);
or UO_252 (O_252,N_4619,N_4578);
and UO_253 (O_253,N_4614,N_4585);
nor UO_254 (O_254,N_4701,N_4694);
nor UO_255 (O_255,N_4611,N_4774);
or UO_256 (O_256,N_4804,N_4822);
or UO_257 (O_257,N_4650,N_4699);
and UO_258 (O_258,N_4728,N_4733);
nor UO_259 (O_259,N_4510,N_4719);
nor UO_260 (O_260,N_4950,N_4710);
nor UO_261 (O_261,N_4518,N_4908);
nor UO_262 (O_262,N_4885,N_4688);
nand UO_263 (O_263,N_4517,N_4798);
nand UO_264 (O_264,N_4590,N_4680);
nor UO_265 (O_265,N_4821,N_4984);
nor UO_266 (O_266,N_4730,N_4620);
and UO_267 (O_267,N_4686,N_4973);
xor UO_268 (O_268,N_4790,N_4996);
nor UO_269 (O_269,N_4624,N_4949);
nor UO_270 (O_270,N_4768,N_4765);
xor UO_271 (O_271,N_4938,N_4941);
nor UO_272 (O_272,N_4808,N_4616);
and UO_273 (O_273,N_4837,N_4954);
and UO_274 (O_274,N_4696,N_4673);
nand UO_275 (O_275,N_4509,N_4566);
or UO_276 (O_276,N_4651,N_4795);
nor UO_277 (O_277,N_4655,N_4803);
and UO_278 (O_278,N_4787,N_4539);
and UO_279 (O_279,N_4771,N_4908);
or UO_280 (O_280,N_4845,N_4916);
and UO_281 (O_281,N_4647,N_4531);
nand UO_282 (O_282,N_4820,N_4904);
nand UO_283 (O_283,N_4650,N_4545);
nand UO_284 (O_284,N_4942,N_4653);
or UO_285 (O_285,N_4606,N_4720);
nor UO_286 (O_286,N_4990,N_4685);
or UO_287 (O_287,N_4533,N_4676);
nor UO_288 (O_288,N_4645,N_4547);
nor UO_289 (O_289,N_4677,N_4874);
or UO_290 (O_290,N_4648,N_4697);
and UO_291 (O_291,N_4964,N_4963);
xnor UO_292 (O_292,N_4943,N_4636);
nor UO_293 (O_293,N_4525,N_4535);
nand UO_294 (O_294,N_4795,N_4550);
and UO_295 (O_295,N_4818,N_4964);
nand UO_296 (O_296,N_4581,N_4975);
nor UO_297 (O_297,N_4773,N_4926);
and UO_298 (O_298,N_4610,N_4630);
nor UO_299 (O_299,N_4841,N_4750);
or UO_300 (O_300,N_4554,N_4670);
and UO_301 (O_301,N_4928,N_4590);
or UO_302 (O_302,N_4541,N_4509);
nand UO_303 (O_303,N_4728,N_4717);
xnor UO_304 (O_304,N_4607,N_4849);
and UO_305 (O_305,N_4760,N_4645);
nand UO_306 (O_306,N_4891,N_4826);
nand UO_307 (O_307,N_4721,N_4621);
and UO_308 (O_308,N_4566,N_4514);
nor UO_309 (O_309,N_4595,N_4932);
and UO_310 (O_310,N_4830,N_4525);
or UO_311 (O_311,N_4954,N_4613);
and UO_312 (O_312,N_4661,N_4813);
or UO_313 (O_313,N_4878,N_4901);
and UO_314 (O_314,N_4854,N_4660);
and UO_315 (O_315,N_4512,N_4708);
and UO_316 (O_316,N_4586,N_4746);
and UO_317 (O_317,N_4567,N_4675);
nor UO_318 (O_318,N_4895,N_4516);
nand UO_319 (O_319,N_4535,N_4585);
and UO_320 (O_320,N_4598,N_4982);
nand UO_321 (O_321,N_4537,N_4543);
or UO_322 (O_322,N_4644,N_4554);
or UO_323 (O_323,N_4570,N_4594);
and UO_324 (O_324,N_4846,N_4737);
nor UO_325 (O_325,N_4691,N_4948);
xor UO_326 (O_326,N_4805,N_4958);
or UO_327 (O_327,N_4587,N_4656);
and UO_328 (O_328,N_4980,N_4673);
nand UO_329 (O_329,N_4512,N_4594);
or UO_330 (O_330,N_4866,N_4979);
nand UO_331 (O_331,N_4975,N_4709);
and UO_332 (O_332,N_4984,N_4698);
nand UO_333 (O_333,N_4978,N_4713);
and UO_334 (O_334,N_4950,N_4861);
nand UO_335 (O_335,N_4982,N_4757);
nand UO_336 (O_336,N_4821,N_4530);
or UO_337 (O_337,N_4882,N_4552);
and UO_338 (O_338,N_4564,N_4907);
nand UO_339 (O_339,N_4682,N_4837);
or UO_340 (O_340,N_4615,N_4546);
and UO_341 (O_341,N_4603,N_4633);
nor UO_342 (O_342,N_4912,N_4713);
or UO_343 (O_343,N_4692,N_4900);
nand UO_344 (O_344,N_4895,N_4540);
nor UO_345 (O_345,N_4552,N_4755);
or UO_346 (O_346,N_4780,N_4815);
and UO_347 (O_347,N_4690,N_4985);
nand UO_348 (O_348,N_4606,N_4879);
xnor UO_349 (O_349,N_4657,N_4717);
or UO_350 (O_350,N_4758,N_4592);
nor UO_351 (O_351,N_4518,N_4923);
and UO_352 (O_352,N_4533,N_4807);
nor UO_353 (O_353,N_4806,N_4760);
nand UO_354 (O_354,N_4566,N_4862);
nand UO_355 (O_355,N_4576,N_4736);
or UO_356 (O_356,N_4626,N_4525);
nor UO_357 (O_357,N_4834,N_4797);
or UO_358 (O_358,N_4898,N_4601);
or UO_359 (O_359,N_4987,N_4571);
nor UO_360 (O_360,N_4629,N_4861);
nand UO_361 (O_361,N_4654,N_4741);
or UO_362 (O_362,N_4654,N_4838);
or UO_363 (O_363,N_4523,N_4694);
nand UO_364 (O_364,N_4924,N_4863);
nor UO_365 (O_365,N_4984,N_4790);
and UO_366 (O_366,N_4837,N_4740);
nand UO_367 (O_367,N_4635,N_4649);
or UO_368 (O_368,N_4761,N_4810);
or UO_369 (O_369,N_4630,N_4816);
or UO_370 (O_370,N_4791,N_4792);
and UO_371 (O_371,N_4872,N_4736);
nand UO_372 (O_372,N_4667,N_4863);
nor UO_373 (O_373,N_4549,N_4952);
and UO_374 (O_374,N_4888,N_4910);
xor UO_375 (O_375,N_4988,N_4767);
and UO_376 (O_376,N_4961,N_4747);
nor UO_377 (O_377,N_4918,N_4798);
nor UO_378 (O_378,N_4596,N_4717);
or UO_379 (O_379,N_4570,N_4535);
nand UO_380 (O_380,N_4876,N_4929);
nor UO_381 (O_381,N_4847,N_4946);
xnor UO_382 (O_382,N_4760,N_4872);
or UO_383 (O_383,N_4991,N_4883);
or UO_384 (O_384,N_4996,N_4666);
nand UO_385 (O_385,N_4587,N_4591);
and UO_386 (O_386,N_4867,N_4914);
or UO_387 (O_387,N_4938,N_4705);
and UO_388 (O_388,N_4818,N_4862);
and UO_389 (O_389,N_4721,N_4685);
nand UO_390 (O_390,N_4647,N_4605);
xor UO_391 (O_391,N_4704,N_4526);
and UO_392 (O_392,N_4962,N_4775);
nor UO_393 (O_393,N_4917,N_4834);
xnor UO_394 (O_394,N_4615,N_4792);
or UO_395 (O_395,N_4595,N_4545);
nor UO_396 (O_396,N_4933,N_4726);
or UO_397 (O_397,N_4589,N_4920);
and UO_398 (O_398,N_4675,N_4962);
nor UO_399 (O_399,N_4757,N_4603);
and UO_400 (O_400,N_4602,N_4783);
xor UO_401 (O_401,N_4727,N_4720);
nand UO_402 (O_402,N_4963,N_4931);
nor UO_403 (O_403,N_4863,N_4622);
or UO_404 (O_404,N_4714,N_4845);
and UO_405 (O_405,N_4736,N_4835);
nand UO_406 (O_406,N_4920,N_4944);
and UO_407 (O_407,N_4551,N_4680);
nand UO_408 (O_408,N_4506,N_4500);
or UO_409 (O_409,N_4699,N_4975);
or UO_410 (O_410,N_4568,N_4539);
and UO_411 (O_411,N_4700,N_4686);
nor UO_412 (O_412,N_4781,N_4571);
nand UO_413 (O_413,N_4989,N_4709);
xor UO_414 (O_414,N_4685,N_4824);
nor UO_415 (O_415,N_4866,N_4897);
nor UO_416 (O_416,N_4521,N_4733);
and UO_417 (O_417,N_4704,N_4901);
nand UO_418 (O_418,N_4576,N_4532);
nor UO_419 (O_419,N_4893,N_4631);
or UO_420 (O_420,N_4885,N_4740);
nand UO_421 (O_421,N_4667,N_4919);
or UO_422 (O_422,N_4696,N_4991);
and UO_423 (O_423,N_4903,N_4889);
and UO_424 (O_424,N_4815,N_4587);
nand UO_425 (O_425,N_4930,N_4684);
nor UO_426 (O_426,N_4622,N_4667);
nand UO_427 (O_427,N_4604,N_4974);
and UO_428 (O_428,N_4960,N_4842);
nor UO_429 (O_429,N_4838,N_4713);
or UO_430 (O_430,N_4915,N_4508);
or UO_431 (O_431,N_4809,N_4759);
nor UO_432 (O_432,N_4555,N_4510);
xor UO_433 (O_433,N_4696,N_4597);
or UO_434 (O_434,N_4865,N_4622);
or UO_435 (O_435,N_4970,N_4781);
and UO_436 (O_436,N_4834,N_4728);
and UO_437 (O_437,N_4978,N_4692);
and UO_438 (O_438,N_4509,N_4797);
or UO_439 (O_439,N_4836,N_4579);
nor UO_440 (O_440,N_4543,N_4862);
and UO_441 (O_441,N_4863,N_4662);
xor UO_442 (O_442,N_4763,N_4974);
or UO_443 (O_443,N_4997,N_4642);
or UO_444 (O_444,N_4900,N_4567);
nand UO_445 (O_445,N_4573,N_4589);
nand UO_446 (O_446,N_4841,N_4729);
and UO_447 (O_447,N_4643,N_4637);
nor UO_448 (O_448,N_4639,N_4946);
or UO_449 (O_449,N_4818,N_4592);
nand UO_450 (O_450,N_4828,N_4999);
xnor UO_451 (O_451,N_4515,N_4760);
nand UO_452 (O_452,N_4657,N_4940);
nor UO_453 (O_453,N_4635,N_4614);
or UO_454 (O_454,N_4555,N_4601);
and UO_455 (O_455,N_4676,N_4566);
nor UO_456 (O_456,N_4642,N_4778);
nor UO_457 (O_457,N_4768,N_4995);
nand UO_458 (O_458,N_4513,N_4963);
nor UO_459 (O_459,N_4938,N_4525);
nor UO_460 (O_460,N_4805,N_4707);
or UO_461 (O_461,N_4733,N_4907);
and UO_462 (O_462,N_4818,N_4839);
or UO_463 (O_463,N_4639,N_4844);
nand UO_464 (O_464,N_4732,N_4524);
and UO_465 (O_465,N_4788,N_4947);
and UO_466 (O_466,N_4981,N_4893);
nand UO_467 (O_467,N_4755,N_4595);
or UO_468 (O_468,N_4704,N_4535);
nand UO_469 (O_469,N_4934,N_4561);
or UO_470 (O_470,N_4756,N_4567);
and UO_471 (O_471,N_4875,N_4547);
nand UO_472 (O_472,N_4938,N_4634);
or UO_473 (O_473,N_4785,N_4512);
and UO_474 (O_474,N_4655,N_4899);
nor UO_475 (O_475,N_4868,N_4799);
nor UO_476 (O_476,N_4519,N_4880);
nand UO_477 (O_477,N_4567,N_4936);
nand UO_478 (O_478,N_4735,N_4894);
and UO_479 (O_479,N_4825,N_4959);
or UO_480 (O_480,N_4614,N_4514);
and UO_481 (O_481,N_4856,N_4514);
or UO_482 (O_482,N_4916,N_4646);
or UO_483 (O_483,N_4824,N_4981);
or UO_484 (O_484,N_4925,N_4697);
nor UO_485 (O_485,N_4895,N_4662);
nor UO_486 (O_486,N_4560,N_4829);
or UO_487 (O_487,N_4873,N_4915);
nand UO_488 (O_488,N_4660,N_4509);
or UO_489 (O_489,N_4544,N_4839);
nand UO_490 (O_490,N_4887,N_4902);
nor UO_491 (O_491,N_4645,N_4847);
or UO_492 (O_492,N_4720,N_4573);
or UO_493 (O_493,N_4716,N_4788);
and UO_494 (O_494,N_4834,N_4687);
xnor UO_495 (O_495,N_4608,N_4579);
and UO_496 (O_496,N_4946,N_4760);
nor UO_497 (O_497,N_4758,N_4878);
and UO_498 (O_498,N_4728,N_4590);
nand UO_499 (O_499,N_4941,N_4670);
and UO_500 (O_500,N_4948,N_4847);
nand UO_501 (O_501,N_4999,N_4742);
nand UO_502 (O_502,N_4652,N_4744);
or UO_503 (O_503,N_4855,N_4712);
or UO_504 (O_504,N_4552,N_4831);
nand UO_505 (O_505,N_4575,N_4506);
or UO_506 (O_506,N_4887,N_4699);
nand UO_507 (O_507,N_4664,N_4752);
nand UO_508 (O_508,N_4921,N_4513);
nand UO_509 (O_509,N_4664,N_4950);
and UO_510 (O_510,N_4505,N_4631);
or UO_511 (O_511,N_4623,N_4792);
nor UO_512 (O_512,N_4771,N_4921);
nand UO_513 (O_513,N_4502,N_4825);
nand UO_514 (O_514,N_4727,N_4608);
and UO_515 (O_515,N_4942,N_4752);
xor UO_516 (O_516,N_4726,N_4685);
or UO_517 (O_517,N_4930,N_4548);
and UO_518 (O_518,N_4752,N_4529);
nor UO_519 (O_519,N_4627,N_4599);
nand UO_520 (O_520,N_4804,N_4518);
and UO_521 (O_521,N_4560,N_4982);
nand UO_522 (O_522,N_4778,N_4761);
or UO_523 (O_523,N_4946,N_4794);
or UO_524 (O_524,N_4761,N_4842);
nor UO_525 (O_525,N_4795,N_4796);
and UO_526 (O_526,N_4746,N_4981);
and UO_527 (O_527,N_4539,N_4859);
nand UO_528 (O_528,N_4963,N_4549);
or UO_529 (O_529,N_4895,N_4780);
nand UO_530 (O_530,N_4735,N_4800);
or UO_531 (O_531,N_4622,N_4950);
nor UO_532 (O_532,N_4823,N_4673);
nand UO_533 (O_533,N_4532,N_4607);
and UO_534 (O_534,N_4867,N_4656);
and UO_535 (O_535,N_4599,N_4573);
xor UO_536 (O_536,N_4764,N_4831);
xnor UO_537 (O_537,N_4529,N_4563);
nor UO_538 (O_538,N_4651,N_4816);
and UO_539 (O_539,N_4962,N_4696);
xnor UO_540 (O_540,N_4711,N_4739);
nor UO_541 (O_541,N_4512,N_4707);
xor UO_542 (O_542,N_4540,N_4501);
or UO_543 (O_543,N_4840,N_4742);
and UO_544 (O_544,N_4661,N_4543);
nor UO_545 (O_545,N_4645,N_4821);
or UO_546 (O_546,N_4668,N_4591);
and UO_547 (O_547,N_4611,N_4888);
nand UO_548 (O_548,N_4513,N_4955);
nand UO_549 (O_549,N_4585,N_4793);
nand UO_550 (O_550,N_4935,N_4504);
and UO_551 (O_551,N_4663,N_4666);
or UO_552 (O_552,N_4586,N_4736);
nor UO_553 (O_553,N_4809,N_4575);
nor UO_554 (O_554,N_4686,N_4919);
nand UO_555 (O_555,N_4973,N_4876);
nor UO_556 (O_556,N_4622,N_4901);
nand UO_557 (O_557,N_4841,N_4853);
or UO_558 (O_558,N_4522,N_4645);
or UO_559 (O_559,N_4769,N_4753);
and UO_560 (O_560,N_4509,N_4559);
or UO_561 (O_561,N_4638,N_4648);
nand UO_562 (O_562,N_4960,N_4765);
nand UO_563 (O_563,N_4852,N_4835);
nand UO_564 (O_564,N_4960,N_4774);
or UO_565 (O_565,N_4687,N_4910);
and UO_566 (O_566,N_4546,N_4614);
or UO_567 (O_567,N_4925,N_4689);
and UO_568 (O_568,N_4999,N_4518);
nand UO_569 (O_569,N_4921,N_4854);
and UO_570 (O_570,N_4700,N_4918);
and UO_571 (O_571,N_4935,N_4622);
or UO_572 (O_572,N_4983,N_4621);
nand UO_573 (O_573,N_4901,N_4990);
nor UO_574 (O_574,N_4932,N_4712);
or UO_575 (O_575,N_4623,N_4640);
nor UO_576 (O_576,N_4801,N_4533);
nor UO_577 (O_577,N_4625,N_4593);
nand UO_578 (O_578,N_4509,N_4567);
or UO_579 (O_579,N_4752,N_4585);
nand UO_580 (O_580,N_4979,N_4936);
or UO_581 (O_581,N_4808,N_4733);
nand UO_582 (O_582,N_4648,N_4662);
or UO_583 (O_583,N_4570,N_4694);
nand UO_584 (O_584,N_4819,N_4987);
nand UO_585 (O_585,N_4769,N_4521);
and UO_586 (O_586,N_4964,N_4939);
or UO_587 (O_587,N_4818,N_4777);
nand UO_588 (O_588,N_4814,N_4798);
or UO_589 (O_589,N_4902,N_4950);
nor UO_590 (O_590,N_4511,N_4502);
and UO_591 (O_591,N_4875,N_4970);
nor UO_592 (O_592,N_4516,N_4595);
or UO_593 (O_593,N_4727,N_4822);
and UO_594 (O_594,N_4720,N_4636);
nor UO_595 (O_595,N_4529,N_4703);
and UO_596 (O_596,N_4807,N_4875);
nand UO_597 (O_597,N_4619,N_4867);
xnor UO_598 (O_598,N_4925,N_4596);
or UO_599 (O_599,N_4688,N_4537);
nor UO_600 (O_600,N_4817,N_4909);
nand UO_601 (O_601,N_4650,N_4995);
and UO_602 (O_602,N_4623,N_4530);
nand UO_603 (O_603,N_4771,N_4663);
nor UO_604 (O_604,N_4661,N_4778);
nand UO_605 (O_605,N_4521,N_4836);
nor UO_606 (O_606,N_4793,N_4822);
nor UO_607 (O_607,N_4954,N_4768);
nand UO_608 (O_608,N_4669,N_4615);
or UO_609 (O_609,N_4940,N_4798);
or UO_610 (O_610,N_4663,N_4853);
and UO_611 (O_611,N_4778,N_4540);
nand UO_612 (O_612,N_4944,N_4657);
nand UO_613 (O_613,N_4663,N_4800);
nand UO_614 (O_614,N_4938,N_4927);
nor UO_615 (O_615,N_4959,N_4969);
nor UO_616 (O_616,N_4551,N_4945);
and UO_617 (O_617,N_4711,N_4669);
or UO_618 (O_618,N_4874,N_4581);
nand UO_619 (O_619,N_4828,N_4776);
xnor UO_620 (O_620,N_4614,N_4963);
xnor UO_621 (O_621,N_4574,N_4700);
nor UO_622 (O_622,N_4889,N_4791);
or UO_623 (O_623,N_4820,N_4722);
or UO_624 (O_624,N_4687,N_4949);
nor UO_625 (O_625,N_4752,N_4559);
or UO_626 (O_626,N_4863,N_4590);
xor UO_627 (O_627,N_4787,N_4530);
nand UO_628 (O_628,N_4833,N_4759);
or UO_629 (O_629,N_4814,N_4819);
nand UO_630 (O_630,N_4969,N_4532);
or UO_631 (O_631,N_4729,N_4611);
or UO_632 (O_632,N_4531,N_4775);
xnor UO_633 (O_633,N_4633,N_4764);
or UO_634 (O_634,N_4994,N_4631);
and UO_635 (O_635,N_4681,N_4559);
nor UO_636 (O_636,N_4950,N_4627);
nor UO_637 (O_637,N_4989,N_4514);
nor UO_638 (O_638,N_4893,N_4501);
or UO_639 (O_639,N_4831,N_4793);
or UO_640 (O_640,N_4844,N_4630);
xnor UO_641 (O_641,N_4844,N_4682);
nor UO_642 (O_642,N_4871,N_4915);
nor UO_643 (O_643,N_4636,N_4645);
xnor UO_644 (O_644,N_4678,N_4535);
nand UO_645 (O_645,N_4627,N_4908);
nor UO_646 (O_646,N_4805,N_4538);
xnor UO_647 (O_647,N_4893,N_4846);
and UO_648 (O_648,N_4544,N_4883);
and UO_649 (O_649,N_4840,N_4690);
or UO_650 (O_650,N_4955,N_4580);
nand UO_651 (O_651,N_4668,N_4735);
nand UO_652 (O_652,N_4754,N_4875);
and UO_653 (O_653,N_4610,N_4571);
or UO_654 (O_654,N_4798,N_4653);
nand UO_655 (O_655,N_4703,N_4893);
nand UO_656 (O_656,N_4716,N_4620);
xor UO_657 (O_657,N_4934,N_4665);
or UO_658 (O_658,N_4917,N_4833);
and UO_659 (O_659,N_4872,N_4707);
nand UO_660 (O_660,N_4606,N_4506);
nor UO_661 (O_661,N_4988,N_4522);
or UO_662 (O_662,N_4663,N_4968);
nor UO_663 (O_663,N_4954,N_4587);
nand UO_664 (O_664,N_4766,N_4863);
nand UO_665 (O_665,N_4924,N_4521);
and UO_666 (O_666,N_4910,N_4742);
and UO_667 (O_667,N_4699,N_4819);
or UO_668 (O_668,N_4574,N_4878);
nor UO_669 (O_669,N_4726,N_4521);
or UO_670 (O_670,N_4996,N_4998);
or UO_671 (O_671,N_4510,N_4724);
or UO_672 (O_672,N_4676,N_4582);
nand UO_673 (O_673,N_4821,N_4784);
nand UO_674 (O_674,N_4737,N_4540);
nand UO_675 (O_675,N_4599,N_4622);
or UO_676 (O_676,N_4940,N_4946);
nor UO_677 (O_677,N_4719,N_4639);
and UO_678 (O_678,N_4869,N_4925);
and UO_679 (O_679,N_4504,N_4602);
or UO_680 (O_680,N_4622,N_4859);
or UO_681 (O_681,N_4920,N_4845);
nand UO_682 (O_682,N_4653,N_4881);
or UO_683 (O_683,N_4908,N_4959);
nand UO_684 (O_684,N_4807,N_4639);
xor UO_685 (O_685,N_4911,N_4923);
nand UO_686 (O_686,N_4877,N_4790);
or UO_687 (O_687,N_4534,N_4805);
or UO_688 (O_688,N_4619,N_4884);
or UO_689 (O_689,N_4873,N_4616);
nand UO_690 (O_690,N_4760,N_4706);
or UO_691 (O_691,N_4731,N_4703);
or UO_692 (O_692,N_4706,N_4651);
nand UO_693 (O_693,N_4781,N_4501);
and UO_694 (O_694,N_4712,N_4801);
nand UO_695 (O_695,N_4741,N_4603);
nor UO_696 (O_696,N_4697,N_4618);
or UO_697 (O_697,N_4763,N_4588);
xor UO_698 (O_698,N_4575,N_4598);
nand UO_699 (O_699,N_4529,N_4680);
or UO_700 (O_700,N_4728,N_4668);
and UO_701 (O_701,N_4850,N_4967);
nor UO_702 (O_702,N_4750,N_4645);
xnor UO_703 (O_703,N_4709,N_4710);
nand UO_704 (O_704,N_4543,N_4863);
nand UO_705 (O_705,N_4962,N_4843);
nand UO_706 (O_706,N_4778,N_4968);
nand UO_707 (O_707,N_4850,N_4979);
nand UO_708 (O_708,N_4695,N_4619);
xnor UO_709 (O_709,N_4790,N_4595);
nand UO_710 (O_710,N_4557,N_4683);
nor UO_711 (O_711,N_4806,N_4961);
nand UO_712 (O_712,N_4857,N_4820);
nor UO_713 (O_713,N_4523,N_4643);
nand UO_714 (O_714,N_4662,N_4782);
nor UO_715 (O_715,N_4832,N_4669);
and UO_716 (O_716,N_4737,N_4866);
and UO_717 (O_717,N_4590,N_4552);
nand UO_718 (O_718,N_4876,N_4861);
and UO_719 (O_719,N_4696,N_4899);
and UO_720 (O_720,N_4745,N_4507);
nand UO_721 (O_721,N_4934,N_4674);
and UO_722 (O_722,N_4661,N_4577);
and UO_723 (O_723,N_4539,N_4601);
or UO_724 (O_724,N_4728,N_4633);
xor UO_725 (O_725,N_4917,N_4604);
xnor UO_726 (O_726,N_4941,N_4547);
nand UO_727 (O_727,N_4791,N_4613);
or UO_728 (O_728,N_4508,N_4581);
nand UO_729 (O_729,N_4799,N_4649);
nand UO_730 (O_730,N_4761,N_4734);
nand UO_731 (O_731,N_4979,N_4734);
nand UO_732 (O_732,N_4908,N_4886);
nand UO_733 (O_733,N_4639,N_4584);
nand UO_734 (O_734,N_4698,N_4535);
nand UO_735 (O_735,N_4676,N_4797);
nand UO_736 (O_736,N_4854,N_4688);
or UO_737 (O_737,N_4652,N_4630);
or UO_738 (O_738,N_4732,N_4671);
and UO_739 (O_739,N_4845,N_4582);
nor UO_740 (O_740,N_4787,N_4733);
nor UO_741 (O_741,N_4838,N_4657);
nand UO_742 (O_742,N_4820,N_4992);
nor UO_743 (O_743,N_4736,N_4625);
or UO_744 (O_744,N_4655,N_4987);
or UO_745 (O_745,N_4781,N_4897);
nor UO_746 (O_746,N_4957,N_4608);
or UO_747 (O_747,N_4717,N_4892);
nor UO_748 (O_748,N_4571,N_4662);
nor UO_749 (O_749,N_4752,N_4765);
nand UO_750 (O_750,N_4681,N_4705);
nand UO_751 (O_751,N_4768,N_4640);
and UO_752 (O_752,N_4905,N_4964);
nand UO_753 (O_753,N_4583,N_4557);
nor UO_754 (O_754,N_4503,N_4880);
nand UO_755 (O_755,N_4762,N_4582);
and UO_756 (O_756,N_4546,N_4550);
or UO_757 (O_757,N_4789,N_4740);
or UO_758 (O_758,N_4642,N_4509);
nand UO_759 (O_759,N_4541,N_4875);
nor UO_760 (O_760,N_4897,N_4630);
and UO_761 (O_761,N_4509,N_4825);
nor UO_762 (O_762,N_4710,N_4581);
nor UO_763 (O_763,N_4820,N_4520);
and UO_764 (O_764,N_4747,N_4933);
xnor UO_765 (O_765,N_4889,N_4861);
and UO_766 (O_766,N_4747,N_4764);
and UO_767 (O_767,N_4723,N_4502);
or UO_768 (O_768,N_4533,N_4795);
nand UO_769 (O_769,N_4965,N_4554);
nor UO_770 (O_770,N_4724,N_4808);
and UO_771 (O_771,N_4775,N_4932);
nor UO_772 (O_772,N_4602,N_4722);
nand UO_773 (O_773,N_4587,N_4694);
nand UO_774 (O_774,N_4680,N_4740);
nand UO_775 (O_775,N_4859,N_4861);
or UO_776 (O_776,N_4841,N_4893);
or UO_777 (O_777,N_4519,N_4827);
nand UO_778 (O_778,N_4767,N_4561);
xnor UO_779 (O_779,N_4868,N_4852);
nor UO_780 (O_780,N_4998,N_4884);
and UO_781 (O_781,N_4894,N_4709);
nor UO_782 (O_782,N_4697,N_4559);
nor UO_783 (O_783,N_4667,N_4658);
nand UO_784 (O_784,N_4898,N_4979);
nand UO_785 (O_785,N_4728,N_4956);
nor UO_786 (O_786,N_4789,N_4504);
and UO_787 (O_787,N_4677,N_4574);
nand UO_788 (O_788,N_4715,N_4739);
nand UO_789 (O_789,N_4980,N_4929);
nand UO_790 (O_790,N_4785,N_4807);
nor UO_791 (O_791,N_4752,N_4855);
nand UO_792 (O_792,N_4527,N_4621);
nor UO_793 (O_793,N_4798,N_4530);
nand UO_794 (O_794,N_4747,N_4578);
nor UO_795 (O_795,N_4768,N_4731);
nand UO_796 (O_796,N_4691,N_4944);
and UO_797 (O_797,N_4665,N_4761);
nor UO_798 (O_798,N_4544,N_4873);
nor UO_799 (O_799,N_4877,N_4832);
and UO_800 (O_800,N_4937,N_4505);
nand UO_801 (O_801,N_4894,N_4715);
or UO_802 (O_802,N_4868,N_4782);
and UO_803 (O_803,N_4871,N_4875);
and UO_804 (O_804,N_4746,N_4627);
nor UO_805 (O_805,N_4947,N_4639);
xor UO_806 (O_806,N_4946,N_4594);
xnor UO_807 (O_807,N_4916,N_4716);
nor UO_808 (O_808,N_4902,N_4841);
and UO_809 (O_809,N_4860,N_4698);
and UO_810 (O_810,N_4655,N_4805);
xnor UO_811 (O_811,N_4632,N_4739);
and UO_812 (O_812,N_4707,N_4566);
or UO_813 (O_813,N_4871,N_4587);
nand UO_814 (O_814,N_4792,N_4815);
xor UO_815 (O_815,N_4742,N_4717);
or UO_816 (O_816,N_4935,N_4661);
nor UO_817 (O_817,N_4722,N_4567);
nor UO_818 (O_818,N_4537,N_4728);
and UO_819 (O_819,N_4544,N_4644);
or UO_820 (O_820,N_4889,N_4621);
nand UO_821 (O_821,N_4756,N_4641);
and UO_822 (O_822,N_4980,N_4988);
xnor UO_823 (O_823,N_4699,N_4584);
nor UO_824 (O_824,N_4897,N_4922);
or UO_825 (O_825,N_4552,N_4704);
nand UO_826 (O_826,N_4729,N_4556);
nor UO_827 (O_827,N_4554,N_4783);
or UO_828 (O_828,N_4524,N_4875);
or UO_829 (O_829,N_4818,N_4889);
and UO_830 (O_830,N_4609,N_4520);
nand UO_831 (O_831,N_4920,N_4568);
nand UO_832 (O_832,N_4795,N_4516);
and UO_833 (O_833,N_4899,N_4949);
nand UO_834 (O_834,N_4815,N_4675);
nor UO_835 (O_835,N_4884,N_4900);
nor UO_836 (O_836,N_4924,N_4710);
nand UO_837 (O_837,N_4533,N_4703);
nand UO_838 (O_838,N_4655,N_4809);
xnor UO_839 (O_839,N_4707,N_4646);
and UO_840 (O_840,N_4871,N_4849);
or UO_841 (O_841,N_4720,N_4906);
nor UO_842 (O_842,N_4773,N_4590);
nand UO_843 (O_843,N_4545,N_4505);
or UO_844 (O_844,N_4577,N_4574);
nand UO_845 (O_845,N_4602,N_4716);
and UO_846 (O_846,N_4504,N_4856);
or UO_847 (O_847,N_4800,N_4991);
or UO_848 (O_848,N_4831,N_4878);
nor UO_849 (O_849,N_4794,N_4544);
or UO_850 (O_850,N_4883,N_4861);
or UO_851 (O_851,N_4958,N_4948);
or UO_852 (O_852,N_4808,N_4935);
nand UO_853 (O_853,N_4726,N_4858);
nand UO_854 (O_854,N_4586,N_4989);
and UO_855 (O_855,N_4748,N_4705);
or UO_856 (O_856,N_4835,N_4934);
and UO_857 (O_857,N_4938,N_4741);
xnor UO_858 (O_858,N_4941,N_4922);
or UO_859 (O_859,N_4699,N_4646);
nand UO_860 (O_860,N_4901,N_4797);
and UO_861 (O_861,N_4868,N_4828);
nand UO_862 (O_862,N_4808,N_4985);
and UO_863 (O_863,N_4906,N_4573);
nand UO_864 (O_864,N_4557,N_4879);
nand UO_865 (O_865,N_4748,N_4976);
or UO_866 (O_866,N_4771,N_4970);
or UO_867 (O_867,N_4911,N_4692);
nor UO_868 (O_868,N_4584,N_4619);
and UO_869 (O_869,N_4742,N_4507);
nor UO_870 (O_870,N_4940,N_4873);
and UO_871 (O_871,N_4952,N_4873);
and UO_872 (O_872,N_4860,N_4938);
nor UO_873 (O_873,N_4705,N_4920);
xnor UO_874 (O_874,N_4656,N_4593);
or UO_875 (O_875,N_4522,N_4903);
nor UO_876 (O_876,N_4666,N_4768);
nor UO_877 (O_877,N_4748,N_4656);
or UO_878 (O_878,N_4957,N_4651);
and UO_879 (O_879,N_4603,N_4959);
nand UO_880 (O_880,N_4566,N_4786);
xnor UO_881 (O_881,N_4742,N_4696);
nand UO_882 (O_882,N_4606,N_4819);
and UO_883 (O_883,N_4506,N_4634);
and UO_884 (O_884,N_4643,N_4741);
nor UO_885 (O_885,N_4745,N_4638);
nand UO_886 (O_886,N_4518,N_4608);
nor UO_887 (O_887,N_4648,N_4615);
nor UO_888 (O_888,N_4731,N_4702);
and UO_889 (O_889,N_4575,N_4782);
nor UO_890 (O_890,N_4641,N_4549);
or UO_891 (O_891,N_4917,N_4809);
nand UO_892 (O_892,N_4703,N_4925);
nor UO_893 (O_893,N_4522,N_4614);
or UO_894 (O_894,N_4847,N_4995);
nand UO_895 (O_895,N_4551,N_4976);
nand UO_896 (O_896,N_4896,N_4910);
nand UO_897 (O_897,N_4591,N_4801);
xor UO_898 (O_898,N_4724,N_4803);
xor UO_899 (O_899,N_4625,N_4967);
nor UO_900 (O_900,N_4547,N_4870);
nand UO_901 (O_901,N_4559,N_4746);
nor UO_902 (O_902,N_4801,N_4521);
xnor UO_903 (O_903,N_4636,N_4935);
or UO_904 (O_904,N_4646,N_4908);
or UO_905 (O_905,N_4906,N_4972);
nand UO_906 (O_906,N_4555,N_4607);
and UO_907 (O_907,N_4775,N_4897);
nand UO_908 (O_908,N_4990,N_4708);
xnor UO_909 (O_909,N_4859,N_4987);
or UO_910 (O_910,N_4630,N_4952);
nor UO_911 (O_911,N_4845,N_4902);
nor UO_912 (O_912,N_4690,N_4862);
and UO_913 (O_913,N_4588,N_4923);
nand UO_914 (O_914,N_4602,N_4618);
or UO_915 (O_915,N_4771,N_4525);
xnor UO_916 (O_916,N_4918,N_4799);
nand UO_917 (O_917,N_4680,N_4561);
and UO_918 (O_918,N_4924,N_4571);
nor UO_919 (O_919,N_4568,N_4676);
nor UO_920 (O_920,N_4992,N_4712);
nand UO_921 (O_921,N_4739,N_4714);
nand UO_922 (O_922,N_4598,N_4527);
or UO_923 (O_923,N_4959,N_4955);
or UO_924 (O_924,N_4692,N_4681);
or UO_925 (O_925,N_4908,N_4656);
nor UO_926 (O_926,N_4763,N_4732);
nor UO_927 (O_927,N_4861,N_4960);
xor UO_928 (O_928,N_4502,N_4982);
or UO_929 (O_929,N_4900,N_4506);
or UO_930 (O_930,N_4578,N_4776);
and UO_931 (O_931,N_4804,N_4693);
nand UO_932 (O_932,N_4639,N_4538);
or UO_933 (O_933,N_4673,N_4549);
or UO_934 (O_934,N_4986,N_4533);
or UO_935 (O_935,N_4990,N_4738);
or UO_936 (O_936,N_4796,N_4606);
nand UO_937 (O_937,N_4770,N_4500);
nor UO_938 (O_938,N_4969,N_4556);
nor UO_939 (O_939,N_4910,N_4895);
and UO_940 (O_940,N_4943,N_4680);
nor UO_941 (O_941,N_4935,N_4800);
or UO_942 (O_942,N_4694,N_4568);
and UO_943 (O_943,N_4533,N_4786);
or UO_944 (O_944,N_4689,N_4535);
nor UO_945 (O_945,N_4752,N_4971);
or UO_946 (O_946,N_4692,N_4977);
nor UO_947 (O_947,N_4579,N_4907);
nand UO_948 (O_948,N_4970,N_4761);
nand UO_949 (O_949,N_4894,N_4746);
nor UO_950 (O_950,N_4923,N_4661);
and UO_951 (O_951,N_4899,N_4730);
nand UO_952 (O_952,N_4729,N_4717);
and UO_953 (O_953,N_4527,N_4657);
nand UO_954 (O_954,N_4714,N_4992);
or UO_955 (O_955,N_4778,N_4754);
nand UO_956 (O_956,N_4982,N_4890);
nor UO_957 (O_957,N_4870,N_4593);
and UO_958 (O_958,N_4653,N_4765);
or UO_959 (O_959,N_4555,N_4880);
and UO_960 (O_960,N_4651,N_4705);
nor UO_961 (O_961,N_4888,N_4635);
or UO_962 (O_962,N_4810,N_4621);
or UO_963 (O_963,N_4815,N_4904);
nand UO_964 (O_964,N_4872,N_4721);
nand UO_965 (O_965,N_4956,N_4891);
and UO_966 (O_966,N_4898,N_4982);
or UO_967 (O_967,N_4514,N_4985);
xor UO_968 (O_968,N_4890,N_4664);
or UO_969 (O_969,N_4565,N_4621);
nand UO_970 (O_970,N_4590,N_4970);
and UO_971 (O_971,N_4840,N_4787);
xnor UO_972 (O_972,N_4913,N_4789);
nand UO_973 (O_973,N_4563,N_4963);
nor UO_974 (O_974,N_4824,N_4817);
nor UO_975 (O_975,N_4847,N_4775);
nand UO_976 (O_976,N_4931,N_4725);
or UO_977 (O_977,N_4684,N_4844);
and UO_978 (O_978,N_4688,N_4825);
nor UO_979 (O_979,N_4693,N_4699);
or UO_980 (O_980,N_4617,N_4604);
and UO_981 (O_981,N_4685,N_4604);
nor UO_982 (O_982,N_4768,N_4966);
or UO_983 (O_983,N_4819,N_4874);
nand UO_984 (O_984,N_4580,N_4995);
nand UO_985 (O_985,N_4648,N_4749);
and UO_986 (O_986,N_4935,N_4785);
xnor UO_987 (O_987,N_4548,N_4737);
and UO_988 (O_988,N_4782,N_4690);
nor UO_989 (O_989,N_4894,N_4674);
or UO_990 (O_990,N_4993,N_4761);
nor UO_991 (O_991,N_4547,N_4774);
and UO_992 (O_992,N_4751,N_4634);
nand UO_993 (O_993,N_4656,N_4835);
nor UO_994 (O_994,N_4566,N_4925);
xnor UO_995 (O_995,N_4868,N_4945);
or UO_996 (O_996,N_4620,N_4841);
nor UO_997 (O_997,N_4871,N_4531);
or UO_998 (O_998,N_4800,N_4525);
nand UO_999 (O_999,N_4711,N_4866);
endmodule